// Benchmark "adder" written by ABC on Wed Jul 13 18:48:41 2022

module adder ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] ,
    \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] ,
    \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] ,
    \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] ,
    \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] ,
    \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] ,
    \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] , \b[60] ,
    \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] , \b[68] ,
    \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] , \b[76] ,
    \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] , \b[84] ,
    \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] ,
    \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127] , cOut  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] ,
    \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] ,
    \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] ,
    \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] ,
    \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] ,
    \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] ,
    \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] ,
    \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] ,
    \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] ,
    \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] ,
    \b[76] , \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] ,
    \b[84] , \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] ,
    \b[92] , \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] , cOut;
  wire new_new_n386__, new_new_n387__, new_new_n389__, new_new_n390__,
    new_new_n391__, new_new_n392__, new_new_n393__, new_new_n395__,
    new_new_n396__, new_new_n397__, new_new_n398__, new_new_n399__,
    new_new_n400__, new_new_n401__, new_new_n403__, new_new_n404__,
    new_new_n405__, new_new_n406__, new_new_n407__, new_new_n408__,
    new_new_n409__, new_new_n411__, new_new_n412__, new_new_n413__,
    new_new_n414__, new_new_n415__, new_new_n416__, new_new_n417__,
    new_new_n419__, new_new_n420__, new_new_n421__, new_new_n422__,
    new_new_n423__, new_new_n424__, new_new_n425__, new_new_n427__,
    new_new_n428__, new_new_n429__, new_new_n430__, new_new_n431__,
    new_new_n432__, new_new_n433__, new_new_n435__, new_new_n436__,
    new_new_n437__, new_new_n438__, new_new_n439__, new_new_n440__,
    new_new_n441__, new_new_n443__, new_new_n444__, new_new_n445__,
    new_new_n446__, new_new_n447__, new_new_n448__, new_new_n449__,
    new_new_n451__, new_new_n452__, new_new_n453__, new_new_n454__,
    new_new_n455__, new_new_n456__, new_new_n457__, new_new_n459__,
    new_new_n460__, new_new_n461__, new_new_n462__, new_new_n463__,
    new_new_n464__, new_new_n465__, new_new_n467__, new_new_n468__,
    new_new_n469__, new_new_n470__, new_new_n471__, new_new_n472__,
    new_new_n473__, new_new_n475__, new_new_n476__, new_new_n477__,
    new_new_n478__, new_new_n479__, new_new_n480__, new_new_n481__,
    new_new_n483__, new_new_n484__, new_new_n485__, new_new_n486__,
    new_new_n487__, new_new_n488__, new_new_n489__, new_new_n491__,
    new_new_n492__, new_new_n493__, new_new_n494__, new_new_n495__,
    new_new_n496__, new_new_n497__, new_new_n499__, new_new_n500__,
    new_new_n501__, new_new_n502__, new_new_n503__, new_new_n504__,
    new_new_n505__, new_new_n507__, new_new_n508__, new_new_n509__,
    new_new_n510__, new_new_n511__, new_new_n512__, new_new_n513__,
    new_new_n515__, new_new_n516__, new_new_n517__, new_new_n518__,
    new_new_n519__, new_new_n520__, new_new_n521__, new_new_n523__,
    new_new_n524__, new_new_n525__, new_new_n526__, new_new_n527__,
    new_new_n528__, new_new_n529__, new_new_n531__, new_new_n532__,
    new_new_n533__, new_new_n534__, new_new_n535__, new_new_n536__,
    new_new_n537__, new_new_n539__, new_new_n540__, new_new_n541__,
    new_new_n542__, new_new_n543__, new_new_n544__, new_new_n545__,
    new_new_n547__, new_new_n548__, new_new_n549__, new_new_n550__,
    new_new_n551__, new_new_n552__, new_new_n553__, new_new_n555__,
    new_new_n556__, new_new_n557__, new_new_n558__, new_new_n559__,
    new_new_n560__, new_new_n561__, new_new_n563__, new_new_n564__,
    new_new_n565__, new_new_n566__, new_new_n567__, new_new_n568__,
    new_new_n569__, new_new_n571__, new_new_n572__, new_new_n573__,
    new_new_n574__, new_new_n575__, new_new_n576__, new_new_n577__,
    new_new_n579__, new_new_n580__, new_new_n581__, new_new_n582__,
    new_new_n583__, new_new_n584__, new_new_n585__, new_new_n587__,
    new_new_n588__, new_new_n589__, new_new_n590__, new_new_n591__,
    new_new_n592__, new_new_n593__, new_new_n595__, new_new_n596__,
    new_new_n597__, new_new_n598__, new_new_n599__, new_new_n600__,
    new_new_n601__, new_new_n603__, new_new_n604__, new_new_n605__,
    new_new_n606__, new_new_n607__, new_new_n608__, new_new_n609__,
    new_new_n611__, new_new_n612__, new_new_n613__, new_new_n614__,
    new_new_n615__, new_new_n616__, new_new_n617__, new_new_n619__,
    new_new_n620__, new_new_n621__, new_new_n622__, new_new_n623__,
    new_new_n624__, new_new_n625__, new_new_n627__, new_new_n628__,
    new_new_n629__, new_new_n630__, new_new_n631__, new_new_n632__,
    new_new_n633__, new_new_n635__, new_new_n636__, new_new_n637__,
    new_new_n638__, new_new_n639__, new_new_n640__, new_new_n641__,
    new_new_n643__, new_new_n644__, new_new_n645__, new_new_n646__,
    new_new_n647__, new_new_n648__, new_new_n649__, new_new_n651__,
    new_new_n652__, new_new_n653__, new_new_n654__, new_new_n655__,
    new_new_n656__, new_new_n657__, new_new_n659__, new_new_n660__,
    new_new_n661__, new_new_n662__, new_new_n663__, new_new_n664__,
    new_new_n665__, new_new_n667__, new_new_n668__, new_new_n669__,
    new_new_n670__, new_new_n671__, new_new_n672__, new_new_n673__,
    new_new_n675__, new_new_n676__, new_new_n677__, new_new_n678__,
    new_new_n679__, new_new_n680__, new_new_n681__, new_new_n683__,
    new_new_n684__, new_new_n685__, new_new_n686__, new_new_n687__,
    new_new_n688__, new_new_n689__, new_new_n691__, new_new_n692__,
    new_new_n693__, new_new_n694__, new_new_n695__, new_new_n696__,
    new_new_n697__, new_new_n699__, new_new_n700__, new_new_n701__,
    new_new_n702__, new_new_n703__, new_new_n704__, new_new_n705__,
    new_new_n707__, new_new_n708__, new_new_n709__, new_new_n710__,
    new_new_n711__, new_new_n712__, new_new_n713__, new_new_n715__,
    new_new_n716__, new_new_n717__, new_new_n718__, new_new_n719__,
    new_new_n720__, new_new_n721__, new_new_n723__, new_new_n724__,
    new_new_n725__, new_new_n726__, new_new_n727__, new_new_n728__,
    new_new_n729__, new_new_n731__, new_new_n732__, new_new_n733__,
    new_new_n734__, new_new_n735__, new_new_n736__, new_new_n737__,
    new_new_n739__, new_new_n740__, new_new_n741__, new_new_n742__,
    new_new_n743__, new_new_n744__, new_new_n745__, new_new_n747__,
    new_new_n748__, new_new_n749__, new_new_n750__, new_new_n751__,
    new_new_n752__, new_new_n753__, new_new_n755__, new_new_n756__,
    new_new_n757__, new_new_n758__, new_new_n759__, new_new_n760__,
    new_new_n761__, new_new_n763__, new_new_n764__, new_new_n765__,
    new_new_n766__, new_new_n767__, new_new_n768__, new_new_n769__,
    new_new_n771__, new_new_n772__, new_new_n773__, new_new_n774__,
    new_new_n775__, new_new_n776__, new_new_n777__, new_new_n779__,
    new_new_n780__, new_new_n781__, new_new_n782__, new_new_n783__,
    new_new_n784__, new_new_n785__, new_new_n787__, new_new_n788__,
    new_new_n789__, new_new_n790__, new_new_n791__, new_new_n792__,
    new_new_n793__, new_new_n795__, new_new_n796__, new_new_n797__,
    new_new_n798__, new_new_n799__, new_new_n800__, new_new_n801__,
    new_new_n803__, new_new_n804__, new_new_n805__, new_new_n806__,
    new_new_n807__, new_new_n808__, new_new_n809__, new_new_n811__,
    new_new_n812__, new_new_n813__, new_new_n814__, new_new_n815__,
    new_new_n816__, new_new_n817__, new_new_n819__, new_new_n820__,
    new_new_n821__, new_new_n822__, new_new_n823__, new_new_n824__,
    new_new_n825__, new_new_n827__, new_new_n828__, new_new_n829__,
    new_new_n830__, new_new_n831__, new_new_n832__, new_new_n833__,
    new_new_n835__, new_new_n836__, new_new_n837__, new_new_n838__,
    new_new_n839__, new_new_n840__, new_new_n841__, new_new_n843__,
    new_new_n844__, new_new_n845__, new_new_n846__, new_new_n847__,
    new_new_n848__, new_new_n849__, new_new_n851__, new_new_n852__,
    new_new_n853__, new_new_n854__, new_new_n855__, new_new_n856__,
    new_new_n857__, new_new_n859__, new_new_n860__, new_new_n861__,
    new_new_n862__, new_new_n863__, new_new_n864__, new_new_n865__,
    new_new_n867__, new_new_n868__, new_new_n869__, new_new_n870__,
    new_new_n871__, new_new_n872__, new_new_n873__, new_new_n875__,
    new_new_n876__, new_new_n877__, new_new_n878__, new_new_n879__,
    new_new_n880__, new_new_n881__, new_new_n883__, new_new_n884__,
    new_new_n885__, new_new_n886__, new_new_n887__, new_new_n888__,
    new_new_n889__, new_new_n891__, new_new_n892__, new_new_n893__,
    new_new_n894__, new_new_n895__, new_new_n896__, new_new_n897__,
    new_new_n899__, new_new_n900__, new_new_n901__, new_new_n902__,
    new_new_n903__, new_new_n904__, new_new_n905__, new_new_n907__,
    new_new_n908__, new_new_n909__, new_new_n910__, new_new_n911__,
    new_new_n912__, new_new_n913__, new_new_n915__, new_new_n916__,
    new_new_n917__, new_new_n918__, new_new_n919__, new_new_n920__,
    new_new_n921__, new_new_n923__, new_new_n924__, new_new_n925__,
    new_new_n926__, new_new_n927__, new_new_n928__, new_new_n929__,
    new_new_n931__, new_new_n932__, new_new_n933__, new_new_n934__,
    new_new_n935__, new_new_n936__, new_new_n937__, new_new_n939__,
    new_new_n940__, new_new_n941__, new_new_n942__, new_new_n943__,
    new_new_n944__, new_new_n945__, new_new_n947__, new_new_n948__,
    new_new_n949__, new_new_n950__, new_new_n951__, new_new_n952__,
    new_new_n953__, new_new_n955__, new_new_n956__, new_new_n957__,
    new_new_n958__, new_new_n959__, new_new_n960__, new_new_n961__,
    new_new_n963__, new_new_n964__, new_new_n965__, new_new_n966__,
    new_new_n967__, new_new_n968__, new_new_n969__, new_new_n971__,
    new_new_n972__, new_new_n973__, new_new_n974__, new_new_n975__,
    new_new_n976__, new_new_n977__, new_new_n979__, new_new_n980__,
    new_new_n981__, new_new_n982__, new_new_n983__, new_new_n984__,
    new_new_n985__, new_new_n987__, new_new_n988__, new_new_n989__,
    new_new_n990__, new_new_n991__, new_new_n992__, new_new_n993__,
    new_new_n995__, new_new_n996__, new_new_n997__, new_new_n998__,
    new_new_n999__, new_new_n1000__, new_new_n1001__, new_new_n1003__,
    new_new_n1004__, new_new_n1005__, new_new_n1006__, new_new_n1007__,
    new_new_n1008__, new_new_n1009__, new_new_n1011__, new_new_n1012__,
    new_new_n1013__, new_new_n1014__, new_new_n1015__, new_new_n1016__,
    new_new_n1017__, new_new_n1019__, new_new_n1020__, new_new_n1021__,
    new_new_n1022__, new_new_n1023__, new_new_n1024__, new_new_n1025__,
    new_new_n1027__, new_new_n1028__, new_new_n1029__, new_new_n1030__,
    new_new_n1031__, new_new_n1032__, new_new_n1033__, new_new_n1035__,
    new_new_n1036__, new_new_n1037__, new_new_n1038__, new_new_n1039__,
    new_new_n1040__, new_new_n1041__, new_new_n1043__, new_new_n1044__,
    new_new_n1045__, new_new_n1046__, new_new_n1047__, new_new_n1048__,
    new_new_n1049__, new_new_n1051__, new_new_n1052__, new_new_n1053__,
    new_new_n1054__, new_new_n1055__, new_new_n1056__, new_new_n1057__,
    new_new_n1059__, new_new_n1060__, new_new_n1061__, new_new_n1062__,
    new_new_n1063__, new_new_n1064__, new_new_n1065__, new_new_n1067__,
    new_new_n1068__, new_new_n1069__, new_new_n1070__, new_new_n1071__,
    new_new_n1072__, new_new_n1073__, new_new_n1075__, new_new_n1076__,
    new_new_n1077__, new_new_n1078__, new_new_n1079__, new_new_n1080__,
    new_new_n1081__, new_new_n1083__, new_new_n1084__, new_new_n1085__,
    new_new_n1086__, new_new_n1087__, new_new_n1088__, new_new_n1089__,
    new_new_n1091__, new_new_n1092__, new_new_n1093__, new_new_n1094__,
    new_new_n1095__, new_new_n1096__, new_new_n1097__, new_new_n1099__,
    new_new_n1100__, new_new_n1101__, new_new_n1102__, new_new_n1103__,
    new_new_n1104__, new_new_n1105__, new_new_n1107__, new_new_n1108__,
    new_new_n1109__, new_new_n1110__, new_new_n1111__, new_new_n1112__,
    new_new_n1113__, new_new_n1115__, new_new_n1116__, new_new_n1117__,
    new_new_n1118__, new_new_n1119__, new_new_n1120__, new_new_n1121__,
    new_new_n1123__, new_new_n1124__, new_new_n1125__, new_new_n1126__,
    new_new_n1127__, new_new_n1128__, new_new_n1129__, new_new_n1131__,
    new_new_n1132__, new_new_n1133__, new_new_n1134__, new_new_n1135__,
    new_new_n1136__, new_new_n1137__, new_new_n1139__, new_new_n1140__,
    new_new_n1141__, new_new_n1142__, new_new_n1143__, new_new_n1144__,
    new_new_n1145__, new_new_n1147__, new_new_n1148__, new_new_n1149__,
    new_new_n1150__, new_new_n1151__, new_new_n1152__, new_new_n1153__,
    new_new_n1155__, new_new_n1156__, new_new_n1157__, new_new_n1158__,
    new_new_n1159__, new_new_n1160__, new_new_n1161__, new_new_n1163__,
    new_new_n1164__, new_new_n1165__, new_new_n1166__, new_new_n1167__,
    new_new_n1168__, new_new_n1169__, new_new_n1171__, new_new_n1172__,
    new_new_n1173__, new_new_n1174__, new_new_n1175__, new_new_n1176__,
    new_new_n1177__, new_new_n1179__, new_new_n1180__, new_new_n1181__,
    new_new_n1182__, new_new_n1183__, new_new_n1184__, new_new_n1185__,
    new_new_n1187__, new_new_n1188__, new_new_n1189__, new_new_n1190__,
    new_new_n1191__, new_new_n1192__, new_new_n1193__, new_new_n1195__,
    new_new_n1196__, new_new_n1197__, new_new_n1198__, new_new_n1199__,
    new_new_n1200__, new_new_n1201__, new_new_n1203__, new_new_n1204__,
    new_new_n1205__, new_new_n1206__, new_new_n1207__, new_new_n1208__,
    new_new_n1209__, new_new_n1211__, new_new_n1212__, new_new_n1213__,
    new_new_n1214__, new_new_n1215__, new_new_n1216__, new_new_n1217__,
    new_new_n1219__, new_new_n1220__, new_new_n1221__, new_new_n1222__,
    new_new_n1223__, new_new_n1224__, new_new_n1225__, new_new_n1227__,
    new_new_n1228__, new_new_n1229__, new_new_n1230__, new_new_n1231__,
    new_new_n1232__, new_new_n1233__, new_new_n1235__, new_new_n1236__,
    new_new_n1237__, new_new_n1238__, new_new_n1239__, new_new_n1240__,
    new_new_n1241__, new_new_n1243__, new_new_n1244__, new_new_n1245__,
    new_new_n1246__, new_new_n1247__, new_new_n1248__, new_new_n1249__,
    new_new_n1251__, new_new_n1252__, new_new_n1253__, new_new_n1254__,
    new_new_n1255__, new_new_n1256__, new_new_n1257__, new_new_n1259__,
    new_new_n1260__, new_new_n1261__, new_new_n1262__, new_new_n1263__,
    new_new_n1264__, new_new_n1265__, new_new_n1267__, new_new_n1268__,
    new_new_n1269__, new_new_n1270__, new_new_n1271__, new_new_n1272__,
    new_new_n1273__, new_new_n1275__, new_new_n1276__, new_new_n1277__,
    new_new_n1278__, new_new_n1279__, new_new_n1280__, new_new_n1281__,
    new_new_n1283__, new_new_n1284__, new_new_n1285__, new_new_n1286__,
    new_new_n1287__, new_new_n1288__, new_new_n1289__, new_new_n1291__,
    new_new_n1292__, new_new_n1293__, new_new_n1294__, new_new_n1295__,
    new_new_n1296__, new_new_n1297__, new_new_n1299__, new_new_n1300__,
    new_new_n1301__, new_new_n1302__, new_new_n1303__, new_new_n1304__,
    new_new_n1305__, new_new_n1307__, new_new_n1308__, new_new_n1309__,
    new_new_n1310__, new_new_n1311__, new_new_n1312__, new_new_n1313__,
    new_new_n1315__, new_new_n1316__, new_new_n1317__, new_new_n1318__,
    new_new_n1319__, new_new_n1320__, new_new_n1321__, new_new_n1323__,
    new_new_n1324__, new_new_n1325__, new_new_n1326__, new_new_n1327__,
    new_new_n1328__, new_new_n1329__, new_new_n1331__, new_new_n1332__,
    new_new_n1333__, new_new_n1334__, new_new_n1335__, new_new_n1336__,
    new_new_n1337__, new_new_n1339__, new_new_n1340__, new_new_n1341__,
    new_new_n1342__, new_new_n1343__, new_new_n1344__, new_new_n1345__,
    new_new_n1347__, new_new_n1348__, new_new_n1349__, new_new_n1350__,
    new_new_n1351__, new_new_n1352__, new_new_n1353__, new_new_n1355__,
    new_new_n1356__, new_new_n1357__, new_new_n1358__, new_new_n1359__,
    new_new_n1360__, new_new_n1361__, new_new_n1363__, new_new_n1364__,
    new_new_n1365__, new_new_n1366__, new_new_n1367__, new_new_n1368__,
    new_new_n1369__, new_new_n1371__, new_new_n1372__, new_new_n1373__,
    new_new_n1374__, new_new_n1375__, new_new_n1376__, new_new_n1377__,
    new_new_n1379__, new_new_n1380__, new_new_n1381__, new_new_n1382__,
    new_new_n1383__, new_new_n1384__, new_new_n1385__, new_new_n1387__,
    new_new_n1388__, new_new_n1389__, new_new_n1390__, new_new_n1391__,
    new_new_n1392__, new_new_n1393__, new_new_n1395__, new_new_n1396__,
    new_new_n1397__, new_new_n1398__, new_new_n1399__, new_new_n1400__,
    new_new_n1401__, new_new_n1403__;
  assign new_new_n386__ = \a[0]  & \b[0] ;
  assign new_new_n387__ = ~\a[0]  & ~\b[0] ;
  assign \f[0]  = ~new_new_n386__ & ~new_new_n387__;
  assign new_new_n389__ = \a[1]  & \b[1] ;
  assign new_new_n390__ = ~\a[1]  & ~\b[1] ;
  assign new_new_n391__ = ~new_new_n389__ & ~new_new_n390__;
  assign new_new_n392__ = new_new_n386__ & ~new_new_n391__;
  assign new_new_n393__ = ~new_new_n386__ & new_new_n391__;
  assign \f[1]  = new_new_n392__ | new_new_n393__;
  assign new_new_n395__ = \a[2]  & \b[2] ;
  assign new_new_n396__ = ~\a[2]  & ~\b[2] ;
  assign new_new_n397__ = ~new_new_n395__ & ~new_new_n396__;
  assign new_new_n398__ = ~new_new_n386__ & ~new_new_n389__;
  assign new_new_n399__ = ~new_new_n390__ & ~new_new_n398__;
  assign new_new_n400__ = new_new_n397__ & ~new_new_n399__;
  assign new_new_n401__ = ~new_new_n397__ & new_new_n399__;
  assign \f[2]  = new_new_n400__ | new_new_n401__;
  assign new_new_n403__ = ~new_new_n395__ & ~new_new_n399__;
  assign new_new_n404__ = ~new_new_n396__ & ~new_new_n403__;
  assign new_new_n405__ = \b[3]  & new_new_n404__;
  assign new_new_n406__ = ~\b[3]  & ~new_new_n404__;
  assign new_new_n407__ = ~new_new_n405__ & ~new_new_n406__;
  assign new_new_n408__ = \a[3]  & new_new_n407__;
  assign new_new_n409__ = ~\a[3]  & ~new_new_n407__;
  assign \f[3]  = ~new_new_n408__ & ~new_new_n409__;
  assign new_new_n411__ = \a[4]  & \b[4] ;
  assign new_new_n412__ = ~\a[4]  & ~\b[4] ;
  assign new_new_n413__ = ~new_new_n411__ & ~new_new_n412__;
  assign new_new_n414__ = ~\a[3]  & ~new_new_n405__;
  assign new_new_n415__ = ~new_new_n406__ & ~new_new_n414__;
  assign new_new_n416__ = ~new_new_n413__ & new_new_n415__;
  assign new_new_n417__ = new_new_n413__ & ~new_new_n415__;
  assign \f[4]  = new_new_n416__ | new_new_n417__;
  assign new_new_n419__ = ~new_new_n411__ & ~new_new_n415__;
  assign new_new_n420__ = ~new_new_n412__ & ~new_new_n419__;
  assign new_new_n421__ = ~\a[5]  & ~\b[5] ;
  assign new_new_n422__ = \a[5]  & \b[5] ;
  assign new_new_n423__ = ~new_new_n421__ & ~new_new_n422__;
  assign new_new_n424__ = new_new_n420__ & ~new_new_n423__;
  assign new_new_n425__ = ~new_new_n420__ & new_new_n423__;
  assign \f[5]  = new_new_n424__ | new_new_n425__;
  assign new_new_n427__ = ~\a[6]  & ~\b[6] ;
  assign new_new_n428__ = \a[6]  & \b[6] ;
  assign new_new_n429__ = ~new_new_n427__ & ~new_new_n428__;
  assign new_new_n430__ = ~new_new_n420__ & ~new_new_n422__;
  assign new_new_n431__ = ~new_new_n421__ & ~new_new_n430__;
  assign new_new_n432__ = ~new_new_n429__ & new_new_n431__;
  assign new_new_n433__ = new_new_n429__ & ~new_new_n431__;
  assign \f[6]  = new_new_n432__ | new_new_n433__;
  assign new_new_n435__ = ~\a[7]  & ~\b[7] ;
  assign new_new_n436__ = \a[7]  & \b[7] ;
  assign new_new_n437__ = ~new_new_n435__ & ~new_new_n436__;
  assign new_new_n438__ = ~new_new_n428__ & ~new_new_n431__;
  assign new_new_n439__ = ~new_new_n427__ & ~new_new_n438__;
  assign new_new_n440__ = ~new_new_n437__ & new_new_n439__;
  assign new_new_n441__ = new_new_n437__ & ~new_new_n439__;
  assign \f[7]  = new_new_n440__ | new_new_n441__;
  assign new_new_n443__ = ~\a[8]  & ~\b[8] ;
  assign new_new_n444__ = \a[8]  & \b[8] ;
  assign new_new_n445__ = ~new_new_n443__ & ~new_new_n444__;
  assign new_new_n446__ = ~new_new_n436__ & ~new_new_n439__;
  assign new_new_n447__ = ~new_new_n435__ & ~new_new_n446__;
  assign new_new_n448__ = ~new_new_n445__ & new_new_n447__;
  assign new_new_n449__ = new_new_n445__ & ~new_new_n447__;
  assign \f[8]  = new_new_n448__ | new_new_n449__;
  assign new_new_n451__ = ~\a[9]  & ~\b[9] ;
  assign new_new_n452__ = \a[9]  & \b[9] ;
  assign new_new_n453__ = ~new_new_n451__ & ~new_new_n452__;
  assign new_new_n454__ = ~new_new_n444__ & ~new_new_n447__;
  assign new_new_n455__ = ~new_new_n443__ & ~new_new_n454__;
  assign new_new_n456__ = ~new_new_n453__ & new_new_n455__;
  assign new_new_n457__ = new_new_n453__ & ~new_new_n455__;
  assign \f[9]  = new_new_n456__ | new_new_n457__;
  assign new_new_n459__ = ~\a[10]  & ~\b[10] ;
  assign new_new_n460__ = \a[10]  & \b[10] ;
  assign new_new_n461__ = ~new_new_n459__ & ~new_new_n460__;
  assign new_new_n462__ = ~new_new_n452__ & ~new_new_n455__;
  assign new_new_n463__ = ~new_new_n451__ & ~new_new_n462__;
  assign new_new_n464__ = ~new_new_n461__ & new_new_n463__;
  assign new_new_n465__ = new_new_n461__ & ~new_new_n463__;
  assign \f[10]  = new_new_n464__ | new_new_n465__;
  assign new_new_n467__ = ~new_new_n460__ & ~new_new_n463__;
  assign new_new_n468__ = ~new_new_n459__ & ~new_new_n467__;
  assign new_new_n469__ = ~\b[11]  & ~new_new_n468__;
  assign new_new_n470__ = \b[11]  & new_new_n468__;
  assign new_new_n471__ = ~new_new_n469__ & ~new_new_n470__;
  assign new_new_n472__ = \a[11]  & ~new_new_n471__;
  assign new_new_n473__ = ~\a[11]  & new_new_n471__;
  assign \f[11]  = new_new_n472__ | new_new_n473__;
  assign new_new_n475__ = ~\a[11]  & ~new_new_n470__;
  assign new_new_n476__ = ~new_new_n469__ & ~new_new_n475__;
  assign new_new_n477__ = ~\a[12]  & ~\b[12] ;
  assign new_new_n478__ = \a[12]  & \b[12] ;
  assign new_new_n479__ = ~new_new_n477__ & ~new_new_n478__;
  assign new_new_n480__ = ~new_new_n476__ & new_new_n479__;
  assign new_new_n481__ = new_new_n476__ & ~new_new_n479__;
  assign \f[12]  = new_new_n480__ | new_new_n481__;
  assign new_new_n483__ = ~new_new_n476__ & ~new_new_n478__;
  assign new_new_n484__ = ~new_new_n477__ & ~new_new_n483__;
  assign new_new_n485__ = ~\b[13]  & ~new_new_n484__;
  assign new_new_n486__ = \b[13]  & new_new_n484__;
  assign new_new_n487__ = ~new_new_n485__ & ~new_new_n486__;
  assign new_new_n488__ = \a[13]  & ~new_new_n487__;
  assign new_new_n489__ = ~\a[13]  & new_new_n487__;
  assign \f[13]  = new_new_n488__ | new_new_n489__;
  assign new_new_n491__ = ~\a[13]  & ~new_new_n486__;
  assign new_new_n492__ = ~new_new_n485__ & ~new_new_n491__;
  assign new_new_n493__ = ~\a[14]  & ~\b[14] ;
  assign new_new_n494__ = \a[14]  & \b[14] ;
  assign new_new_n495__ = ~new_new_n493__ & ~new_new_n494__;
  assign new_new_n496__ = ~new_new_n492__ & new_new_n495__;
  assign new_new_n497__ = new_new_n492__ & ~new_new_n495__;
  assign \f[14]  = new_new_n496__ | new_new_n497__;
  assign new_new_n499__ = ~new_new_n492__ & ~new_new_n494__;
  assign new_new_n500__ = ~new_new_n493__ & ~new_new_n499__;
  assign new_new_n501__ = ~\b[15]  & ~new_new_n500__;
  assign new_new_n502__ = \b[15]  & new_new_n500__;
  assign new_new_n503__ = ~new_new_n501__ & ~new_new_n502__;
  assign new_new_n504__ = \a[15]  & ~new_new_n503__;
  assign new_new_n505__ = ~\a[15]  & new_new_n503__;
  assign \f[15]  = new_new_n504__ | new_new_n505__;
  assign new_new_n507__ = ~\a[15]  & ~new_new_n502__;
  assign new_new_n508__ = ~new_new_n501__ & ~new_new_n507__;
  assign new_new_n509__ = ~\a[16]  & ~\b[16] ;
  assign new_new_n510__ = \a[16]  & \b[16] ;
  assign new_new_n511__ = ~new_new_n509__ & ~new_new_n510__;
  assign new_new_n512__ = ~new_new_n508__ & new_new_n511__;
  assign new_new_n513__ = new_new_n508__ & ~new_new_n511__;
  assign \f[16]  = new_new_n512__ | new_new_n513__;
  assign new_new_n515__ = ~new_new_n508__ & ~new_new_n510__;
  assign new_new_n516__ = ~new_new_n509__ & ~new_new_n515__;
  assign new_new_n517__ = ~\b[17]  & ~new_new_n516__;
  assign new_new_n518__ = \b[17]  & new_new_n516__;
  assign new_new_n519__ = ~new_new_n517__ & ~new_new_n518__;
  assign new_new_n520__ = \a[17]  & ~new_new_n519__;
  assign new_new_n521__ = ~\a[17]  & new_new_n519__;
  assign \f[17]  = new_new_n520__ | new_new_n521__;
  assign new_new_n523__ = ~\a[17]  & ~new_new_n518__;
  assign new_new_n524__ = ~new_new_n517__ & ~new_new_n523__;
  assign new_new_n525__ = ~\a[18]  & ~\b[18] ;
  assign new_new_n526__ = \a[18]  & \b[18] ;
  assign new_new_n527__ = ~new_new_n525__ & ~new_new_n526__;
  assign new_new_n528__ = ~new_new_n524__ & new_new_n527__;
  assign new_new_n529__ = new_new_n524__ & ~new_new_n527__;
  assign \f[18]  = new_new_n528__ | new_new_n529__;
  assign new_new_n531__ = ~new_new_n524__ & ~new_new_n526__;
  assign new_new_n532__ = ~new_new_n525__ & ~new_new_n531__;
  assign new_new_n533__ = ~\b[19]  & ~new_new_n532__;
  assign new_new_n534__ = \b[19]  & new_new_n532__;
  assign new_new_n535__ = ~new_new_n533__ & ~new_new_n534__;
  assign new_new_n536__ = \a[19]  & ~new_new_n535__;
  assign new_new_n537__ = ~\a[19]  & new_new_n535__;
  assign \f[19]  = new_new_n536__ | new_new_n537__;
  assign new_new_n539__ = ~\a[19]  & ~new_new_n534__;
  assign new_new_n540__ = ~new_new_n533__ & ~new_new_n539__;
  assign new_new_n541__ = ~\a[20]  & ~\b[20] ;
  assign new_new_n542__ = \a[20]  & \b[20] ;
  assign new_new_n543__ = ~new_new_n541__ & ~new_new_n542__;
  assign new_new_n544__ = ~new_new_n540__ & new_new_n543__;
  assign new_new_n545__ = new_new_n540__ & ~new_new_n543__;
  assign \f[20]  = new_new_n544__ | new_new_n545__;
  assign new_new_n547__ = ~new_new_n540__ & ~new_new_n542__;
  assign new_new_n548__ = ~new_new_n541__ & ~new_new_n547__;
  assign new_new_n549__ = ~\b[21]  & ~new_new_n548__;
  assign new_new_n550__ = \b[21]  & new_new_n548__;
  assign new_new_n551__ = ~new_new_n549__ & ~new_new_n550__;
  assign new_new_n552__ = \a[21]  & ~new_new_n551__;
  assign new_new_n553__ = ~\a[21]  & new_new_n551__;
  assign \f[21]  = new_new_n552__ | new_new_n553__;
  assign new_new_n555__ = ~\a[21]  & ~new_new_n550__;
  assign new_new_n556__ = ~new_new_n549__ & ~new_new_n555__;
  assign new_new_n557__ = ~\a[22]  & ~\b[22] ;
  assign new_new_n558__ = \a[22]  & \b[22] ;
  assign new_new_n559__ = ~new_new_n557__ & ~new_new_n558__;
  assign new_new_n560__ = ~new_new_n556__ & new_new_n559__;
  assign new_new_n561__ = new_new_n556__ & ~new_new_n559__;
  assign \f[22]  = new_new_n560__ | new_new_n561__;
  assign new_new_n563__ = ~new_new_n556__ & ~new_new_n558__;
  assign new_new_n564__ = ~new_new_n557__ & ~new_new_n563__;
  assign new_new_n565__ = ~\b[23]  & ~new_new_n564__;
  assign new_new_n566__ = \b[23]  & new_new_n564__;
  assign new_new_n567__ = ~new_new_n565__ & ~new_new_n566__;
  assign new_new_n568__ = \a[23]  & ~new_new_n567__;
  assign new_new_n569__ = ~\a[23]  & new_new_n567__;
  assign \f[23]  = new_new_n568__ | new_new_n569__;
  assign new_new_n571__ = ~\a[23]  & ~new_new_n566__;
  assign new_new_n572__ = ~new_new_n565__ & ~new_new_n571__;
  assign new_new_n573__ = ~\a[24]  & ~\b[24] ;
  assign new_new_n574__ = \a[24]  & \b[24] ;
  assign new_new_n575__ = ~new_new_n573__ & ~new_new_n574__;
  assign new_new_n576__ = ~new_new_n572__ & new_new_n575__;
  assign new_new_n577__ = new_new_n572__ & ~new_new_n575__;
  assign \f[24]  = new_new_n576__ | new_new_n577__;
  assign new_new_n579__ = ~new_new_n572__ & ~new_new_n574__;
  assign new_new_n580__ = ~new_new_n573__ & ~new_new_n579__;
  assign new_new_n581__ = ~\b[25]  & ~new_new_n580__;
  assign new_new_n582__ = \b[25]  & new_new_n580__;
  assign new_new_n583__ = ~new_new_n581__ & ~new_new_n582__;
  assign new_new_n584__ = \a[25]  & ~new_new_n583__;
  assign new_new_n585__ = ~\a[25]  & new_new_n583__;
  assign \f[25]  = new_new_n584__ | new_new_n585__;
  assign new_new_n587__ = ~\a[25]  & ~new_new_n582__;
  assign new_new_n588__ = ~new_new_n581__ & ~new_new_n587__;
  assign new_new_n589__ = ~\a[26]  & ~\b[26] ;
  assign new_new_n590__ = \a[26]  & \b[26] ;
  assign new_new_n591__ = ~new_new_n589__ & ~new_new_n590__;
  assign new_new_n592__ = ~new_new_n588__ & new_new_n591__;
  assign new_new_n593__ = new_new_n588__ & ~new_new_n591__;
  assign \f[26]  = new_new_n592__ | new_new_n593__;
  assign new_new_n595__ = ~new_new_n588__ & ~new_new_n590__;
  assign new_new_n596__ = ~new_new_n589__ & ~new_new_n595__;
  assign new_new_n597__ = ~\b[27]  & ~new_new_n596__;
  assign new_new_n598__ = \b[27]  & new_new_n596__;
  assign new_new_n599__ = ~new_new_n597__ & ~new_new_n598__;
  assign new_new_n600__ = \a[27]  & ~new_new_n599__;
  assign new_new_n601__ = ~\a[27]  & new_new_n599__;
  assign \f[27]  = new_new_n600__ | new_new_n601__;
  assign new_new_n603__ = ~\a[27]  & ~new_new_n598__;
  assign new_new_n604__ = ~new_new_n597__ & ~new_new_n603__;
  assign new_new_n605__ = ~\a[28]  & ~\b[28] ;
  assign new_new_n606__ = \a[28]  & \b[28] ;
  assign new_new_n607__ = ~new_new_n605__ & ~new_new_n606__;
  assign new_new_n608__ = ~new_new_n604__ & new_new_n607__;
  assign new_new_n609__ = new_new_n604__ & ~new_new_n607__;
  assign \f[28]  = new_new_n608__ | new_new_n609__;
  assign new_new_n611__ = ~new_new_n604__ & ~new_new_n606__;
  assign new_new_n612__ = ~new_new_n605__ & ~new_new_n611__;
  assign new_new_n613__ = ~\b[29]  & ~new_new_n612__;
  assign new_new_n614__ = \b[29]  & new_new_n612__;
  assign new_new_n615__ = ~new_new_n613__ & ~new_new_n614__;
  assign new_new_n616__ = \a[29]  & ~new_new_n615__;
  assign new_new_n617__ = ~\a[29]  & new_new_n615__;
  assign \f[29]  = new_new_n616__ | new_new_n617__;
  assign new_new_n619__ = ~\a[29]  & ~new_new_n614__;
  assign new_new_n620__ = ~new_new_n613__ & ~new_new_n619__;
  assign new_new_n621__ = ~\a[30]  & ~\b[30] ;
  assign new_new_n622__ = \a[30]  & \b[30] ;
  assign new_new_n623__ = ~new_new_n621__ & ~new_new_n622__;
  assign new_new_n624__ = ~new_new_n620__ & new_new_n623__;
  assign new_new_n625__ = new_new_n620__ & ~new_new_n623__;
  assign \f[30]  = new_new_n624__ | new_new_n625__;
  assign new_new_n627__ = ~new_new_n620__ & ~new_new_n622__;
  assign new_new_n628__ = ~new_new_n621__ & ~new_new_n627__;
  assign new_new_n629__ = ~\b[31]  & ~new_new_n628__;
  assign new_new_n630__ = \b[31]  & new_new_n628__;
  assign new_new_n631__ = ~new_new_n629__ & ~new_new_n630__;
  assign new_new_n632__ = \a[31]  & ~new_new_n631__;
  assign new_new_n633__ = ~\a[31]  & new_new_n631__;
  assign \f[31]  = new_new_n632__ | new_new_n633__;
  assign new_new_n635__ = ~\a[31]  & ~new_new_n630__;
  assign new_new_n636__ = ~new_new_n629__ & ~new_new_n635__;
  assign new_new_n637__ = ~\a[32]  & ~\b[32] ;
  assign new_new_n638__ = \a[32]  & \b[32] ;
  assign new_new_n639__ = ~new_new_n637__ & ~new_new_n638__;
  assign new_new_n640__ = ~new_new_n636__ & new_new_n639__;
  assign new_new_n641__ = new_new_n636__ & ~new_new_n639__;
  assign \f[32]  = new_new_n640__ | new_new_n641__;
  assign new_new_n643__ = ~new_new_n636__ & ~new_new_n638__;
  assign new_new_n644__ = ~new_new_n637__ & ~new_new_n643__;
  assign new_new_n645__ = ~\b[33]  & ~new_new_n644__;
  assign new_new_n646__ = \b[33]  & new_new_n644__;
  assign new_new_n647__ = ~new_new_n645__ & ~new_new_n646__;
  assign new_new_n648__ = \a[33]  & ~new_new_n647__;
  assign new_new_n649__ = ~\a[33]  & new_new_n647__;
  assign \f[33]  = new_new_n648__ | new_new_n649__;
  assign new_new_n651__ = ~\a[33]  & ~new_new_n646__;
  assign new_new_n652__ = ~new_new_n645__ & ~new_new_n651__;
  assign new_new_n653__ = ~\a[34]  & ~\b[34] ;
  assign new_new_n654__ = \a[34]  & \b[34] ;
  assign new_new_n655__ = ~new_new_n653__ & ~new_new_n654__;
  assign new_new_n656__ = ~new_new_n652__ & new_new_n655__;
  assign new_new_n657__ = new_new_n652__ & ~new_new_n655__;
  assign \f[34]  = new_new_n656__ | new_new_n657__;
  assign new_new_n659__ = ~new_new_n652__ & ~new_new_n654__;
  assign new_new_n660__ = ~new_new_n653__ & ~new_new_n659__;
  assign new_new_n661__ = ~\b[35]  & ~new_new_n660__;
  assign new_new_n662__ = \b[35]  & new_new_n660__;
  assign new_new_n663__ = ~new_new_n661__ & ~new_new_n662__;
  assign new_new_n664__ = \a[35]  & ~new_new_n663__;
  assign new_new_n665__ = ~\a[35]  & new_new_n663__;
  assign \f[35]  = new_new_n664__ | new_new_n665__;
  assign new_new_n667__ = ~\a[35]  & ~new_new_n662__;
  assign new_new_n668__ = ~new_new_n661__ & ~new_new_n667__;
  assign new_new_n669__ = ~\a[36]  & ~\b[36] ;
  assign new_new_n670__ = \a[36]  & \b[36] ;
  assign new_new_n671__ = ~new_new_n669__ & ~new_new_n670__;
  assign new_new_n672__ = ~new_new_n668__ & new_new_n671__;
  assign new_new_n673__ = new_new_n668__ & ~new_new_n671__;
  assign \f[36]  = new_new_n672__ | new_new_n673__;
  assign new_new_n675__ = ~new_new_n668__ & ~new_new_n670__;
  assign new_new_n676__ = ~new_new_n669__ & ~new_new_n675__;
  assign new_new_n677__ = ~\b[37]  & ~new_new_n676__;
  assign new_new_n678__ = \b[37]  & new_new_n676__;
  assign new_new_n679__ = ~new_new_n677__ & ~new_new_n678__;
  assign new_new_n680__ = \a[37]  & ~new_new_n679__;
  assign new_new_n681__ = ~\a[37]  & new_new_n679__;
  assign \f[37]  = new_new_n680__ | new_new_n681__;
  assign new_new_n683__ = ~\a[37]  & ~new_new_n678__;
  assign new_new_n684__ = ~new_new_n677__ & ~new_new_n683__;
  assign new_new_n685__ = ~\a[38]  & ~\b[38] ;
  assign new_new_n686__ = \a[38]  & \b[38] ;
  assign new_new_n687__ = ~new_new_n685__ & ~new_new_n686__;
  assign new_new_n688__ = ~new_new_n684__ & new_new_n687__;
  assign new_new_n689__ = new_new_n684__ & ~new_new_n687__;
  assign \f[38]  = new_new_n688__ | new_new_n689__;
  assign new_new_n691__ = ~new_new_n684__ & ~new_new_n686__;
  assign new_new_n692__ = ~new_new_n685__ & ~new_new_n691__;
  assign new_new_n693__ = ~\b[39]  & ~new_new_n692__;
  assign new_new_n694__ = \b[39]  & new_new_n692__;
  assign new_new_n695__ = ~new_new_n693__ & ~new_new_n694__;
  assign new_new_n696__ = \a[39]  & ~new_new_n695__;
  assign new_new_n697__ = ~\a[39]  & new_new_n695__;
  assign \f[39]  = new_new_n696__ | new_new_n697__;
  assign new_new_n699__ = ~\a[39]  & ~new_new_n694__;
  assign new_new_n700__ = ~new_new_n693__ & ~new_new_n699__;
  assign new_new_n701__ = ~\a[40]  & ~\b[40] ;
  assign new_new_n702__ = \a[40]  & \b[40] ;
  assign new_new_n703__ = ~new_new_n701__ & ~new_new_n702__;
  assign new_new_n704__ = ~new_new_n700__ & new_new_n703__;
  assign new_new_n705__ = new_new_n700__ & ~new_new_n703__;
  assign \f[40]  = new_new_n704__ | new_new_n705__;
  assign new_new_n707__ = ~new_new_n700__ & ~new_new_n702__;
  assign new_new_n708__ = ~new_new_n701__ & ~new_new_n707__;
  assign new_new_n709__ = ~\b[41]  & ~new_new_n708__;
  assign new_new_n710__ = \b[41]  & new_new_n708__;
  assign new_new_n711__ = ~new_new_n709__ & ~new_new_n710__;
  assign new_new_n712__ = \a[41]  & ~new_new_n711__;
  assign new_new_n713__ = ~\a[41]  & new_new_n711__;
  assign \f[41]  = new_new_n712__ | new_new_n713__;
  assign new_new_n715__ = ~\a[41]  & ~new_new_n710__;
  assign new_new_n716__ = ~new_new_n709__ & ~new_new_n715__;
  assign new_new_n717__ = ~\a[42]  & ~\b[42] ;
  assign new_new_n718__ = \a[42]  & \b[42] ;
  assign new_new_n719__ = ~new_new_n717__ & ~new_new_n718__;
  assign new_new_n720__ = ~new_new_n716__ & new_new_n719__;
  assign new_new_n721__ = new_new_n716__ & ~new_new_n719__;
  assign \f[42]  = new_new_n720__ | new_new_n721__;
  assign new_new_n723__ = ~new_new_n716__ & ~new_new_n718__;
  assign new_new_n724__ = ~new_new_n717__ & ~new_new_n723__;
  assign new_new_n725__ = ~\b[43]  & ~new_new_n724__;
  assign new_new_n726__ = \b[43]  & new_new_n724__;
  assign new_new_n727__ = ~new_new_n725__ & ~new_new_n726__;
  assign new_new_n728__ = \a[43]  & ~new_new_n727__;
  assign new_new_n729__ = ~\a[43]  & new_new_n727__;
  assign \f[43]  = new_new_n728__ | new_new_n729__;
  assign new_new_n731__ = ~\a[43]  & ~new_new_n726__;
  assign new_new_n732__ = ~new_new_n725__ & ~new_new_n731__;
  assign new_new_n733__ = ~\a[44]  & ~\b[44] ;
  assign new_new_n734__ = \a[44]  & \b[44] ;
  assign new_new_n735__ = ~new_new_n733__ & ~new_new_n734__;
  assign new_new_n736__ = ~new_new_n732__ & new_new_n735__;
  assign new_new_n737__ = new_new_n732__ & ~new_new_n735__;
  assign \f[44]  = new_new_n736__ | new_new_n737__;
  assign new_new_n739__ = ~new_new_n732__ & ~new_new_n734__;
  assign new_new_n740__ = ~new_new_n733__ & ~new_new_n739__;
  assign new_new_n741__ = ~\b[45]  & ~new_new_n740__;
  assign new_new_n742__ = \b[45]  & new_new_n740__;
  assign new_new_n743__ = ~new_new_n741__ & ~new_new_n742__;
  assign new_new_n744__ = \a[45]  & ~new_new_n743__;
  assign new_new_n745__ = ~\a[45]  & new_new_n743__;
  assign \f[45]  = new_new_n744__ | new_new_n745__;
  assign new_new_n747__ = ~\a[45]  & ~new_new_n742__;
  assign new_new_n748__ = ~new_new_n741__ & ~new_new_n747__;
  assign new_new_n749__ = ~\a[46]  & ~\b[46] ;
  assign new_new_n750__ = \a[46]  & \b[46] ;
  assign new_new_n751__ = ~new_new_n749__ & ~new_new_n750__;
  assign new_new_n752__ = ~new_new_n748__ & new_new_n751__;
  assign new_new_n753__ = new_new_n748__ & ~new_new_n751__;
  assign \f[46]  = new_new_n752__ | new_new_n753__;
  assign new_new_n755__ = ~new_new_n748__ & ~new_new_n750__;
  assign new_new_n756__ = ~new_new_n749__ & ~new_new_n755__;
  assign new_new_n757__ = ~\b[47]  & ~new_new_n756__;
  assign new_new_n758__ = \b[47]  & new_new_n756__;
  assign new_new_n759__ = ~new_new_n757__ & ~new_new_n758__;
  assign new_new_n760__ = \a[47]  & ~new_new_n759__;
  assign new_new_n761__ = ~\a[47]  & new_new_n759__;
  assign \f[47]  = new_new_n760__ | new_new_n761__;
  assign new_new_n763__ = ~\a[47]  & ~new_new_n758__;
  assign new_new_n764__ = ~new_new_n757__ & ~new_new_n763__;
  assign new_new_n765__ = ~\a[48]  & ~\b[48] ;
  assign new_new_n766__ = \a[48]  & \b[48] ;
  assign new_new_n767__ = ~new_new_n765__ & ~new_new_n766__;
  assign new_new_n768__ = ~new_new_n764__ & new_new_n767__;
  assign new_new_n769__ = new_new_n764__ & ~new_new_n767__;
  assign \f[48]  = new_new_n768__ | new_new_n769__;
  assign new_new_n771__ = ~new_new_n764__ & ~new_new_n766__;
  assign new_new_n772__ = ~new_new_n765__ & ~new_new_n771__;
  assign new_new_n773__ = ~\b[49]  & ~new_new_n772__;
  assign new_new_n774__ = \b[49]  & new_new_n772__;
  assign new_new_n775__ = ~new_new_n773__ & ~new_new_n774__;
  assign new_new_n776__ = \a[49]  & ~new_new_n775__;
  assign new_new_n777__ = ~\a[49]  & new_new_n775__;
  assign \f[49]  = new_new_n776__ | new_new_n777__;
  assign new_new_n779__ = ~\a[49]  & ~new_new_n774__;
  assign new_new_n780__ = ~new_new_n773__ & ~new_new_n779__;
  assign new_new_n781__ = ~\a[50]  & ~\b[50] ;
  assign new_new_n782__ = \a[50]  & \b[50] ;
  assign new_new_n783__ = ~new_new_n781__ & ~new_new_n782__;
  assign new_new_n784__ = ~new_new_n780__ & new_new_n783__;
  assign new_new_n785__ = new_new_n780__ & ~new_new_n783__;
  assign \f[50]  = new_new_n784__ | new_new_n785__;
  assign new_new_n787__ = ~new_new_n780__ & ~new_new_n782__;
  assign new_new_n788__ = ~new_new_n781__ & ~new_new_n787__;
  assign new_new_n789__ = ~\b[51]  & ~new_new_n788__;
  assign new_new_n790__ = \b[51]  & new_new_n788__;
  assign new_new_n791__ = ~new_new_n789__ & ~new_new_n790__;
  assign new_new_n792__ = \a[51]  & ~new_new_n791__;
  assign new_new_n793__ = ~\a[51]  & new_new_n791__;
  assign \f[51]  = new_new_n792__ | new_new_n793__;
  assign new_new_n795__ = ~\a[51]  & ~new_new_n790__;
  assign new_new_n796__ = ~new_new_n789__ & ~new_new_n795__;
  assign new_new_n797__ = ~\a[52]  & ~\b[52] ;
  assign new_new_n798__ = \a[52]  & \b[52] ;
  assign new_new_n799__ = ~new_new_n797__ & ~new_new_n798__;
  assign new_new_n800__ = ~new_new_n796__ & new_new_n799__;
  assign new_new_n801__ = new_new_n796__ & ~new_new_n799__;
  assign \f[52]  = new_new_n800__ | new_new_n801__;
  assign new_new_n803__ = ~new_new_n796__ & ~new_new_n798__;
  assign new_new_n804__ = ~new_new_n797__ & ~new_new_n803__;
  assign new_new_n805__ = ~\b[53]  & ~new_new_n804__;
  assign new_new_n806__ = \b[53]  & new_new_n804__;
  assign new_new_n807__ = ~new_new_n805__ & ~new_new_n806__;
  assign new_new_n808__ = \a[53]  & ~new_new_n807__;
  assign new_new_n809__ = ~\a[53]  & new_new_n807__;
  assign \f[53]  = new_new_n808__ | new_new_n809__;
  assign new_new_n811__ = ~\a[53]  & ~new_new_n806__;
  assign new_new_n812__ = ~new_new_n805__ & ~new_new_n811__;
  assign new_new_n813__ = ~\a[54]  & ~\b[54] ;
  assign new_new_n814__ = \a[54]  & \b[54] ;
  assign new_new_n815__ = ~new_new_n813__ & ~new_new_n814__;
  assign new_new_n816__ = ~new_new_n812__ & new_new_n815__;
  assign new_new_n817__ = new_new_n812__ & ~new_new_n815__;
  assign \f[54]  = new_new_n816__ | new_new_n817__;
  assign new_new_n819__ = ~new_new_n812__ & ~new_new_n814__;
  assign new_new_n820__ = ~new_new_n813__ & ~new_new_n819__;
  assign new_new_n821__ = ~\b[55]  & ~new_new_n820__;
  assign new_new_n822__ = \b[55]  & new_new_n820__;
  assign new_new_n823__ = ~new_new_n821__ & ~new_new_n822__;
  assign new_new_n824__ = \a[55]  & ~new_new_n823__;
  assign new_new_n825__ = ~\a[55]  & new_new_n823__;
  assign \f[55]  = new_new_n824__ | new_new_n825__;
  assign new_new_n827__ = ~\a[55]  & ~new_new_n822__;
  assign new_new_n828__ = ~new_new_n821__ & ~new_new_n827__;
  assign new_new_n829__ = ~\a[56]  & ~\b[56] ;
  assign new_new_n830__ = \a[56]  & \b[56] ;
  assign new_new_n831__ = ~new_new_n829__ & ~new_new_n830__;
  assign new_new_n832__ = ~new_new_n828__ & new_new_n831__;
  assign new_new_n833__ = new_new_n828__ & ~new_new_n831__;
  assign \f[56]  = new_new_n832__ | new_new_n833__;
  assign new_new_n835__ = ~new_new_n828__ & ~new_new_n830__;
  assign new_new_n836__ = ~new_new_n829__ & ~new_new_n835__;
  assign new_new_n837__ = ~\b[57]  & ~new_new_n836__;
  assign new_new_n838__ = \b[57]  & new_new_n836__;
  assign new_new_n839__ = ~new_new_n837__ & ~new_new_n838__;
  assign new_new_n840__ = \a[57]  & ~new_new_n839__;
  assign new_new_n841__ = ~\a[57]  & new_new_n839__;
  assign \f[57]  = new_new_n840__ | new_new_n841__;
  assign new_new_n843__ = ~\a[57]  & ~new_new_n838__;
  assign new_new_n844__ = ~new_new_n837__ & ~new_new_n843__;
  assign new_new_n845__ = ~\a[58]  & ~\b[58] ;
  assign new_new_n846__ = \a[58]  & \b[58] ;
  assign new_new_n847__ = ~new_new_n845__ & ~new_new_n846__;
  assign new_new_n848__ = ~new_new_n844__ & new_new_n847__;
  assign new_new_n849__ = new_new_n844__ & ~new_new_n847__;
  assign \f[58]  = new_new_n848__ | new_new_n849__;
  assign new_new_n851__ = ~new_new_n844__ & ~new_new_n846__;
  assign new_new_n852__ = ~new_new_n845__ & ~new_new_n851__;
  assign new_new_n853__ = ~\b[59]  & ~new_new_n852__;
  assign new_new_n854__ = \b[59]  & new_new_n852__;
  assign new_new_n855__ = ~new_new_n853__ & ~new_new_n854__;
  assign new_new_n856__ = \a[59]  & ~new_new_n855__;
  assign new_new_n857__ = ~\a[59]  & new_new_n855__;
  assign \f[59]  = new_new_n856__ | new_new_n857__;
  assign new_new_n859__ = ~\a[59]  & ~new_new_n854__;
  assign new_new_n860__ = ~new_new_n853__ & ~new_new_n859__;
  assign new_new_n861__ = ~\a[60]  & ~\b[60] ;
  assign new_new_n862__ = \a[60]  & \b[60] ;
  assign new_new_n863__ = ~new_new_n861__ & ~new_new_n862__;
  assign new_new_n864__ = ~new_new_n860__ & new_new_n863__;
  assign new_new_n865__ = new_new_n860__ & ~new_new_n863__;
  assign \f[60]  = new_new_n864__ | new_new_n865__;
  assign new_new_n867__ = ~new_new_n860__ & ~new_new_n862__;
  assign new_new_n868__ = ~new_new_n861__ & ~new_new_n867__;
  assign new_new_n869__ = ~\b[61]  & ~new_new_n868__;
  assign new_new_n870__ = \b[61]  & new_new_n868__;
  assign new_new_n871__ = ~new_new_n869__ & ~new_new_n870__;
  assign new_new_n872__ = \a[61]  & ~new_new_n871__;
  assign new_new_n873__ = ~\a[61]  & new_new_n871__;
  assign \f[61]  = new_new_n872__ | new_new_n873__;
  assign new_new_n875__ = ~\a[61]  & ~new_new_n870__;
  assign new_new_n876__ = ~new_new_n869__ & ~new_new_n875__;
  assign new_new_n877__ = ~\a[62]  & ~\b[62] ;
  assign new_new_n878__ = \a[62]  & \b[62] ;
  assign new_new_n879__ = ~new_new_n877__ & ~new_new_n878__;
  assign new_new_n880__ = ~new_new_n876__ & new_new_n879__;
  assign new_new_n881__ = new_new_n876__ & ~new_new_n879__;
  assign \f[62]  = new_new_n880__ | new_new_n881__;
  assign new_new_n883__ = ~new_new_n876__ & ~new_new_n878__;
  assign new_new_n884__ = ~new_new_n877__ & ~new_new_n883__;
  assign new_new_n885__ = ~\b[63]  & ~new_new_n884__;
  assign new_new_n886__ = \b[63]  & new_new_n884__;
  assign new_new_n887__ = ~new_new_n885__ & ~new_new_n886__;
  assign new_new_n888__ = \a[63]  & ~new_new_n887__;
  assign new_new_n889__ = ~\a[63]  & new_new_n887__;
  assign \f[63]  = new_new_n888__ | new_new_n889__;
  assign new_new_n891__ = ~\a[63]  & ~new_new_n886__;
  assign new_new_n892__ = ~new_new_n885__ & ~new_new_n891__;
  assign new_new_n893__ = ~\a[64]  & ~\b[64] ;
  assign new_new_n894__ = \a[64]  & \b[64] ;
  assign new_new_n895__ = ~new_new_n893__ & ~new_new_n894__;
  assign new_new_n896__ = ~new_new_n892__ & new_new_n895__;
  assign new_new_n897__ = new_new_n892__ & ~new_new_n895__;
  assign \f[64]  = new_new_n896__ | new_new_n897__;
  assign new_new_n899__ = ~new_new_n892__ & ~new_new_n894__;
  assign new_new_n900__ = ~new_new_n893__ & ~new_new_n899__;
  assign new_new_n901__ = ~\b[65]  & ~new_new_n900__;
  assign new_new_n902__ = \b[65]  & new_new_n900__;
  assign new_new_n903__ = ~new_new_n901__ & ~new_new_n902__;
  assign new_new_n904__ = \a[65]  & ~new_new_n903__;
  assign new_new_n905__ = ~\a[65]  & new_new_n903__;
  assign \f[65]  = new_new_n904__ | new_new_n905__;
  assign new_new_n907__ = ~\a[65]  & ~new_new_n902__;
  assign new_new_n908__ = ~new_new_n901__ & ~new_new_n907__;
  assign new_new_n909__ = ~\a[66]  & ~\b[66] ;
  assign new_new_n910__ = \a[66]  & \b[66] ;
  assign new_new_n911__ = ~new_new_n909__ & ~new_new_n910__;
  assign new_new_n912__ = ~new_new_n908__ & new_new_n911__;
  assign new_new_n913__ = new_new_n908__ & ~new_new_n911__;
  assign \f[66]  = new_new_n912__ | new_new_n913__;
  assign new_new_n915__ = ~new_new_n908__ & ~new_new_n910__;
  assign new_new_n916__ = ~new_new_n909__ & ~new_new_n915__;
  assign new_new_n917__ = ~\b[67]  & ~new_new_n916__;
  assign new_new_n918__ = \b[67]  & new_new_n916__;
  assign new_new_n919__ = ~new_new_n917__ & ~new_new_n918__;
  assign new_new_n920__ = \a[67]  & ~new_new_n919__;
  assign new_new_n921__ = ~\a[67]  & new_new_n919__;
  assign \f[67]  = new_new_n920__ | new_new_n921__;
  assign new_new_n923__ = ~\a[67]  & ~new_new_n918__;
  assign new_new_n924__ = ~new_new_n917__ & ~new_new_n923__;
  assign new_new_n925__ = ~\a[68]  & ~\b[68] ;
  assign new_new_n926__ = \a[68]  & \b[68] ;
  assign new_new_n927__ = ~new_new_n925__ & ~new_new_n926__;
  assign new_new_n928__ = ~new_new_n924__ & new_new_n927__;
  assign new_new_n929__ = new_new_n924__ & ~new_new_n927__;
  assign \f[68]  = new_new_n928__ | new_new_n929__;
  assign new_new_n931__ = ~new_new_n924__ & ~new_new_n926__;
  assign new_new_n932__ = ~new_new_n925__ & ~new_new_n931__;
  assign new_new_n933__ = ~\b[69]  & ~new_new_n932__;
  assign new_new_n934__ = \b[69]  & new_new_n932__;
  assign new_new_n935__ = ~new_new_n933__ & ~new_new_n934__;
  assign new_new_n936__ = \a[69]  & ~new_new_n935__;
  assign new_new_n937__ = ~\a[69]  & new_new_n935__;
  assign \f[69]  = new_new_n936__ | new_new_n937__;
  assign new_new_n939__ = ~\a[69]  & ~new_new_n934__;
  assign new_new_n940__ = ~new_new_n933__ & ~new_new_n939__;
  assign new_new_n941__ = ~\a[70]  & ~\b[70] ;
  assign new_new_n942__ = \a[70]  & \b[70] ;
  assign new_new_n943__ = ~new_new_n941__ & ~new_new_n942__;
  assign new_new_n944__ = ~new_new_n940__ & new_new_n943__;
  assign new_new_n945__ = new_new_n940__ & ~new_new_n943__;
  assign \f[70]  = new_new_n944__ | new_new_n945__;
  assign new_new_n947__ = ~new_new_n940__ & ~new_new_n942__;
  assign new_new_n948__ = ~new_new_n941__ & ~new_new_n947__;
  assign new_new_n949__ = ~\b[71]  & ~new_new_n948__;
  assign new_new_n950__ = \b[71]  & new_new_n948__;
  assign new_new_n951__ = ~new_new_n949__ & ~new_new_n950__;
  assign new_new_n952__ = \a[71]  & ~new_new_n951__;
  assign new_new_n953__ = ~\a[71]  & new_new_n951__;
  assign \f[71]  = new_new_n952__ | new_new_n953__;
  assign new_new_n955__ = ~\a[71]  & ~new_new_n950__;
  assign new_new_n956__ = ~new_new_n949__ & ~new_new_n955__;
  assign new_new_n957__ = ~\a[72]  & ~\b[72] ;
  assign new_new_n958__ = \a[72]  & \b[72] ;
  assign new_new_n959__ = ~new_new_n957__ & ~new_new_n958__;
  assign new_new_n960__ = ~new_new_n956__ & new_new_n959__;
  assign new_new_n961__ = new_new_n956__ & ~new_new_n959__;
  assign \f[72]  = new_new_n960__ | new_new_n961__;
  assign new_new_n963__ = ~new_new_n956__ & ~new_new_n958__;
  assign new_new_n964__ = ~new_new_n957__ & ~new_new_n963__;
  assign new_new_n965__ = ~\b[73]  & ~new_new_n964__;
  assign new_new_n966__ = \b[73]  & new_new_n964__;
  assign new_new_n967__ = ~new_new_n965__ & ~new_new_n966__;
  assign new_new_n968__ = \a[73]  & ~new_new_n967__;
  assign new_new_n969__ = ~\a[73]  & new_new_n967__;
  assign \f[73]  = new_new_n968__ | new_new_n969__;
  assign new_new_n971__ = ~\a[73]  & ~new_new_n966__;
  assign new_new_n972__ = ~new_new_n965__ & ~new_new_n971__;
  assign new_new_n973__ = ~\a[74]  & ~\b[74] ;
  assign new_new_n974__ = \a[74]  & \b[74] ;
  assign new_new_n975__ = ~new_new_n973__ & ~new_new_n974__;
  assign new_new_n976__ = ~new_new_n972__ & new_new_n975__;
  assign new_new_n977__ = new_new_n972__ & ~new_new_n975__;
  assign \f[74]  = new_new_n976__ | new_new_n977__;
  assign new_new_n979__ = ~new_new_n972__ & ~new_new_n974__;
  assign new_new_n980__ = ~new_new_n973__ & ~new_new_n979__;
  assign new_new_n981__ = ~\b[75]  & ~new_new_n980__;
  assign new_new_n982__ = \b[75]  & new_new_n980__;
  assign new_new_n983__ = ~new_new_n981__ & ~new_new_n982__;
  assign new_new_n984__ = \a[75]  & ~new_new_n983__;
  assign new_new_n985__ = ~\a[75]  & new_new_n983__;
  assign \f[75]  = new_new_n984__ | new_new_n985__;
  assign new_new_n987__ = ~\a[75]  & ~new_new_n982__;
  assign new_new_n988__ = ~new_new_n981__ & ~new_new_n987__;
  assign new_new_n989__ = ~\a[76]  & ~\b[76] ;
  assign new_new_n990__ = \a[76]  & \b[76] ;
  assign new_new_n991__ = ~new_new_n989__ & ~new_new_n990__;
  assign new_new_n992__ = ~new_new_n988__ & new_new_n991__;
  assign new_new_n993__ = new_new_n988__ & ~new_new_n991__;
  assign \f[76]  = new_new_n992__ | new_new_n993__;
  assign new_new_n995__ = ~new_new_n988__ & ~new_new_n990__;
  assign new_new_n996__ = ~new_new_n989__ & ~new_new_n995__;
  assign new_new_n997__ = ~\b[77]  & ~new_new_n996__;
  assign new_new_n998__ = \b[77]  & new_new_n996__;
  assign new_new_n999__ = ~new_new_n997__ & ~new_new_n998__;
  assign new_new_n1000__ = \a[77]  & ~new_new_n999__;
  assign new_new_n1001__ = ~\a[77]  & new_new_n999__;
  assign \f[77]  = new_new_n1000__ | new_new_n1001__;
  assign new_new_n1003__ = ~\a[77]  & ~new_new_n998__;
  assign new_new_n1004__ = ~new_new_n997__ & ~new_new_n1003__;
  assign new_new_n1005__ = ~\a[78]  & ~\b[78] ;
  assign new_new_n1006__ = \a[78]  & \b[78] ;
  assign new_new_n1007__ = ~new_new_n1005__ & ~new_new_n1006__;
  assign new_new_n1008__ = ~new_new_n1004__ & new_new_n1007__;
  assign new_new_n1009__ = new_new_n1004__ & ~new_new_n1007__;
  assign \f[78]  = new_new_n1008__ | new_new_n1009__;
  assign new_new_n1011__ = ~new_new_n1004__ & ~new_new_n1006__;
  assign new_new_n1012__ = ~new_new_n1005__ & ~new_new_n1011__;
  assign new_new_n1013__ = ~\b[79]  & ~new_new_n1012__;
  assign new_new_n1014__ = \b[79]  & new_new_n1012__;
  assign new_new_n1015__ = ~new_new_n1013__ & ~new_new_n1014__;
  assign new_new_n1016__ = \a[79]  & ~new_new_n1015__;
  assign new_new_n1017__ = ~\a[79]  & new_new_n1015__;
  assign \f[79]  = new_new_n1016__ | new_new_n1017__;
  assign new_new_n1019__ = ~\a[79]  & ~new_new_n1014__;
  assign new_new_n1020__ = ~new_new_n1013__ & ~new_new_n1019__;
  assign new_new_n1021__ = ~\a[80]  & ~\b[80] ;
  assign new_new_n1022__ = \a[80]  & \b[80] ;
  assign new_new_n1023__ = ~new_new_n1021__ & ~new_new_n1022__;
  assign new_new_n1024__ = ~new_new_n1020__ & new_new_n1023__;
  assign new_new_n1025__ = new_new_n1020__ & ~new_new_n1023__;
  assign \f[80]  = new_new_n1024__ | new_new_n1025__;
  assign new_new_n1027__ = ~new_new_n1020__ & ~new_new_n1022__;
  assign new_new_n1028__ = ~new_new_n1021__ & ~new_new_n1027__;
  assign new_new_n1029__ = ~\b[81]  & ~new_new_n1028__;
  assign new_new_n1030__ = \b[81]  & new_new_n1028__;
  assign new_new_n1031__ = ~new_new_n1029__ & ~new_new_n1030__;
  assign new_new_n1032__ = \a[81]  & ~new_new_n1031__;
  assign new_new_n1033__ = ~\a[81]  & new_new_n1031__;
  assign \f[81]  = new_new_n1032__ | new_new_n1033__;
  assign new_new_n1035__ = ~\a[81]  & ~new_new_n1030__;
  assign new_new_n1036__ = ~new_new_n1029__ & ~new_new_n1035__;
  assign new_new_n1037__ = ~\a[82]  & ~\b[82] ;
  assign new_new_n1038__ = \a[82]  & \b[82] ;
  assign new_new_n1039__ = ~new_new_n1037__ & ~new_new_n1038__;
  assign new_new_n1040__ = ~new_new_n1036__ & new_new_n1039__;
  assign new_new_n1041__ = new_new_n1036__ & ~new_new_n1039__;
  assign \f[82]  = new_new_n1040__ | new_new_n1041__;
  assign new_new_n1043__ = ~new_new_n1036__ & ~new_new_n1038__;
  assign new_new_n1044__ = ~new_new_n1037__ & ~new_new_n1043__;
  assign new_new_n1045__ = ~\b[83]  & ~new_new_n1044__;
  assign new_new_n1046__ = \b[83]  & new_new_n1044__;
  assign new_new_n1047__ = ~new_new_n1045__ & ~new_new_n1046__;
  assign new_new_n1048__ = \a[83]  & ~new_new_n1047__;
  assign new_new_n1049__ = ~\a[83]  & new_new_n1047__;
  assign \f[83]  = new_new_n1048__ | new_new_n1049__;
  assign new_new_n1051__ = ~\a[83]  & ~new_new_n1046__;
  assign new_new_n1052__ = ~new_new_n1045__ & ~new_new_n1051__;
  assign new_new_n1053__ = ~\a[84]  & ~\b[84] ;
  assign new_new_n1054__ = \a[84]  & \b[84] ;
  assign new_new_n1055__ = ~new_new_n1053__ & ~new_new_n1054__;
  assign new_new_n1056__ = ~new_new_n1052__ & new_new_n1055__;
  assign new_new_n1057__ = new_new_n1052__ & ~new_new_n1055__;
  assign \f[84]  = new_new_n1056__ | new_new_n1057__;
  assign new_new_n1059__ = ~new_new_n1052__ & ~new_new_n1054__;
  assign new_new_n1060__ = ~new_new_n1053__ & ~new_new_n1059__;
  assign new_new_n1061__ = ~\b[85]  & ~new_new_n1060__;
  assign new_new_n1062__ = \b[85]  & new_new_n1060__;
  assign new_new_n1063__ = ~new_new_n1061__ & ~new_new_n1062__;
  assign new_new_n1064__ = \a[85]  & ~new_new_n1063__;
  assign new_new_n1065__ = ~\a[85]  & new_new_n1063__;
  assign \f[85]  = new_new_n1064__ | new_new_n1065__;
  assign new_new_n1067__ = ~\a[85]  & ~new_new_n1062__;
  assign new_new_n1068__ = ~new_new_n1061__ & ~new_new_n1067__;
  assign new_new_n1069__ = ~\a[86]  & ~\b[86] ;
  assign new_new_n1070__ = \a[86]  & \b[86] ;
  assign new_new_n1071__ = ~new_new_n1069__ & ~new_new_n1070__;
  assign new_new_n1072__ = ~new_new_n1068__ & new_new_n1071__;
  assign new_new_n1073__ = new_new_n1068__ & ~new_new_n1071__;
  assign \f[86]  = new_new_n1072__ | new_new_n1073__;
  assign new_new_n1075__ = ~new_new_n1068__ & ~new_new_n1070__;
  assign new_new_n1076__ = ~new_new_n1069__ & ~new_new_n1075__;
  assign new_new_n1077__ = ~\b[87]  & ~new_new_n1076__;
  assign new_new_n1078__ = \b[87]  & new_new_n1076__;
  assign new_new_n1079__ = ~new_new_n1077__ & ~new_new_n1078__;
  assign new_new_n1080__ = \a[87]  & ~new_new_n1079__;
  assign new_new_n1081__ = ~\a[87]  & new_new_n1079__;
  assign \f[87]  = new_new_n1080__ | new_new_n1081__;
  assign new_new_n1083__ = ~\a[87]  & ~new_new_n1078__;
  assign new_new_n1084__ = ~new_new_n1077__ & ~new_new_n1083__;
  assign new_new_n1085__ = ~\a[88]  & ~\b[88] ;
  assign new_new_n1086__ = \a[88]  & \b[88] ;
  assign new_new_n1087__ = ~new_new_n1085__ & ~new_new_n1086__;
  assign new_new_n1088__ = ~new_new_n1084__ & new_new_n1087__;
  assign new_new_n1089__ = new_new_n1084__ & ~new_new_n1087__;
  assign \f[88]  = new_new_n1088__ | new_new_n1089__;
  assign new_new_n1091__ = ~new_new_n1084__ & ~new_new_n1086__;
  assign new_new_n1092__ = ~new_new_n1085__ & ~new_new_n1091__;
  assign new_new_n1093__ = ~\b[89]  & ~new_new_n1092__;
  assign new_new_n1094__ = \b[89]  & new_new_n1092__;
  assign new_new_n1095__ = ~new_new_n1093__ & ~new_new_n1094__;
  assign new_new_n1096__ = \a[89]  & ~new_new_n1095__;
  assign new_new_n1097__ = ~\a[89]  & new_new_n1095__;
  assign \f[89]  = new_new_n1096__ | new_new_n1097__;
  assign new_new_n1099__ = ~\a[89]  & ~new_new_n1094__;
  assign new_new_n1100__ = ~new_new_n1093__ & ~new_new_n1099__;
  assign new_new_n1101__ = ~\a[90]  & ~\b[90] ;
  assign new_new_n1102__ = \a[90]  & \b[90] ;
  assign new_new_n1103__ = ~new_new_n1101__ & ~new_new_n1102__;
  assign new_new_n1104__ = ~new_new_n1100__ & new_new_n1103__;
  assign new_new_n1105__ = new_new_n1100__ & ~new_new_n1103__;
  assign \f[90]  = new_new_n1104__ | new_new_n1105__;
  assign new_new_n1107__ = ~new_new_n1100__ & ~new_new_n1102__;
  assign new_new_n1108__ = ~new_new_n1101__ & ~new_new_n1107__;
  assign new_new_n1109__ = ~\b[91]  & ~new_new_n1108__;
  assign new_new_n1110__ = \b[91]  & new_new_n1108__;
  assign new_new_n1111__ = ~new_new_n1109__ & ~new_new_n1110__;
  assign new_new_n1112__ = \a[91]  & ~new_new_n1111__;
  assign new_new_n1113__ = ~\a[91]  & new_new_n1111__;
  assign \f[91]  = new_new_n1112__ | new_new_n1113__;
  assign new_new_n1115__ = ~\a[91]  & ~new_new_n1110__;
  assign new_new_n1116__ = ~new_new_n1109__ & ~new_new_n1115__;
  assign new_new_n1117__ = ~\a[92]  & ~\b[92] ;
  assign new_new_n1118__ = \a[92]  & \b[92] ;
  assign new_new_n1119__ = ~new_new_n1117__ & ~new_new_n1118__;
  assign new_new_n1120__ = ~new_new_n1116__ & new_new_n1119__;
  assign new_new_n1121__ = new_new_n1116__ & ~new_new_n1119__;
  assign \f[92]  = new_new_n1120__ | new_new_n1121__;
  assign new_new_n1123__ = ~new_new_n1116__ & ~new_new_n1118__;
  assign new_new_n1124__ = ~new_new_n1117__ & ~new_new_n1123__;
  assign new_new_n1125__ = ~\b[93]  & ~new_new_n1124__;
  assign new_new_n1126__ = \b[93]  & new_new_n1124__;
  assign new_new_n1127__ = ~new_new_n1125__ & ~new_new_n1126__;
  assign new_new_n1128__ = \a[93]  & ~new_new_n1127__;
  assign new_new_n1129__ = ~\a[93]  & new_new_n1127__;
  assign \f[93]  = new_new_n1128__ | new_new_n1129__;
  assign new_new_n1131__ = ~\a[93]  & ~new_new_n1126__;
  assign new_new_n1132__ = ~new_new_n1125__ & ~new_new_n1131__;
  assign new_new_n1133__ = ~\a[94]  & ~\b[94] ;
  assign new_new_n1134__ = \a[94]  & \b[94] ;
  assign new_new_n1135__ = ~new_new_n1133__ & ~new_new_n1134__;
  assign new_new_n1136__ = ~new_new_n1132__ & new_new_n1135__;
  assign new_new_n1137__ = new_new_n1132__ & ~new_new_n1135__;
  assign \f[94]  = new_new_n1136__ | new_new_n1137__;
  assign new_new_n1139__ = ~new_new_n1132__ & ~new_new_n1134__;
  assign new_new_n1140__ = ~new_new_n1133__ & ~new_new_n1139__;
  assign new_new_n1141__ = ~\b[95]  & ~new_new_n1140__;
  assign new_new_n1142__ = \b[95]  & new_new_n1140__;
  assign new_new_n1143__ = ~new_new_n1141__ & ~new_new_n1142__;
  assign new_new_n1144__ = \a[95]  & ~new_new_n1143__;
  assign new_new_n1145__ = ~\a[95]  & new_new_n1143__;
  assign \f[95]  = new_new_n1144__ | new_new_n1145__;
  assign new_new_n1147__ = ~\a[95]  & ~new_new_n1142__;
  assign new_new_n1148__ = ~new_new_n1141__ & ~new_new_n1147__;
  assign new_new_n1149__ = ~\a[96]  & ~\b[96] ;
  assign new_new_n1150__ = \a[96]  & \b[96] ;
  assign new_new_n1151__ = ~new_new_n1149__ & ~new_new_n1150__;
  assign new_new_n1152__ = ~new_new_n1148__ & new_new_n1151__;
  assign new_new_n1153__ = new_new_n1148__ & ~new_new_n1151__;
  assign \f[96]  = new_new_n1152__ | new_new_n1153__;
  assign new_new_n1155__ = ~new_new_n1148__ & ~new_new_n1150__;
  assign new_new_n1156__ = ~new_new_n1149__ & ~new_new_n1155__;
  assign new_new_n1157__ = ~\b[97]  & ~new_new_n1156__;
  assign new_new_n1158__ = \b[97]  & new_new_n1156__;
  assign new_new_n1159__ = ~new_new_n1157__ & ~new_new_n1158__;
  assign new_new_n1160__ = \a[97]  & ~new_new_n1159__;
  assign new_new_n1161__ = ~\a[97]  & new_new_n1159__;
  assign \f[97]  = new_new_n1160__ | new_new_n1161__;
  assign new_new_n1163__ = ~\a[97]  & ~new_new_n1158__;
  assign new_new_n1164__ = ~new_new_n1157__ & ~new_new_n1163__;
  assign new_new_n1165__ = ~\a[98]  & ~\b[98] ;
  assign new_new_n1166__ = \a[98]  & \b[98] ;
  assign new_new_n1167__ = ~new_new_n1165__ & ~new_new_n1166__;
  assign new_new_n1168__ = ~new_new_n1164__ & new_new_n1167__;
  assign new_new_n1169__ = new_new_n1164__ & ~new_new_n1167__;
  assign \f[98]  = new_new_n1168__ | new_new_n1169__;
  assign new_new_n1171__ = ~new_new_n1164__ & ~new_new_n1166__;
  assign new_new_n1172__ = ~new_new_n1165__ & ~new_new_n1171__;
  assign new_new_n1173__ = ~\b[99]  & ~new_new_n1172__;
  assign new_new_n1174__ = \b[99]  & new_new_n1172__;
  assign new_new_n1175__ = ~new_new_n1173__ & ~new_new_n1174__;
  assign new_new_n1176__ = \a[99]  & ~new_new_n1175__;
  assign new_new_n1177__ = ~\a[99]  & new_new_n1175__;
  assign \f[99]  = new_new_n1176__ | new_new_n1177__;
  assign new_new_n1179__ = ~\a[99]  & ~new_new_n1174__;
  assign new_new_n1180__ = ~new_new_n1173__ & ~new_new_n1179__;
  assign new_new_n1181__ = ~\a[100]  & ~\b[100] ;
  assign new_new_n1182__ = \a[100]  & \b[100] ;
  assign new_new_n1183__ = ~new_new_n1181__ & ~new_new_n1182__;
  assign new_new_n1184__ = ~new_new_n1180__ & new_new_n1183__;
  assign new_new_n1185__ = new_new_n1180__ & ~new_new_n1183__;
  assign \f[100]  = new_new_n1184__ | new_new_n1185__;
  assign new_new_n1187__ = ~new_new_n1180__ & ~new_new_n1182__;
  assign new_new_n1188__ = ~new_new_n1181__ & ~new_new_n1187__;
  assign new_new_n1189__ = ~\b[101]  & ~new_new_n1188__;
  assign new_new_n1190__ = \b[101]  & new_new_n1188__;
  assign new_new_n1191__ = ~new_new_n1189__ & ~new_new_n1190__;
  assign new_new_n1192__ = \a[101]  & ~new_new_n1191__;
  assign new_new_n1193__ = ~\a[101]  & new_new_n1191__;
  assign \f[101]  = new_new_n1192__ | new_new_n1193__;
  assign new_new_n1195__ = ~\a[101]  & ~new_new_n1190__;
  assign new_new_n1196__ = ~new_new_n1189__ & ~new_new_n1195__;
  assign new_new_n1197__ = ~\a[102]  & ~\b[102] ;
  assign new_new_n1198__ = \a[102]  & \b[102] ;
  assign new_new_n1199__ = ~new_new_n1197__ & ~new_new_n1198__;
  assign new_new_n1200__ = ~new_new_n1196__ & new_new_n1199__;
  assign new_new_n1201__ = new_new_n1196__ & ~new_new_n1199__;
  assign \f[102]  = new_new_n1200__ | new_new_n1201__;
  assign new_new_n1203__ = ~new_new_n1196__ & ~new_new_n1198__;
  assign new_new_n1204__ = ~new_new_n1197__ & ~new_new_n1203__;
  assign new_new_n1205__ = ~\b[103]  & ~new_new_n1204__;
  assign new_new_n1206__ = \b[103]  & new_new_n1204__;
  assign new_new_n1207__ = ~new_new_n1205__ & ~new_new_n1206__;
  assign new_new_n1208__ = \a[103]  & ~new_new_n1207__;
  assign new_new_n1209__ = ~\a[103]  & new_new_n1207__;
  assign \f[103]  = new_new_n1208__ | new_new_n1209__;
  assign new_new_n1211__ = ~\a[103]  & ~new_new_n1206__;
  assign new_new_n1212__ = ~new_new_n1205__ & ~new_new_n1211__;
  assign new_new_n1213__ = ~\a[104]  & ~\b[104] ;
  assign new_new_n1214__ = \a[104]  & \b[104] ;
  assign new_new_n1215__ = ~new_new_n1213__ & ~new_new_n1214__;
  assign new_new_n1216__ = ~new_new_n1212__ & new_new_n1215__;
  assign new_new_n1217__ = new_new_n1212__ & ~new_new_n1215__;
  assign \f[104]  = new_new_n1216__ | new_new_n1217__;
  assign new_new_n1219__ = ~new_new_n1212__ & ~new_new_n1214__;
  assign new_new_n1220__ = ~new_new_n1213__ & ~new_new_n1219__;
  assign new_new_n1221__ = ~\b[105]  & ~new_new_n1220__;
  assign new_new_n1222__ = \b[105]  & new_new_n1220__;
  assign new_new_n1223__ = ~new_new_n1221__ & ~new_new_n1222__;
  assign new_new_n1224__ = \a[105]  & ~new_new_n1223__;
  assign new_new_n1225__ = ~\a[105]  & new_new_n1223__;
  assign \f[105]  = new_new_n1224__ | new_new_n1225__;
  assign new_new_n1227__ = ~\a[105]  & ~new_new_n1222__;
  assign new_new_n1228__ = ~new_new_n1221__ & ~new_new_n1227__;
  assign new_new_n1229__ = ~\a[106]  & ~\b[106] ;
  assign new_new_n1230__ = \a[106]  & \b[106] ;
  assign new_new_n1231__ = ~new_new_n1229__ & ~new_new_n1230__;
  assign new_new_n1232__ = ~new_new_n1228__ & new_new_n1231__;
  assign new_new_n1233__ = new_new_n1228__ & ~new_new_n1231__;
  assign \f[106]  = new_new_n1232__ | new_new_n1233__;
  assign new_new_n1235__ = ~new_new_n1228__ & ~new_new_n1230__;
  assign new_new_n1236__ = ~new_new_n1229__ & ~new_new_n1235__;
  assign new_new_n1237__ = ~\b[107]  & ~new_new_n1236__;
  assign new_new_n1238__ = \b[107]  & new_new_n1236__;
  assign new_new_n1239__ = ~new_new_n1237__ & ~new_new_n1238__;
  assign new_new_n1240__ = \a[107]  & ~new_new_n1239__;
  assign new_new_n1241__ = ~\a[107]  & new_new_n1239__;
  assign \f[107]  = new_new_n1240__ | new_new_n1241__;
  assign new_new_n1243__ = ~\a[107]  & ~new_new_n1238__;
  assign new_new_n1244__ = ~new_new_n1237__ & ~new_new_n1243__;
  assign new_new_n1245__ = ~\a[108]  & ~\b[108] ;
  assign new_new_n1246__ = \a[108]  & \b[108] ;
  assign new_new_n1247__ = ~new_new_n1245__ & ~new_new_n1246__;
  assign new_new_n1248__ = ~new_new_n1244__ & new_new_n1247__;
  assign new_new_n1249__ = new_new_n1244__ & ~new_new_n1247__;
  assign \f[108]  = new_new_n1248__ | new_new_n1249__;
  assign new_new_n1251__ = ~new_new_n1244__ & ~new_new_n1246__;
  assign new_new_n1252__ = ~new_new_n1245__ & ~new_new_n1251__;
  assign new_new_n1253__ = ~\b[109]  & ~new_new_n1252__;
  assign new_new_n1254__ = \b[109]  & new_new_n1252__;
  assign new_new_n1255__ = ~new_new_n1253__ & ~new_new_n1254__;
  assign new_new_n1256__ = \a[109]  & ~new_new_n1255__;
  assign new_new_n1257__ = ~\a[109]  & new_new_n1255__;
  assign \f[109]  = new_new_n1256__ | new_new_n1257__;
  assign new_new_n1259__ = ~\a[109]  & ~new_new_n1254__;
  assign new_new_n1260__ = ~new_new_n1253__ & ~new_new_n1259__;
  assign new_new_n1261__ = ~\a[110]  & ~\b[110] ;
  assign new_new_n1262__ = \a[110]  & \b[110] ;
  assign new_new_n1263__ = ~new_new_n1261__ & ~new_new_n1262__;
  assign new_new_n1264__ = ~new_new_n1260__ & new_new_n1263__;
  assign new_new_n1265__ = new_new_n1260__ & ~new_new_n1263__;
  assign \f[110]  = new_new_n1264__ | new_new_n1265__;
  assign new_new_n1267__ = ~new_new_n1260__ & ~new_new_n1262__;
  assign new_new_n1268__ = ~new_new_n1261__ & ~new_new_n1267__;
  assign new_new_n1269__ = ~\b[111]  & ~new_new_n1268__;
  assign new_new_n1270__ = \b[111]  & new_new_n1268__;
  assign new_new_n1271__ = ~new_new_n1269__ & ~new_new_n1270__;
  assign new_new_n1272__ = \a[111]  & ~new_new_n1271__;
  assign new_new_n1273__ = ~\a[111]  & new_new_n1271__;
  assign \f[111]  = new_new_n1272__ | new_new_n1273__;
  assign new_new_n1275__ = ~\a[111]  & ~new_new_n1270__;
  assign new_new_n1276__ = ~new_new_n1269__ & ~new_new_n1275__;
  assign new_new_n1277__ = ~\a[112]  & ~\b[112] ;
  assign new_new_n1278__ = \a[112]  & \b[112] ;
  assign new_new_n1279__ = ~new_new_n1277__ & ~new_new_n1278__;
  assign new_new_n1280__ = ~new_new_n1276__ & new_new_n1279__;
  assign new_new_n1281__ = new_new_n1276__ & ~new_new_n1279__;
  assign \f[112]  = new_new_n1280__ | new_new_n1281__;
  assign new_new_n1283__ = ~new_new_n1276__ & ~new_new_n1278__;
  assign new_new_n1284__ = ~new_new_n1277__ & ~new_new_n1283__;
  assign new_new_n1285__ = ~\b[113]  & ~new_new_n1284__;
  assign new_new_n1286__ = \b[113]  & new_new_n1284__;
  assign new_new_n1287__ = ~new_new_n1285__ & ~new_new_n1286__;
  assign new_new_n1288__ = \a[113]  & ~new_new_n1287__;
  assign new_new_n1289__ = ~\a[113]  & new_new_n1287__;
  assign \f[113]  = new_new_n1288__ | new_new_n1289__;
  assign new_new_n1291__ = ~\a[113]  & ~new_new_n1286__;
  assign new_new_n1292__ = ~new_new_n1285__ & ~new_new_n1291__;
  assign new_new_n1293__ = ~\a[114]  & ~\b[114] ;
  assign new_new_n1294__ = \a[114]  & \b[114] ;
  assign new_new_n1295__ = ~new_new_n1293__ & ~new_new_n1294__;
  assign new_new_n1296__ = ~new_new_n1292__ & new_new_n1295__;
  assign new_new_n1297__ = new_new_n1292__ & ~new_new_n1295__;
  assign \f[114]  = new_new_n1296__ | new_new_n1297__;
  assign new_new_n1299__ = ~new_new_n1292__ & ~new_new_n1294__;
  assign new_new_n1300__ = ~new_new_n1293__ & ~new_new_n1299__;
  assign new_new_n1301__ = ~\b[115]  & ~new_new_n1300__;
  assign new_new_n1302__ = \b[115]  & new_new_n1300__;
  assign new_new_n1303__ = ~new_new_n1301__ & ~new_new_n1302__;
  assign new_new_n1304__ = \a[115]  & ~new_new_n1303__;
  assign new_new_n1305__ = ~\a[115]  & new_new_n1303__;
  assign \f[115]  = new_new_n1304__ | new_new_n1305__;
  assign new_new_n1307__ = ~\a[115]  & ~new_new_n1302__;
  assign new_new_n1308__ = ~new_new_n1301__ & ~new_new_n1307__;
  assign new_new_n1309__ = ~\a[116]  & ~\b[116] ;
  assign new_new_n1310__ = \a[116]  & \b[116] ;
  assign new_new_n1311__ = ~new_new_n1309__ & ~new_new_n1310__;
  assign new_new_n1312__ = ~new_new_n1308__ & new_new_n1311__;
  assign new_new_n1313__ = new_new_n1308__ & ~new_new_n1311__;
  assign \f[116]  = new_new_n1312__ | new_new_n1313__;
  assign new_new_n1315__ = ~new_new_n1308__ & ~new_new_n1310__;
  assign new_new_n1316__ = ~new_new_n1309__ & ~new_new_n1315__;
  assign new_new_n1317__ = ~\b[117]  & ~new_new_n1316__;
  assign new_new_n1318__ = \b[117]  & new_new_n1316__;
  assign new_new_n1319__ = ~new_new_n1317__ & ~new_new_n1318__;
  assign new_new_n1320__ = \a[117]  & ~new_new_n1319__;
  assign new_new_n1321__ = ~\a[117]  & new_new_n1319__;
  assign \f[117]  = new_new_n1320__ | new_new_n1321__;
  assign new_new_n1323__ = ~\a[117]  & ~new_new_n1318__;
  assign new_new_n1324__ = ~new_new_n1317__ & ~new_new_n1323__;
  assign new_new_n1325__ = ~\a[118]  & ~\b[118] ;
  assign new_new_n1326__ = \a[118]  & \b[118] ;
  assign new_new_n1327__ = ~new_new_n1325__ & ~new_new_n1326__;
  assign new_new_n1328__ = ~new_new_n1324__ & new_new_n1327__;
  assign new_new_n1329__ = new_new_n1324__ & ~new_new_n1327__;
  assign \f[118]  = new_new_n1328__ | new_new_n1329__;
  assign new_new_n1331__ = ~new_new_n1324__ & ~new_new_n1326__;
  assign new_new_n1332__ = ~new_new_n1325__ & ~new_new_n1331__;
  assign new_new_n1333__ = ~\b[119]  & ~new_new_n1332__;
  assign new_new_n1334__ = \b[119]  & new_new_n1332__;
  assign new_new_n1335__ = ~new_new_n1333__ & ~new_new_n1334__;
  assign new_new_n1336__ = \a[119]  & ~new_new_n1335__;
  assign new_new_n1337__ = ~\a[119]  & new_new_n1335__;
  assign \f[119]  = new_new_n1336__ | new_new_n1337__;
  assign new_new_n1339__ = ~\a[119]  & ~new_new_n1334__;
  assign new_new_n1340__ = ~new_new_n1333__ & ~new_new_n1339__;
  assign new_new_n1341__ = ~\a[120]  & ~\b[120] ;
  assign new_new_n1342__ = \a[120]  & \b[120] ;
  assign new_new_n1343__ = ~new_new_n1341__ & ~new_new_n1342__;
  assign new_new_n1344__ = ~new_new_n1340__ & new_new_n1343__;
  assign new_new_n1345__ = new_new_n1340__ & ~new_new_n1343__;
  assign \f[120]  = new_new_n1344__ | new_new_n1345__;
  assign new_new_n1347__ = ~new_new_n1340__ & ~new_new_n1342__;
  assign new_new_n1348__ = ~new_new_n1341__ & ~new_new_n1347__;
  assign new_new_n1349__ = ~\b[121]  & ~new_new_n1348__;
  assign new_new_n1350__ = \b[121]  & new_new_n1348__;
  assign new_new_n1351__ = ~new_new_n1349__ & ~new_new_n1350__;
  assign new_new_n1352__ = \a[121]  & ~new_new_n1351__;
  assign new_new_n1353__ = ~\a[121]  & new_new_n1351__;
  assign \f[121]  = new_new_n1352__ | new_new_n1353__;
  assign new_new_n1355__ = ~\a[121]  & ~new_new_n1350__;
  assign new_new_n1356__ = ~new_new_n1349__ & ~new_new_n1355__;
  assign new_new_n1357__ = ~\a[122]  & ~\b[122] ;
  assign new_new_n1358__ = \a[122]  & \b[122] ;
  assign new_new_n1359__ = ~new_new_n1357__ & ~new_new_n1358__;
  assign new_new_n1360__ = ~new_new_n1356__ & new_new_n1359__;
  assign new_new_n1361__ = new_new_n1356__ & ~new_new_n1359__;
  assign \f[122]  = new_new_n1360__ | new_new_n1361__;
  assign new_new_n1363__ = ~new_new_n1356__ & ~new_new_n1358__;
  assign new_new_n1364__ = ~new_new_n1357__ & ~new_new_n1363__;
  assign new_new_n1365__ = ~\b[123]  & ~new_new_n1364__;
  assign new_new_n1366__ = \b[123]  & new_new_n1364__;
  assign new_new_n1367__ = ~new_new_n1365__ & ~new_new_n1366__;
  assign new_new_n1368__ = \a[123]  & ~new_new_n1367__;
  assign new_new_n1369__ = ~\a[123]  & new_new_n1367__;
  assign \f[123]  = new_new_n1368__ | new_new_n1369__;
  assign new_new_n1371__ = ~\a[123]  & ~new_new_n1366__;
  assign new_new_n1372__ = ~new_new_n1365__ & ~new_new_n1371__;
  assign new_new_n1373__ = ~\a[124]  & ~\b[124] ;
  assign new_new_n1374__ = \a[124]  & \b[124] ;
  assign new_new_n1375__ = ~new_new_n1373__ & ~new_new_n1374__;
  assign new_new_n1376__ = ~new_new_n1372__ & new_new_n1375__;
  assign new_new_n1377__ = new_new_n1372__ & ~new_new_n1375__;
  assign \f[124]  = new_new_n1376__ | new_new_n1377__;
  assign new_new_n1379__ = ~new_new_n1372__ & ~new_new_n1374__;
  assign new_new_n1380__ = ~new_new_n1373__ & ~new_new_n1379__;
  assign new_new_n1381__ = ~\b[125]  & ~new_new_n1380__;
  assign new_new_n1382__ = \b[125]  & new_new_n1380__;
  assign new_new_n1383__ = ~new_new_n1381__ & ~new_new_n1382__;
  assign new_new_n1384__ = \a[125]  & ~new_new_n1383__;
  assign new_new_n1385__ = ~\a[125]  & new_new_n1383__;
  assign \f[125]  = new_new_n1384__ | new_new_n1385__;
  assign new_new_n1387__ = ~\a[125]  & ~new_new_n1382__;
  assign new_new_n1388__ = ~new_new_n1381__ & ~new_new_n1387__;
  assign new_new_n1389__ = \a[126]  & \b[126] ;
  assign new_new_n1390__ = ~\a[126]  & ~\b[126] ;
  assign new_new_n1391__ = ~new_new_n1389__ & ~new_new_n1390__;
  assign new_new_n1392__ = new_new_n1388__ & ~new_new_n1391__;
  assign new_new_n1393__ = ~new_new_n1388__ & new_new_n1391__;
  assign \f[126]  = new_new_n1392__ | new_new_n1393__;
  assign new_new_n1395__ = \a[127]  & \b[127] ;
  assign new_new_n1396__ = ~\a[127]  & ~\b[127] ;
  assign new_new_n1397__ = ~new_new_n1395__ & ~new_new_n1396__;
  assign new_new_n1398__ = ~new_new_n1388__ & ~new_new_n1389__;
  assign new_new_n1399__ = ~new_new_n1390__ & ~new_new_n1398__;
  assign new_new_n1400__ = new_new_n1397__ & ~new_new_n1399__;
  assign new_new_n1401__ = ~new_new_n1397__ & new_new_n1399__;
  assign \f[127]  = new_new_n1400__ | new_new_n1401__;
  assign new_new_n1403__ = ~new_new_n1395__ & ~new_new_n1399__;
  assign cOut = ~new_new_n1396__ & ~new_new_n1403__;
endmodule


