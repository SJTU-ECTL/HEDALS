// Benchmark "sin" written by ABC on Wed Jul 13 18:49:26 2022

module sin ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24;
  wire new_new_n50__, new_new_n51__, new_new_n52__, new_new_n53__,
    new_new_n54__, new_new_n55__, new_new_n56__, new_new_n57__,
    new_new_n58__, new_new_n59__, new_new_n60__, new_new_n61__,
    new_new_n62__, new_new_n63__, new_new_n64__, new_new_n65__,
    new_new_n66__, new_new_n67__, new_new_n68__, new_new_n69__,
    new_new_n70__, new_new_n71__, new_new_n72__, new_new_n73__,
    new_new_n74__, new_new_n75__, new_new_n76__, new_new_n77__,
    new_new_n78__, new_new_n79__, new_new_n80__, new_new_n81__,
    new_new_n82__, new_new_n83__, new_new_n84__, new_new_n85__,
    new_new_n86__, new_new_n87__, new_new_n88__, new_new_n89__,
    new_new_n90__, new_new_n91__, new_new_n92__, new_new_n93__,
    new_new_n94__, new_new_n95__, new_new_n96__, new_new_n97__,
    new_new_n98__, new_new_n99__, new_new_n100__, new_new_n101__,
    new_new_n102__, new_new_n103__, new_new_n104__, new_new_n105__,
    new_new_n106__, new_new_n107__, new_new_n108__, new_new_n109__,
    new_new_n110__, new_new_n111__, new_new_n112__, new_new_n113__,
    new_new_n114__, new_new_n115__, new_new_n116__, new_new_n117__,
    new_new_n118__, new_new_n119__, new_new_n120__, new_new_n121__,
    new_new_n122__, new_new_n123__, new_new_n124__, new_new_n125__,
    new_new_n126__, new_new_n127__, new_new_n128__, new_new_n129__,
    new_new_n130__, new_new_n131__, new_new_n132__, new_new_n133__,
    new_new_n134__, new_new_n135__, new_new_n136__, new_new_n137__,
    new_new_n138__, new_new_n139__, new_new_n140__, new_new_n141__,
    new_new_n142__, new_new_n143__, new_new_n144__, new_new_n145__,
    new_new_n146__, new_new_n147__, new_new_n148__, new_new_n149__,
    new_new_n150__, new_new_n151__, new_new_n152__, new_new_n153__,
    new_new_n154__, new_new_n155__, new_new_n156__, new_new_n157__,
    new_new_n158__, new_new_n159__, new_new_n160__, new_new_n161__,
    new_new_n162__, new_new_n163__, new_new_n164__, new_new_n165__,
    new_new_n166__, new_new_n167__, new_new_n168__, new_new_n169__,
    new_new_n170__, new_new_n171__, new_new_n172__, new_new_n173__,
    new_new_n174__, new_new_n175__, new_new_n176__, new_new_n177__,
    new_new_n178__, new_new_n179__, new_new_n180__, new_new_n181__,
    new_new_n182__, new_new_n183__, new_new_n184__, new_new_n185__,
    new_new_n186__, new_new_n187__, new_new_n188__, new_new_n189__,
    new_new_n190__, new_new_n191__, new_new_n192__, new_new_n193__,
    new_new_n194__, new_new_n195__, new_new_n196__, new_new_n197__,
    new_new_n198__, new_new_n199__, new_new_n200__, new_new_n201__,
    new_new_n202__, new_new_n203__, new_new_n204__, new_new_n205__,
    new_new_n206__, new_new_n207__, new_new_n208__, new_new_n209__,
    new_new_n210__, new_new_n211__, new_new_n212__, new_new_n213__,
    new_new_n214__, new_new_n215__, new_new_n216__, new_new_n217__,
    new_new_n218__, new_new_n219__, new_new_n220__, new_new_n221__,
    new_new_n222__, new_new_n223__, new_new_n224__, new_new_n225__,
    new_new_n226__, new_new_n227__, new_new_n228__, new_new_n229__,
    new_new_n230__, new_new_n231__, new_new_n232__, new_new_n233__,
    new_new_n234__, new_new_n235__, new_new_n236__, new_new_n237__,
    new_new_n238__, new_new_n239__, new_new_n240__, new_new_n241__,
    new_new_n242__, new_new_n243__, new_new_n244__, new_new_n245__,
    new_new_n246__, new_new_n247__, new_new_n248__, new_new_n249__,
    new_new_n250__, new_new_n251__, new_new_n252__, new_new_n253__,
    new_new_n254__, new_new_n255__, new_new_n256__, new_new_n257__,
    new_new_n258__, new_new_n259__, new_new_n260__, new_new_n261__,
    new_new_n262__, new_new_n263__, new_new_n264__, new_new_n265__,
    new_new_n266__, new_new_n267__, new_new_n268__, new_new_n269__,
    new_new_n270__, new_new_n271__, new_new_n272__, new_new_n273__,
    new_new_n274__, new_new_n275__, new_new_n276__, new_new_n277__,
    new_new_n278__, new_new_n279__, new_new_n280__, new_new_n281__,
    new_new_n282__, new_new_n283__, new_new_n284__, new_new_n285__,
    new_new_n286__, new_new_n287__, new_new_n288__, new_new_n289__,
    new_new_n290__, new_new_n291__, new_new_n292__, new_new_n293__,
    new_new_n294__, new_new_n295__, new_new_n296__, new_new_n297__,
    new_new_n298__, new_new_n299__, new_new_n300__, new_new_n301__,
    new_new_n302__, new_new_n303__, new_new_n304__, new_new_n305__,
    new_new_n306__, new_new_n307__, new_new_n308__, new_new_n309__,
    new_new_n310__, new_new_n311__, new_new_n312__, new_new_n313__,
    new_new_n314__, new_new_n315__, new_new_n316__, new_new_n317__,
    new_new_n318__, new_new_n319__, new_new_n320__, new_new_n321__,
    new_new_n322__, new_new_n323__, new_new_n324__, new_new_n325__,
    new_new_n326__, new_new_n327__, new_new_n328__, new_new_n329__,
    new_new_n330__, new_new_n331__, new_new_n332__, new_new_n333__,
    new_new_n334__, new_new_n335__, new_new_n336__, new_new_n337__,
    new_new_n338__, new_new_n339__, new_new_n340__, new_new_n341__,
    new_new_n342__, new_new_n343__, new_new_n344__, new_new_n345__,
    new_new_n346__, new_new_n347__, new_new_n348__, new_new_n349__,
    new_new_n350__, new_new_n351__, new_new_n352__, new_new_n353__,
    new_new_n354__, new_new_n355__, new_new_n356__, new_new_n357__,
    new_new_n358__, new_new_n359__, new_new_n360__, new_new_n361__,
    new_new_n362__, new_new_n363__, new_new_n364__, new_new_n365__,
    new_new_n366__, new_new_n367__, new_new_n368__, new_new_n369__,
    new_new_n370__, new_new_n371__, new_new_n372__, new_new_n373__,
    new_new_n374__, new_new_n375__, new_new_n376__, new_new_n377__,
    new_new_n378__, new_new_n379__, new_new_n380__, new_new_n381__,
    new_new_n382__, new_new_n383__, new_new_n384__, new_new_n385__,
    new_new_n386__, new_new_n387__, new_new_n388__, new_new_n389__,
    new_new_n390__, new_new_n391__, new_new_n392__, new_new_n393__,
    new_new_n394__, new_new_n395__, new_new_n396__, new_new_n397__,
    new_new_n398__, new_new_n399__, new_new_n400__, new_new_n401__,
    new_new_n402__, new_new_n403__, new_new_n404__, new_new_n405__,
    new_new_n406__, new_new_n407__, new_new_n408__, new_new_n409__,
    new_new_n410__, new_new_n411__, new_new_n412__, new_new_n413__,
    new_new_n414__, new_new_n415__, new_new_n416__, new_new_n417__,
    new_new_n418__, new_new_n419__, new_new_n420__, new_new_n421__,
    new_new_n422__, new_new_n423__, new_new_n424__, new_new_n425__,
    new_new_n426__, new_new_n427__, new_new_n428__, new_new_n429__,
    new_new_n430__, new_new_n431__, new_new_n432__, new_new_n433__,
    new_new_n434__, new_new_n435__, new_new_n436__, new_new_n437__,
    new_new_n438__, new_new_n439__, new_new_n440__, new_new_n441__,
    new_new_n442__, new_new_n443__, new_new_n444__, new_new_n445__,
    new_new_n446__, new_new_n447__, new_new_n448__, new_new_n449__,
    new_new_n450__, new_new_n451__, new_new_n452__, new_new_n453__,
    new_new_n454__, new_new_n455__, new_new_n456__, new_new_n457__,
    new_new_n458__, new_new_n459__, new_new_n460__, new_new_n461__,
    new_new_n462__, new_new_n463__, new_new_n464__, new_new_n465__,
    new_new_n466__, new_new_n467__, new_new_n468__, new_new_n469__,
    new_new_n470__, new_new_n471__, new_new_n472__, new_new_n473__,
    new_new_n474__, new_new_n475__, new_new_n476__, new_new_n477__,
    new_new_n478__, new_new_n479__, new_new_n480__, new_new_n481__,
    new_new_n482__, new_new_n483__, new_new_n484__, new_new_n485__,
    new_new_n486__, new_new_n487__, new_new_n488__, new_new_n489__,
    new_new_n490__, new_new_n491__, new_new_n492__, new_new_n493__,
    new_new_n494__, new_new_n495__, new_new_n496__, new_new_n497__,
    new_new_n498__, new_new_n499__, new_new_n500__, new_new_n501__,
    new_new_n502__, new_new_n503__, new_new_n504__, new_new_n505__,
    new_new_n506__, new_new_n507__, new_new_n508__, new_new_n509__,
    new_new_n510__, new_new_n511__, new_new_n512__, new_new_n513__,
    new_new_n514__, new_new_n515__, new_new_n516__, new_new_n517__,
    new_new_n518__, new_new_n519__, new_new_n520__, new_new_n521__,
    new_new_n522__, new_new_n523__, new_new_n524__, new_new_n525__,
    new_new_n526__, new_new_n527__, new_new_n528__, new_new_n529__,
    new_new_n530__, new_new_n531__, new_new_n532__, new_new_n533__,
    new_new_n534__, new_new_n535__, new_new_n536__, new_new_n537__,
    new_new_n538__, new_new_n539__, new_new_n540__, new_new_n541__,
    new_new_n542__, new_new_n543__, new_new_n544__, new_new_n545__,
    new_new_n546__, new_new_n547__, new_new_n548__, new_new_n549__,
    new_new_n550__, new_new_n551__, new_new_n552__, new_new_n553__,
    new_new_n554__, new_new_n555__, new_new_n556__, new_new_n557__,
    new_new_n558__, new_new_n559__, new_new_n560__, new_new_n561__,
    new_new_n562__, new_new_n563__, new_new_n564__, new_new_n565__,
    new_new_n566__, new_new_n567__, new_new_n568__, new_new_n569__,
    new_new_n570__, new_new_n571__, new_new_n572__, new_new_n573__,
    new_new_n574__, new_new_n575__, new_new_n576__, new_new_n577__,
    new_new_n578__, new_new_n579__, new_new_n580__, new_new_n581__,
    new_new_n582__, new_new_n583__, new_new_n584__, new_new_n585__,
    new_new_n586__, new_new_n587__, new_new_n588__, new_new_n589__,
    new_new_n590__, new_new_n591__, new_new_n592__, new_new_n593__,
    new_new_n594__, new_new_n595__, new_new_n596__, new_new_n597__,
    new_new_n598__, new_new_n599__, new_new_n600__, new_new_n601__,
    new_new_n602__, new_new_n603__, new_new_n604__, new_new_n605__,
    new_new_n606__, new_new_n607__, new_new_n608__, new_new_n609__,
    new_new_n610__, new_new_n611__, new_new_n612__, new_new_n613__,
    new_new_n614__, new_new_n615__, new_new_n616__, new_new_n617__,
    new_new_n618__, new_new_n619__, new_new_n620__, new_new_n621__,
    new_new_n622__, new_new_n623__, new_new_n624__, new_new_n625__,
    new_new_n626__, new_new_n627__, new_new_n628__, new_new_n629__,
    new_new_n630__, new_new_n631__, new_new_n632__, new_new_n633__,
    new_new_n634__, new_new_n635__, new_new_n636__, new_new_n637__,
    new_new_n638__, new_new_n639__, new_new_n640__, new_new_n641__,
    new_new_n642__, new_new_n643__, new_new_n644__, new_new_n645__,
    new_new_n646__, new_new_n647__, new_new_n648__, new_new_n649__,
    new_new_n650__, new_new_n651__, new_new_n652__, new_new_n653__,
    new_new_n654__, new_new_n655__, new_new_n656__, new_new_n657__,
    new_new_n658__, new_new_n659__, new_new_n660__, new_new_n661__,
    new_new_n662__, new_new_n663__, new_new_n664__, new_new_n665__,
    new_new_n666__, new_new_n667__, new_new_n668__, new_new_n669__,
    new_new_n670__, new_new_n671__, new_new_n672__, new_new_n673__,
    new_new_n674__, new_new_n675__, new_new_n676__, new_new_n677__,
    new_new_n678__, new_new_n679__, new_new_n680__, new_new_n681__,
    new_new_n682__, new_new_n683__, new_new_n684__, new_new_n685__,
    new_new_n686__, new_new_n687__, new_new_n688__, new_new_n689__,
    new_new_n690__, new_new_n691__, new_new_n692__, new_new_n693__,
    new_new_n694__, new_new_n695__, new_new_n696__, new_new_n697__,
    new_new_n698__, new_new_n699__, new_new_n700__, new_new_n701__,
    new_new_n702__, new_new_n703__, new_new_n704__, new_new_n705__,
    new_new_n706__, new_new_n707__, new_new_n708__, new_new_n709__,
    new_new_n710__, new_new_n711__, new_new_n712__, new_new_n713__,
    new_new_n714__, new_new_n715__, new_new_n716__, new_new_n717__,
    new_new_n718__, new_new_n719__, new_new_n720__, new_new_n721__,
    new_new_n722__, new_new_n723__, new_new_n724__, new_new_n725__,
    new_new_n726__, new_new_n727__, new_new_n728__, new_new_n729__,
    new_new_n730__, new_new_n731__, new_new_n732__, new_new_n733__,
    new_new_n734__, new_new_n735__, new_new_n736__, new_new_n737__,
    new_new_n738__, new_new_n739__, new_new_n740__, new_new_n741__,
    new_new_n742__, new_new_n743__, new_new_n744__, new_new_n745__,
    new_new_n746__, new_new_n747__, new_new_n748__, new_new_n749__,
    new_new_n750__, new_new_n751__, new_new_n752__, new_new_n753__,
    new_new_n754__, new_new_n755__, new_new_n756__, new_new_n757__,
    new_new_n758__, new_new_n759__, new_new_n760__, new_new_n761__,
    new_new_n762__, new_new_n763__, new_new_n764__, new_new_n765__,
    new_new_n766__, new_new_n767__, new_new_n768__, new_new_n769__,
    new_new_n770__, new_new_n771__, new_new_n772__, new_new_n773__,
    new_new_n774__, new_new_n775__, new_new_n776__, new_new_n777__,
    new_new_n778__, new_new_n779__, new_new_n780__, new_new_n781__,
    new_new_n782__, new_new_n783__, new_new_n784__, new_new_n785__,
    new_new_n786__, new_new_n787__, new_new_n788__, new_new_n789__,
    new_new_n790__, new_new_n791__, new_new_n792__, new_new_n793__,
    new_new_n794__, new_new_n795__, new_new_n796__, new_new_n797__,
    new_new_n798__, new_new_n799__, new_new_n800__, new_new_n801__,
    new_new_n802__, new_new_n803__, new_new_n804__, new_new_n805__,
    new_new_n806__, new_new_n807__, new_new_n808__, new_new_n809__,
    new_new_n810__, new_new_n811__, new_new_n812__, new_new_n813__,
    new_new_n814__, new_new_n815__, new_new_n816__, new_new_n817__,
    new_new_n818__, new_new_n819__, new_new_n820__, new_new_n821__,
    new_new_n822__, new_new_n823__, new_new_n824__, new_new_n825__,
    new_new_n826__, new_new_n827__, new_new_n828__, new_new_n829__,
    new_new_n830__, new_new_n831__, new_new_n832__, new_new_n833__,
    new_new_n834__, new_new_n835__, new_new_n836__, new_new_n837__,
    new_new_n838__, new_new_n839__, new_new_n840__, new_new_n841__,
    new_new_n842__, new_new_n843__, new_new_n844__, new_new_n845__,
    new_new_n846__, new_new_n847__, new_new_n848__, new_new_n849__,
    new_new_n850__, new_new_n851__, new_new_n852__, new_new_n853__,
    new_new_n854__, new_new_n855__, new_new_n856__, new_new_n857__,
    new_new_n858__, new_new_n859__, new_new_n860__, new_new_n861__,
    new_new_n862__, new_new_n863__, new_new_n864__, new_new_n865__,
    new_new_n866__, new_new_n867__, new_new_n868__, new_new_n869__,
    new_new_n870__, new_new_n871__, new_new_n872__, new_new_n873__,
    new_new_n874__, new_new_n875__, new_new_n876__, new_new_n877__,
    new_new_n878__, new_new_n879__, new_new_n880__, new_new_n881__,
    new_new_n882__, new_new_n883__, new_new_n884__, new_new_n885__,
    new_new_n886__, new_new_n887__, new_new_n888__, new_new_n889__,
    new_new_n890__, new_new_n891__, new_new_n892__, new_new_n893__,
    new_new_n894__, new_new_n895__, new_new_n896__, new_new_n897__,
    new_new_n898__, new_new_n899__, new_new_n900__, new_new_n901__,
    new_new_n902__, new_new_n903__, new_new_n904__, new_new_n905__,
    new_new_n906__, new_new_n907__, new_new_n908__, new_new_n909__,
    new_new_n910__, new_new_n911__, new_new_n912__, new_new_n913__,
    new_new_n914__, new_new_n915__, new_new_n916__, new_new_n917__,
    new_new_n918__, new_new_n919__, new_new_n920__, new_new_n921__,
    new_new_n922__, new_new_n923__, new_new_n924__, new_new_n925__,
    new_new_n926__, new_new_n927__, new_new_n928__, new_new_n929__,
    new_new_n930__, new_new_n931__, new_new_n932__, new_new_n933__,
    new_new_n934__, new_new_n935__, new_new_n936__, new_new_n937__,
    new_new_n938__, new_new_n939__, new_new_n940__, new_new_n941__,
    new_new_n942__, new_new_n943__, new_new_n944__, new_new_n945__,
    new_new_n946__, new_new_n947__, new_new_n948__, new_new_n949__,
    new_new_n950__, new_new_n951__, new_new_n952__, new_new_n953__,
    new_new_n954__, new_new_n955__, new_new_n956__, new_new_n957__,
    new_new_n958__, new_new_n959__, new_new_n960__, new_new_n961__,
    new_new_n962__, new_new_n963__, new_new_n964__, new_new_n965__,
    new_new_n966__, new_new_n967__, new_new_n968__, new_new_n969__,
    new_new_n970__, new_new_n971__, new_new_n972__, new_new_n973__,
    new_new_n974__, new_new_n975__, new_new_n976__, new_new_n977__,
    new_new_n978__, new_new_n979__, new_new_n980__, new_new_n981__,
    new_new_n982__, new_new_n983__, new_new_n984__, new_new_n985__,
    new_new_n986__, new_new_n987__, new_new_n988__, new_new_n989__,
    new_new_n990__, new_new_n991__, new_new_n992__, new_new_n993__,
    new_new_n994__, new_new_n995__, new_new_n996__, new_new_n997__,
    new_new_n998__, new_new_n999__, new_new_n1000__, new_new_n1001__,
    new_new_n1002__, new_new_n1003__, new_new_n1004__, new_new_n1005__,
    new_new_n1006__, new_new_n1007__, new_new_n1008__, new_new_n1009__,
    new_new_n1010__, new_new_n1011__, new_new_n1012__, new_new_n1013__,
    new_new_n1014__, new_new_n1015__, new_new_n1016__, new_new_n1017__,
    new_new_n1018__, new_new_n1019__, new_new_n1020__, new_new_n1021__,
    new_new_n1022__, new_new_n1023__, new_new_n1024__, new_new_n1025__,
    new_new_n1026__, new_new_n1027__, new_new_n1028__, new_new_n1029__,
    new_new_n1030__, new_new_n1031__, new_new_n1032__, new_new_n1033__,
    new_new_n1034__, new_new_n1035__, new_new_n1036__, new_new_n1037__,
    new_new_n1038__, new_new_n1039__, new_new_n1040__, new_new_n1041__,
    new_new_n1042__, new_new_n1043__, new_new_n1044__, new_new_n1045__,
    new_new_n1046__, new_new_n1047__, new_new_n1048__, new_new_n1049__,
    new_new_n1050__, new_new_n1051__, new_new_n1052__, new_new_n1053__,
    new_new_n1054__, new_new_n1055__, new_new_n1056__, new_new_n1057__,
    new_new_n1058__, new_new_n1059__, new_new_n1060__, new_new_n1061__,
    new_new_n1062__, new_new_n1063__, new_new_n1064__, new_new_n1065__,
    new_new_n1066__, new_new_n1067__, new_new_n1068__, new_new_n1069__,
    new_new_n1070__, new_new_n1071__, new_new_n1072__, new_new_n1073__,
    new_new_n1074__, new_new_n1075__, new_new_n1076__, new_new_n1077__,
    new_new_n1078__, new_new_n1079__, new_new_n1080__, new_new_n1081__,
    new_new_n1082__, new_new_n1083__, new_new_n1084__, new_new_n1085__,
    new_new_n1086__, new_new_n1087__, new_new_n1088__, new_new_n1089__,
    new_new_n1090__, new_new_n1091__, new_new_n1092__, new_new_n1093__,
    new_new_n1094__, new_new_n1095__, new_new_n1096__, new_new_n1097__,
    new_new_n1098__, new_new_n1099__, new_new_n1100__, new_new_n1101__,
    new_new_n1102__, new_new_n1103__, new_new_n1104__, new_new_n1105__,
    new_new_n1106__, new_new_n1107__, new_new_n1108__, new_new_n1109__,
    new_new_n1110__, new_new_n1111__, new_new_n1112__, new_new_n1113__,
    new_new_n1114__, new_new_n1115__, new_new_n1116__, new_new_n1117__,
    new_new_n1118__, new_new_n1119__, new_new_n1120__, new_new_n1121__,
    new_new_n1122__, new_new_n1123__, new_new_n1124__, new_new_n1125__,
    new_new_n1126__, new_new_n1127__, new_new_n1128__, new_new_n1129__,
    new_new_n1130__, new_new_n1131__, new_new_n1132__, new_new_n1133__,
    new_new_n1134__, new_new_n1135__, new_new_n1136__, new_new_n1137__,
    new_new_n1138__, new_new_n1139__, new_new_n1140__, new_new_n1141__,
    new_new_n1142__, new_new_n1143__, new_new_n1144__, new_new_n1145__,
    new_new_n1146__, new_new_n1147__, new_new_n1148__, new_new_n1149__,
    new_new_n1150__, new_new_n1151__, new_new_n1152__, new_new_n1153__,
    new_new_n1154__, new_new_n1155__, new_new_n1156__, new_new_n1157__,
    new_new_n1158__, new_new_n1159__, new_new_n1160__, new_new_n1161__,
    new_new_n1162__, new_new_n1163__, new_new_n1164__, new_new_n1165__,
    new_new_n1166__, new_new_n1167__, new_new_n1168__, new_new_n1169__,
    new_new_n1170__, new_new_n1171__, new_new_n1172__, new_new_n1173__,
    new_new_n1174__, new_new_n1175__, new_new_n1176__, new_new_n1177__,
    new_new_n1178__, new_new_n1179__, new_new_n1180__, new_new_n1181__,
    new_new_n1182__, new_new_n1183__, new_new_n1184__, new_new_n1185__,
    new_new_n1186__, new_new_n1187__, new_new_n1188__, new_new_n1189__,
    new_new_n1190__, new_new_n1191__, new_new_n1192__, new_new_n1193__,
    new_new_n1194__, new_new_n1195__, new_new_n1196__, new_new_n1197__,
    new_new_n1198__, new_new_n1199__, new_new_n1200__, new_new_n1201__,
    new_new_n1202__, new_new_n1203__, new_new_n1204__, new_new_n1205__,
    new_new_n1206__, new_new_n1207__, new_new_n1208__, new_new_n1209__,
    new_new_n1210__, new_new_n1211__, new_new_n1212__, new_new_n1213__,
    new_new_n1214__, new_new_n1215__, new_new_n1216__, new_new_n1217__,
    new_new_n1218__, new_new_n1219__, new_new_n1220__, new_new_n1221__,
    new_new_n1222__, new_new_n1223__, new_new_n1224__, new_new_n1225__,
    new_new_n1226__, new_new_n1227__, new_new_n1228__, new_new_n1229__,
    new_new_n1230__, new_new_n1231__, new_new_n1232__, new_new_n1233__,
    new_new_n1234__, new_new_n1235__, new_new_n1236__, new_new_n1237__,
    new_new_n1238__, new_new_n1239__, new_new_n1240__, new_new_n1241__,
    new_new_n1242__, new_new_n1243__, new_new_n1244__, new_new_n1245__,
    new_new_n1246__, new_new_n1247__, new_new_n1248__, new_new_n1249__,
    new_new_n1250__, new_new_n1251__, new_new_n1252__, new_new_n1253__,
    new_new_n1254__, new_new_n1255__, new_new_n1256__, new_new_n1257__,
    new_new_n1258__, new_new_n1259__, new_new_n1260__, new_new_n1261__,
    new_new_n1262__, new_new_n1263__, new_new_n1264__, new_new_n1265__,
    new_new_n1266__, new_new_n1267__, new_new_n1268__, new_new_n1269__,
    new_new_n1270__, new_new_n1271__, new_new_n1272__, new_new_n1273__,
    new_new_n1274__, new_new_n1275__, new_new_n1276__, new_new_n1277__,
    new_new_n1278__, new_new_n1279__, new_new_n1280__, new_new_n1281__,
    new_new_n1282__, new_new_n1283__, new_new_n1284__, new_new_n1285__,
    new_new_n1286__, new_new_n1287__, new_new_n1288__, new_new_n1289__,
    new_new_n1290__, new_new_n1291__, new_new_n1292__, new_new_n1293__,
    new_new_n1294__, new_new_n1295__, new_new_n1296__, new_new_n1297__,
    new_new_n1298__, new_new_n1299__, new_new_n1300__, new_new_n1301__,
    new_new_n1302__, new_new_n1303__, new_new_n1304__, new_new_n1305__,
    new_new_n1306__, new_new_n1307__, new_new_n1308__, new_new_n1309__,
    new_new_n1310__, new_new_n1311__, new_new_n1312__, new_new_n1313__,
    new_new_n1314__, new_new_n1315__, new_new_n1316__, new_new_n1317__,
    new_new_n1318__, new_new_n1319__, new_new_n1320__, new_new_n1321__,
    new_new_n1322__, new_new_n1323__, new_new_n1324__, new_new_n1325__,
    new_new_n1326__, new_new_n1327__, new_new_n1328__, new_new_n1329__,
    new_new_n1330__, new_new_n1331__, new_new_n1332__, new_new_n1333__,
    new_new_n1334__, new_new_n1335__, new_new_n1336__, new_new_n1337__,
    new_new_n1338__, new_new_n1339__, new_new_n1340__, new_new_n1341__,
    new_new_n1342__, new_new_n1343__, new_new_n1344__, new_new_n1345__,
    new_new_n1346__, new_new_n1347__, new_new_n1348__, new_new_n1349__,
    new_new_n1350__, new_new_n1351__, new_new_n1352__, new_new_n1353__,
    new_new_n1354__, new_new_n1355__, new_new_n1356__, new_new_n1357__,
    new_new_n1358__, new_new_n1359__, new_new_n1360__, new_new_n1361__,
    new_new_n1362__, new_new_n1363__, new_new_n1364__, new_new_n1365__,
    new_new_n1366__, new_new_n1367__, new_new_n1368__, new_new_n1369__,
    new_new_n1370__, new_new_n1371__, new_new_n1372__, new_new_n1373__,
    new_new_n1374__, new_new_n1375__, new_new_n1376__, new_new_n1377__,
    new_new_n1378__, new_new_n1379__, new_new_n1380__, new_new_n1381__,
    new_new_n1382__, new_new_n1383__, new_new_n1384__, new_new_n1385__,
    new_new_n1386__, new_new_n1387__, new_new_n1388__, new_new_n1389__,
    new_new_n1390__, new_new_n1391__, new_new_n1392__, new_new_n1393__,
    new_new_n1394__, new_new_n1395__, new_new_n1396__, new_new_n1397__,
    new_new_n1398__, new_new_n1399__, new_new_n1400__, new_new_n1401__,
    new_new_n1402__, new_new_n1403__, new_new_n1404__, new_new_n1405__,
    new_new_n1406__, new_new_n1407__, new_new_n1408__, new_new_n1409__,
    new_new_n1410__, new_new_n1411__, new_new_n1412__, new_new_n1413__,
    new_new_n1414__, new_new_n1415__, new_new_n1416__, new_new_n1417__,
    new_new_n1418__, new_new_n1419__, new_new_n1420__, new_new_n1421__,
    new_new_n1422__, new_new_n1423__, new_new_n1424__, new_new_n1425__,
    new_new_n1426__, new_new_n1427__, new_new_n1428__, new_new_n1429__,
    new_new_n1430__, new_new_n1431__, new_new_n1432__, new_new_n1433__,
    new_new_n1434__, new_new_n1435__, new_new_n1436__, new_new_n1437__,
    new_new_n1438__, new_new_n1439__, new_new_n1440__, new_new_n1441__,
    new_new_n1442__, new_new_n1443__, new_new_n1444__, new_new_n1445__,
    new_new_n1446__, new_new_n1447__, new_new_n1448__, new_new_n1449__,
    new_new_n1450__, new_new_n1451__, new_new_n1452__, new_new_n1453__,
    new_new_n1454__, new_new_n1455__, new_new_n1456__, new_new_n1457__,
    new_new_n1458__, new_new_n1459__, new_new_n1460__, new_new_n1461__,
    new_new_n1462__, new_new_n1463__, new_new_n1464__, new_new_n1465__,
    new_new_n1466__, new_new_n1467__, new_new_n1468__, new_new_n1469__,
    new_new_n1470__, new_new_n1471__, new_new_n1472__, new_new_n1473__,
    new_new_n1474__, new_new_n1475__, new_new_n1476__, new_new_n1477__,
    new_new_n1478__, new_new_n1479__, new_new_n1480__, new_new_n1481__,
    new_new_n1482__, new_new_n1483__, new_new_n1484__, new_new_n1485__,
    new_new_n1486__, new_new_n1487__, new_new_n1488__, new_new_n1489__,
    new_new_n1490__, new_new_n1491__, new_new_n1492__, new_new_n1493__,
    new_new_n1494__, new_new_n1495__, new_new_n1496__, new_new_n1497__,
    new_new_n1498__, new_new_n1499__, new_new_n1500__, new_new_n1501__,
    new_new_n1502__, new_new_n1503__, new_new_n1504__, new_new_n1505__,
    new_new_n1506__, new_new_n1507__, new_new_n1508__, new_new_n1509__,
    new_new_n1510__, new_new_n1511__, new_new_n1512__, new_new_n1513__,
    new_new_n1514__, new_new_n1515__, new_new_n1516__, new_new_n1517__,
    new_new_n1518__, new_new_n1519__, new_new_n1520__, new_new_n1521__,
    new_new_n1522__, new_new_n1523__, new_new_n1524__, new_new_n1525__,
    new_new_n1526__, new_new_n1527__, new_new_n1528__, new_new_n1529__,
    new_new_n1530__, new_new_n1531__, new_new_n1532__, new_new_n1533__,
    new_new_n1534__, new_new_n1535__, new_new_n1536__, new_new_n1537__,
    new_new_n1538__, new_new_n1539__, new_new_n1540__, new_new_n1541__,
    new_new_n1542__, new_new_n1543__, new_new_n1544__, new_new_n1545__,
    new_new_n1546__, new_new_n1547__, new_new_n1548__, new_new_n1549__,
    new_new_n1550__, new_new_n1551__, new_new_n1552__, new_new_n1553__,
    new_new_n1554__, new_new_n1555__, new_new_n1556__, new_new_n1557__,
    new_new_n1558__, new_new_n1559__, new_new_n1560__, new_new_n1561__,
    new_new_n1562__, new_new_n1563__, new_new_n1564__, new_new_n1565__,
    new_new_n1566__, new_new_n1567__, new_new_n1568__, new_new_n1569__,
    new_new_n1570__, new_new_n1571__, new_new_n1572__, new_new_n1573__,
    new_new_n1574__, new_new_n1575__, new_new_n1576__, new_new_n1577__,
    new_new_n1578__, new_new_n1579__, new_new_n1580__, new_new_n1581__,
    new_new_n1582__, new_new_n1583__, new_new_n1584__, new_new_n1585__,
    new_new_n1586__, new_new_n1587__, new_new_n1588__, new_new_n1589__,
    new_new_n1590__, new_new_n1591__, new_new_n1592__, new_new_n1593__,
    new_new_n1594__, new_new_n1595__, new_new_n1596__, new_new_n1597__,
    new_new_n1598__, new_new_n1599__, new_new_n1600__, new_new_n1601__,
    new_new_n1602__, new_new_n1603__, new_new_n1604__, new_new_n1605__,
    new_new_n1606__, new_new_n1607__, new_new_n1608__, new_new_n1609__,
    new_new_n1610__, new_new_n1611__, new_new_n1612__, new_new_n1613__,
    new_new_n1614__, new_new_n1615__, new_new_n1616__, new_new_n1617__,
    new_new_n1618__, new_new_n1619__, new_new_n1620__, new_new_n1621__,
    new_new_n1622__, new_new_n1623__, new_new_n1624__, new_new_n1625__,
    new_new_n1626__, new_new_n1627__, new_new_n1628__, new_new_n1629__,
    new_new_n1630__, new_new_n1631__, new_new_n1632__, new_new_n1633__,
    new_new_n1634__, new_new_n1635__, new_new_n1636__, new_new_n1637__,
    new_new_n1638__, new_new_n1639__, new_new_n1640__, new_new_n1641__,
    new_new_n1642__, new_new_n1643__, new_new_n1644__, new_new_n1645__,
    new_new_n1646__, new_new_n1647__, new_new_n1648__, new_new_n1649__,
    new_new_n1650__, new_new_n1651__, new_new_n1652__, new_new_n1653__,
    new_new_n1654__, new_new_n1655__, new_new_n1656__, new_new_n1657__,
    new_new_n1658__, new_new_n1659__, new_new_n1660__, new_new_n1661__,
    new_new_n1662__, new_new_n1663__, new_new_n1664__, new_new_n1665__,
    new_new_n1666__, new_new_n1667__, new_new_n1668__, new_new_n1669__,
    new_new_n1670__, new_new_n1671__, new_new_n1672__, new_new_n1673__,
    new_new_n1674__, new_new_n1675__, new_new_n1676__, new_new_n1677__,
    new_new_n1678__, new_new_n1679__, new_new_n1680__, new_new_n1681__,
    new_new_n1682__, new_new_n1683__, new_new_n1684__, new_new_n1685__,
    new_new_n1686__, new_new_n1687__, new_new_n1688__, new_new_n1689__,
    new_new_n1690__, new_new_n1691__, new_new_n1692__, new_new_n1693__,
    new_new_n1694__, new_new_n1695__, new_new_n1696__, new_new_n1697__,
    new_new_n1698__, new_new_n1699__, new_new_n1700__, new_new_n1701__,
    new_new_n1702__, new_new_n1703__, new_new_n1704__, new_new_n1705__,
    new_new_n1706__, new_new_n1707__, new_new_n1708__, new_new_n1709__,
    new_new_n1710__, new_new_n1711__, new_new_n1712__, new_new_n1713__,
    new_new_n1714__, new_new_n1715__, new_new_n1716__, new_new_n1717__,
    new_new_n1718__, new_new_n1719__, new_new_n1720__, new_new_n1721__,
    new_new_n1722__, new_new_n1723__, new_new_n1724__, new_new_n1725__,
    new_new_n1726__, new_new_n1727__, new_new_n1728__, new_new_n1729__,
    new_new_n1730__, new_new_n1731__, new_new_n1732__, new_new_n1733__,
    new_new_n1734__, new_new_n1735__, new_new_n1736__, new_new_n1737__,
    new_new_n1738__, new_new_n1739__, new_new_n1740__, new_new_n1741__,
    new_new_n1742__, new_new_n1743__, new_new_n1744__, new_new_n1745__,
    new_new_n1746__, new_new_n1747__, new_new_n1748__, new_new_n1749__,
    new_new_n1750__, new_new_n1751__, new_new_n1752__, new_new_n1753__,
    new_new_n1754__, new_new_n1755__, new_new_n1756__, new_new_n1757__,
    new_new_n1758__, new_new_n1759__, new_new_n1760__, new_new_n1761__,
    new_new_n1762__, new_new_n1763__, new_new_n1764__, new_new_n1765__,
    new_new_n1766__, new_new_n1767__, new_new_n1768__, new_new_n1769__,
    new_new_n1770__, new_new_n1771__, new_new_n1772__, new_new_n1773__,
    new_new_n1774__, new_new_n1775__, new_new_n1776__, new_new_n1777__,
    new_new_n1778__, new_new_n1779__, new_new_n1780__, new_new_n1781__,
    new_new_n1782__, new_new_n1783__, new_new_n1784__, new_new_n1785__,
    new_new_n1786__, new_new_n1787__, new_new_n1788__, new_new_n1789__,
    new_new_n1790__, new_new_n1791__, new_new_n1792__, new_new_n1793__,
    new_new_n1794__, new_new_n1795__, new_new_n1796__, new_new_n1797__,
    new_new_n1798__, new_new_n1799__, new_new_n1800__, new_new_n1801__,
    new_new_n1802__, new_new_n1803__, new_new_n1804__, new_new_n1805__,
    new_new_n1806__, new_new_n1807__, new_new_n1808__, new_new_n1809__,
    new_new_n1810__, new_new_n1811__, new_new_n1812__, new_new_n1813__,
    new_new_n1814__, new_new_n1815__, new_new_n1816__, new_new_n1817__,
    new_new_n1818__, new_new_n1819__, new_new_n1820__, new_new_n1821__,
    new_new_n1822__, new_new_n1823__, new_new_n1824__, new_new_n1825__,
    new_new_n1826__, new_new_n1827__, new_new_n1828__, new_new_n1829__,
    new_new_n1830__, new_new_n1831__, new_new_n1832__, new_new_n1833__,
    new_new_n1834__, new_new_n1835__, new_new_n1836__, new_new_n1837__,
    new_new_n1838__, new_new_n1839__, new_new_n1840__, new_new_n1841__,
    new_new_n1842__, new_new_n1843__, new_new_n1844__, new_new_n1845__,
    new_new_n1846__, new_new_n1847__, new_new_n1848__, new_new_n1849__,
    new_new_n1850__, new_new_n1851__, new_new_n1852__, new_new_n1853__,
    new_new_n1854__, new_new_n1855__, new_new_n1856__, new_new_n1857__,
    new_new_n1858__, new_new_n1859__, new_new_n1860__, new_new_n1861__,
    new_new_n1862__, new_new_n1863__, new_new_n1864__, new_new_n1865__,
    new_new_n1866__, new_new_n1867__, new_new_n1868__, new_new_n1869__,
    new_new_n1870__, new_new_n1871__, new_new_n1872__, new_new_n1873__,
    new_new_n1874__, new_new_n1875__, new_new_n1876__, new_new_n1877__,
    new_new_n1878__, new_new_n1879__, new_new_n1880__, new_new_n1881__,
    new_new_n1882__, new_new_n1883__, new_new_n1884__, new_new_n1885__,
    new_new_n1886__, new_new_n1887__, new_new_n1888__, new_new_n1889__,
    new_new_n1890__, new_new_n1891__, new_new_n1892__, new_new_n1893__,
    new_new_n1894__, new_new_n1895__, new_new_n1896__, new_new_n1897__,
    new_new_n1898__, new_new_n1899__, new_new_n1900__, new_new_n1901__,
    new_new_n1902__, new_new_n1903__, new_new_n1904__, new_new_n1905__,
    new_new_n1906__, new_new_n1907__, new_new_n1908__, new_new_n1909__,
    new_new_n1910__, new_new_n1911__, new_new_n1912__, new_new_n1913__,
    new_new_n1914__, new_new_n1915__, new_new_n1916__, new_new_n1917__,
    new_new_n1918__, new_new_n1919__, new_new_n1920__, new_new_n1921__,
    new_new_n1922__, new_new_n1923__, new_new_n1924__, new_new_n1925__,
    new_new_n1926__, new_new_n1927__, new_new_n1928__, new_new_n1929__,
    new_new_n1930__, new_new_n1931__, new_new_n1932__, new_new_n1933__,
    new_new_n1934__, new_new_n1935__, new_new_n1936__, new_new_n1937__,
    new_new_n1938__, new_new_n1939__, new_new_n1940__, new_new_n1941__,
    new_new_n1942__, new_new_n1943__, new_new_n1944__, new_new_n1945__,
    new_new_n1946__, new_new_n1947__, new_new_n1948__, new_new_n1949__,
    new_new_n1950__, new_new_n1951__, new_new_n1952__, new_new_n1953__,
    new_new_n1954__, new_new_n1955__, new_new_n1956__, new_new_n1957__,
    new_new_n1958__, new_new_n1959__, new_new_n1960__, new_new_n1961__,
    new_new_n1962__, new_new_n1963__, new_new_n1964__, new_new_n1965__,
    new_new_n1966__, new_new_n1967__, new_new_n1968__, new_new_n1969__,
    new_new_n1970__, new_new_n1971__, new_new_n1972__, new_new_n1973__,
    new_new_n1974__, new_new_n1975__, new_new_n1976__, new_new_n1977__,
    new_new_n1978__, new_new_n1979__, new_new_n1980__, new_new_n1981__,
    new_new_n1982__, new_new_n1983__, new_new_n1984__, new_new_n1985__,
    new_new_n1986__, new_new_n1987__, new_new_n1988__, new_new_n1989__,
    new_new_n1990__, new_new_n1991__, new_new_n1992__, new_new_n1993__,
    new_new_n1994__, new_new_n1995__, new_new_n1996__, new_new_n1997__,
    new_new_n1998__, new_new_n1999__, new_new_n2000__, new_new_n2001__,
    new_new_n2002__, new_new_n2003__, new_new_n2004__, new_new_n2005__,
    new_new_n2006__, new_new_n2007__, new_new_n2008__, new_new_n2009__,
    new_new_n2010__, new_new_n2011__, new_new_n2012__, new_new_n2013__,
    new_new_n2014__, new_new_n2015__, new_new_n2016__, new_new_n2017__,
    new_new_n2018__, new_new_n2019__, new_new_n2020__, new_new_n2021__,
    new_new_n2022__, new_new_n2023__, new_new_n2024__, new_new_n2025__,
    new_new_n2026__, new_new_n2027__, new_new_n2028__, new_new_n2029__,
    new_new_n2030__, new_new_n2031__, new_new_n2032__, new_new_n2033__,
    new_new_n2034__, new_new_n2035__, new_new_n2036__, new_new_n2037__,
    new_new_n2038__, new_new_n2039__, new_new_n2040__, new_new_n2041__,
    new_new_n2042__, new_new_n2043__, new_new_n2044__, new_new_n2045__,
    new_new_n2046__, new_new_n2047__, new_new_n2048__, new_new_n2049__,
    new_new_n2050__, new_new_n2051__, new_new_n2052__, new_new_n2053__,
    new_new_n2054__, new_new_n2055__, new_new_n2056__, new_new_n2057__,
    new_new_n2058__, new_new_n2059__, new_new_n2060__, new_new_n2061__,
    new_new_n2062__, new_new_n2063__, new_new_n2064__, new_new_n2065__,
    new_new_n2066__, new_new_n2067__, new_new_n2068__, new_new_n2069__,
    new_new_n2070__, new_new_n2071__, new_new_n2072__, new_new_n2073__,
    new_new_n2074__, new_new_n2075__, new_new_n2076__, new_new_n2077__,
    new_new_n2078__, new_new_n2079__, new_new_n2080__, new_new_n2081__,
    new_new_n2082__, new_new_n2083__, new_new_n2084__, new_new_n2085__,
    new_new_n2086__, new_new_n2087__, new_new_n2088__, new_new_n2089__,
    new_new_n2090__, new_new_n2091__, new_new_n2092__, new_new_n2093__,
    new_new_n2094__, new_new_n2095__, new_new_n2096__, new_new_n2097__,
    new_new_n2098__, new_new_n2099__, new_new_n2100__, new_new_n2101__,
    new_new_n2102__, new_new_n2103__, new_new_n2104__, new_new_n2105__,
    new_new_n2106__, new_new_n2107__, new_new_n2108__, new_new_n2109__,
    new_new_n2110__, new_new_n2111__, new_new_n2112__, new_new_n2113__,
    new_new_n2114__, new_new_n2115__, new_new_n2116__, new_new_n2117__,
    new_new_n2118__, new_new_n2119__, new_new_n2120__, new_new_n2121__,
    new_new_n2122__, new_new_n2123__, new_new_n2124__, new_new_n2125__,
    new_new_n2126__, new_new_n2127__, new_new_n2128__, new_new_n2129__,
    new_new_n2130__, new_new_n2131__, new_new_n2132__, new_new_n2133__,
    new_new_n2134__, new_new_n2135__, new_new_n2136__, new_new_n2137__,
    new_new_n2138__, new_new_n2139__, new_new_n2140__, new_new_n2141__,
    new_new_n2142__, new_new_n2143__, new_new_n2144__, new_new_n2145__,
    new_new_n2146__, new_new_n2147__, new_new_n2148__, new_new_n2149__,
    new_new_n2150__, new_new_n2151__, new_new_n2152__, new_new_n2153__,
    new_new_n2154__, new_new_n2155__, new_new_n2156__, new_new_n2157__,
    new_new_n2158__, new_new_n2159__, new_new_n2160__, new_new_n2161__,
    new_new_n2162__, new_new_n2163__, new_new_n2164__, new_new_n2165__,
    new_new_n2166__, new_new_n2167__, new_new_n2168__, new_new_n2169__,
    new_new_n2170__, new_new_n2171__, new_new_n2172__, new_new_n2173__,
    new_new_n2174__, new_new_n2175__, new_new_n2176__, new_new_n2177__,
    new_new_n2178__, new_new_n2179__, new_new_n2180__, new_new_n2181__,
    new_new_n2182__, new_new_n2183__, new_new_n2184__, new_new_n2185__,
    new_new_n2186__, new_new_n2187__, new_new_n2188__, new_new_n2189__,
    new_new_n2190__, new_new_n2191__, new_new_n2192__, new_new_n2193__,
    new_new_n2194__, new_new_n2195__, new_new_n2196__, new_new_n2197__,
    new_new_n2198__, new_new_n2199__, new_new_n2200__, new_new_n2201__,
    new_new_n2202__, new_new_n2203__, new_new_n2204__, new_new_n2205__,
    new_new_n2206__, new_new_n2207__, new_new_n2208__, new_new_n2209__,
    new_new_n2210__, new_new_n2211__, new_new_n2212__, new_new_n2213__,
    new_new_n2214__, new_new_n2215__, new_new_n2216__, new_new_n2217__,
    new_new_n2218__, new_new_n2219__, new_new_n2220__, new_new_n2221__,
    new_new_n2222__, new_new_n2223__, new_new_n2224__, new_new_n2225__,
    new_new_n2226__, new_new_n2227__, new_new_n2228__, new_new_n2229__,
    new_new_n2230__, new_new_n2231__, new_new_n2232__, new_new_n2233__,
    new_new_n2234__, new_new_n2235__, new_new_n2236__, new_new_n2237__,
    new_new_n2238__, new_new_n2239__, new_new_n2240__, new_new_n2241__,
    new_new_n2242__, new_new_n2243__, new_new_n2244__, new_new_n2245__,
    new_new_n2246__, new_new_n2247__, new_new_n2248__, new_new_n2249__,
    new_new_n2250__, new_new_n2251__, new_new_n2252__, new_new_n2253__,
    new_new_n2254__, new_new_n2255__, new_new_n2256__, new_new_n2257__,
    new_new_n2258__, new_new_n2259__, new_new_n2260__, new_new_n2261__,
    new_new_n2262__, new_new_n2263__, new_new_n2264__, new_new_n2265__,
    new_new_n2266__, new_new_n2267__, new_new_n2268__, new_new_n2269__,
    new_new_n2270__, new_new_n2271__, new_new_n2272__, new_new_n2273__,
    new_new_n2274__, new_new_n2275__, new_new_n2276__, new_new_n2277__,
    new_new_n2278__, new_new_n2279__, new_new_n2280__, new_new_n2281__,
    new_new_n2282__, new_new_n2283__, new_new_n2284__, new_new_n2285__,
    new_new_n2286__, new_new_n2287__, new_new_n2288__, new_new_n2289__,
    new_new_n2290__, new_new_n2291__, new_new_n2292__, new_new_n2293__,
    new_new_n2294__, new_new_n2295__, new_new_n2296__, new_new_n2297__,
    new_new_n2298__, new_new_n2299__, new_new_n2300__, new_new_n2301__,
    new_new_n2302__, new_new_n2303__, new_new_n2304__, new_new_n2305__,
    new_new_n2306__, new_new_n2307__, new_new_n2308__, new_new_n2309__,
    new_new_n2310__, new_new_n2311__, new_new_n2312__, new_new_n2313__,
    new_new_n2314__, new_new_n2315__, new_new_n2316__, new_new_n2317__,
    new_new_n2318__, new_new_n2319__, new_new_n2320__, new_new_n2321__,
    new_new_n2322__, new_new_n2323__, new_new_n2324__, new_new_n2325__,
    new_new_n2326__, new_new_n2327__, new_new_n2328__, new_new_n2329__,
    new_new_n2330__, new_new_n2331__, new_new_n2332__, new_new_n2333__,
    new_new_n2334__, new_new_n2335__, new_new_n2336__, new_new_n2337__,
    new_new_n2338__, new_new_n2339__, new_new_n2340__, new_new_n2341__,
    new_new_n2342__, new_new_n2343__, new_new_n2344__, new_new_n2345__,
    new_new_n2346__, new_new_n2347__, new_new_n2348__, new_new_n2349__,
    new_new_n2350__, new_new_n2351__, new_new_n2352__, new_new_n2353__,
    new_new_n2354__, new_new_n2355__, new_new_n2356__, new_new_n2357__,
    new_new_n2358__, new_new_n2359__, new_new_n2360__, new_new_n2361__,
    new_new_n2362__, new_new_n2363__, new_new_n2364__, new_new_n2365__,
    new_new_n2366__, new_new_n2367__, new_new_n2368__, new_new_n2369__,
    new_new_n2370__, new_new_n2371__, new_new_n2372__, new_new_n2373__,
    new_new_n2374__, new_new_n2375__, new_new_n2376__, new_new_n2377__,
    new_new_n2378__, new_new_n2379__, new_new_n2380__, new_new_n2381__,
    new_new_n2382__, new_new_n2383__, new_new_n2384__, new_new_n2385__,
    new_new_n2386__, new_new_n2387__, new_new_n2388__, new_new_n2389__,
    new_new_n2390__, new_new_n2391__, new_new_n2392__, new_new_n2393__,
    new_new_n2394__, new_new_n2395__, new_new_n2396__, new_new_n2397__,
    new_new_n2398__, new_new_n2399__, new_new_n2400__, new_new_n2401__,
    new_new_n2402__, new_new_n2403__, new_new_n2404__, new_new_n2405__,
    new_new_n2406__, new_new_n2407__, new_new_n2408__, new_new_n2409__,
    new_new_n2410__, new_new_n2411__, new_new_n2412__, new_new_n2413__,
    new_new_n2414__, new_new_n2415__, new_new_n2416__, new_new_n2417__,
    new_new_n2418__, new_new_n2419__, new_new_n2420__, new_new_n2421__,
    new_new_n2422__, new_new_n2423__, new_new_n2424__, new_new_n2425__,
    new_new_n2426__, new_new_n2427__, new_new_n2428__, new_new_n2429__,
    new_new_n2430__, new_new_n2431__, new_new_n2432__, new_new_n2433__,
    new_new_n2434__, new_new_n2435__, new_new_n2436__, new_new_n2437__,
    new_new_n2438__, new_new_n2439__, new_new_n2440__, new_new_n2441__,
    new_new_n2442__, new_new_n2443__, new_new_n2444__, new_new_n2445__,
    new_new_n2446__, new_new_n2447__, new_new_n2448__, new_new_n2449__,
    new_new_n2450__, new_new_n2451__, new_new_n2452__, new_new_n2453__,
    new_new_n2454__, new_new_n2455__, new_new_n2456__, new_new_n2457__,
    new_new_n2458__, new_new_n2459__, new_new_n2460__, new_new_n2461__,
    new_new_n2462__, new_new_n2463__, new_new_n2464__, new_new_n2465__,
    new_new_n2466__, new_new_n2467__, new_new_n2468__, new_new_n2469__,
    new_new_n2470__, new_new_n2471__, new_new_n2472__, new_new_n2473__,
    new_new_n2474__, new_new_n2475__, new_new_n2476__, new_new_n2477__,
    new_new_n2478__, new_new_n2479__, new_new_n2480__, new_new_n2481__,
    new_new_n2482__, new_new_n2483__, new_new_n2484__, new_new_n2485__,
    new_new_n2486__, new_new_n2487__, new_new_n2488__, new_new_n2489__,
    new_new_n2490__, new_new_n2491__, new_new_n2492__, new_new_n2493__,
    new_new_n2494__, new_new_n2495__, new_new_n2496__, new_new_n2497__,
    new_new_n2498__, new_new_n2499__, new_new_n2500__, new_new_n2501__,
    new_new_n2502__, new_new_n2503__, new_new_n2504__, new_new_n2505__,
    new_new_n2506__, new_new_n2507__, new_new_n2508__, new_new_n2509__,
    new_new_n2510__, new_new_n2511__, new_new_n2512__, new_new_n2513__,
    new_new_n2514__, new_new_n2515__, new_new_n2516__, new_new_n2517__,
    new_new_n2518__, new_new_n2519__, new_new_n2520__, new_new_n2521__,
    new_new_n2522__, new_new_n2523__, new_new_n2524__, new_new_n2525__,
    new_new_n2526__, new_new_n2527__, new_new_n2528__, new_new_n2529__,
    new_new_n2530__, new_new_n2531__, new_new_n2532__, new_new_n2533__,
    new_new_n2534__, new_new_n2535__, new_new_n2536__, new_new_n2537__,
    new_new_n2538__, new_new_n2539__, new_new_n2540__, new_new_n2541__,
    new_new_n2542__, new_new_n2543__, new_new_n2544__, new_new_n2545__,
    new_new_n2546__, new_new_n2547__, new_new_n2548__, new_new_n2549__,
    new_new_n2550__, new_new_n2551__, new_new_n2552__, new_new_n2553__,
    new_new_n2554__, new_new_n2555__, new_new_n2556__, new_new_n2557__,
    new_new_n2558__, new_new_n2559__, new_new_n2560__, new_new_n2561__,
    new_new_n2562__, new_new_n2563__, new_new_n2564__, new_new_n2565__,
    new_new_n2566__, new_new_n2567__, new_new_n2568__, new_new_n2569__,
    new_new_n2570__, new_new_n2571__, new_new_n2572__, new_new_n2573__,
    new_new_n2574__, new_new_n2575__, new_new_n2576__, new_new_n2577__,
    new_new_n2578__, new_new_n2579__, new_new_n2580__, new_new_n2581__,
    new_new_n2582__, new_new_n2583__, new_new_n2584__, new_new_n2585__,
    new_new_n2586__, new_new_n2587__, new_new_n2588__, new_new_n2589__,
    new_new_n2590__, new_new_n2591__, new_new_n2592__, new_new_n2593__,
    new_new_n2594__, new_new_n2595__, new_new_n2596__, new_new_n2597__,
    new_new_n2598__, new_new_n2599__, new_new_n2600__, new_new_n2601__,
    new_new_n2602__, new_new_n2603__, new_new_n2604__, new_new_n2605__,
    new_new_n2606__, new_new_n2607__, new_new_n2608__, new_new_n2609__,
    new_new_n2610__, new_new_n2611__, new_new_n2612__, new_new_n2613__,
    new_new_n2614__, new_new_n2615__, new_new_n2616__, new_new_n2617__,
    new_new_n2618__, new_new_n2619__, new_new_n2620__, new_new_n2621__,
    new_new_n2622__, new_new_n2623__, new_new_n2624__, new_new_n2625__,
    new_new_n2626__, new_new_n2627__, new_new_n2628__, new_new_n2629__,
    new_new_n2630__, new_new_n2631__, new_new_n2632__, new_new_n2633__,
    new_new_n2634__, new_new_n2635__, new_new_n2636__, new_new_n2637__,
    new_new_n2638__, new_new_n2639__, new_new_n2640__, new_new_n2641__,
    new_new_n2642__, new_new_n2643__, new_new_n2644__, new_new_n2645__,
    new_new_n2646__, new_new_n2647__, new_new_n2648__, new_new_n2649__,
    new_new_n2650__, new_new_n2651__, new_new_n2652__, new_new_n2653__,
    new_new_n2654__, new_new_n2655__, new_new_n2656__, new_new_n2657__,
    new_new_n2658__, new_new_n2659__, new_new_n2660__, new_new_n2661__,
    new_new_n2662__, new_new_n2663__, new_new_n2664__, new_new_n2665__,
    new_new_n2666__, new_new_n2667__, new_new_n2668__, new_new_n2669__,
    new_new_n2670__, new_new_n2671__, new_new_n2672__, new_new_n2673__,
    new_new_n2674__, new_new_n2675__, new_new_n2676__, new_new_n2677__,
    new_new_n2678__, new_new_n2679__, new_new_n2680__, new_new_n2681__,
    new_new_n2682__, new_new_n2683__, new_new_n2684__, new_new_n2685__,
    new_new_n2686__, new_new_n2687__, new_new_n2688__, new_new_n2689__,
    new_new_n2690__, new_new_n2691__, new_new_n2692__, new_new_n2693__,
    new_new_n2694__, new_new_n2695__, new_new_n2696__, new_new_n2697__,
    new_new_n2698__, new_new_n2699__, new_new_n2700__, new_new_n2701__,
    new_new_n2702__, new_new_n2703__, new_new_n2704__, new_new_n2705__,
    new_new_n2706__, new_new_n2707__, new_new_n2708__, new_new_n2709__,
    new_new_n2710__, new_new_n2711__, new_new_n2712__, new_new_n2713__,
    new_new_n2714__, new_new_n2715__, new_new_n2716__, new_new_n2717__,
    new_new_n2718__, new_new_n2719__, new_new_n2720__, new_new_n2721__,
    new_new_n2722__, new_new_n2723__, new_new_n2724__, new_new_n2725__,
    new_new_n2726__, new_new_n2727__, new_new_n2728__, new_new_n2729__,
    new_new_n2730__, new_new_n2731__, new_new_n2732__, new_new_n2733__,
    new_new_n2734__, new_new_n2735__, new_new_n2736__, new_new_n2737__,
    new_new_n2738__, new_new_n2739__, new_new_n2740__, new_new_n2741__,
    new_new_n2742__, new_new_n2743__, new_new_n2744__, new_new_n2745__,
    new_new_n2746__, new_new_n2747__, new_new_n2748__, new_new_n2749__,
    new_new_n2750__, new_new_n2751__, new_new_n2752__, new_new_n2753__,
    new_new_n2754__, new_new_n2755__, new_new_n2756__, new_new_n2757__,
    new_new_n2758__, new_new_n2759__, new_new_n2760__, new_new_n2761__,
    new_new_n2762__, new_new_n2763__, new_new_n2764__, new_new_n2765__,
    new_new_n2766__, new_new_n2767__, new_new_n2768__, new_new_n2769__,
    new_new_n2770__, new_new_n2771__, new_new_n2772__, new_new_n2773__,
    new_new_n2774__, new_new_n2775__, new_new_n2776__, new_new_n2777__,
    new_new_n2778__, new_new_n2779__, new_new_n2780__, new_new_n2781__,
    new_new_n2782__, new_new_n2783__, new_new_n2784__, new_new_n2785__,
    new_new_n2786__, new_new_n2787__, new_new_n2788__, new_new_n2789__,
    new_new_n2790__, new_new_n2791__, new_new_n2792__, new_new_n2793__,
    new_new_n2794__, new_new_n2795__, new_new_n2796__, new_new_n2797__,
    new_new_n2798__, new_new_n2799__, new_new_n2800__, new_new_n2801__,
    new_new_n2802__, new_new_n2803__, new_new_n2804__, new_new_n2805__,
    new_new_n2806__, new_new_n2807__, new_new_n2808__, new_new_n2809__,
    new_new_n2810__, new_new_n2811__, new_new_n2812__, new_new_n2813__,
    new_new_n2814__, new_new_n2815__, new_new_n2816__, new_new_n2817__,
    new_new_n2818__, new_new_n2819__, new_new_n2820__, new_new_n2821__,
    new_new_n2822__, new_new_n2823__, new_new_n2824__, new_new_n2825__,
    new_new_n2826__, new_new_n2827__, new_new_n2828__, new_new_n2829__,
    new_new_n2830__, new_new_n2831__, new_new_n2832__, new_new_n2833__,
    new_new_n2834__, new_new_n2835__, new_new_n2836__, new_new_n2837__,
    new_new_n2838__, new_new_n2839__, new_new_n2840__, new_new_n2841__,
    new_new_n2842__, new_new_n2843__, new_new_n2844__, new_new_n2845__,
    new_new_n2846__, new_new_n2847__, new_new_n2848__, new_new_n2849__,
    new_new_n2850__, new_new_n2851__, new_new_n2852__, new_new_n2853__,
    new_new_n2854__, new_new_n2855__, new_new_n2856__, new_new_n2857__,
    new_new_n2858__, new_new_n2859__, new_new_n2860__, new_new_n2861__,
    new_new_n2862__, new_new_n2863__, new_new_n2864__, new_new_n2865__,
    new_new_n2866__, new_new_n2867__, new_new_n2868__, new_new_n2869__,
    new_new_n2870__, new_new_n2871__, new_new_n2872__, new_new_n2873__,
    new_new_n2874__, new_new_n2875__, new_new_n2876__, new_new_n2877__,
    new_new_n2878__, new_new_n2879__, new_new_n2880__, new_new_n2881__,
    new_new_n2882__, new_new_n2883__, new_new_n2884__, new_new_n2885__,
    new_new_n2886__, new_new_n2887__, new_new_n2888__, new_new_n2889__,
    new_new_n2890__, new_new_n2891__, new_new_n2892__, new_new_n2893__,
    new_new_n2894__, new_new_n2895__, new_new_n2896__, new_new_n2897__,
    new_new_n2898__, new_new_n2899__, new_new_n2900__, new_new_n2901__,
    new_new_n2902__, new_new_n2903__, new_new_n2904__, new_new_n2905__,
    new_new_n2906__, new_new_n2907__, new_new_n2908__, new_new_n2909__,
    new_new_n2910__, new_new_n2911__, new_new_n2912__, new_new_n2913__,
    new_new_n2914__, new_new_n2915__, new_new_n2916__, new_new_n2917__,
    new_new_n2918__, new_new_n2919__, new_new_n2920__, new_new_n2921__,
    new_new_n2922__, new_new_n2923__, new_new_n2924__, new_new_n2925__,
    new_new_n2926__, new_new_n2927__, new_new_n2928__, new_new_n2929__,
    new_new_n2930__, new_new_n2931__, new_new_n2932__, new_new_n2933__,
    new_new_n2934__, new_new_n2935__, new_new_n2936__, new_new_n2937__,
    new_new_n2938__, new_new_n2939__, new_new_n2940__, new_new_n2941__,
    new_new_n2942__, new_new_n2943__, new_new_n2944__, new_new_n2945__,
    new_new_n2946__, new_new_n2947__, new_new_n2948__, new_new_n2949__,
    new_new_n2950__, new_new_n2951__, new_new_n2952__, new_new_n2953__,
    new_new_n2954__, new_new_n2955__, new_new_n2956__, new_new_n2957__,
    new_new_n2958__, new_new_n2959__, new_new_n2960__, new_new_n2961__,
    new_new_n2962__, new_new_n2963__, new_new_n2964__, new_new_n2965__,
    new_new_n2966__, new_new_n2967__, new_new_n2968__, new_new_n2969__,
    new_new_n2970__, new_new_n2971__, new_new_n2972__, new_new_n2973__,
    new_new_n2974__, new_new_n2975__, new_new_n2976__, new_new_n2977__,
    new_new_n2978__, new_new_n2979__, new_new_n2980__, new_new_n2981__,
    new_new_n2982__, new_new_n2983__, new_new_n2984__, new_new_n2985__,
    new_new_n2986__, new_new_n2987__, new_new_n2988__, new_new_n2989__,
    new_new_n2990__, new_new_n2991__, new_new_n2992__, new_new_n2993__,
    new_new_n2994__, new_new_n2995__, new_new_n2996__, new_new_n2997__,
    new_new_n2998__, new_new_n2999__, new_new_n3000__, new_new_n3001__,
    new_new_n3002__, new_new_n3003__, new_new_n3004__, new_new_n3005__,
    new_new_n3006__, new_new_n3007__, new_new_n3008__, new_new_n3009__,
    new_new_n3010__, new_new_n3011__, new_new_n3012__, new_new_n3013__,
    new_new_n3014__, new_new_n3015__, new_new_n3016__, new_new_n3017__,
    new_new_n3018__, new_new_n3019__, new_new_n3020__, new_new_n3021__,
    new_new_n3022__, new_new_n3023__, new_new_n3024__, new_new_n3025__,
    new_new_n3026__, new_new_n3027__, new_new_n3028__, new_new_n3029__,
    new_new_n3030__, new_new_n3031__, new_new_n3032__, new_new_n3033__,
    new_new_n3034__, new_new_n3035__, new_new_n3036__, new_new_n3037__,
    new_new_n3038__, new_new_n3039__, new_new_n3040__, new_new_n3041__,
    new_new_n3042__, new_new_n3043__, new_new_n3044__, new_new_n3045__,
    new_new_n3046__, new_new_n3047__, new_new_n3048__, new_new_n3049__,
    new_new_n3050__, new_new_n3051__, new_new_n3052__, new_new_n3053__,
    new_new_n3054__, new_new_n3055__, new_new_n3056__, new_new_n3057__,
    new_new_n3058__, new_new_n3059__, new_new_n3060__, new_new_n3061__,
    new_new_n3062__, new_new_n3063__, new_new_n3064__, new_new_n3065__,
    new_new_n3066__, new_new_n3067__, new_new_n3068__, new_new_n3069__,
    new_new_n3070__, new_new_n3071__, new_new_n3072__, new_new_n3073__,
    new_new_n3074__, new_new_n3075__, new_new_n3076__, new_new_n3077__,
    new_new_n3078__, new_new_n3079__, new_new_n3080__, new_new_n3081__,
    new_new_n3082__, new_new_n3083__, new_new_n3084__, new_new_n3085__,
    new_new_n3086__, new_new_n3087__, new_new_n3088__, new_new_n3089__,
    new_new_n3090__, new_new_n3091__, new_new_n3092__, new_new_n3093__,
    new_new_n3094__, new_new_n3095__, new_new_n3096__, new_new_n3097__,
    new_new_n3098__, new_new_n3099__, new_new_n3100__, new_new_n3101__,
    new_new_n3102__, new_new_n3103__, new_new_n3104__, new_new_n3105__,
    new_new_n3106__, new_new_n3107__, new_new_n3108__, new_new_n3109__,
    new_new_n3110__, new_new_n3111__, new_new_n3112__, new_new_n3113__,
    new_new_n3114__, new_new_n3115__, new_new_n3116__, new_new_n3117__,
    new_new_n3118__, new_new_n3119__, new_new_n3120__, new_new_n3121__,
    new_new_n3122__, new_new_n3123__, new_new_n3124__, new_new_n3125__,
    new_new_n3126__, new_new_n3127__, new_new_n3128__, new_new_n3129__,
    new_new_n3130__, new_new_n3131__, new_new_n3132__, new_new_n3133__,
    new_new_n3134__, new_new_n3135__, new_new_n3136__, new_new_n3137__,
    new_new_n3138__, new_new_n3139__, new_new_n3140__, new_new_n3141__,
    new_new_n3142__, new_new_n3143__, new_new_n3144__, new_new_n3145__,
    new_new_n3146__, new_new_n3147__, new_new_n3148__, new_new_n3149__,
    new_new_n3150__, new_new_n3151__, new_new_n3152__, new_new_n3153__,
    new_new_n3154__, new_new_n3155__, new_new_n3156__, new_new_n3157__,
    new_new_n3158__, new_new_n3159__, new_new_n3160__, new_new_n3161__,
    new_new_n3162__, new_new_n3163__, new_new_n3164__, new_new_n3165__,
    new_new_n3166__, new_new_n3167__, new_new_n3168__, new_new_n3169__,
    new_new_n3170__, new_new_n3171__, new_new_n3172__, new_new_n3173__,
    new_new_n3174__, new_new_n3175__, new_new_n3176__, new_new_n3177__,
    new_new_n3178__, new_new_n3179__, new_new_n3180__, new_new_n3181__,
    new_new_n3182__, new_new_n3183__, new_new_n3184__, new_new_n3185__,
    new_new_n3186__, new_new_n3187__, new_new_n3188__, new_new_n3189__,
    new_new_n3190__, new_new_n3191__, new_new_n3192__, new_new_n3193__,
    new_new_n3194__, new_new_n3195__, new_new_n3196__, new_new_n3197__,
    new_new_n3198__, new_new_n3199__, new_new_n3200__, new_new_n3201__,
    new_new_n3202__, new_new_n3203__, new_new_n3204__, new_new_n3205__,
    new_new_n3206__, new_new_n3207__, new_new_n3208__, new_new_n3209__,
    new_new_n3210__, new_new_n3211__, new_new_n3212__, new_new_n3213__,
    new_new_n3214__, new_new_n3215__, new_new_n3216__, new_new_n3217__,
    new_new_n3218__, new_new_n3219__, new_new_n3220__, new_new_n3221__,
    new_new_n3222__, new_new_n3223__, new_new_n3224__, new_new_n3225__,
    new_new_n3226__, new_new_n3227__, new_new_n3228__, new_new_n3229__,
    new_new_n3230__, new_new_n3231__, new_new_n3232__, new_new_n3233__,
    new_new_n3234__, new_new_n3235__, new_new_n3236__, new_new_n3237__,
    new_new_n3238__, new_new_n3239__, new_new_n3240__, new_new_n3241__,
    new_new_n3242__, new_new_n3243__, new_new_n3244__, new_new_n3245__,
    new_new_n3246__, new_new_n3247__, new_new_n3248__, new_new_n3249__,
    new_new_n3250__, new_new_n3251__, new_new_n3252__, new_new_n3253__,
    new_new_n3254__, new_new_n3255__, new_new_n3256__, new_new_n3257__,
    new_new_n3258__, new_new_n3259__, new_new_n3260__, new_new_n3261__,
    new_new_n3262__, new_new_n3263__, new_new_n3264__, new_new_n3265__,
    new_new_n3266__, new_new_n3267__, new_new_n3268__, new_new_n3269__,
    new_new_n3270__, new_new_n3271__, new_new_n3272__, new_new_n3273__,
    new_new_n3274__, new_new_n3275__, new_new_n3276__, new_new_n3277__,
    new_new_n3278__, new_new_n3279__, new_new_n3280__, new_new_n3281__,
    new_new_n3282__, new_new_n3283__, new_new_n3284__, new_new_n3285__,
    new_new_n3286__, new_new_n3287__, new_new_n3288__, new_new_n3289__,
    new_new_n3290__, new_new_n3291__, new_new_n3292__, new_new_n3293__,
    new_new_n3294__, new_new_n3295__, new_new_n3296__, new_new_n3297__,
    new_new_n3298__, new_new_n3299__, new_new_n3300__, new_new_n3301__,
    new_new_n3302__, new_new_n3303__, new_new_n3304__, new_new_n3305__,
    new_new_n3306__, new_new_n3307__, new_new_n3308__, new_new_n3309__,
    new_new_n3310__, new_new_n3311__, new_new_n3312__, new_new_n3313__,
    new_new_n3314__, new_new_n3315__, new_new_n3316__, new_new_n3317__,
    new_new_n3318__, new_new_n3319__, new_new_n3320__, new_new_n3321__,
    new_new_n3322__, new_new_n3323__, new_new_n3324__, new_new_n3325__,
    new_new_n3326__, new_new_n3327__, new_new_n3328__, new_new_n3329__,
    new_new_n3330__, new_new_n3331__, new_new_n3332__, new_new_n3333__,
    new_new_n3334__, new_new_n3335__, new_new_n3336__, new_new_n3337__,
    new_new_n3338__, new_new_n3339__, new_new_n3340__, new_new_n3341__,
    new_new_n3342__, new_new_n3343__, new_new_n3344__, new_new_n3345__,
    new_new_n3346__, new_new_n3347__, new_new_n3348__, new_new_n3349__,
    new_new_n3350__, new_new_n3351__, new_new_n3352__, new_new_n3353__,
    new_new_n3354__, new_new_n3355__, new_new_n3356__, new_new_n3357__,
    new_new_n3358__, new_new_n3359__, new_new_n3360__, new_new_n3361__,
    new_new_n3362__, new_new_n3363__, new_new_n3364__, new_new_n3365__,
    new_new_n3366__, new_new_n3367__, new_new_n3368__, new_new_n3369__,
    new_new_n3370__, new_new_n3371__, new_new_n3372__, new_new_n3373__,
    new_new_n3374__, new_new_n3375__, new_new_n3376__, new_new_n3377__,
    new_new_n3378__, new_new_n3379__, new_new_n3380__, new_new_n3381__,
    new_new_n3382__, new_new_n3383__, new_new_n3384__, new_new_n3385__,
    new_new_n3386__, new_new_n3387__, new_new_n3388__, new_new_n3389__,
    new_new_n3390__, new_new_n3391__, new_new_n3392__, new_new_n3393__,
    new_new_n3394__, new_new_n3395__, new_new_n3396__, new_new_n3397__,
    new_new_n3398__, new_new_n3399__, new_new_n3400__, new_new_n3401__,
    new_new_n3402__, new_new_n3403__, new_new_n3404__, new_new_n3405__,
    new_new_n3406__, new_new_n3407__, new_new_n3408__, new_new_n3409__,
    new_new_n3410__, new_new_n3411__, new_new_n3412__, new_new_n3413__,
    new_new_n3414__, new_new_n3415__, new_new_n3416__, new_new_n3417__,
    new_new_n3418__, new_new_n3419__, new_new_n3420__, new_new_n3421__,
    new_new_n3422__, new_new_n3423__, new_new_n3424__, new_new_n3425__,
    new_new_n3426__, new_new_n3427__, new_new_n3428__, new_new_n3429__,
    new_new_n3430__, new_new_n3431__, new_new_n3432__, new_new_n3433__,
    new_new_n3434__, new_new_n3435__, new_new_n3436__, new_new_n3437__,
    new_new_n3438__, new_new_n3439__, new_new_n3440__, new_new_n3441__,
    new_new_n3442__, new_new_n3443__, new_new_n3444__, new_new_n3445__,
    new_new_n3446__, new_new_n3447__, new_new_n3448__, new_new_n3449__,
    new_new_n3450__, new_new_n3451__, new_new_n3452__, new_new_n3453__,
    new_new_n3454__, new_new_n3455__, new_new_n3456__, new_new_n3457__,
    new_new_n3458__, new_new_n3459__, new_new_n3460__, new_new_n3461__,
    new_new_n3462__, new_new_n3463__, new_new_n3464__, new_new_n3465__,
    new_new_n3466__, new_new_n3467__, new_new_n3468__, new_new_n3469__,
    new_new_n3470__, new_new_n3471__, new_new_n3472__, new_new_n3473__,
    new_new_n3474__, new_new_n3475__, new_new_n3476__, new_new_n3477__,
    new_new_n3478__, new_new_n3479__, new_new_n3480__, new_new_n3481__,
    new_new_n3482__, new_new_n3483__, new_new_n3484__, new_new_n3485__,
    new_new_n3486__, new_new_n3487__, new_new_n3488__, new_new_n3489__,
    new_new_n3490__, new_new_n3491__, new_new_n3492__, new_new_n3493__,
    new_new_n3494__, new_new_n3495__, new_new_n3496__, new_new_n3497__,
    new_new_n3498__, new_new_n3499__, new_new_n3500__, new_new_n3501__,
    new_new_n3502__, new_new_n3503__, new_new_n3504__, new_new_n3505__,
    new_new_n3506__, new_new_n3507__, new_new_n3508__, new_new_n3509__,
    new_new_n3510__, new_new_n3511__, new_new_n3512__, new_new_n3513__,
    new_new_n3514__, new_new_n3515__, new_new_n3516__, new_new_n3517__,
    new_new_n3518__, new_new_n3519__, new_new_n3520__, new_new_n3521__,
    new_new_n3522__, new_new_n3523__, new_new_n3524__, new_new_n3525__,
    new_new_n3526__, new_new_n3527__, new_new_n3528__, new_new_n3529__,
    new_new_n3530__, new_new_n3531__, new_new_n3532__, new_new_n3533__,
    new_new_n3534__, new_new_n3535__, new_new_n3536__, new_new_n3537__,
    new_new_n3538__, new_new_n3539__, new_new_n3540__, new_new_n3541__,
    new_new_n3542__, new_new_n3543__, new_new_n3544__, new_new_n3545__,
    new_new_n3546__, new_new_n3547__, new_new_n3548__, new_new_n3549__,
    new_new_n3550__, new_new_n3551__, new_new_n3552__, new_new_n3553__,
    new_new_n3554__, new_new_n3555__, new_new_n3556__, new_new_n3557__,
    new_new_n3558__, new_new_n3559__, new_new_n3560__, new_new_n3561__,
    new_new_n3562__, new_new_n3563__, new_new_n3564__, new_new_n3565__,
    new_new_n3566__, new_new_n3567__, new_new_n3568__, new_new_n3569__,
    new_new_n3570__, new_new_n3571__, new_new_n3572__, new_new_n3573__,
    new_new_n3574__, new_new_n3575__, new_new_n3576__, new_new_n3577__,
    new_new_n3578__, new_new_n3579__, new_new_n3580__, new_new_n3581__,
    new_new_n3582__, new_new_n3583__, new_new_n3584__, new_new_n3585__,
    new_new_n3586__, new_new_n3587__, new_new_n3588__, new_new_n3589__,
    new_new_n3590__, new_new_n3591__, new_new_n3592__, new_new_n3593__,
    new_new_n3594__, new_new_n3595__, new_new_n3596__, new_new_n3597__,
    new_new_n3598__, new_new_n3599__, new_new_n3600__, new_new_n3601__,
    new_new_n3602__, new_new_n3603__, new_new_n3604__, new_new_n3605__,
    new_new_n3606__, new_new_n3607__, new_new_n3608__, new_new_n3609__,
    new_new_n3610__, new_new_n3611__, new_new_n3612__, new_new_n3613__,
    new_new_n3614__, new_new_n3615__, new_new_n3616__, new_new_n3617__,
    new_new_n3618__, new_new_n3619__, new_new_n3620__, new_new_n3621__,
    new_new_n3622__, new_new_n3623__, new_new_n3624__, new_new_n3625__,
    new_new_n3626__, new_new_n3627__, new_new_n3628__, new_new_n3629__,
    new_new_n3630__, new_new_n3631__, new_new_n3632__, new_new_n3633__,
    new_new_n3634__, new_new_n3635__, new_new_n3636__, new_new_n3637__,
    new_new_n3638__, new_new_n3639__, new_new_n3640__, new_new_n3641__,
    new_new_n3642__, new_new_n3643__, new_new_n3644__, new_new_n3645__,
    new_new_n3646__, new_new_n3647__, new_new_n3648__, new_new_n3649__,
    new_new_n3650__, new_new_n3651__, new_new_n3652__, new_new_n3653__,
    new_new_n3654__, new_new_n3655__, new_new_n3656__, new_new_n3657__,
    new_new_n3658__, new_new_n3659__, new_new_n3660__, new_new_n3661__,
    new_new_n3662__, new_new_n3663__, new_new_n3664__, new_new_n3665__,
    new_new_n3666__, new_new_n3667__, new_new_n3668__, new_new_n3669__,
    new_new_n3670__, new_new_n3671__, new_new_n3672__, new_new_n3673__,
    new_new_n3674__, new_new_n3675__, new_new_n3676__, new_new_n3677__,
    new_new_n3678__, new_new_n3679__, new_new_n3680__, new_new_n3681__,
    new_new_n3682__, new_new_n3683__, new_new_n3684__, new_new_n3685__,
    new_new_n3686__, new_new_n3687__, new_new_n3688__, new_new_n3689__,
    new_new_n3690__, new_new_n3691__, new_new_n3692__, new_new_n3693__,
    new_new_n3694__, new_new_n3695__, new_new_n3696__, new_new_n3697__,
    new_new_n3698__, new_new_n3699__, new_new_n3700__, new_new_n3701__,
    new_new_n3702__, new_new_n3703__, new_new_n3704__, new_new_n3705__,
    new_new_n3706__, new_new_n3707__, new_new_n3708__, new_new_n3709__,
    new_new_n3710__, new_new_n3711__, new_new_n3712__, new_new_n3713__,
    new_new_n3714__, new_new_n3715__, new_new_n3716__, new_new_n3717__,
    new_new_n3718__, new_new_n3719__, new_new_n3720__, new_new_n3721__,
    new_new_n3722__, new_new_n3723__, new_new_n3724__, new_new_n3725__,
    new_new_n3726__, new_new_n3727__, new_new_n3728__, new_new_n3729__,
    new_new_n3730__, new_new_n3731__, new_new_n3732__, new_new_n3733__,
    new_new_n3734__, new_new_n3735__, new_new_n3736__, new_new_n3737__,
    new_new_n3738__, new_new_n3739__, new_new_n3740__, new_new_n3741__,
    new_new_n3742__, new_new_n3743__, new_new_n3744__, new_new_n3745__,
    new_new_n3746__, new_new_n3747__, new_new_n3748__, new_new_n3749__,
    new_new_n3750__, new_new_n3751__, new_new_n3752__, new_new_n3753__,
    new_new_n3754__, new_new_n3755__, new_new_n3756__, new_new_n3757__,
    new_new_n3758__, new_new_n3759__, new_new_n3760__, new_new_n3761__,
    new_new_n3762__, new_new_n3763__, new_new_n3764__, new_new_n3765__,
    new_new_n3766__, new_new_n3767__, new_new_n3768__, new_new_n3769__,
    new_new_n3770__, new_new_n3771__, new_new_n3772__, new_new_n3773__,
    new_new_n3774__, new_new_n3775__, new_new_n3776__, new_new_n3777__,
    new_new_n3778__, new_new_n3779__, new_new_n3780__, new_new_n3781__,
    new_new_n3782__, new_new_n3783__, new_new_n3784__, new_new_n3785__,
    new_new_n3786__, new_new_n3787__, new_new_n3788__, new_new_n3789__,
    new_new_n3790__, new_new_n3791__, new_new_n3792__, new_new_n3793__,
    new_new_n3794__, new_new_n3795__, new_new_n3796__, new_new_n3797__,
    new_new_n3798__, new_new_n3799__, new_new_n3800__, new_new_n3801__,
    new_new_n3802__, new_new_n3803__, new_new_n3804__, new_new_n3805__,
    new_new_n3806__, new_new_n3807__, new_new_n3808__, new_new_n3809__,
    new_new_n3810__, new_new_n3811__, new_new_n3812__, new_new_n3813__,
    new_new_n3814__, new_new_n3815__, new_new_n3816__, new_new_n3817__,
    new_new_n3818__, new_new_n3819__, new_new_n3820__, new_new_n3821__,
    new_new_n3822__, new_new_n3823__, new_new_n3824__, new_new_n3825__,
    new_new_n3826__, new_new_n3827__, new_new_n3828__, new_new_n3829__,
    new_new_n3830__, new_new_n3831__, new_new_n3832__, new_new_n3833__,
    new_new_n3834__, new_new_n3835__, new_new_n3836__, new_new_n3837__,
    new_new_n3838__, new_new_n3839__, new_new_n3840__, new_new_n3841__,
    new_new_n3842__, new_new_n3843__, new_new_n3844__, new_new_n3845__,
    new_new_n3846__, new_new_n3847__, new_new_n3848__, new_new_n3849__,
    new_new_n3850__, new_new_n3851__, new_new_n3852__, new_new_n3853__,
    new_new_n3854__, new_new_n3855__, new_new_n3856__, new_new_n3857__,
    new_new_n3858__, new_new_n3859__, new_new_n3860__, new_new_n3861__,
    new_new_n3862__, new_new_n3863__, new_new_n3864__, new_new_n3865__,
    new_new_n3866__, new_new_n3867__, new_new_n3868__, new_new_n3869__,
    new_new_n3870__, new_new_n3871__, new_new_n3872__, new_new_n3873__,
    new_new_n3874__, new_new_n3875__, new_new_n3876__, new_new_n3877__,
    new_new_n3878__, new_new_n3879__, new_new_n3880__, new_new_n3881__,
    new_new_n3882__, new_new_n3883__, new_new_n3884__, new_new_n3885__,
    new_new_n3886__, new_new_n3887__, new_new_n3888__, new_new_n3889__,
    new_new_n3890__, new_new_n3891__, new_new_n3892__, new_new_n3893__,
    new_new_n3894__, new_new_n3895__, new_new_n3896__, new_new_n3897__,
    new_new_n3898__, new_new_n3899__, new_new_n3900__, new_new_n3901__,
    new_new_n3902__, new_new_n3903__, new_new_n3904__, new_new_n3905__,
    new_new_n3906__, new_new_n3907__, new_new_n3908__, new_new_n3909__,
    new_new_n3910__, new_new_n3911__, new_new_n3912__, new_new_n3913__,
    new_new_n3914__, new_new_n3915__, new_new_n3916__, new_new_n3917__,
    new_new_n3918__, new_new_n3919__, new_new_n3920__, new_new_n3921__,
    new_new_n3922__, new_new_n3923__, new_new_n3924__, new_new_n3925__,
    new_new_n3926__, new_new_n3927__, new_new_n3928__, new_new_n3929__,
    new_new_n3930__, new_new_n3931__, new_new_n3932__, new_new_n3933__,
    new_new_n3934__, new_new_n3935__, new_new_n3936__, new_new_n3937__,
    new_new_n3938__, new_new_n3939__, new_new_n3940__, new_new_n3941__,
    new_new_n3942__, new_new_n3943__, new_new_n3944__, new_new_n3945__,
    new_new_n3946__, new_new_n3947__, new_new_n3948__, new_new_n3949__,
    new_new_n3950__, new_new_n3951__, new_new_n3952__, new_new_n3953__,
    new_new_n3954__, new_new_n3955__, new_new_n3956__, new_new_n3957__,
    new_new_n3958__, new_new_n3959__, new_new_n3960__, new_new_n3961__,
    new_new_n3962__, new_new_n3963__, new_new_n3964__, new_new_n3965__,
    new_new_n3966__, new_new_n3967__, new_new_n3968__, new_new_n3969__,
    new_new_n3970__, new_new_n3971__, new_new_n3972__, new_new_n3973__,
    new_new_n3974__, new_new_n3975__, new_new_n3976__, new_new_n3977__,
    new_new_n3978__, new_new_n3979__, new_new_n3980__, new_new_n3981__,
    new_new_n3982__, new_new_n3983__, new_new_n3984__, new_new_n3985__,
    new_new_n3986__, new_new_n3987__, new_new_n3988__, new_new_n3989__,
    new_new_n3990__, new_new_n3991__, new_new_n3992__, new_new_n3993__,
    new_new_n3994__, new_new_n3995__, new_new_n3996__, new_new_n3997__,
    new_new_n3998__, new_new_n3999__, new_new_n4000__, new_new_n4001__,
    new_new_n4002__, new_new_n4003__, new_new_n4004__, new_new_n4005__,
    new_new_n4006__, new_new_n4007__, new_new_n4008__, new_new_n4009__,
    new_new_n4010__, new_new_n4011__, new_new_n4012__, new_new_n4013__,
    new_new_n4014__, new_new_n4015__, new_new_n4016__, new_new_n4017__,
    new_new_n4018__, new_new_n4019__, new_new_n4020__, new_new_n4021__,
    new_new_n4022__, new_new_n4023__, new_new_n4024__, new_new_n4025__,
    new_new_n4026__, new_new_n4027__, new_new_n4028__, new_new_n4029__,
    new_new_n4030__, new_new_n4031__, new_new_n4032__, new_new_n4033__,
    new_new_n4034__, new_new_n4035__, new_new_n4036__, new_new_n4037__,
    new_new_n4038__, new_new_n4039__, new_new_n4040__, new_new_n4041__,
    new_new_n4042__, new_new_n4043__, new_new_n4044__, new_new_n4045__,
    new_new_n4046__, new_new_n4047__, new_new_n4048__, new_new_n4049__,
    new_new_n4050__, new_new_n4051__, new_new_n4052__, new_new_n4053__,
    new_new_n4054__, new_new_n4055__, new_new_n4056__, new_new_n4057__,
    new_new_n4058__, new_new_n4059__, new_new_n4060__, new_new_n4061__,
    new_new_n4062__, new_new_n4063__, new_new_n4064__, new_new_n4065__,
    new_new_n4066__, new_new_n4067__, new_new_n4068__, new_new_n4069__,
    new_new_n4070__, new_new_n4071__, new_new_n4072__, new_new_n4073__,
    new_new_n4074__, new_new_n4075__, new_new_n4076__, new_new_n4077__,
    new_new_n4078__, new_new_n4079__, new_new_n4080__, new_new_n4081__,
    new_new_n4082__, new_new_n4083__, new_new_n4084__, new_new_n4085__,
    new_new_n4086__, new_new_n4087__, new_new_n4088__, new_new_n4089__,
    new_new_n4090__, new_new_n4091__, new_new_n4092__, new_new_n4093__,
    new_new_n4094__, new_new_n4095__, new_new_n4096__, new_new_n4097__,
    new_new_n4098__, new_new_n4099__, new_new_n4100__, new_new_n4101__,
    new_new_n4102__, new_new_n4103__, new_new_n4104__, new_new_n4105__,
    new_new_n4106__, new_new_n4107__, new_new_n4108__, new_new_n4109__,
    new_new_n4110__, new_new_n4111__, new_new_n4112__, new_new_n4113__,
    new_new_n4114__, new_new_n4115__, new_new_n4116__, new_new_n4117__,
    new_new_n4118__, new_new_n4119__, new_new_n4120__, new_new_n4121__,
    new_new_n4122__, new_new_n4123__, new_new_n4124__, new_new_n4125__,
    new_new_n4126__, new_new_n4127__, new_new_n4128__, new_new_n4129__,
    new_new_n4130__, new_new_n4131__, new_new_n4132__, new_new_n4133__,
    new_new_n4134__, new_new_n4135__, new_new_n4136__, new_new_n4137__,
    new_new_n4138__, new_new_n4139__, new_new_n4140__, new_new_n4141__,
    new_new_n4142__, new_new_n4143__, new_new_n4144__, new_new_n4145__,
    new_new_n4146__, new_new_n4147__, new_new_n4148__, new_new_n4149__,
    new_new_n4150__, new_new_n4151__, new_new_n4152__, new_new_n4153__,
    new_new_n4154__, new_new_n4155__, new_new_n4156__, new_new_n4157__,
    new_new_n4158__, new_new_n4159__, new_new_n4160__, new_new_n4161__,
    new_new_n4162__, new_new_n4163__, new_new_n4164__, new_new_n4165__,
    new_new_n4166__, new_new_n4167__, new_new_n4168__, new_new_n4169__,
    new_new_n4170__, new_new_n4171__, new_new_n4172__, new_new_n4173__,
    new_new_n4174__, new_new_n4175__, new_new_n4176__, new_new_n4177__,
    new_new_n4178__, new_new_n4179__, new_new_n4180__, new_new_n4181__,
    new_new_n4182__, new_new_n4183__, new_new_n4184__, new_new_n4185__,
    new_new_n4186__, new_new_n4187__, new_new_n4188__, new_new_n4189__,
    new_new_n4190__, new_new_n4191__, new_new_n4192__, new_new_n4193__,
    new_new_n4194__, new_new_n4195__, new_new_n4196__, new_new_n4197__,
    new_new_n4198__, new_new_n4199__, new_new_n4200__, new_new_n4201__,
    new_new_n4202__, new_new_n4203__, new_new_n4204__, new_new_n4205__,
    new_new_n4206__, new_new_n4207__, new_new_n4208__, new_new_n4209__,
    new_new_n4210__, new_new_n4211__, new_new_n4212__, new_new_n4213__,
    new_new_n4214__, new_new_n4215__, new_new_n4216__, new_new_n4217__,
    new_new_n4218__, new_new_n4219__, new_new_n4220__, new_new_n4221__,
    new_new_n4222__, new_new_n4223__, new_new_n4224__, new_new_n4225__,
    new_new_n4226__, new_new_n4227__, new_new_n4228__, new_new_n4229__,
    new_new_n4230__, new_new_n4231__, new_new_n4232__, new_new_n4233__,
    new_new_n4234__, new_new_n4235__, new_new_n4236__, new_new_n4237__,
    new_new_n4238__, new_new_n4239__, new_new_n4240__, new_new_n4241__,
    new_new_n4242__, new_new_n4243__, new_new_n4244__, new_new_n4245__,
    new_new_n4246__, new_new_n4247__, new_new_n4248__, new_new_n4249__,
    new_new_n4250__, new_new_n4251__, new_new_n4252__, new_new_n4253__,
    new_new_n4254__, new_new_n4255__, new_new_n4256__, new_new_n4257__,
    new_new_n4258__, new_new_n4259__, new_new_n4260__, new_new_n4261__,
    new_new_n4262__, new_new_n4263__, new_new_n4264__, new_new_n4265__,
    new_new_n4266__, new_new_n4267__, new_new_n4268__, new_new_n4269__,
    new_new_n4270__, new_new_n4271__, new_new_n4272__, new_new_n4273__,
    new_new_n4274__, new_new_n4275__, new_new_n4276__, new_new_n4277__,
    new_new_n4278__, new_new_n4279__, new_new_n4280__, new_new_n4281__,
    new_new_n4282__, new_new_n4283__, new_new_n4284__, new_new_n4285__,
    new_new_n4286__, new_new_n4287__, new_new_n4288__, new_new_n4289__,
    new_new_n4290__, new_new_n4291__, new_new_n4292__, new_new_n4293__,
    new_new_n4294__, new_new_n4295__, new_new_n4296__, new_new_n4297__,
    new_new_n4298__, new_new_n4299__, new_new_n4300__, new_new_n4301__,
    new_new_n4302__, new_new_n4303__, new_new_n4304__, new_new_n4305__,
    new_new_n4306__, new_new_n4307__, new_new_n4308__, new_new_n4309__,
    new_new_n4310__, new_new_n4311__, new_new_n4312__, new_new_n4313__,
    new_new_n4314__, new_new_n4315__, new_new_n4316__, new_new_n4317__,
    new_new_n4318__, new_new_n4319__, new_new_n4320__, new_new_n4321__,
    new_new_n4322__, new_new_n4323__, new_new_n4324__, new_new_n4325__,
    new_new_n4326__, new_new_n4327__, new_new_n4328__, new_new_n4329__,
    new_new_n4330__, new_new_n4331__, new_new_n4332__, new_new_n4333__,
    new_new_n4334__, new_new_n4335__, new_new_n4336__, new_new_n4337__,
    new_new_n4338__, new_new_n4339__, new_new_n4340__, new_new_n4341__,
    new_new_n4342__, new_new_n4343__, new_new_n4344__, new_new_n4345__,
    new_new_n4346__, new_new_n4347__, new_new_n4348__, new_new_n4349__,
    new_new_n4350__, new_new_n4351__, new_new_n4352__, new_new_n4353__,
    new_new_n4354__, new_new_n4355__, new_new_n4356__, new_new_n4357__,
    new_new_n4358__, new_new_n4359__, new_new_n4360__, new_new_n4361__,
    new_new_n4362__, new_new_n4363__, new_new_n4364__, new_new_n4365__,
    new_new_n4366__, new_new_n4367__, new_new_n4368__, new_new_n4369__,
    new_new_n4370__, new_new_n4371__, new_new_n4372__, new_new_n4373__,
    new_new_n4374__, new_new_n4375__, new_new_n4376__, new_new_n4377__,
    new_new_n4378__, new_new_n4379__, new_new_n4380__, new_new_n4381__,
    new_new_n4382__, new_new_n4383__, new_new_n4384__, new_new_n4385__,
    new_new_n4386__, new_new_n4387__, new_new_n4388__, new_new_n4389__,
    new_new_n4390__, new_new_n4391__, new_new_n4392__, new_new_n4393__,
    new_new_n4394__, new_new_n4395__, new_new_n4396__, new_new_n4397__,
    new_new_n4398__, new_new_n4399__, new_new_n4400__, new_new_n4401__,
    new_new_n4402__, new_new_n4403__, new_new_n4404__, new_new_n4405__,
    new_new_n4406__, new_new_n4407__, new_new_n4408__, new_new_n4409__,
    new_new_n4410__, new_new_n4411__, new_new_n4412__, new_new_n4413__,
    new_new_n4414__, new_new_n4415__, new_new_n4416__, new_new_n4417__,
    new_new_n4418__, new_new_n4419__, new_new_n4420__, new_new_n4421__,
    new_new_n4422__, new_new_n4423__, new_new_n4424__, new_new_n4425__,
    new_new_n4426__, new_new_n4427__, new_new_n4428__, new_new_n4429__,
    new_new_n4430__, new_new_n4431__, new_new_n4432__, new_new_n4433__,
    new_new_n4434__, new_new_n4435__, new_new_n4436__, new_new_n4437__,
    new_new_n4438__, new_new_n4439__, new_new_n4440__, new_new_n4441__,
    new_new_n4442__, new_new_n4443__, new_new_n4444__, new_new_n4445__,
    new_new_n4446__, new_new_n4447__, new_new_n4448__, new_new_n4449__,
    new_new_n4450__, new_new_n4451__, new_new_n4452__, new_new_n4453__,
    new_new_n4454__, new_new_n4455__, new_new_n4456__, new_new_n4457__,
    new_new_n4458__, new_new_n4459__, new_new_n4460__, new_new_n4461__,
    new_new_n4462__, new_new_n4463__, new_new_n4464__, new_new_n4465__,
    new_new_n4466__, new_new_n4467__, new_new_n4468__, new_new_n4469__,
    new_new_n4470__, new_new_n4471__, new_new_n4472__, new_new_n4473__,
    new_new_n4474__, new_new_n4475__, new_new_n4476__, new_new_n4477__,
    new_new_n4478__, new_new_n4479__, new_new_n4480__, new_new_n4481__,
    new_new_n4482__, new_new_n4483__, new_new_n4484__, new_new_n4485__,
    new_new_n4486__, new_new_n4487__, new_new_n4488__, new_new_n4489__,
    new_new_n4490__, new_new_n4491__, new_new_n4492__, new_new_n4493__,
    new_new_n4494__, new_new_n4495__, new_new_n4496__, new_new_n4497__,
    new_new_n4498__, new_new_n4499__, new_new_n4500__, new_new_n4501__,
    new_new_n4502__, new_new_n4503__, new_new_n4504__, new_new_n4505__,
    new_new_n4506__, new_new_n4507__, new_new_n4508__, new_new_n4509__,
    new_new_n4510__, new_new_n4511__, new_new_n4512__, new_new_n4513__,
    new_new_n4514__, new_new_n4515__, new_new_n4516__, new_new_n4517__,
    new_new_n4518__, new_new_n4519__, new_new_n4520__, new_new_n4521__,
    new_new_n4522__, new_new_n4523__, new_new_n4524__, new_new_n4525__,
    new_new_n4526__, new_new_n4527__, new_new_n4528__, new_new_n4529__,
    new_new_n4530__, new_new_n4531__, new_new_n4532__, new_new_n4533__,
    new_new_n4534__, new_new_n4535__, new_new_n4536__, new_new_n4537__,
    new_new_n4538__, new_new_n4539__, new_new_n4540__, new_new_n4541__,
    new_new_n4542__, new_new_n4543__, new_new_n4544__, new_new_n4545__,
    new_new_n4546__, new_new_n4547__, new_new_n4548__, new_new_n4549__,
    new_new_n4550__, new_new_n4551__, new_new_n4552__, new_new_n4553__,
    new_new_n4554__, new_new_n4555__, new_new_n4556__, new_new_n4557__,
    new_new_n4558__, new_new_n4559__, new_new_n4560__, new_new_n4561__,
    new_new_n4562__, new_new_n4563__, new_new_n4564__, new_new_n4565__,
    new_new_n4566__, new_new_n4567__, new_new_n4568__, new_new_n4569__,
    new_new_n4570__, new_new_n4571__, new_new_n4572__, new_new_n4573__,
    new_new_n4574__, new_new_n4575__, new_new_n4576__, new_new_n4577__,
    new_new_n4578__, new_new_n4579__, new_new_n4580__, new_new_n4581__,
    new_new_n4582__, new_new_n4583__, new_new_n4584__, new_new_n4585__,
    new_new_n4586__, new_new_n4587__, new_new_n4588__, new_new_n4589__,
    new_new_n4590__, new_new_n4591__, new_new_n4592__, new_new_n4593__,
    new_new_n4594__, new_new_n4595__, new_new_n4596__, new_new_n4597__,
    new_new_n4598__, new_new_n4599__, new_new_n4600__, new_new_n4601__,
    new_new_n4602__, new_new_n4603__, new_new_n4604__, new_new_n4605__,
    new_new_n4606__, new_new_n4607__, new_new_n4608__, new_new_n4609__,
    new_new_n4610__, new_new_n4611__, new_new_n4612__, new_new_n4613__,
    new_new_n4614__, new_new_n4615__, new_new_n4616__, new_new_n4617__,
    new_new_n4618__, new_new_n4619__, new_new_n4620__, new_new_n4621__,
    new_new_n4622__, new_new_n4623__, new_new_n4624__, new_new_n4625__,
    new_new_n4626__, new_new_n4627__, new_new_n4628__, new_new_n4629__,
    new_new_n4630__, new_new_n4631__, new_new_n4632__, new_new_n4633__,
    new_new_n4634__, new_new_n4635__, new_new_n4636__, new_new_n4637__,
    new_new_n4638__, new_new_n4639__, new_new_n4640__, new_new_n4641__,
    new_new_n4642__, new_new_n4643__, new_new_n4644__, new_new_n4645__,
    new_new_n4646__, new_new_n4647__, new_new_n4648__, new_new_n4649__,
    new_new_n4650__, new_new_n4651__, new_new_n4652__, new_new_n4653__,
    new_new_n4654__, new_new_n4655__, new_new_n4656__, new_new_n4657__,
    new_new_n4658__, new_new_n4659__, new_new_n4660__, new_new_n4661__,
    new_new_n4662__, new_new_n4663__, new_new_n4664__, new_new_n4665__,
    new_new_n4666__, new_new_n4667__, new_new_n4668__, new_new_n4669__,
    new_new_n4670__, new_new_n4671__, new_new_n4672__, new_new_n4673__,
    new_new_n4674__, new_new_n4675__, new_new_n4676__, new_new_n4677__,
    new_new_n4678__, new_new_n4679__, new_new_n4680__, new_new_n4681__,
    new_new_n4682__, new_new_n4683__, new_new_n4684__, new_new_n4685__,
    new_new_n4686__, new_new_n4687__, new_new_n4688__, new_new_n4689__,
    new_new_n4690__, new_new_n4691__, new_new_n4692__, new_new_n4693__,
    new_new_n4695__, new_new_n4696__, new_new_n4697__, new_new_n4698__,
    new_new_n4699__, new_new_n4700__, new_new_n4701__, new_new_n4702__,
    new_new_n4703__, new_new_n4704__, new_new_n4705__, new_new_n4706__,
    new_new_n4707__, new_new_n4708__, new_new_n4709__, new_new_n4710__,
    new_new_n4711__, new_new_n4712__, new_new_n4713__, new_new_n4714__,
    new_new_n4715__, new_new_n4716__, new_new_n4717__, new_new_n4718__,
    new_new_n4719__, new_new_n4720__, new_new_n4721__, new_new_n4722__,
    new_new_n4723__, new_new_n4724__, new_new_n4725__, new_new_n4726__,
    new_new_n4727__, new_new_n4728__, new_new_n4729__, new_new_n4730__,
    new_new_n4731__, new_new_n4732__, new_new_n4733__, new_new_n4734__,
    new_new_n4735__, new_new_n4736__, new_new_n4737__, new_new_n4738__,
    new_new_n4739__, new_new_n4740__, new_new_n4741__, new_new_n4742__,
    new_new_n4743__, new_new_n4744__, new_new_n4745__, new_new_n4746__,
    new_new_n4747__, new_new_n4748__, new_new_n4749__, new_new_n4750__,
    new_new_n4751__, new_new_n4752__, new_new_n4753__, new_new_n4754__,
    new_new_n4755__, new_new_n4756__, new_new_n4757__, new_new_n4758__,
    new_new_n4759__, new_new_n4760__, new_new_n4761__, new_new_n4762__,
    new_new_n4763__, new_new_n4764__, new_new_n4765__, new_new_n4766__,
    new_new_n4767__, new_new_n4768__, new_new_n4769__, new_new_n4770__,
    new_new_n4771__, new_new_n4772__, new_new_n4773__, new_new_n4774__,
    new_new_n4775__, new_new_n4776__, new_new_n4777__, new_new_n4778__,
    new_new_n4779__, new_new_n4780__, new_new_n4781__, new_new_n4782__,
    new_new_n4783__, new_new_n4784__, new_new_n4785__, new_new_n4786__,
    new_new_n4787__, new_new_n4788__, new_new_n4789__, new_new_n4790__,
    new_new_n4791__, new_new_n4792__, new_new_n4793__, new_new_n4794__,
    new_new_n4795__, new_new_n4796__, new_new_n4797__, new_new_n4798__,
    new_new_n4799__, new_new_n4800__, new_new_n4801__, new_new_n4802__,
    new_new_n4803__, new_new_n4804__, new_new_n4805__, new_new_n4806__,
    new_new_n4807__, new_new_n4808__, new_new_n4809__, new_new_n4810__,
    new_new_n4811__, new_new_n4812__, new_new_n4813__, new_new_n4814__,
    new_new_n4815__, new_new_n4816__, new_new_n4817__, new_new_n4818__,
    new_new_n4819__, new_new_n4820__, new_new_n4821__, new_new_n4822__,
    new_new_n4823__, new_new_n4824__, new_new_n4825__, new_new_n4826__,
    new_new_n4827__, new_new_n4828__, new_new_n4829__, new_new_n4830__,
    new_new_n4831__, new_new_n4832__, new_new_n4833__, new_new_n4834__,
    new_new_n4835__, new_new_n4836__, new_new_n4837__, new_new_n4838__,
    new_new_n4839__, new_new_n4840__, new_new_n4841__, new_new_n4842__,
    new_new_n4843__, new_new_n4844__, new_new_n4845__, new_new_n4846__,
    new_new_n4847__, new_new_n4848__, new_new_n4849__, new_new_n4850__,
    new_new_n4851__, new_new_n4852__, new_new_n4853__, new_new_n4854__,
    new_new_n4855__, new_new_n4856__, new_new_n4857__, new_new_n4858__,
    new_new_n4859__, new_new_n4860__, new_new_n4861__, new_new_n4862__,
    new_new_n4863__, new_new_n4864__, new_new_n4865__, new_new_n4866__,
    new_new_n4867__, new_new_n4868__, new_new_n4869__, new_new_n4870__,
    new_new_n4871__, new_new_n4872__, new_new_n4873__, new_new_n4874__,
    new_new_n4875__, new_new_n4876__, new_new_n4877__, new_new_n4878__,
    new_new_n4879__, new_new_n4880__, new_new_n4881__, new_new_n4882__,
    new_new_n4883__, new_new_n4884__, new_new_n4885__, new_new_n4886__,
    new_new_n4887__, new_new_n4888__, new_new_n4889__, new_new_n4890__,
    new_new_n4891__, new_new_n4892__, new_new_n4893__, new_new_n4894__,
    new_new_n4895__, new_new_n4896__, new_new_n4897__, new_new_n4898__,
    new_new_n4899__, new_new_n4900__, new_new_n4901__, new_new_n4902__,
    new_new_n4903__, new_new_n4904__, new_new_n4905__, new_new_n4906__,
    new_new_n4907__, new_new_n4908__, new_new_n4909__, new_new_n4910__,
    new_new_n4911__, new_new_n4912__, new_new_n4913__, new_new_n4915__,
    new_new_n4916__, new_new_n4917__, new_new_n4918__, new_new_n4919__,
    new_new_n4920__, new_new_n4921__, new_new_n4922__, new_new_n4923__,
    new_new_n4924__, new_new_n4925__, new_new_n4926__, new_new_n4927__,
    new_new_n4928__, new_new_n4929__, new_new_n4930__, new_new_n4931__,
    new_new_n4932__, new_new_n4933__, new_new_n4934__, new_new_n4935__,
    new_new_n4936__, new_new_n4937__, new_new_n4938__, new_new_n4939__,
    new_new_n4940__, new_new_n4941__, new_new_n4942__, new_new_n4943__,
    new_new_n4944__, new_new_n4945__, new_new_n4946__, new_new_n4947__,
    new_new_n4948__, new_new_n4949__, new_new_n4950__, new_new_n4951__,
    new_new_n4952__, new_new_n4953__, new_new_n4954__, new_new_n4955__,
    new_new_n4956__, new_new_n4957__, new_new_n4958__, new_new_n4959__,
    new_new_n4960__, new_new_n4961__, new_new_n4962__, new_new_n4963__,
    new_new_n4964__, new_new_n4965__, new_new_n4966__, new_new_n4967__,
    new_new_n4968__, new_new_n4969__, new_new_n4970__, new_new_n4971__,
    new_new_n4972__, new_new_n4973__, new_new_n4974__, new_new_n4975__,
    new_new_n4976__, new_new_n4977__, new_new_n4978__, new_new_n4979__,
    new_new_n4980__, new_new_n4981__, new_new_n4982__, new_new_n4983__,
    new_new_n4984__, new_new_n4985__, new_new_n4986__, new_new_n4987__,
    new_new_n4988__, new_new_n4989__, new_new_n4990__, new_new_n4991__,
    new_new_n4992__, new_new_n4993__, new_new_n4994__, new_new_n4995__,
    new_new_n4996__, new_new_n4997__, new_new_n4998__, new_new_n4999__,
    new_new_n5000__, new_new_n5001__, new_new_n5002__, new_new_n5003__,
    new_new_n5004__, new_new_n5005__, new_new_n5006__, new_new_n5007__,
    new_new_n5008__, new_new_n5009__, new_new_n5010__, new_new_n5011__,
    new_new_n5012__, new_new_n5013__, new_new_n5014__, new_new_n5015__,
    new_new_n5016__, new_new_n5017__, new_new_n5018__, new_new_n5019__,
    new_new_n5020__, new_new_n5021__, new_new_n5022__, new_new_n5023__,
    new_new_n5024__, new_new_n5025__, new_new_n5026__, new_new_n5027__,
    new_new_n5028__, new_new_n5029__, new_new_n5030__, new_new_n5031__,
    new_new_n5032__, new_new_n5033__, new_new_n5034__, new_new_n5035__,
    new_new_n5036__, new_new_n5037__, new_new_n5038__, new_new_n5039__,
    new_new_n5040__, new_new_n5041__, new_new_n5042__, new_new_n5043__,
    new_new_n5044__, new_new_n5045__, new_new_n5046__, new_new_n5047__,
    new_new_n5048__, new_new_n5049__, new_new_n5050__, new_new_n5051__,
    new_new_n5052__, new_new_n5053__, new_new_n5054__, new_new_n5055__,
    new_new_n5056__, new_new_n5057__, new_new_n5058__, new_new_n5059__,
    new_new_n5060__, new_new_n5061__, new_new_n5062__, new_new_n5063__,
    new_new_n5064__, new_new_n5065__, new_new_n5066__, new_new_n5067__,
    new_new_n5068__, new_new_n5069__, new_new_n5070__, new_new_n5071__,
    new_new_n5072__, new_new_n5073__, new_new_n5074__, new_new_n5075__,
    new_new_n5076__, new_new_n5077__, new_new_n5078__, new_new_n5079__,
    new_new_n5080__, new_new_n5081__, new_new_n5082__, new_new_n5083__,
    new_new_n5084__, new_new_n5085__, new_new_n5086__, new_new_n5087__,
    new_new_n5088__, new_new_n5089__, new_new_n5090__, new_new_n5091__,
    new_new_n5092__, new_new_n5093__, new_new_n5094__, new_new_n5095__,
    new_new_n5096__, new_new_n5097__, new_new_n5098__, new_new_n5099__,
    new_new_n5100__, new_new_n5101__, new_new_n5102__, new_new_n5103__,
    new_new_n5104__, new_new_n5105__, new_new_n5106__, new_new_n5107__,
    new_new_n5108__, new_new_n5109__, new_new_n5110__, new_new_n5112__,
    new_new_n5113__, new_new_n5114__, new_new_n5115__, new_new_n5116__,
    new_new_n5117__, new_new_n5118__, new_new_n5119__, new_new_n5120__,
    new_new_n5121__, new_new_n5122__, new_new_n5123__, new_new_n5124__,
    new_new_n5125__, new_new_n5126__, new_new_n5127__, new_new_n5128__,
    new_new_n5129__, new_new_n5130__, new_new_n5131__, new_new_n5132__,
    new_new_n5133__, new_new_n5134__, new_new_n5135__, new_new_n5136__,
    new_new_n5137__, new_new_n5138__, new_new_n5139__, new_new_n5140__,
    new_new_n5141__, new_new_n5142__, new_new_n5143__, new_new_n5144__,
    new_new_n5145__, new_new_n5146__, new_new_n5147__, new_new_n5148__,
    new_new_n5149__, new_new_n5150__, new_new_n5151__, new_new_n5152__,
    new_new_n5153__, new_new_n5154__, new_new_n5155__, new_new_n5156__,
    new_new_n5157__, new_new_n5158__, new_new_n5159__, new_new_n5160__,
    new_new_n5161__, new_new_n5162__, new_new_n5163__, new_new_n5164__,
    new_new_n5165__, new_new_n5166__, new_new_n5167__, new_new_n5168__,
    new_new_n5169__, new_new_n5170__, new_new_n5171__, new_new_n5172__,
    new_new_n5173__, new_new_n5174__, new_new_n5175__, new_new_n5176__,
    new_new_n5177__, new_new_n5178__, new_new_n5179__, new_new_n5180__,
    new_new_n5181__, new_new_n5182__, new_new_n5183__, new_new_n5184__,
    new_new_n5185__, new_new_n5186__, new_new_n5187__, new_new_n5188__,
    new_new_n5189__, new_new_n5190__, new_new_n5191__, new_new_n5192__,
    new_new_n5193__, new_new_n5194__, new_new_n5195__, new_new_n5196__,
    new_new_n5197__, new_new_n5198__, new_new_n5199__, new_new_n5200__,
    new_new_n5201__, new_new_n5202__, new_new_n5203__, new_new_n5204__,
    new_new_n5205__, new_new_n5206__, new_new_n5207__, new_new_n5208__,
    new_new_n5209__, new_new_n5210__, new_new_n5211__, new_new_n5212__,
    new_new_n5213__, new_new_n5214__, new_new_n5215__, new_new_n5216__,
    new_new_n5217__, new_new_n5218__, new_new_n5219__, new_new_n5220__,
    new_new_n5221__, new_new_n5222__, new_new_n5223__, new_new_n5224__,
    new_new_n5225__, new_new_n5226__, new_new_n5227__, new_new_n5228__,
    new_new_n5229__, new_new_n5230__, new_new_n5231__, new_new_n5232__,
    new_new_n5233__, new_new_n5234__, new_new_n5235__, new_new_n5236__,
    new_new_n5237__, new_new_n5238__, new_new_n5239__, new_new_n5240__,
    new_new_n5241__, new_new_n5242__, new_new_n5243__, new_new_n5244__,
    new_new_n5245__, new_new_n5246__, new_new_n5247__, new_new_n5248__,
    new_new_n5249__, new_new_n5250__, new_new_n5251__, new_new_n5252__,
    new_new_n5253__, new_new_n5254__, new_new_n5255__, new_new_n5256__,
    new_new_n5257__, new_new_n5258__, new_new_n5259__, new_new_n5260__,
    new_new_n5261__, new_new_n5262__, new_new_n5263__, new_new_n5264__,
    new_new_n5265__, new_new_n5266__, new_new_n5267__, new_new_n5268__,
    new_new_n5269__, new_new_n5270__, new_new_n5271__, new_new_n5272__,
    new_new_n5273__, new_new_n5274__, new_new_n5275__, new_new_n5276__,
    new_new_n5277__, new_new_n5278__, new_new_n5279__, new_new_n5280__,
    new_new_n5281__, new_new_n5282__, new_new_n5283__, new_new_n5284__,
    new_new_n5285__, new_new_n5286__, new_new_n5287__, new_new_n5288__,
    new_new_n5289__, new_new_n5290__, new_new_n5291__, new_new_n5292__,
    new_new_n5294__, new_new_n5295__, new_new_n5296__, new_new_n5297__,
    new_new_n5298__, new_new_n5299__, new_new_n5300__, new_new_n5301__,
    new_new_n5302__, new_new_n5303__, new_new_n5304__, new_new_n5305__,
    new_new_n5306__, new_new_n5307__, new_new_n5308__, new_new_n5309__,
    new_new_n5310__, new_new_n5311__, new_new_n5312__, new_new_n5313__,
    new_new_n5314__, new_new_n5315__, new_new_n5316__, new_new_n5317__,
    new_new_n5318__, new_new_n5319__, new_new_n5320__, new_new_n5321__,
    new_new_n5322__, new_new_n5323__, new_new_n5324__, new_new_n5325__,
    new_new_n5326__, new_new_n5327__, new_new_n5328__, new_new_n5329__,
    new_new_n5330__, new_new_n5331__, new_new_n5332__, new_new_n5333__,
    new_new_n5334__, new_new_n5335__, new_new_n5336__, new_new_n5337__,
    new_new_n5338__, new_new_n5339__, new_new_n5340__, new_new_n5341__,
    new_new_n5342__, new_new_n5343__, new_new_n5344__, new_new_n5345__,
    new_new_n5346__, new_new_n5347__, new_new_n5348__, new_new_n5349__,
    new_new_n5350__, new_new_n5351__, new_new_n5352__, new_new_n5353__,
    new_new_n5354__, new_new_n5355__, new_new_n5356__, new_new_n5357__,
    new_new_n5358__, new_new_n5359__, new_new_n5360__, new_new_n5361__,
    new_new_n5362__, new_new_n5363__, new_new_n5364__, new_new_n5365__,
    new_new_n5366__, new_new_n5367__, new_new_n5368__, new_new_n5369__,
    new_new_n5370__, new_new_n5371__, new_new_n5372__, new_new_n5373__,
    new_new_n5374__, new_new_n5375__, new_new_n5376__, new_new_n5377__,
    new_new_n5378__, new_new_n5379__, new_new_n5380__, new_new_n5381__,
    new_new_n5382__, new_new_n5383__, new_new_n5384__, new_new_n5385__,
    new_new_n5386__, new_new_n5387__, new_new_n5388__, new_new_n5389__,
    new_new_n5390__, new_new_n5391__, new_new_n5392__, new_new_n5393__,
    new_new_n5394__, new_new_n5395__, new_new_n5396__, new_new_n5397__,
    new_new_n5398__, new_new_n5399__, new_new_n5400__, new_new_n5401__,
    new_new_n5402__, new_new_n5403__, new_new_n5404__, new_new_n5405__,
    new_new_n5406__, new_new_n5407__, new_new_n5408__, new_new_n5409__,
    new_new_n5410__, new_new_n5411__, new_new_n5412__, new_new_n5413__,
    new_new_n5414__, new_new_n5415__, new_new_n5416__, new_new_n5417__,
    new_new_n5418__, new_new_n5419__, new_new_n5420__, new_new_n5421__,
    new_new_n5422__, new_new_n5423__, new_new_n5424__, new_new_n5425__,
    new_new_n5426__, new_new_n5427__, new_new_n5428__, new_new_n5429__,
    new_new_n5430__, new_new_n5431__, new_new_n5432__, new_new_n5433__,
    new_new_n5434__, new_new_n5435__, new_new_n5436__, new_new_n5437__,
    new_new_n5438__, new_new_n5439__, new_new_n5440__, new_new_n5441__,
    new_new_n5442__, new_new_n5443__, new_new_n5444__, new_new_n5445__,
    new_new_n5446__, new_new_n5447__, new_new_n5448__, new_new_n5449__,
    new_new_n5450__, new_new_n5451__, new_new_n5452__, new_new_n5454__,
    new_new_n5455__, new_new_n5456__, new_new_n5457__, new_new_n5458__,
    new_new_n5459__, new_new_n5460__, new_new_n5461__, new_new_n5462__,
    new_new_n5463__, new_new_n5464__, new_new_n5465__, new_new_n5466__,
    new_new_n5467__, new_new_n5468__, new_new_n5469__, new_new_n5470__,
    new_new_n5471__, new_new_n5472__, new_new_n5473__, new_new_n5474__,
    new_new_n5475__, new_new_n5476__, new_new_n5477__, new_new_n5478__,
    new_new_n5479__, new_new_n5480__, new_new_n5481__, new_new_n5482__,
    new_new_n5483__, new_new_n5484__, new_new_n5485__, new_new_n5486__,
    new_new_n5487__, new_new_n5488__, new_new_n5489__, new_new_n5490__,
    new_new_n5491__, new_new_n5492__, new_new_n5493__, new_new_n5494__,
    new_new_n5495__, new_new_n5496__, new_new_n5497__, new_new_n5498__,
    new_new_n5499__, new_new_n5500__, new_new_n5501__, new_new_n5502__,
    new_new_n5503__, new_new_n5504__, new_new_n5505__, new_new_n5506__,
    new_new_n5507__, new_new_n5508__, new_new_n5509__, new_new_n5510__,
    new_new_n5511__, new_new_n5512__, new_new_n5513__, new_new_n5514__,
    new_new_n5515__, new_new_n5516__, new_new_n5517__, new_new_n5518__,
    new_new_n5519__, new_new_n5520__, new_new_n5521__, new_new_n5522__,
    new_new_n5523__, new_new_n5524__, new_new_n5525__, new_new_n5526__,
    new_new_n5527__, new_new_n5528__, new_new_n5529__, new_new_n5530__,
    new_new_n5531__, new_new_n5532__, new_new_n5533__, new_new_n5534__,
    new_new_n5535__, new_new_n5536__, new_new_n5537__, new_new_n5538__,
    new_new_n5539__, new_new_n5540__, new_new_n5541__, new_new_n5542__,
    new_new_n5543__, new_new_n5544__, new_new_n5545__, new_new_n5546__,
    new_new_n5547__, new_new_n5548__, new_new_n5549__, new_new_n5550__,
    new_new_n5551__, new_new_n5552__, new_new_n5553__, new_new_n5554__,
    new_new_n5555__, new_new_n5556__, new_new_n5557__, new_new_n5558__,
    new_new_n5559__, new_new_n5560__, new_new_n5561__, new_new_n5562__,
    new_new_n5563__, new_new_n5564__, new_new_n5565__, new_new_n5566__,
    new_new_n5567__, new_new_n5568__, new_new_n5569__, new_new_n5570__,
    new_new_n5571__, new_new_n5572__, new_new_n5573__, new_new_n5574__,
    new_new_n5575__, new_new_n5576__, new_new_n5577__, new_new_n5578__,
    new_new_n5579__, new_new_n5580__, new_new_n5581__, new_new_n5582__,
    new_new_n5583__, new_new_n5584__, new_new_n5585__, new_new_n5586__,
    new_new_n5587__, new_new_n5588__, new_new_n5589__, new_new_n5590__,
    new_new_n5591__, new_new_n5592__, new_new_n5593__, new_new_n5594__,
    new_new_n5595__, new_new_n5596__, new_new_n5597__, new_new_n5598__,
    new_new_n5599__, new_new_n5600__, new_new_n5601__, new_new_n5602__,
    new_new_n5603__, new_new_n5604__, new_new_n5605__, new_new_n5606__,
    new_new_n5607__, new_new_n5608__, new_new_n5609__, new_new_n5610__,
    new_new_n5611__, new_new_n5612__, new_new_n5613__, new_new_n5614__,
    new_new_n5615__, new_new_n5616__, new_new_n5617__, new_new_n5618__,
    new_new_n5619__, new_new_n5620__, new_new_n5621__, new_new_n5622__,
    new_new_n5623__, new_new_n5624__, new_new_n5625__, new_new_n5626__,
    new_new_n5627__, new_new_n5628__, new_new_n5629__, new_new_n5630__,
    new_new_n5631__, new_new_n5632__, new_new_n5633__, new_new_n5634__,
    new_new_n5635__, new_new_n5636__, new_new_n5637__, new_new_n5638__,
    new_new_n5639__, new_new_n5640__, new_new_n5641__, new_new_n5642__,
    new_new_n5643__, new_new_n5644__, new_new_n5645__, new_new_n5647__,
    new_new_n5648__, new_new_n5649__, new_new_n5650__, new_new_n5651__,
    new_new_n5652__, new_new_n5653__, new_new_n5654__, new_new_n5655__,
    new_new_n5656__, new_new_n5657__, new_new_n5658__, new_new_n5659__,
    new_new_n5660__, new_new_n5661__, new_new_n5662__, new_new_n5663__,
    new_new_n5664__, new_new_n5665__, new_new_n5666__, new_new_n5667__,
    new_new_n5668__, new_new_n5669__, new_new_n5670__, new_new_n5671__,
    new_new_n5672__, new_new_n5673__, new_new_n5674__, new_new_n5675__,
    new_new_n5676__, new_new_n5677__, new_new_n5678__, new_new_n5679__,
    new_new_n5680__, new_new_n5681__, new_new_n5682__, new_new_n5683__,
    new_new_n5684__, new_new_n5685__, new_new_n5686__, new_new_n5687__,
    new_new_n5688__, new_new_n5689__, new_new_n5690__, new_new_n5691__,
    new_new_n5692__, new_new_n5693__, new_new_n5694__, new_new_n5695__,
    new_new_n5696__, new_new_n5697__, new_new_n5698__, new_new_n5699__,
    new_new_n5700__, new_new_n5701__, new_new_n5702__, new_new_n5703__,
    new_new_n5704__, new_new_n5705__, new_new_n5706__, new_new_n5707__,
    new_new_n5708__, new_new_n5709__, new_new_n5710__, new_new_n5711__,
    new_new_n5712__, new_new_n5713__, new_new_n5714__, new_new_n5715__,
    new_new_n5716__, new_new_n5717__, new_new_n5718__, new_new_n5719__,
    new_new_n5720__, new_new_n5721__, new_new_n5722__, new_new_n5723__,
    new_new_n5724__, new_new_n5725__, new_new_n5726__, new_new_n5727__,
    new_new_n5728__, new_new_n5729__, new_new_n5730__, new_new_n5731__,
    new_new_n5732__, new_new_n5733__, new_new_n5734__, new_new_n5735__,
    new_new_n5736__, new_new_n5737__, new_new_n5738__, new_new_n5739__,
    new_new_n5740__, new_new_n5741__, new_new_n5742__, new_new_n5743__,
    new_new_n5744__, new_new_n5745__, new_new_n5746__, new_new_n5747__,
    new_new_n5748__, new_new_n5749__, new_new_n5750__, new_new_n5751__,
    new_new_n5752__, new_new_n5753__, new_new_n5754__, new_new_n5755__,
    new_new_n5756__, new_new_n5757__, new_new_n5758__, new_new_n5759__,
    new_new_n5760__, new_new_n5761__, new_new_n5762__, new_new_n5763__,
    new_new_n5764__, new_new_n5765__, new_new_n5766__, new_new_n5767__,
    new_new_n5768__, new_new_n5769__, new_new_n5770__, new_new_n5771__,
    new_new_n5772__, new_new_n5773__, new_new_n5774__, new_new_n5775__,
    new_new_n5776__, new_new_n5777__, new_new_n5778__, new_new_n5779__,
    new_new_n5780__, new_new_n5781__, new_new_n5782__, new_new_n5783__,
    new_new_n5784__, new_new_n5785__, new_new_n5786__, new_new_n5787__,
    new_new_n5788__, new_new_n5789__, new_new_n5790__, new_new_n5791__,
    new_new_n5792__, new_new_n5793__, new_new_n5794__, new_new_n5795__,
    new_new_n5796__, new_new_n5797__, new_new_n5798__, new_new_n5799__,
    new_new_n5800__, new_new_n5801__, new_new_n5802__, new_new_n5803__,
    new_new_n5804__, new_new_n5805__, new_new_n5806__, new_new_n5807__,
    new_new_n5808__, new_new_n5809__, new_new_n5810__, new_new_n5811__,
    new_new_n5812__, new_new_n5813__, new_new_n5814__, new_new_n5815__,
    new_new_n5816__, new_new_n5817__, new_new_n5818__, new_new_n5820__,
    new_new_n5821__, new_new_n5822__, new_new_n5823__, new_new_n5824__,
    new_new_n5825__, new_new_n5826__, new_new_n5827__, new_new_n5828__,
    new_new_n5829__, new_new_n5830__, new_new_n5831__, new_new_n5832__,
    new_new_n5833__, new_new_n5834__, new_new_n5835__, new_new_n5836__,
    new_new_n5837__, new_new_n5838__, new_new_n5839__, new_new_n5840__,
    new_new_n5841__, new_new_n5842__, new_new_n5843__, new_new_n5844__,
    new_new_n5845__, new_new_n5846__, new_new_n5847__, new_new_n5848__,
    new_new_n5849__, new_new_n5850__, new_new_n5851__, new_new_n5852__,
    new_new_n5853__, new_new_n5854__, new_new_n5855__, new_new_n5856__,
    new_new_n5857__, new_new_n5858__, new_new_n5859__, new_new_n5860__,
    new_new_n5861__, new_new_n5862__, new_new_n5863__, new_new_n5864__,
    new_new_n5865__, new_new_n5866__, new_new_n5867__, new_new_n5868__,
    new_new_n5869__, new_new_n5870__, new_new_n5871__, new_new_n5872__,
    new_new_n5873__, new_new_n5874__, new_new_n5875__, new_new_n5876__,
    new_new_n5877__, new_new_n5878__, new_new_n5879__, new_new_n5880__,
    new_new_n5881__, new_new_n5882__, new_new_n5883__, new_new_n5884__,
    new_new_n5885__, new_new_n5886__, new_new_n5887__, new_new_n5888__,
    new_new_n5889__, new_new_n5890__, new_new_n5891__, new_new_n5892__,
    new_new_n5893__, new_new_n5894__, new_new_n5895__, new_new_n5896__,
    new_new_n5897__, new_new_n5898__, new_new_n5899__, new_new_n5900__,
    new_new_n5901__, new_new_n5902__, new_new_n5903__, new_new_n5904__,
    new_new_n5905__, new_new_n5906__, new_new_n5907__, new_new_n5908__,
    new_new_n5909__, new_new_n5910__, new_new_n5911__, new_new_n5912__,
    new_new_n5913__, new_new_n5914__, new_new_n5915__, new_new_n5916__,
    new_new_n5917__, new_new_n5918__, new_new_n5919__, new_new_n5920__,
    new_new_n5921__, new_new_n5922__, new_new_n5923__, new_new_n5924__,
    new_new_n5925__, new_new_n5926__, new_new_n5927__, new_new_n5928__,
    new_new_n5929__, new_new_n5930__, new_new_n5931__, new_new_n5932__,
    new_new_n5933__, new_new_n5934__, new_new_n5935__, new_new_n5936__,
    new_new_n5937__, new_new_n5938__, new_new_n5939__, new_new_n5940__,
    new_new_n5941__, new_new_n5942__, new_new_n5943__, new_new_n5944__,
    new_new_n5945__, new_new_n5946__, new_new_n5947__, new_new_n5948__,
    new_new_n5949__, new_new_n5950__, new_new_n5951__, new_new_n5952__,
    new_new_n5953__, new_new_n5954__, new_new_n5955__, new_new_n5956__,
    new_new_n5957__, new_new_n5958__, new_new_n5959__, new_new_n5960__,
    new_new_n5961__, new_new_n5962__, new_new_n5963__, new_new_n5964__,
    new_new_n5965__, new_new_n5966__, new_new_n5967__, new_new_n5968__,
    new_new_n5969__, new_new_n5971__, new_new_n5972__, new_new_n5973__,
    new_new_n5974__, new_new_n5975__, new_new_n5976__, new_new_n5977__,
    new_new_n5978__, new_new_n5979__, new_new_n5980__, new_new_n5981__,
    new_new_n5982__, new_new_n5983__, new_new_n5984__, new_new_n5985__,
    new_new_n5986__, new_new_n5987__, new_new_n5988__, new_new_n5989__,
    new_new_n5990__, new_new_n5991__, new_new_n5992__, new_new_n5993__,
    new_new_n5994__, new_new_n5995__, new_new_n5996__, new_new_n5997__,
    new_new_n5998__, new_new_n5999__, new_new_n6000__, new_new_n6001__,
    new_new_n6002__, new_new_n6003__, new_new_n6004__, new_new_n6005__,
    new_new_n6006__, new_new_n6007__, new_new_n6008__, new_new_n6009__,
    new_new_n6010__, new_new_n6011__, new_new_n6012__, new_new_n6013__,
    new_new_n6014__, new_new_n6015__, new_new_n6016__, new_new_n6017__,
    new_new_n6018__, new_new_n6019__, new_new_n6020__, new_new_n6021__,
    new_new_n6022__, new_new_n6023__, new_new_n6024__, new_new_n6025__,
    new_new_n6026__, new_new_n6027__, new_new_n6028__, new_new_n6029__,
    new_new_n6030__, new_new_n6031__, new_new_n6032__, new_new_n6033__,
    new_new_n6034__, new_new_n6035__, new_new_n6036__, new_new_n6037__,
    new_new_n6038__, new_new_n6039__, new_new_n6040__, new_new_n6041__,
    new_new_n6042__, new_new_n6043__, new_new_n6044__, new_new_n6045__,
    new_new_n6046__, new_new_n6047__, new_new_n6048__, new_new_n6049__,
    new_new_n6050__, new_new_n6051__, new_new_n6052__, new_new_n6053__,
    new_new_n6054__, new_new_n6055__, new_new_n6056__, new_new_n6057__,
    new_new_n6058__, new_new_n6059__, new_new_n6060__, new_new_n6061__,
    new_new_n6062__, new_new_n6063__, new_new_n6064__, new_new_n6065__,
    new_new_n6066__, new_new_n6067__, new_new_n6068__, new_new_n6069__,
    new_new_n6070__, new_new_n6071__, new_new_n6072__, new_new_n6073__,
    new_new_n6074__, new_new_n6075__, new_new_n6076__, new_new_n6077__,
    new_new_n6078__, new_new_n6079__, new_new_n6080__, new_new_n6081__,
    new_new_n6082__, new_new_n6083__, new_new_n6084__, new_new_n6085__,
    new_new_n6086__, new_new_n6087__, new_new_n6088__, new_new_n6089__,
    new_new_n6090__, new_new_n6091__, new_new_n6092__, new_new_n6093__,
    new_new_n6094__, new_new_n6095__, new_new_n6096__, new_new_n6097__,
    new_new_n6098__, new_new_n6099__, new_new_n6100__, new_new_n6101__,
    new_new_n6102__, new_new_n6103__, new_new_n6104__, new_new_n6105__,
    new_new_n6106__, new_new_n6107__, new_new_n6108__, new_new_n6109__,
    new_new_n6110__, new_new_n6111__, new_new_n6112__, new_new_n6113__,
    new_new_n6114__, new_new_n6115__, new_new_n6116__, new_new_n6117__,
    new_new_n6118__, new_new_n6119__, new_new_n6120__, new_new_n6121__,
    new_new_n6122__, new_new_n6123__, new_new_n6124__, new_new_n6125__,
    new_new_n6126__, new_new_n6127__, new_new_n6129__, new_new_n6130__,
    new_new_n6131__, new_new_n6132__, new_new_n6133__, new_new_n6134__,
    new_new_n6135__, new_new_n6136__, new_new_n6137__, new_new_n6138__,
    new_new_n6139__, new_new_n6140__, new_new_n6141__, new_new_n6142__,
    new_new_n6143__, new_new_n6144__, new_new_n6145__, new_new_n6146__,
    new_new_n6147__, new_new_n6148__, new_new_n6149__, new_new_n6150__,
    new_new_n6151__, new_new_n6152__, new_new_n6153__, new_new_n6154__,
    new_new_n6155__, new_new_n6156__, new_new_n6157__, new_new_n6158__,
    new_new_n6159__, new_new_n6160__, new_new_n6161__, new_new_n6162__,
    new_new_n6163__, new_new_n6164__, new_new_n6165__, new_new_n6166__,
    new_new_n6167__, new_new_n6168__, new_new_n6169__, new_new_n6170__,
    new_new_n6171__, new_new_n6172__, new_new_n6173__, new_new_n6174__,
    new_new_n6175__, new_new_n6176__, new_new_n6177__, new_new_n6178__,
    new_new_n6179__, new_new_n6180__, new_new_n6181__, new_new_n6182__,
    new_new_n6183__, new_new_n6184__, new_new_n6185__, new_new_n6186__,
    new_new_n6187__, new_new_n6188__, new_new_n6189__, new_new_n6190__,
    new_new_n6191__, new_new_n6192__, new_new_n6193__, new_new_n6194__,
    new_new_n6195__, new_new_n6196__, new_new_n6197__, new_new_n6198__,
    new_new_n6199__, new_new_n6200__, new_new_n6201__, new_new_n6202__,
    new_new_n6203__, new_new_n6204__, new_new_n6205__, new_new_n6206__,
    new_new_n6207__, new_new_n6208__, new_new_n6209__, new_new_n6210__,
    new_new_n6211__, new_new_n6212__, new_new_n6213__, new_new_n6214__,
    new_new_n6215__, new_new_n6216__, new_new_n6217__, new_new_n6218__,
    new_new_n6219__, new_new_n6220__, new_new_n6221__, new_new_n6222__,
    new_new_n6223__, new_new_n6224__, new_new_n6225__, new_new_n6226__,
    new_new_n6227__, new_new_n6228__, new_new_n6229__, new_new_n6230__,
    new_new_n6231__, new_new_n6232__, new_new_n6233__, new_new_n6234__,
    new_new_n6235__, new_new_n6236__, new_new_n6237__, new_new_n6238__,
    new_new_n6239__, new_new_n6240__, new_new_n6241__, new_new_n6242__,
    new_new_n6243__, new_new_n6244__, new_new_n6245__, new_new_n6246__,
    new_new_n6247__, new_new_n6248__, new_new_n6249__, new_new_n6250__,
    new_new_n6251__, new_new_n6252__, new_new_n6253__, new_new_n6254__,
    new_new_n6255__, new_new_n6256__, new_new_n6257__, new_new_n6258__,
    new_new_n6259__, new_new_n6260__, new_new_n6261__, new_new_n6262__,
    new_new_n6263__, new_new_n6264__, new_new_n6265__, new_new_n6266__,
    new_new_n6267__, new_new_n6268__, new_new_n6269__, new_new_n6270__,
    new_new_n6271__, new_new_n6273__, new_new_n6274__, new_new_n6275__,
    new_new_n6276__, new_new_n6277__, new_new_n6278__, new_new_n6279__,
    new_new_n6280__, new_new_n6281__, new_new_n6282__, new_new_n6283__,
    new_new_n6284__, new_new_n6285__, new_new_n6286__, new_new_n6287__,
    new_new_n6288__, new_new_n6289__, new_new_n6290__, new_new_n6291__,
    new_new_n6292__, new_new_n6293__, new_new_n6294__, new_new_n6295__,
    new_new_n6296__, new_new_n6297__, new_new_n6298__, new_new_n6299__,
    new_new_n6300__, new_new_n6301__, new_new_n6302__, new_new_n6303__,
    new_new_n6304__, new_new_n6305__, new_new_n6306__, new_new_n6307__,
    new_new_n6308__, new_new_n6309__, new_new_n6310__, new_new_n6311__,
    new_new_n6312__, new_new_n6313__, new_new_n6314__, new_new_n6315__,
    new_new_n6316__, new_new_n6317__, new_new_n6318__, new_new_n6319__,
    new_new_n6320__, new_new_n6321__, new_new_n6322__, new_new_n6323__,
    new_new_n6324__, new_new_n6325__, new_new_n6326__, new_new_n6327__,
    new_new_n6328__, new_new_n6329__, new_new_n6330__, new_new_n6331__,
    new_new_n6332__, new_new_n6333__, new_new_n6334__, new_new_n6335__,
    new_new_n6336__, new_new_n6337__, new_new_n6338__, new_new_n6339__,
    new_new_n6340__, new_new_n6341__, new_new_n6342__, new_new_n6343__,
    new_new_n6344__, new_new_n6345__, new_new_n6346__, new_new_n6347__,
    new_new_n6348__, new_new_n6349__, new_new_n6350__, new_new_n6351__,
    new_new_n6352__, new_new_n6353__, new_new_n6354__, new_new_n6355__,
    new_new_n6356__, new_new_n6357__, new_new_n6358__, new_new_n6359__,
    new_new_n6360__, new_new_n6361__, new_new_n6362__, new_new_n6363__,
    new_new_n6364__, new_new_n6365__, new_new_n6366__, new_new_n6367__,
    new_new_n6368__, new_new_n6369__, new_new_n6370__, new_new_n6371__,
    new_new_n6372__, new_new_n6373__, new_new_n6374__, new_new_n6375__,
    new_new_n6376__, new_new_n6377__, new_new_n6378__, new_new_n6379__,
    new_new_n6380__, new_new_n6381__, new_new_n6382__, new_new_n6383__,
    new_new_n6384__, new_new_n6385__, new_new_n6386__, new_new_n6387__,
    new_new_n6388__, new_new_n6389__, new_new_n6390__, new_new_n6391__,
    new_new_n6392__, new_new_n6393__, new_new_n6394__, new_new_n6395__,
    new_new_n6396__, new_new_n6397__, new_new_n6398__, new_new_n6399__,
    new_new_n6401__, new_new_n6402__, new_new_n6403__, new_new_n6404__,
    new_new_n6405__, new_new_n6406__, new_new_n6407__, new_new_n6408__,
    new_new_n6409__, new_new_n6410__, new_new_n6411__, new_new_n6412__,
    new_new_n6413__, new_new_n6414__, new_new_n6415__, new_new_n6416__,
    new_new_n6417__, new_new_n6418__, new_new_n6419__, new_new_n6420__,
    new_new_n6421__, new_new_n6422__, new_new_n6423__, new_new_n6424__,
    new_new_n6425__, new_new_n6426__, new_new_n6427__, new_new_n6428__,
    new_new_n6429__, new_new_n6430__, new_new_n6431__, new_new_n6432__,
    new_new_n6433__, new_new_n6434__, new_new_n6435__, new_new_n6436__,
    new_new_n6437__, new_new_n6438__, new_new_n6439__, new_new_n6440__,
    new_new_n6441__, new_new_n6442__, new_new_n6443__, new_new_n6444__,
    new_new_n6445__, new_new_n6446__, new_new_n6447__, new_new_n6448__,
    new_new_n6449__, new_new_n6450__, new_new_n6451__, new_new_n6452__,
    new_new_n6453__, new_new_n6454__, new_new_n6455__, new_new_n6456__,
    new_new_n6457__, new_new_n6458__, new_new_n6459__, new_new_n6460__,
    new_new_n6461__, new_new_n6462__, new_new_n6463__, new_new_n6464__,
    new_new_n6465__, new_new_n6466__, new_new_n6467__, new_new_n6468__,
    new_new_n6469__, new_new_n6470__, new_new_n6471__, new_new_n6472__,
    new_new_n6473__, new_new_n6474__, new_new_n6475__, new_new_n6476__,
    new_new_n6477__, new_new_n6478__, new_new_n6479__, new_new_n6480__,
    new_new_n6481__, new_new_n6482__, new_new_n6483__, new_new_n6484__,
    new_new_n6485__, new_new_n6486__, new_new_n6487__, new_new_n6488__,
    new_new_n6489__, new_new_n6490__, new_new_n6491__, new_new_n6492__,
    new_new_n6493__, new_new_n6494__, new_new_n6495__, new_new_n6496__,
    new_new_n6497__, new_new_n6498__, new_new_n6500__, new_new_n6501__,
    new_new_n6502__, new_new_n6503__, new_new_n6504__, new_new_n6505__,
    new_new_n6506__, new_new_n6507__, new_new_n6508__, new_new_n6509__,
    new_new_n6510__, new_new_n6511__, new_new_n6512__, new_new_n6513__,
    new_new_n6514__, new_new_n6515__, new_new_n6516__, new_new_n6517__,
    new_new_n6518__, new_new_n6519__, new_new_n6520__, new_new_n6521__,
    new_new_n6522__, new_new_n6523__, new_new_n6524__, new_new_n6525__,
    new_new_n6526__, new_new_n6527__, new_new_n6528__, new_new_n6529__,
    new_new_n6530__, new_new_n6531__, new_new_n6532__, new_new_n6533__,
    new_new_n6534__, new_new_n6535__, new_new_n6536__, new_new_n6537__,
    new_new_n6538__, new_new_n6539__, new_new_n6540__, new_new_n6541__,
    new_new_n6542__, new_new_n6543__, new_new_n6544__, new_new_n6545__,
    new_new_n6546__, new_new_n6547__, new_new_n6548__, new_new_n6549__,
    new_new_n6550__, new_new_n6551__, new_new_n6552__, new_new_n6553__,
    new_new_n6554__, new_new_n6555__, new_new_n6556__, new_new_n6557__,
    new_new_n6558__, new_new_n6559__, new_new_n6560__, new_new_n6561__,
    new_new_n6562__, new_new_n6563__, new_new_n6564__, new_new_n6565__,
    new_new_n6566__, new_new_n6567__, new_new_n6568__, new_new_n6569__,
    new_new_n6570__, new_new_n6571__, new_new_n6572__, new_new_n6573__,
    new_new_n6574__, new_new_n6575__, new_new_n6576__, new_new_n6577__,
    new_new_n6578__, new_new_n6579__, new_new_n6580__, new_new_n6581__,
    new_new_n6582__, new_new_n6583__, new_new_n6584__, new_new_n6585__,
    new_new_n6586__, new_new_n6587__, new_new_n6588__, new_new_n6589__,
    new_new_n6590__, new_new_n6591__, new_new_n6592__, new_new_n6593__,
    new_new_n6594__, new_new_n6595__, new_new_n6596__, new_new_n6597__,
    new_new_n6598__, new_new_n6599__, new_new_n6600__, new_new_n6601__,
    new_new_n6602__, new_new_n6603__, new_new_n6604__, new_new_n6605__,
    new_new_n6606__, new_new_n6607__, new_new_n6608__, new_new_n6609__,
    new_new_n6611__, new_new_n6612__, new_new_n6613__, new_new_n6614__,
    new_new_n6615__, new_new_n6616__, new_new_n6617__, new_new_n6618__,
    new_new_n6619__, new_new_n6620__, new_new_n6621__, new_new_n6622__,
    new_new_n6623__, new_new_n6624__, new_new_n6625__, new_new_n6626__,
    new_new_n6627__, new_new_n6628__, new_new_n6629__, new_new_n6630__,
    new_new_n6631__, new_new_n6632__, new_new_n6633__, new_new_n6634__,
    new_new_n6635__, new_new_n6636__, new_new_n6637__, new_new_n6638__,
    new_new_n6639__, new_new_n6640__, new_new_n6641__, new_new_n6642__,
    new_new_n6643__, new_new_n6644__, new_new_n6645__, new_new_n6646__,
    new_new_n6647__, new_new_n6648__, new_new_n6649__, new_new_n6650__,
    new_new_n6651__, new_new_n6652__, new_new_n6653__, new_new_n6654__,
    new_new_n6655__, new_new_n6656__, new_new_n6657__, new_new_n6658__,
    new_new_n6659__, new_new_n6660__, new_new_n6661__, new_new_n6662__,
    new_new_n6663__, new_new_n6664__, new_new_n6665__, new_new_n6666__,
    new_new_n6667__, new_new_n6668__, new_new_n6669__, new_new_n6670__,
    new_new_n6671__, new_new_n6672__, new_new_n6673__, new_new_n6674__,
    new_new_n6675__, new_new_n6676__, new_new_n6677__, new_new_n6678__,
    new_new_n6679__, new_new_n6680__, new_new_n6681__, new_new_n6682__,
    new_new_n6683__, new_new_n6684__, new_new_n6685__, new_new_n6686__,
    new_new_n6687__, new_new_n6688__, new_new_n6689__, new_new_n6690__,
    new_new_n6691__, new_new_n6692__, new_new_n6693__, new_new_n6694__,
    new_new_n6695__, new_new_n6696__, new_new_n6697__, new_new_n6698__,
    new_new_n6699__, new_new_n6700__, new_new_n6701__, new_new_n6702__,
    new_new_n6703__, new_new_n6704__, new_new_n6705__, new_new_n6706__,
    new_new_n6707__, new_new_n6708__, new_new_n6709__, new_new_n6710__,
    new_new_n6711__, new_new_n6712__, new_new_n6713__, new_new_n6714__,
    new_new_n6716__, new_new_n6717__, new_new_n6718__, new_new_n6719__,
    new_new_n6720__, new_new_n6721__, new_new_n6722__, new_new_n6723__,
    new_new_n6724__, new_new_n6725__, new_new_n6726__, new_new_n6727__,
    new_new_n6728__, new_new_n6729__, new_new_n6730__, new_new_n6731__,
    new_new_n6732__, new_new_n6733__, new_new_n6734__, new_new_n6735__,
    new_new_n6736__, new_new_n6737__, new_new_n6738__, new_new_n6739__,
    new_new_n6740__, new_new_n6741__, new_new_n6742__, new_new_n6743__,
    new_new_n6744__, new_new_n6745__, new_new_n6746__, new_new_n6747__,
    new_new_n6748__, new_new_n6749__, new_new_n6750__, new_new_n6751__,
    new_new_n6752__, new_new_n6753__, new_new_n6754__, new_new_n6755__,
    new_new_n6756__, new_new_n6757__, new_new_n6758__, new_new_n6759__,
    new_new_n6760__, new_new_n6761__, new_new_n6762__, new_new_n6763__,
    new_new_n6764__, new_new_n6765__, new_new_n6766__, new_new_n6767__,
    new_new_n6768__, new_new_n6769__, new_new_n6770__, new_new_n6771__,
    new_new_n6772__, new_new_n6773__, new_new_n6774__, new_new_n6775__,
    new_new_n6776__, new_new_n6777__, new_new_n6778__, new_new_n6779__,
    new_new_n6780__, new_new_n6781__, new_new_n6783__, new_new_n6784__,
    new_new_n6785__, new_new_n6786__, new_new_n6787__, new_new_n6788__,
    new_new_n6789__, new_new_n6790__, new_new_n6791__, new_new_n6792__,
    new_new_n6793__, new_new_n6794__, new_new_n6795__, new_new_n6796__,
    new_new_n6797__, new_new_n6798__, new_new_n6799__, new_new_n6800__,
    new_new_n6801__, new_new_n6802__, new_new_n6803__, new_new_n6804__,
    new_new_n6805__, new_new_n6806__, new_new_n6807__, new_new_n6808__,
    new_new_n6809__, new_new_n6810__, new_new_n6811__, new_new_n6812__,
    new_new_n6813__, new_new_n6814__, new_new_n6815__, new_new_n6816__,
    new_new_n6817__, new_new_n6818__, new_new_n6819__, new_new_n6820__,
    new_new_n6821__, new_new_n6822__, new_new_n6823__, new_new_n6824__,
    new_new_n6825__, new_new_n6826__, new_new_n6827__, new_new_n6828__,
    new_new_n6829__, new_new_n6830__, new_new_n6831__, new_new_n6832__,
    new_new_n6833__, new_new_n6834__, new_new_n6835__, new_new_n6836__,
    new_new_n6837__, new_new_n6838__, new_new_n6839__, new_new_n6840__,
    new_new_n6841__, new_new_n6842__, new_new_n6843__, new_new_n6844__,
    new_new_n6845__, new_new_n6846__, new_new_n6847__, new_new_n6848__,
    new_new_n6849__, new_new_n6850__, new_new_n6851__, new_new_n6852__,
    new_new_n6853__, new_new_n6854__, new_new_n6855__, new_new_n6856__,
    new_new_n6857__, new_new_n6858__, new_new_n6859__, new_new_n6860__,
    new_new_n6861__, new_new_n6862__, new_new_n6863__, new_new_n6864__,
    new_new_n6866__, new_new_n6867__, new_new_n6868__, new_new_n6869__,
    new_new_n6870__, new_new_n6871__, new_new_n6872__, new_new_n6873__,
    new_new_n6874__, new_new_n6875__, new_new_n6876__, new_new_n6877__,
    new_new_n6878__, new_new_n6879__, new_new_n6880__, new_new_n6881__,
    new_new_n6882__, new_new_n6883__, new_new_n6884__, new_new_n6885__,
    new_new_n6886__, new_new_n6887__, new_new_n6888__, new_new_n6889__,
    new_new_n6890__, new_new_n6891__, new_new_n6892__, new_new_n6893__,
    new_new_n6894__, new_new_n6895__, new_new_n6896__, new_new_n6897__,
    new_new_n6898__, new_new_n6899__, new_new_n6900__, new_new_n6901__,
    new_new_n6902__, new_new_n6903__, new_new_n6904__, new_new_n6905__,
    new_new_n6906__, new_new_n6907__, new_new_n6908__, new_new_n6909__,
    new_new_n6910__, new_new_n6911__, new_new_n6912__, new_new_n6913__,
    new_new_n6914__, new_new_n6915__, new_new_n6916__, new_new_n6917__,
    new_new_n6918__, new_new_n6919__, new_new_n6920__, new_new_n6922__,
    new_new_n6923__, new_new_n6924__, new_new_n6925__, new_new_n6926__,
    new_new_n6927__, new_new_n6928__, new_new_n6929__, new_new_n6930__,
    new_new_n6931__, new_new_n6932__, new_new_n6933__, new_new_n6934__,
    new_new_n6935__, new_new_n6936__, new_new_n6937__, new_new_n6938__,
    new_new_n6939__, new_new_n6940__, new_new_n6941__, new_new_n6942__,
    new_new_n6943__, new_new_n6944__, new_new_n6945__, new_new_n6946__,
    new_new_n6947__, new_new_n6949__, new_new_n6950__, new_new_n6951__,
    new_new_n6952__, new_new_n6953__, new_new_n6954__, new_new_n6955__,
    new_new_n6956__, new_new_n6957__, new_new_n6958__, new_new_n6959__,
    new_new_n6960__, new_new_n6961__, new_new_n6962__, new_new_n6963__,
    new_new_n6964__, new_new_n6965__, new_new_n6966__, new_new_n6967__,
    new_new_n6968__, new_new_n6969__, new_new_n6970__, new_new_n6971__,
    new_new_n6972__, new_new_n6973__, new_new_n6974__, new_new_n6975__,
    new_new_n6976__, new_new_n6977__, new_new_n6978__, new_new_n6979__,
    new_new_n6980__, new_new_n6981__, new_new_n6982__, new_new_n6983__,
    new_new_n6984__, new_new_n6985__, new_new_n6986__, new_new_n6988__,
    new_new_n6989__, new_new_n6990__, new_new_n6991__, new_new_n6992__,
    new_new_n6993__, new_new_n6994__, new_new_n6995__, new_new_n6996__,
    new_new_n6997__, new_new_n6998__, new_new_n6999__, new_new_n7000__,
    new_new_n7001__, new_new_n7002__, new_new_n7003__, new_new_n7004__,
    new_new_n7005__, new_new_n7006__, new_new_n7007__, new_new_n7008__,
    new_new_n7009__, new_new_n7010__, new_new_n7011__, new_new_n7013__,
    new_new_n7014__, new_new_n7015__, new_new_n7016__, new_new_n7017__,
    new_new_n7018__, new_new_n7019__, new_new_n7020__, new_new_n7021__,
    new_new_n7022__, new_new_n7023__, new_new_n7024__, new_new_n7025__,
    new_new_n7026__, new_new_n7027__, new_new_n7028__, new_new_n7029__,
    new_new_n7030__, new_new_n7031__, new_new_n7032__, new_new_n7033__,
    new_new_n7034__, new_new_n7035__, new_new_n7036__, new_new_n7037__,
    new_new_n7038__, new_new_n7040__, new_new_n7041__, new_new_n7042__,
    new_new_n7043__, new_new_n7044__, new_new_n7045__, new_new_n7046__,
    new_new_n7047__, new_new_n7048__, new_new_n7049__, new_new_n7050__,
    new_new_n7051__, new_new_n7052__, new_new_n7053__, new_new_n7054__,
    new_new_n7055__, new_new_n7056__, new_new_n7057__, new_new_n7058__,
    new_new_n7059__, new_new_n7060__, new_new_n7061__, new_new_n7063__,
    new_new_n7064__, new_new_n7065__, new_new_n7066__, new_new_n7067__,
    new_new_n7068__, new_new_n7069__, new_new_n7070__, new_new_n7071__,
    new_new_n7072__, new_new_n7073__, new_new_n7074__, new_new_n7075__,
    new_new_n7076__, new_new_n7077__, new_new_n7078__, new_new_n7080__,
    new_new_n7081__, new_new_n7082__, new_new_n7083__, new_new_n7084__,
    new_new_n7085__, new_new_n7086__, new_new_n7087__, new_new_n7088__,
    new_new_n7089__, new_new_n7091__, new_new_n7092__;
  assign new_new_n50__ = ~pi20 & ~pi21;
  assign new_new_n51__ = pi22 & new_new_n50__;
  assign new_new_n52__ = pi20 & pi21;
  assign new_new_n53__ = ~pi22 & new_new_n52__;
  assign new_new_n54__ = ~new_new_n51__ & ~new_new_n53__;
  assign new_new_n55__ = ~pi19 & ~pi22;
  assign new_new_n56__ = ~pi05 & ~pi06;
  assign new_new_n57__ = ~pi00 & ~pi01;
  assign new_new_n58__ = ~pi02 & ~pi03;
  assign new_new_n59__ = new_new_n57__ & new_new_n58__;
  assign new_new_n60__ = ~pi04 & ~pi07;
  assign new_new_n61__ = new_new_n56__ & new_new_n60__;
  assign new_new_n62__ = new_new_n59__ & new_new_n61__;
  assign new_new_n63__ = ~pi08 & ~pi09;
  assign new_new_n64__ = ~pi10 & new_new_n63__;
  assign new_new_n65__ = ~pi11 & new_new_n64__;
  assign new_new_n66__ = new_new_n62__ & new_new_n65__;
  assign new_new_n67__ = ~pi12 & ~pi13;
  assign new_new_n68__ = ~pi14 & new_new_n67__;
  assign new_new_n69__ = ~pi15 & new_new_n68__;
  assign new_new_n70__ = new_new_n66__ & new_new_n69__;
  assign new_new_n71__ = ~pi17 & pi18;
  assign new_new_n72__ = ~pi16 & new_new_n71__;
  assign new_new_n73__ = new_new_n70__ & ~new_new_n72__;
  assign new_new_n74__ = pi16 & pi17;
  assign new_new_n75__ = ~pi18 & new_new_n74__;
  assign new_new_n76__ = ~new_new_n70__ & ~new_new_n75__;
  assign new_new_n77__ = ~new_new_n73__ & ~new_new_n76__;
  assign new_new_n78__ = new_new_n55__ & new_new_n77__;
  assign new_new_n79__ = pi19 & pi22;
  assign new_new_n80__ = new_new_n72__ & new_new_n79__;
  assign new_new_n81__ = ~new_new_n78__ & ~new_new_n80__;
  assign new_new_n82__ = ~pi22 & ~new_new_n66__;
  assign new_new_n83__ = ~pi22 & ~new_new_n68__;
  assign new_new_n84__ = ~new_new_n82__ & ~new_new_n83__;
  assign new_new_n85__ = pi15 & ~new_new_n84__;
  assign new_new_n86__ = ~pi15 & new_new_n84__;
  assign new_new_n87__ = ~new_new_n85__ & ~new_new_n86__;
  assign new_new_n88__ = ~new_new_n81__ & new_new_n87__;
  assign new_new_n89__ = ~new_new_n54__ & new_new_n88__;
  assign new_new_n90__ = ~pi18 & ~pi19;
  assign new_new_n91__ = ~pi16 & ~pi17;
  assign new_new_n92__ = new_new_n90__ & new_new_n91__;
  assign new_new_n93__ = new_new_n70__ & new_new_n92__;
  assign new_new_n94__ = ~pi22 & ~new_new_n93__;
  assign new_new_n95__ = ~pi20 & pi21;
  assign new_new_n96__ = ~new_new_n94__ & new_new_n95__;
  assign new_new_n97__ = pi20 & ~pi21;
  assign new_new_n98__ = new_new_n94__ & new_new_n97__;
  assign new_new_n99__ = ~new_new_n96__ & ~new_new_n98__;
  assign new_new_n100__ = ~new_new_n87__ & ~new_new_n99__;
  assign new_new_n101__ = pi19 & ~pi22;
  assign new_new_n102__ = pi16 & ~new_new_n70__;
  assign new_new_n103__ = ~pi16 & new_new_n70__;
  assign new_new_n104__ = ~new_new_n102__ & ~new_new_n103__;
  assign new_new_n105__ = new_new_n71__ & new_new_n104__;
  assign new_new_n106__ = new_new_n101__ & new_new_n105__;
  assign new_new_n107__ = pi16 & pi22;
  assign new_new_n108__ = pi17 & new_new_n107__;
  assign new_new_n109__ = new_new_n90__ & new_new_n108__;
  assign new_new_n110__ = ~new_new_n106__ & ~new_new_n109__;
  assign new_new_n111__ = new_new_n100__ & ~new_new_n110__;
  assign new_new_n112__ = ~new_new_n89__ & ~new_new_n111__;
  assign new_new_n113__ = new_new_n55__ & new_new_n105__;
  assign new_new_n114__ = new_new_n75__ & new_new_n79__;
  assign new_new_n115__ = ~new_new_n113__ & ~new_new_n114__;
  assign new_new_n116__ = ~new_new_n54__ & new_new_n87__;
  assign new_new_n117__ = ~new_new_n115__ & new_new_n116__;
  assign new_new_n118__ = ~pi21 & ~pi22;
  assign new_new_n119__ = pi20 & ~new_new_n93__;
  assign new_new_n120__ = ~pi20 & new_new_n93__;
  assign new_new_n121__ = ~new_new_n119__ & ~new_new_n120__;
  assign new_new_n122__ = new_new_n118__ & new_new_n121__;
  assign new_new_n123__ = pi22 & new_new_n52__;
  assign new_new_n124__ = ~new_new_n122__ & ~new_new_n123__;
  assign new_new_n125__ = ~new_new_n87__ & ~new_new_n124__;
  assign new_new_n126__ = pi18 & ~pi19;
  assign new_new_n127__ = ~pi22 & new_new_n126__;
  assign new_new_n128__ = ~pi16 & pi17;
  assign new_new_n129__ = new_new_n70__ & ~new_new_n128__;
  assign new_new_n130__ = pi16 & ~pi17;
  assign new_new_n131__ = ~new_new_n70__ & ~new_new_n130__;
  assign new_new_n132__ = ~new_new_n129__ & ~new_new_n131__;
  assign new_new_n133__ = new_new_n127__ & new_new_n132__;
  assign new_new_n134__ = ~pi18 & new_new_n79__;
  assign new_new_n135__ = new_new_n128__ & new_new_n134__;
  assign new_new_n136__ = ~new_new_n133__ & ~new_new_n135__;
  assign new_new_n137__ = new_new_n125__ & ~new_new_n136__;
  assign new_new_n138__ = pi21 & ~pi22;
  assign new_new_n139__ = new_new_n121__ & new_new_n138__;
  assign new_new_n140__ = pi22 & new_new_n97__;
  assign new_new_n141__ = ~new_new_n139__ & ~new_new_n140__;
  assign new_new_n142__ = pi17 & new_new_n104__;
  assign new_new_n143__ = ~pi22 & new_new_n90__;
  assign new_new_n144__ = new_new_n142__ & new_new_n143__;
  assign new_new_n145__ = pi18 & pi19;
  assign new_new_n146__ = pi22 & new_new_n130__;
  assign new_new_n147__ = new_new_n145__ & new_new_n146__;
  assign new_new_n148__ = ~new_new_n144__ & ~new_new_n147__;
  assign new_new_n149__ = new_new_n87__ & ~new_new_n148__;
  assign new_new_n150__ = ~new_new_n141__ & new_new_n149__;
  assign new_new_n151__ = ~new_new_n137__ & ~new_new_n150__;
  assign new_new_n152__ = ~pi17 & ~pi18;
  assign new_new_n153__ = ~pi19 & new_new_n152__;
  assign new_new_n154__ = ~pi22 & ~new_new_n70__;
  assign new_new_n155__ = ~pi16 & ~new_new_n154__;
  assign new_new_n156__ = new_new_n153__ & new_new_n155__;
  assign new_new_n157__ = pi18 & new_new_n101__;
  assign new_new_n158__ = pi17 & new_new_n102__;
  assign new_new_n159__ = new_new_n157__ & new_new_n158__;
  assign new_new_n160__ = ~new_new_n156__ & ~new_new_n159__;
  assign new_new_n161__ = new_new_n125__ & ~new_new_n160__;
  assign new_new_n162__ = ~new_new_n87__ & ~new_new_n141__;
  assign new_new_n163__ = ~new_new_n160__ & new_new_n162__;
  assign new_new_n164__ = new_new_n127__ & new_new_n142__;
  assign new_new_n165__ = new_new_n130__ & new_new_n134__;
  assign new_new_n166__ = ~new_new_n164__ & ~new_new_n165__;
  assign new_new_n167__ = ~new_new_n87__ & ~new_new_n166__;
  assign new_new_n168__ = ~new_new_n141__ & new_new_n167__;
  assign new_new_n169__ = ~new_new_n163__ & ~new_new_n168__;
  assign new_new_n170__ = ~pi18 & new_new_n101__;
  assign new_new_n171__ = new_new_n132__ & new_new_n170__;
  assign new_new_n172__ = pi22 & new_new_n128__;
  assign new_new_n173__ = new_new_n126__ & new_new_n172__;
  assign new_new_n174__ = ~new_new_n171__ & ~new_new_n173__;
  assign new_new_n175__ = ~new_new_n99__ & ~new_new_n174__;
  assign new_new_n176__ = new_new_n87__ & new_new_n175__;
  assign new_new_n177__ = new_new_n108__ & new_new_n126__;
  assign new_new_n178__ = new_new_n101__ & new_new_n152__;
  assign new_new_n179__ = new_new_n104__ & new_new_n178__;
  assign new_new_n180__ = ~new_new_n177__ & ~new_new_n179__;
  assign new_new_n181__ = ~new_new_n54__ & ~new_new_n87__;
  assign new_new_n182__ = ~new_new_n100__ & ~new_new_n181__;
  assign new_new_n183__ = ~new_new_n180__ & ~new_new_n182__;
  assign new_new_n184__ = ~new_new_n54__ & ~new_new_n110__;
  assign new_new_n185__ = new_new_n87__ & new_new_n184__;
  assign new_new_n186__ = new_new_n125__ & ~new_new_n148__;
  assign new_new_n187__ = new_new_n116__ & ~new_new_n148__;
  assign new_new_n188__ = ~new_new_n136__ & new_new_n162__;
  assign new_new_n189__ = new_new_n180__ & ~new_new_n188__;
  assign new_new_n190__ = ~new_new_n125__ & ~new_new_n162__;
  assign new_new_n191__ = ~new_new_n189__ & ~new_new_n190__;
  assign new_new_n192__ = new_new_n124__ & new_new_n141__;
  assign new_new_n193__ = new_new_n87__ & ~new_new_n192__;
  assign new_new_n194__ = ~new_new_n181__ & ~new_new_n193__;
  assign new_new_n195__ = new_new_n87__ & ~new_new_n141__;
  assign new_new_n196__ = new_new_n110__ & new_new_n160__;
  assign new_new_n197__ = new_new_n195__ & ~new_new_n196__;
  assign new_new_n198__ = new_new_n115__ & ~new_new_n197__;
  assign new_new_n199__ = ~new_new_n194__ & ~new_new_n198__;
  assign new_new_n200__ = new_new_n87__ & ~new_new_n166__;
  assign new_new_n201__ = ~new_new_n99__ & new_new_n200__;
  assign new_new_n202__ = ~new_new_n191__ & ~new_new_n201__;
  assign new_new_n203__ = ~new_new_n199__ & new_new_n202__;
  assign new_new_n204__ = ~new_new_n176__ & ~new_new_n187__;
  assign new_new_n205__ = ~new_new_n183__ & new_new_n204__;
  assign new_new_n206__ = ~new_new_n185__ & ~new_new_n186__;
  assign new_new_n207__ = new_new_n205__ & new_new_n206__;
  assign new_new_n208__ = new_new_n169__ & new_new_n207__;
  assign new_new_n209__ = new_new_n203__ & new_new_n208__;
  assign new_new_n210__ = new_new_n108__ & new_new_n145__;
  assign new_new_n211__ = ~pi22 & new_new_n153__;
  assign new_new_n212__ = new_new_n104__ & new_new_n211__;
  assign new_new_n213__ = ~new_new_n210__ & ~new_new_n212__;
  assign new_new_n214__ = new_new_n148__ & new_new_n213__;
  assign new_new_n215__ = new_new_n100__ & ~new_new_n214__;
  assign new_new_n216__ = new_new_n132__ & new_new_n143__;
  assign new_new_n217__ = new_new_n145__ & new_new_n172__;
  assign new_new_n218__ = ~new_new_n216__ & ~new_new_n217__;
  assign new_new_n219__ = new_new_n116__ & ~new_new_n218__;
  assign new_new_n220__ = ~new_new_n136__ & new_new_n195__;
  assign new_new_n221__ = new_new_n166__ & new_new_n174__;
  assign new_new_n222__ = new_new_n125__ & ~new_new_n221__;
  assign new_new_n223__ = new_new_n87__ & ~new_new_n99__;
  assign new_new_n224__ = ~new_new_n180__ & new_new_n223__;
  assign new_new_n225__ = new_new_n90__ & new_new_n172__;
  assign new_new_n226__ = new_new_n132__ & new_new_n157__;
  assign new_new_n227__ = ~new_new_n225__ & ~new_new_n226__;
  assign new_new_n228__ = ~new_new_n54__ & ~new_new_n227__;
  assign new_new_n229__ = ~new_new_n87__ & new_new_n228__;
  assign new_new_n230__ = ~new_new_n219__ & ~new_new_n224__;
  assign new_new_n231__ = ~new_new_n229__ & new_new_n230__;
  assign new_new_n232__ = ~new_new_n215__ & ~new_new_n220__;
  assign new_new_n233__ = ~new_new_n222__ & new_new_n232__;
  assign new_new_n234__ = new_new_n231__ & new_new_n233__;
  assign new_new_n235__ = pi19 & new_new_n152__;
  assign new_new_n236__ = new_new_n155__ & new_new_n235__;
  assign new_new_n237__ = new_new_n127__ & new_new_n158__;
  assign new_new_n238__ = ~new_new_n236__ & ~new_new_n237__;
  assign new_new_n239__ = new_new_n181__ & ~new_new_n238__;
  assign new_new_n240__ = ~new_new_n180__ & new_new_n195__;
  assign new_new_n241__ = ~new_new_n239__ & ~new_new_n240__;
  assign new_new_n242__ = ~new_new_n87__ & ~new_new_n115__;
  assign new_new_n243__ = ~new_new_n99__ & new_new_n242__;
  assign new_new_n244__ = new_new_n87__ & ~new_new_n124__;
  assign new_new_n245__ = ~new_new_n223__ & ~new_new_n244__;
  assign new_new_n246__ = new_new_n110__ & new_new_n227__;
  assign new_new_n247__ = ~new_new_n245__ & ~new_new_n246__;
  assign new_new_n248__ = ~new_new_n174__ & new_new_n195__;
  assign new_new_n249__ = ~new_new_n87__ & ~new_new_n227__;
  assign new_new_n250__ = ~new_new_n99__ & new_new_n249__;
  assign new_new_n251__ = ~new_new_n81__ & ~new_new_n87__;
  assign new_new_n252__ = ~new_new_n99__ & new_new_n251__;
  assign new_new_n253__ = new_new_n142__ & new_new_n157__;
  assign new_new_n254__ = ~pi19 & new_new_n107__;
  assign new_new_n255__ = new_new_n152__ & new_new_n254__;
  assign new_new_n256__ = ~new_new_n253__ & ~new_new_n255__;
  assign new_new_n257__ = new_new_n162__ & ~new_new_n256__;
  assign new_new_n258__ = ~new_new_n81__ & new_new_n244__;
  assign new_new_n259__ = new_new_n223__ & ~new_new_n238__;
  assign new_new_n260__ = ~new_new_n258__ & ~new_new_n259__;
  assign new_new_n261__ = new_new_n110__ & new_new_n238__;
  assign new_new_n262__ = new_new_n125__ & ~new_new_n261__;
  assign new_new_n263__ = ~new_new_n257__ & ~new_new_n262__;
  assign new_new_n264__ = new_new_n260__ & new_new_n263__;
  assign new_new_n265__ = new_new_n180__ & new_new_n218__;
  assign new_new_n266__ = new_new_n244__ & ~new_new_n265__;
  assign new_new_n267__ = new_new_n223__ & ~new_new_n227__;
  assign new_new_n268__ = new_new_n142__ & new_new_n170__;
  assign new_new_n269__ = new_new_n71__ & new_new_n254__;
  assign new_new_n270__ = ~new_new_n268__ & ~new_new_n269__;
  assign new_new_n271__ = ~new_new_n116__ & ~new_new_n162__;
  assign new_new_n272__ = ~new_new_n270__ & ~new_new_n271__;
  assign new_new_n273__ = new_new_n87__ & ~new_new_n218__;
  assign new_new_n274__ = ~new_new_n141__ & new_new_n273__;
  assign new_new_n275__ = new_new_n136__ & new_new_n256__;
  assign new_new_n276__ = new_new_n181__ & ~new_new_n275__;
  assign new_new_n277__ = new_new_n223__ & ~new_new_n256__;
  assign new_new_n278__ = ~new_new_n110__ & new_new_n181__;
  assign new_new_n279__ = ~new_new_n277__ & ~new_new_n278__;
  assign new_new_n280__ = ~new_new_n267__ & ~new_new_n274__;
  assign new_new_n281__ = ~new_new_n276__ & new_new_n280__;
  assign new_new_n282__ = new_new_n279__ & new_new_n281__;
  assign new_new_n283__ = ~new_new_n272__ & new_new_n282__;
  assign new_new_n284__ = new_new_n264__ & ~new_new_n266__;
  assign new_new_n285__ = new_new_n283__ & new_new_n284__;
  assign new_new_n286__ = ~new_new_n117__ & ~new_new_n250__;
  assign new_new_n287__ = ~new_new_n252__ & new_new_n286__;
  assign new_new_n288__ = new_new_n112__ & ~new_new_n161__;
  assign new_new_n289__ = ~new_new_n243__ & ~new_new_n248__;
  assign new_new_n290__ = new_new_n288__ & new_new_n289__;
  assign new_new_n291__ = new_new_n151__ & new_new_n287__;
  assign new_new_n292__ = new_new_n241__ & ~new_new_n247__;
  assign new_new_n293__ = new_new_n291__ & new_new_n292__;
  assign new_new_n294__ = new_new_n290__ & new_new_n293__;
  assign new_new_n295__ = new_new_n234__ & new_new_n294__;
  assign new_new_n296__ = new_new_n285__ & new_new_n295__;
  assign new_new_n297__ = new_new_n209__ & new_new_n296__;
  assign new_new_n298__ = ~pi22 & ~new_new_n62__;
  assign new_new_n299__ = pi08 & ~new_new_n298__;
  assign new_new_n300__ = ~pi08 & new_new_n298__;
  assign new_new_n301__ = ~new_new_n299__ & ~new_new_n300__;
  assign new_new_n302__ = ~pi04 & new_new_n59__;
  assign new_new_n303__ = ~pi22 & ~new_new_n302__;
  assign new_new_n304__ = ~pi05 & ~new_new_n303__;
  assign new_new_n305__ = ~pi22 & ~new_new_n304__;
  assign new_new_n306__ = ~pi06 & ~new_new_n305__;
  assign new_new_n307__ = pi06 & new_new_n305__;
  assign new_new_n308__ = ~new_new_n306__ & ~new_new_n307__;
  assign new_new_n309__ = pi05 & new_new_n303__;
  assign new_new_n310__ = ~new_new_n304__ & ~new_new_n309__;
  assign new_new_n311__ = new_new_n308__ & new_new_n310__;
  assign new_new_n312__ = ~pi22 & ~new_new_n56__;
  assign new_new_n313__ = ~new_new_n303__ & ~new_new_n312__;
  assign new_new_n314__ = pi07 & ~new_new_n313__;
  assign new_new_n315__ = ~pi07 & new_new_n313__;
  assign new_new_n316__ = ~new_new_n314__ & ~new_new_n315__;
  assign new_new_n317__ = new_new_n311__ & ~new_new_n316__;
  assign new_new_n318__ = ~new_new_n308__ & ~new_new_n310__;
  assign new_new_n319__ = new_new_n316__ & new_new_n318__;
  assign new_new_n320__ = ~new_new_n317__ & ~new_new_n319__;
  assign new_new_n321__ = ~new_new_n110__ & new_new_n125__;
  assign new_new_n322__ = new_new_n162__ & ~new_new_n270__;
  assign new_new_n323__ = ~new_new_n87__ & new_new_n175__;
  assign new_new_n324__ = new_new_n125__ & ~new_new_n180__;
  assign new_new_n325__ = new_new_n100__ & ~new_new_n136__;
  assign new_new_n326__ = ~new_new_n252__ & ~new_new_n325__;
  assign new_new_n327__ = new_new_n87__ & ~new_new_n238__;
  assign new_new_n328__ = ~new_new_n124__ & new_new_n327__;
  assign new_new_n329__ = ~new_new_n323__ & ~new_new_n328__;
  assign new_new_n330__ = ~new_new_n322__ & new_new_n329__;
  assign new_new_n331__ = ~new_new_n324__ & new_new_n326__;
  assign new_new_n332__ = new_new_n330__ & new_new_n331__;
  assign new_new_n333__ = new_new_n166__ & new_new_n180__;
  assign new_new_n334__ = new_new_n181__ & ~new_new_n333__;
  assign new_new_n335__ = ~new_new_n148__ & new_new_n181__;
  assign new_new_n336__ = ~new_new_n141__ & ~new_new_n213__;
  assign new_new_n337__ = new_new_n87__ & new_new_n336__;
  assign new_new_n338__ = ~new_new_n335__ & ~new_new_n337__;
  assign new_new_n339__ = new_new_n162__ & ~new_new_n218__;
  assign new_new_n340__ = ~new_new_n116__ & new_new_n238__;
  assign new_new_n341__ = new_new_n174__ & ~new_new_n195__;
  assign new_new_n342__ = ~new_new_n340__ & ~new_new_n341__;
  assign new_new_n343__ = ~new_new_n100__ & ~new_new_n116__;
  assign new_new_n344__ = new_new_n77__ & new_new_n101__;
  assign new_new_n345__ = pi22 & new_new_n91__;
  assign new_new_n346__ = new_new_n126__ & new_new_n345__;
  assign new_new_n347__ = ~new_new_n344__ & ~new_new_n346__;
  assign new_new_n348__ = new_new_n116__ & ~new_new_n270__;
  assign new_new_n349__ = new_new_n347__ & ~new_new_n348__;
  assign new_new_n350__ = ~new_new_n343__ & ~new_new_n349__;
  assign new_new_n351__ = new_new_n100__ & ~new_new_n238__;
  assign new_new_n352__ = ~new_new_n321__ & ~new_new_n351__;
  assign new_new_n353__ = ~new_new_n334__ & ~new_new_n339__;
  assign new_new_n354__ = new_new_n352__ & new_new_n353__;
  assign new_new_n355__ = new_new_n338__ & ~new_new_n342__;
  assign new_new_n356__ = ~new_new_n350__ & new_new_n355__;
  assign new_new_n357__ = new_new_n332__ & new_new_n354__;
  assign new_new_n358__ = new_new_n356__ & new_new_n357__;
  assign new_new_n359__ = ~new_new_n141__ & ~new_new_n174__;
  assign new_new_n360__ = new_new_n160__ & new_new_n347__;
  assign new_new_n361__ = ~new_new_n124__ & ~new_new_n360__;
  assign new_new_n362__ = ~new_new_n359__ & ~new_new_n361__;
  assign new_new_n363__ = new_new_n87__ & ~new_new_n362__;
  assign new_new_n364__ = new_new_n160__ & ~new_new_n223__;
  assign new_new_n365__ = ~new_new_n195__ & new_new_n347__;
  assign new_new_n366__ = new_new_n270__ & new_new_n365__;
  assign new_new_n367__ = ~new_new_n364__ & ~new_new_n366__;
  assign new_new_n368__ = new_new_n180__ & new_new_n227__;
  assign new_new_n369__ = new_new_n81__ & new_new_n368__;
  assign new_new_n370__ = new_new_n195__ & ~new_new_n369__;
  assign new_new_n371__ = new_new_n115__ & new_new_n166__;
  assign new_new_n372__ = new_new_n223__ & ~new_new_n371__;
  assign new_new_n373__ = new_new_n116__ & ~new_new_n256__;
  assign new_new_n374__ = ~new_new_n188__ & ~new_new_n373__;
  assign new_new_n375__ = ~new_new_n372__ & new_new_n374__;
  assign new_new_n376__ = new_new_n162__ & ~new_new_n221__;
  assign new_new_n377__ = new_new_n125__ & ~new_new_n238__;
  assign new_new_n378__ = ~new_new_n219__ & ~new_new_n377__;
  assign new_new_n379__ = new_new_n195__ & ~new_new_n256__;
  assign new_new_n380__ = ~new_new_n239__ & ~new_new_n376__;
  assign new_new_n381__ = ~new_new_n379__ & new_new_n380__;
  assign new_new_n382__ = new_new_n378__ & new_new_n381__;
  assign new_new_n383__ = new_new_n181__ & ~new_new_n218__;
  assign new_new_n384__ = new_new_n87__ & new_new_n228__;
  assign new_new_n385__ = ~new_new_n383__ & ~new_new_n384__;
  assign new_new_n386__ = new_new_n125__ & ~new_new_n166__;
  assign new_new_n387__ = ~new_new_n370__ & new_new_n385__;
  assign new_new_n388__ = ~new_new_n386__ & new_new_n387__;
  assign new_new_n389__ = ~new_new_n367__ & new_new_n388__;
  assign new_new_n390__ = new_new_n375__ & new_new_n389__;
  assign new_new_n391__ = new_new_n382__ & new_new_n390__;
  assign new_new_n392__ = ~new_new_n54__ & ~new_new_n213__;
  assign new_new_n393__ = ~new_new_n115__ & ~new_new_n141__;
  assign new_new_n394__ = ~new_new_n392__ & ~new_new_n393__;
  assign new_new_n395__ = new_new_n87__ & ~new_new_n394__;
  assign new_new_n396__ = new_new_n54__ & new_new_n110__;
  assign new_new_n397__ = ~new_new_n162__ & ~new_new_n242__;
  assign new_new_n398__ = ~new_new_n396__ & ~new_new_n397__;
  assign new_new_n399__ = ~new_new_n180__ & new_new_n244__;
  assign new_new_n400__ = ~new_new_n224__ & ~new_new_n399__;
  assign new_new_n401__ = ~new_new_n395__ & new_new_n400__;
  assign new_new_n402__ = ~new_new_n398__ & new_new_n401__;
  assign new_new_n403__ = ~new_new_n99__ & new_new_n149__;
  assign new_new_n404__ = new_new_n100__ & ~new_new_n256__;
  assign new_new_n405__ = ~new_new_n267__ & ~new_new_n404__;
  assign new_new_n406__ = ~new_new_n403__ & new_new_n405__;
  assign new_new_n407__ = new_new_n218__ & new_new_n406__;
  assign new_new_n408__ = ~new_new_n99__ & ~new_new_n407__;
  assign new_new_n409__ = ~new_new_n136__ & new_new_n181__;
  assign new_new_n410__ = ~new_new_n81__ & new_new_n181__;
  assign new_new_n411__ = ~new_new_n409__ & ~new_new_n410__;
  assign new_new_n412__ = ~new_new_n110__ & ~new_new_n124__;
  assign new_new_n413__ = new_new_n87__ & new_new_n412__;
  assign new_new_n414__ = new_new_n160__ & new_new_n256__;
  assign new_new_n415__ = ~new_new_n116__ & ~new_new_n125__;
  assign new_new_n416__ = ~new_new_n414__ & ~new_new_n415__;
  assign new_new_n417__ = new_new_n148__ & new_new_n347__;
  assign new_new_n418__ = new_new_n162__ & ~new_new_n417__;
  assign new_new_n419__ = new_new_n411__ & ~new_new_n413__;
  assign new_new_n420__ = ~new_new_n418__ & new_new_n419__;
  assign new_new_n421__ = ~new_new_n416__ & new_new_n420__;
  assign new_new_n422__ = ~new_new_n87__ & ~new_new_n347__;
  assign new_new_n423__ = ~new_new_n124__ & new_new_n422__;
  assign new_new_n424__ = ~new_new_n185__ & ~new_new_n423__;
  assign new_new_n425__ = ~new_new_n363__ & new_new_n424__;
  assign new_new_n426__ = new_new_n402__ & new_new_n425__;
  assign new_new_n427__ = ~new_new_n408__ & new_new_n421__;
  assign new_new_n428__ = new_new_n426__ & new_new_n427__;
  assign new_new_n429__ = new_new_n358__ & new_new_n428__;
  assign new_new_n430__ = new_new_n391__ & new_new_n429__;
  assign new_new_n431__ = ~pi12 & new_new_n66__;
  assign new_new_n432__ = ~pi22 & ~new_new_n431__;
  assign new_new_n433__ = ~pi13 & ~new_new_n432__;
  assign new_new_n434__ = ~pi22 & ~new_new_n433__;
  assign new_new_n435__ = pi14 & ~new_new_n434__;
  assign new_new_n436__ = ~pi14 & new_new_n434__;
  assign new_new_n437__ = ~new_new_n435__ & ~new_new_n436__;
  assign new_new_n438__ = new_new_n81__ & new_new_n227__;
  assign new_new_n439__ = new_new_n195__ & ~new_new_n438__;
  assign new_new_n440__ = new_new_n283__ & ~new_new_n439__;
  assign new_new_n441__ = ~new_new_n149__ & ~new_new_n251__;
  assign new_new_n442__ = ~new_new_n124__ & ~new_new_n441__;
  assign new_new_n443__ = ~new_new_n166__ & new_new_n195__;
  assign new_new_n444__ = ~new_new_n442__ & ~new_new_n443__;
  assign new_new_n445__ = ~new_new_n136__ & new_new_n244__;
  assign new_new_n446__ = ~new_new_n218__ & new_new_n223__;
  assign new_new_n447__ = new_new_n116__ & ~new_new_n166__;
  assign new_new_n448__ = ~new_new_n162__ & ~new_new_n223__;
  assign new_new_n449__ = new_new_n110__ & new_new_n166__;
  assign new_new_n450__ = new_new_n448__ & new_new_n449__;
  assign new_new_n451__ = ~new_new_n110__ & new_new_n162__;
  assign new_new_n452__ = new_new_n81__ & ~new_new_n244__;
  assign new_new_n453__ = ~new_new_n451__ & new_new_n452__;
  assign new_new_n454__ = ~new_new_n450__ & ~new_new_n453__;
  assign new_new_n455__ = ~new_new_n100__ & ~new_new_n125__;
  assign new_new_n456__ = ~new_new_n99__ & ~new_new_n148__;
  assign new_new_n457__ = ~new_new_n87__ & new_new_n456__;
  assign new_new_n458__ = new_new_n227__ & ~new_new_n457__;
  assign new_new_n459__ = ~new_new_n455__ & ~new_new_n458__;
  assign new_new_n460__ = ~new_new_n383__ & ~new_new_n410__;
  assign new_new_n461__ = ~new_new_n325__ & new_new_n460__;
  assign new_new_n462__ = ~new_new_n336__ & ~new_new_n446__;
  assign new_new_n463__ = ~new_new_n447__ & new_new_n462__;
  assign new_new_n464__ = ~new_new_n445__ & new_new_n461__;
  assign new_new_n465__ = new_new_n463__ & new_new_n464__;
  assign new_new_n466__ = new_new_n444__ & new_new_n465__;
  assign new_new_n467__ = ~new_new_n454__ & ~new_new_n459__;
  assign new_new_n468__ = new_new_n466__ & new_new_n467__;
  assign new_new_n469__ = ~new_new_n99__ & new_new_n167__;
  assign new_new_n470__ = ~new_new_n403__ & ~new_new_n469__;
  assign new_new_n471__ = new_new_n195__ & ~new_new_n347__;
  assign new_new_n472__ = new_new_n87__ & ~new_new_n110__;
  assign new_new_n473__ = new_new_n148__ & ~new_new_n472__;
  assign new_new_n474__ = ~new_new_n271__ & ~new_new_n473__;
  assign new_new_n475__ = new_new_n100__ & ~new_new_n218__;
  assign new_new_n476__ = ~new_new_n474__ & ~new_new_n475__;
  assign new_new_n477__ = new_new_n87__ & ~new_new_n213__;
  assign new_new_n478__ = ~new_new_n124__ & new_new_n477__;
  assign new_new_n479__ = ~new_new_n100__ & new_new_n265__;
  assign new_new_n480__ = ~new_new_n116__ & new_new_n174__;
  assign new_new_n481__ = new_new_n270__ & new_new_n480__;
  assign new_new_n482__ = ~new_new_n479__ & ~new_new_n481__;
  assign new_new_n483__ = new_new_n227__ & new_new_n347__;
  assign new_new_n484__ = new_new_n115__ & new_new_n483__;
  assign new_new_n485__ = new_new_n244__ & ~new_new_n484__;
  assign new_new_n486__ = ~new_new_n482__ & ~new_new_n485__;
  assign new_new_n487__ = new_new_n218__ & new_new_n256__;
  assign new_new_n488__ = ~new_new_n162__ & new_new_n487__;
  assign new_new_n489__ = new_new_n180__ & ~new_new_n244__;
  assign new_new_n490__ = new_new_n160__ & new_new_n489__;
  assign new_new_n491__ = ~new_new_n488__ & ~new_new_n490__;
  assign new_new_n492__ = ~new_new_n125__ & new_new_n270__;
  assign new_new_n493__ = ~new_new_n181__ & ~new_new_n223__;
  assign new_new_n494__ = new_new_n218__ & new_new_n347__;
  assign new_new_n495__ = new_new_n493__ & new_new_n494__;
  assign new_new_n496__ = ~new_new_n492__ & ~new_new_n495__;
  assign new_new_n497__ = new_new_n115__ & new_new_n136__;
  assign new_new_n498__ = new_new_n125__ & ~new_new_n497__;
  assign new_new_n499__ = ~new_new_n321__ & ~new_new_n498__;
  assign new_new_n500__ = new_new_n486__ & ~new_new_n496__;
  assign new_new_n501__ = new_new_n499__ & new_new_n500__;
  assign new_new_n502__ = ~new_new_n491__ & new_new_n501__;
  assign new_new_n503__ = ~new_new_n188__ & ~new_new_n478__;
  assign new_new_n504__ = new_new_n241__ & new_new_n503__;
  assign new_new_n505__ = new_new_n502__ & new_new_n504__;
  assign new_new_n506__ = ~new_new_n160__ & new_new_n195__;
  assign new_new_n507__ = new_new_n162__ & ~new_new_n227__;
  assign new_new_n508__ = new_new_n125__ & ~new_new_n214__;
  assign new_new_n509__ = ~new_new_n117__ & ~new_new_n373__;
  assign new_new_n510__ = ~new_new_n201__ & new_new_n509__;
  assign new_new_n511__ = ~new_new_n471__ & ~new_new_n506__;
  assign new_new_n512__ = ~new_new_n507__ & ~new_new_n508__;
  assign new_new_n513__ = new_new_n511__ & new_new_n512__;
  assign new_new_n514__ = new_new_n260__ & new_new_n510__;
  assign new_new_n515__ = new_new_n470__ & new_new_n514__;
  assign new_new_n516__ = new_new_n476__ & new_new_n513__;
  assign new_new_n517__ = new_new_n515__ & new_new_n516__;
  assign new_new_n518__ = new_new_n440__ & new_new_n517__;
  assign new_new_n519__ = new_new_n468__ & new_new_n518__;
  assign new_new_n520__ = new_new_n505__ & new_new_n519__;
  assign new_new_n521__ = ~new_new_n437__ & new_new_n520__;
  assign new_new_n522__ = ~new_new_n116__ & new_new_n218__;
  assign new_new_n523__ = ~new_new_n489__ & ~new_new_n522__;
  assign new_new_n524__ = new_new_n141__ & ~new_new_n223__;
  assign new_new_n525__ = ~new_new_n218__ & ~new_new_n524__;
  assign new_new_n526__ = ~new_new_n322__ & ~new_new_n498__;
  assign new_new_n527__ = ~new_new_n116__ & new_new_n180__;
  assign new_new_n528__ = ~new_new_n200__ & new_new_n527__;
  assign new_new_n529__ = ~new_new_n54__ & ~new_new_n174__;
  assign new_new_n530__ = ~new_new_n174__ & ~new_new_n180__;
  assign new_new_n531__ = new_new_n124__ & ~new_new_n529__;
  assign new_new_n532__ = ~new_new_n530__ & new_new_n531__;
  assign new_new_n533__ = ~new_new_n528__ & ~new_new_n532__;
  assign new_new_n534__ = ~new_new_n186__ & ~new_new_n222__;
  assign new_new_n535__ = ~new_new_n525__ & new_new_n534__;
  assign new_new_n536__ = ~new_new_n523__ & new_new_n526__;
  assign new_new_n537__ = ~new_new_n533__ & new_new_n536__;
  assign new_new_n538__ = new_new_n535__ & new_new_n537__;
  assign new_new_n539__ = ~new_new_n192__ & ~new_new_n238__;
  assign new_new_n540__ = new_new_n88__ & ~new_new_n99__;
  assign new_new_n541__ = ~new_new_n539__ & ~new_new_n540__;
  assign new_new_n542__ = new_new_n87__ & ~new_new_n541__;
  assign new_new_n543__ = new_new_n110__ & new_new_n115__;
  assign new_new_n544__ = new_new_n347__ & new_new_n543__;
  assign new_new_n545__ = new_new_n223__ & ~new_new_n544__;
  assign new_new_n546__ = ~new_new_n174__ & new_new_n244__;
  assign new_new_n547__ = ~new_new_n337__ & ~new_new_n410__;
  assign new_new_n548__ = ~new_new_n377__ & ~new_new_n546__;
  assign new_new_n549__ = new_new_n547__ & new_new_n548__;
  assign new_new_n550__ = ~new_new_n545__ & new_new_n549__;
  assign new_new_n551__ = new_new_n115__ & new_new_n213__;
  assign new_new_n552__ = new_new_n136__ & new_new_n551__;
  assign new_new_n553__ = new_new_n244__ & ~new_new_n552__;
  assign new_new_n554__ = new_new_n110__ & new_new_n213__;
  assign new_new_n555__ = ~new_new_n110__ & new_new_n195__;
  assign new_new_n556__ = ~new_new_n116__ & ~new_new_n555__;
  assign new_new_n557__ = ~new_new_n554__ & ~new_new_n556__;
  assign new_new_n558__ = ~new_new_n124__ & ~new_new_n270__;
  assign new_new_n559__ = new_new_n181__ & ~new_new_n213__;
  assign new_new_n560__ = ~new_new_n174__ & new_new_n181__;
  assign new_new_n561__ = ~new_new_n559__ & ~new_new_n560__;
  assign new_new_n562__ = ~new_new_n384__ & new_new_n561__;
  assign new_new_n563__ = ~new_new_n558__ & new_new_n562__;
  assign new_new_n564__ = new_new_n100__ & ~new_new_n347__;
  assign new_new_n565__ = new_new_n115__ & ~new_new_n564__;
  assign new_new_n566__ = ~new_new_n182__ & ~new_new_n565__;
  assign new_new_n567__ = ~new_new_n258__ & ~new_new_n506__;
  assign new_new_n568__ = ~new_new_n566__ & new_new_n567__;
  assign new_new_n569__ = new_new_n444__ & new_new_n568__;
  assign new_new_n570__ = ~new_new_n87__ & ~new_new_n218__;
  assign new_new_n571__ = ~new_new_n124__ & new_new_n570__;
  assign new_new_n572__ = new_new_n117__ & ~new_new_n552__;
  assign new_new_n573__ = ~new_new_n229__ & ~new_new_n323__;
  assign new_new_n574__ = ~new_new_n456__ & ~new_new_n571__;
  assign new_new_n575__ = new_new_n573__ & new_new_n574__;
  assign new_new_n576__ = ~new_new_n553__ & new_new_n575__;
  assign new_new_n577__ = new_new_n563__ & ~new_new_n572__;
  assign new_new_n578__ = new_new_n576__ & new_new_n577__;
  assign new_new_n579__ = ~new_new_n557__ & new_new_n578__;
  assign new_new_n580__ = new_new_n569__ & new_new_n579__;
  assign new_new_n581__ = new_new_n81__ & new_new_n270__;
  assign new_new_n582__ = new_new_n110__ & new_new_n581__;
  assign new_new_n583__ = new_new_n100__ & ~new_new_n582__;
  assign new_new_n584__ = ~new_new_n150__ & ~new_new_n583__;
  assign new_new_n585__ = new_new_n213__ & new_new_n360__;
  assign new_new_n586__ = new_new_n162__ & ~new_new_n585__;
  assign new_new_n587__ = new_new_n110__ & new_new_n180__;
  assign new_new_n588__ = new_new_n181__ & ~new_new_n587__;
  assign new_new_n589__ = new_new_n136__ & new_new_n270__;
  assign new_new_n590__ = ~new_new_n188__ & ~new_new_n223__;
  assign new_new_n591__ = ~new_new_n589__ & ~new_new_n590__;
  assign new_new_n592__ = ~new_new_n239__ & ~new_new_n475__;
  assign new_new_n593__ = ~new_new_n591__ & new_new_n592__;
  assign new_new_n594__ = new_new_n116__ & ~new_new_n136__;
  assign new_new_n595__ = new_new_n162__ & ~new_new_n238__;
  assign new_new_n596__ = new_new_n125__ & ~new_new_n213__;
  assign new_new_n597__ = ~new_new_n168__ & ~new_new_n594__;
  assign new_new_n598__ = ~new_new_n471__ & ~new_new_n595__;
  assign new_new_n599__ = ~new_new_n596__ & new_new_n598__;
  assign new_new_n600__ = new_new_n597__ & new_new_n599__;
  assign new_new_n601__ = ~new_new_n586__ & ~new_new_n588__;
  assign new_new_n602__ = ~new_new_n542__ & new_new_n601__;
  assign new_new_n603__ = new_new_n584__ & new_new_n602__;
  assign new_new_n604__ = new_new_n550__ & new_new_n593__;
  assign new_new_n605__ = new_new_n600__ & new_new_n604__;
  assign new_new_n606__ = new_new_n538__ & new_new_n603__;
  assign new_new_n607__ = new_new_n605__ & new_new_n606__;
  assign new_new_n608__ = new_new_n580__ & new_new_n607__;
  assign new_new_n609__ = new_new_n430__ & ~new_new_n608__;
  assign new_new_n610__ = ~new_new_n521__ & new_new_n609__;
  assign new_new_n611__ = ~pi08 & new_new_n62__;
  assign new_new_n612__ = ~pi22 & ~new_new_n611__;
  assign new_new_n613__ = ~pi09 & ~new_new_n612__;
  assign new_new_n614__ = pi09 & new_new_n612__;
  assign new_new_n615__ = ~new_new_n613__ & ~new_new_n614__;
  assign new_new_n616__ = new_new_n81__ & new_new_n99__;
  assign new_new_n617__ = ~new_new_n115__ & new_new_n244__;
  assign new_new_n618__ = new_new_n616__ & ~new_new_n617__;
  assign new_new_n619__ = new_new_n100__ & ~new_new_n213__;
  assign new_new_n620__ = new_new_n124__ & new_new_n218__;
  assign new_new_n621__ = ~new_new_n619__ & new_new_n620__;
  assign new_new_n622__ = ~new_new_n618__ & ~new_new_n621__;
  assign new_new_n623__ = new_new_n124__ & new_new_n166__;
  assign new_new_n624__ = new_new_n238__ & new_new_n623__;
  assign new_new_n625__ = new_new_n99__ & new_new_n347__;
  assign new_new_n626__ = new_new_n180__ & new_new_n625__;
  assign new_new_n627__ = ~new_new_n624__ & ~new_new_n626__;
  assign new_new_n628__ = ~new_new_n546__ & ~new_new_n627__;
  assign new_new_n629__ = new_new_n81__ & new_new_n148__;
  assign new_new_n630__ = ~new_new_n87__ & ~new_new_n629__;
  assign new_new_n631__ = ~new_new_n477__ & ~new_new_n630__;
  assign new_new_n632__ = ~new_new_n99__ & ~new_new_n631__;
  assign new_new_n633__ = new_new_n223__ & ~new_new_n629__;
  assign new_new_n634__ = ~new_new_n413__ & ~new_new_n445__;
  assign new_new_n635__ = ~new_new_n633__ & new_new_n634__;
  assign new_new_n636__ = new_new_n499__ & new_new_n635__;
  assign new_new_n637__ = new_new_n628__ & ~new_new_n632__;
  assign new_new_n638__ = new_new_n636__ & new_new_n637__;
  assign new_new_n639__ = new_new_n180__ & new_new_n497__;
  assign new_new_n640__ = ~new_new_n99__ & ~new_new_n639__;
  assign new_new_n641__ = new_new_n238__ & new_new_n270__;
  assign new_new_n642__ = ~new_new_n222__ & new_new_n641__;
  assign new_new_n643__ = ~new_new_n124__ & ~new_new_n642__;
  assign new_new_n644__ = ~new_new_n176__ & ~new_new_n640__;
  assign new_new_n645__ = ~new_new_n643__ & new_new_n644__;
  assign new_new_n646__ = new_new_n124__ & ~new_new_n622__;
  assign new_new_n647__ = new_new_n645__ & new_new_n646__;
  assign new_new_n648__ = new_new_n638__ & new_new_n647__;
  assign new_new_n649__ = new_new_n615__ & ~new_new_n648__;
  assign new_new_n650__ = pi13 & new_new_n432__;
  assign new_new_n651__ = ~new_new_n433__ & ~new_new_n650__;
  assign new_new_n652__ = new_new_n166__ & ~new_new_n251__;
  assign new_new_n653__ = ~new_new_n327__ & new_new_n652__;
  assign new_new_n654__ = new_new_n497__ & new_new_n653__;
  assign new_new_n655__ = ~new_new_n54__ & ~new_new_n654__;
  assign new_new_n656__ = new_new_n110__ & new_new_n256__;
  assign new_new_n657__ = new_new_n100__ & ~new_new_n656__;
  assign new_new_n658__ = new_new_n136__ & new_new_n213__;
  assign new_new_n659__ = new_new_n195__ & ~new_new_n658__;
  assign new_new_n660__ = ~new_new_n339__ & ~new_new_n657__;
  assign new_new_n661__ = ~new_new_n659__ & new_new_n660__;
  assign new_new_n662__ = new_new_n162__ & ~new_new_n213__;
  assign new_new_n663__ = new_new_n81__ & new_new_n218__;
  assign new_new_n664__ = new_new_n87__ & ~new_new_n663__;
  assign new_new_n665__ = new_new_n115__ & new_new_n148__;
  assign new_new_n666__ = ~new_new_n664__ & new_new_n665__;
  assign new_new_n667__ = ~new_new_n141__ & ~new_new_n666__;
  assign new_new_n668__ = new_new_n246__ & new_new_n414__;
  assign new_new_n669__ = ~new_new_n99__ & ~new_new_n668__;
  assign new_new_n670__ = ~new_new_n81__ & ~new_new_n141__;
  assign new_new_n671__ = ~new_new_n87__ & new_new_n670__;
  assign new_new_n672__ = ~new_new_n323__ & ~new_new_n662__;
  assign new_new_n673__ = ~new_new_n671__ & new_new_n672__;
  assign new_new_n674__ = ~new_new_n667__ & ~new_new_n669__;
  assign new_new_n675__ = new_new_n673__ & new_new_n674__;
  assign new_new_n676__ = new_new_n661__ & new_new_n675__;
  assign new_new_n677__ = new_new_n270__ & new_new_n347__;
  assign new_new_n678__ = new_new_n100__ & ~new_new_n677__;
  assign new_new_n679__ = ~new_new_n88__ & new_new_n218__;
  assign new_new_n680__ = new_new_n214__ & new_new_n679__;
  assign new_new_n681__ = ~new_new_n54__ & ~new_new_n680__;
  assign new_new_n682__ = ~new_new_n163__ & ~new_new_n678__;
  assign new_new_n683__ = ~new_new_n681__ & new_new_n682__;
  assign new_new_n684__ = ~new_new_n367__ & new_new_n683__;
  assign new_new_n685__ = ~new_new_n655__ & new_new_n684__;
  assign new_new_n686__ = new_new_n676__ & new_new_n685__;
  assign new_new_n687__ = ~new_new_n651__ & new_new_n686__;
  assign new_new_n688__ = new_new_n651__ & ~new_new_n686__;
  assign new_new_n689__ = ~new_new_n687__ & ~new_new_n688__;
  assign new_new_n690__ = ~new_new_n160__ & new_new_n223__;
  assign new_new_n691__ = ~new_new_n87__ & ~new_new_n256__;
  assign new_new_n692__ = ~new_new_n124__ & new_new_n691__;
  assign new_new_n693__ = new_new_n238__ & ~new_new_n692__;
  assign new_new_n694__ = ~new_new_n190__ & ~new_new_n693__;
  assign new_new_n695__ = ~new_new_n87__ & new_new_n270__;
  assign new_new_n696__ = new_new_n87__ & new_new_n180__;
  assign new_new_n697__ = new_new_n160__ & new_new_n696__;
  assign new_new_n698__ = ~new_new_n124__ & ~new_new_n697__;
  assign new_new_n699__ = ~new_new_n443__ & ~new_new_n698__;
  assign new_new_n700__ = ~new_new_n695__ & ~new_new_n699__;
  assign new_new_n701__ = ~new_new_n347__ & ~new_new_n493__;
  assign new_new_n702__ = ~new_new_n348__ & ~new_new_n690__;
  assign new_new_n703__ = new_new_n112__ & new_new_n702__;
  assign new_new_n704__ = ~new_new_n701__ & new_new_n703__;
  assign new_new_n705__ = ~new_new_n694__ & new_new_n704__;
  assign new_new_n706__ = ~new_new_n700__ & new_new_n705__;
  assign new_new_n707__ = new_new_n505__ & new_new_n706__;
  assign new_new_n708__ = ~new_new_n168__ & ~new_new_n258__;
  assign new_new_n709__ = ~new_new_n124__ & new_new_n149__;
  assign new_new_n710__ = ~new_new_n248__ & ~new_new_n267__;
  assign new_new_n711__ = ~new_new_n596__ & ~new_new_n709__;
  assign new_new_n712__ = new_new_n710__ & new_new_n711__;
  assign new_new_n713__ = new_new_n708__ & new_new_n712__;
  assign new_new_n714__ = ~new_new_n124__ & ~new_new_n166__;
  assign new_new_n715__ = new_new_n174__ & ~new_new_n714__;
  assign new_new_n716__ = new_new_n124__ & ~new_new_n181__;
  assign new_new_n717__ = ~new_new_n162__ & new_new_n716__;
  assign new_new_n718__ = ~new_new_n715__ & ~new_new_n717__;
  assign new_new_n719__ = new_new_n160__ & new_new_n238__;
  assign new_new_n720__ = ~new_new_n116__ & new_new_n719__;
  assign new_new_n721__ = ~new_new_n365__ & ~new_new_n720__;
  assign new_new_n722__ = ~new_new_n383__ & ~new_new_n718__;
  assign new_new_n723__ = ~new_new_n721__ & new_new_n722__;
  assign new_new_n724__ = new_new_n81__ & ~new_new_n100__;
  assign new_new_n725__ = ~new_new_n125__ & new_new_n160__;
  assign new_new_n726__ = ~new_new_n724__ & ~new_new_n725__;
  assign new_new_n727__ = ~new_new_n335__ & ~new_new_n726__;
  assign new_new_n728__ = ~new_new_n161__ & ~new_new_n619__;
  assign new_new_n729__ = ~new_new_n187__ & ~new_new_n328__;
  assign new_new_n730__ = ~new_new_n180__ & new_new_n181__;
  assign new_new_n731__ = ~new_new_n186__ & ~new_new_n413__;
  assign new_new_n732__ = new_new_n244__ & ~new_new_n589__;
  assign new_new_n733__ = new_new_n227__ & ~new_new_n404__;
  assign new_new_n734__ = ~new_new_n455__ & ~new_new_n733__;
  assign new_new_n735__ = new_new_n54__ & new_new_n99__;
  assign new_new_n736__ = new_new_n87__ & ~new_new_n735__;
  assign new_new_n737__ = new_new_n213__ & ~new_new_n529__;
  assign new_new_n738__ = new_new_n736__ & ~new_new_n737__;
  assign new_new_n739__ = ~new_new_n732__ & ~new_new_n738__;
  assign new_new_n740__ = ~new_new_n734__ & new_new_n739__;
  assign new_new_n741__ = ~new_new_n277__ & new_new_n731__;
  assign new_new_n742__ = new_new_n740__ & new_new_n741__;
  assign new_new_n743__ = new_new_n87__ & ~new_new_n270__;
  assign new_new_n744__ = ~new_new_n141__ & new_new_n743__;
  assign new_new_n745__ = ~new_new_n99__ & new_new_n472__;
  assign new_new_n746__ = ~new_new_n744__ & ~new_new_n745__;
  assign new_new_n747__ = ~new_new_n559__ & ~new_new_n730__;
  assign new_new_n748__ = ~new_new_n564__ & new_new_n747__;
  assign new_new_n749__ = ~new_new_n324__ & new_new_n748__;
  assign new_new_n750__ = new_new_n729__ & new_new_n749__;
  assign new_new_n751__ = new_new_n728__ & new_new_n746__;
  assign new_new_n752__ = new_new_n750__ & new_new_n751__;
  assign new_new_n753__ = new_new_n727__ & new_new_n752__;
  assign new_new_n754__ = new_new_n713__ & new_new_n723__;
  assign new_new_n755__ = new_new_n742__ & new_new_n754__;
  assign new_new_n756__ = new_new_n753__ & new_new_n755__;
  assign new_new_n757__ = new_new_n707__ & new_new_n756__;
  assign new_new_n758__ = ~new_new_n608__ & ~new_new_n757__;
  assign new_new_n759__ = new_new_n608__ & new_new_n757__;
  assign new_new_n760__ = ~new_new_n758__ & ~new_new_n759__;
  assign new_new_n761__ = new_new_n689__ & new_new_n760__;
  assign new_new_n762__ = ~pi12 & ~new_new_n82__;
  assign new_new_n763__ = pi12 & new_new_n82__;
  assign new_new_n764__ = ~new_new_n762__ & ~new_new_n763__;
  assign new_new_n765__ = ~new_new_n608__ & ~new_new_n764__;
  assign new_new_n766__ = new_new_n608__ & new_new_n764__;
  assign new_new_n767__ = ~new_new_n765__ & ~new_new_n766__;
  assign new_new_n768__ = ~new_new_n686__ & ~new_new_n764__;
  assign new_new_n769__ = new_new_n686__ & new_new_n764__;
  assign new_new_n770__ = ~new_new_n768__ & ~new_new_n769__;
  assign new_new_n771__ = ~new_new_n760__ & ~new_new_n770__;
  assign new_new_n772__ = new_new_n767__ & new_new_n771__;
  assign new_new_n773__ = ~new_new_n761__ & ~new_new_n772__;
  assign new_new_n774__ = ~new_new_n649__ & ~new_new_n773__;
  assign new_new_n775__ = new_new_n649__ & new_new_n773__;
  assign new_new_n776__ = ~new_new_n774__ & ~new_new_n775__;
  assign new_new_n777__ = ~new_new_n520__ & ~new_new_n608__;
  assign new_new_n778__ = ~new_new_n437__ & ~new_new_n520__;
  assign new_new_n779__ = new_new_n608__ & ~new_new_n778__;
  assign new_new_n780__ = ~new_new_n430__ & ~new_new_n777__;
  assign new_new_n781__ = ~new_new_n779__ & new_new_n780__;
  assign new_new_n782__ = ~new_new_n610__ & ~new_new_n781__;
  assign new_new_n783__ = ~new_new_n776__ & new_new_n782__;
  assign new_new_n784__ = ~new_new_n430__ & ~new_new_n520__;
  assign new_new_n785__ = ~new_new_n608__ & ~new_new_n784__;
  assign new_new_n786__ = ~new_new_n521__ & new_new_n785__;
  assign new_new_n787__ = ~new_new_n781__ & ~new_new_n786__;
  assign new_new_n788__ = new_new_n776__ & ~new_new_n787__;
  assign new_new_n789__ = ~new_new_n783__ & ~new_new_n788__;
  assign new_new_n790__ = ~new_new_n99__ & ~new_new_n677__;
  assign new_new_n791__ = new_new_n676__ & ~new_new_n790__;
  assign new_new_n792__ = new_new_n648__ & new_new_n791__;
  assign new_new_n793__ = new_new_n246__ & new_new_n347__;
  assign new_new_n794__ = new_new_n256__ & new_new_n793__;
  assign new_new_n795__ = ~new_new_n141__ & ~new_new_n794__;
  assign new_new_n796__ = ~new_new_n322__ & ~new_new_n795__;
  assign new_new_n797__ = new_new_n174__ & new_new_n238__;
  assign new_new_n798__ = new_new_n166__ & new_new_n797__;
  assign new_new_n799__ = ~new_new_n87__ & ~new_new_n136__;
  assign new_new_n800__ = new_new_n180__ & ~new_new_n799__;
  assign new_new_n801__ = ~new_new_n743__ & new_new_n800__;
  assign new_new_n802__ = new_new_n798__ & new_new_n801__;
  assign new_new_n803__ = ~new_new_n141__ & ~new_new_n802__;
  assign new_new_n804__ = new_new_n796__ & ~new_new_n803__;
  assign new_new_n805__ = new_new_n686__ & new_new_n804__;
  assign new_new_n806__ = ~pi22 & ~new_new_n64__;
  assign new_new_n807__ = ~new_new_n298__ & ~new_new_n806__;
  assign new_new_n808__ = pi11 & ~new_new_n807__;
  assign new_new_n809__ = ~pi11 & new_new_n807__;
  assign new_new_n810__ = ~new_new_n808__ & ~new_new_n809__;
  assign new_new_n811__ = ~new_new_n805__ & new_new_n810__;
  assign new_new_n812__ = new_new_n792__ & ~new_new_n811__;
  assign new_new_n813__ = ~pi22 & ~new_new_n613__;
  assign new_new_n814__ = pi10 & ~new_new_n813__;
  assign new_new_n815__ = ~pi10 & new_new_n813__;
  assign new_new_n816__ = ~new_new_n814__ & ~new_new_n815__;
  assign new_new_n817__ = new_new_n791__ & new_new_n816__;
  assign new_new_n818__ = ~new_new_n805__ & ~new_new_n816__;
  assign new_new_n819__ = ~new_new_n817__ & ~new_new_n818__;
  assign new_new_n820__ = ~new_new_n812__ & ~new_new_n819__;
  assign new_new_n821__ = new_new_n437__ & new_new_n608__;
  assign new_new_n822__ = ~new_new_n437__ & ~new_new_n608__;
  assign new_new_n823__ = new_new_n430__ & new_new_n520__;
  assign new_new_n824__ = ~new_new_n784__ & ~new_new_n823__;
  assign new_new_n825__ = ~new_new_n821__ & ~new_new_n822__;
  assign new_new_n826__ = new_new_n824__ & new_new_n825__;
  assign new_new_n827__ = new_new_n608__ & ~new_new_n651__;
  assign new_new_n828__ = ~new_new_n608__ & new_new_n651__;
  assign new_new_n829__ = ~new_new_n827__ & ~new_new_n828__;
  assign new_new_n830__ = ~new_new_n430__ & new_new_n651__;
  assign new_new_n831__ = new_new_n430__ & ~new_new_n651__;
  assign new_new_n832__ = ~new_new_n830__ & ~new_new_n831__;
  assign new_new_n833__ = ~new_new_n824__ & new_new_n829__;
  assign new_new_n834__ = ~new_new_n832__ & new_new_n833__;
  assign new_new_n835__ = ~new_new_n826__ & ~new_new_n834__;
  assign new_new_n836__ = new_new_n760__ & ~new_new_n770__;
  assign new_new_n837__ = new_new_n608__ & new_new_n810__;
  assign new_new_n838__ = ~new_new_n608__ & ~new_new_n810__;
  assign new_new_n839__ = ~new_new_n837__ & ~new_new_n838__;
  assign new_new_n840__ = new_new_n686__ & new_new_n810__;
  assign new_new_n841__ = ~new_new_n686__ & ~new_new_n810__;
  assign new_new_n842__ = ~new_new_n840__ & ~new_new_n841__;
  assign new_new_n843__ = ~new_new_n760__ & ~new_new_n842__;
  assign new_new_n844__ = new_new_n839__ & new_new_n843__;
  assign new_new_n845__ = ~new_new_n836__ & ~new_new_n844__;
  assign new_new_n846__ = new_new_n835__ & new_new_n845__;
  assign new_new_n847__ = ~new_new_n835__ & ~new_new_n845__;
  assign new_new_n848__ = ~new_new_n615__ & ~new_new_n791__;
  assign new_new_n849__ = ~new_new_n805__ & ~new_new_n817__;
  assign new_new_n850__ = ~new_new_n848__ & new_new_n849__;
  assign new_new_n851__ = new_new_n648__ & ~new_new_n850__;
  assign new_new_n852__ = new_new_n615__ & new_new_n805__;
  assign new_new_n853__ = ~new_new_n851__ & ~new_new_n852__;
  assign new_new_n854__ = ~new_new_n847__ & ~new_new_n853__;
  assign new_new_n855__ = ~new_new_n846__ & ~new_new_n854__;
  assign new_new_n856__ = ~new_new_n820__ & ~new_new_n855__;
  assign new_new_n857__ = new_new_n820__ & new_new_n855__;
  assign new_new_n858__ = ~new_new_n856__ & ~new_new_n857__;
  assign new_new_n859__ = ~new_new_n248__ & ~new_new_n671__;
  assign new_new_n860__ = new_new_n162__ & ~new_new_n261__;
  assign new_new_n861__ = ~new_new_n227__ & new_new_n244__;
  assign new_new_n862__ = ~new_new_n176__ & ~new_new_n571__;
  assign new_new_n863__ = new_new_n244__ & ~new_new_n270__;
  assign new_new_n864__ = ~new_new_n224__ & ~new_new_n863__;
  assign new_new_n865__ = ~new_new_n337__ & ~new_new_n619__;
  assign new_new_n866__ = ~new_new_n860__ & ~new_new_n861__;
  assign new_new_n867__ = new_new_n862__ & new_new_n866__;
  assign new_new_n868__ = new_new_n864__ & new_new_n865__;
  assign new_new_n869__ = new_new_n867__ & new_new_n868__;
  assign new_new_n870__ = ~new_new_n148__ & new_new_n162__;
  assign new_new_n871__ = ~new_new_n690__ & ~new_new_n870__;
  assign new_new_n872__ = ~new_new_n186__ & ~new_new_n339__;
  assign new_new_n873__ = ~new_new_n117__ & ~new_new_n730__;
  assign new_new_n874__ = ~new_new_n384__ & new_new_n873__;
  assign new_new_n875__ = new_new_n871__ & new_new_n874__;
  assign new_new_n876__ = new_new_n872__ & new_new_n875__;
  assign new_new_n877__ = new_new_n116__ & ~new_new_n160__;
  assign new_new_n878__ = ~new_new_n410__ & ~new_new_n877__;
  assign new_new_n879__ = ~new_new_n325__ & new_new_n878__;
  assign new_new_n880__ = ~new_new_n243__ & new_new_n879__;
  assign new_new_n881__ = ~new_new_n692__ & new_new_n880__;
  assign new_new_n882__ = new_new_n125__ & ~new_new_n551__;
  assign new_new_n883__ = new_new_n54__ & new_new_n141__;
  assign new_new_n884__ = new_new_n87__ & ~new_new_n180__;
  assign new_new_n885__ = ~new_new_n883__ & new_new_n884__;
  assign new_new_n886__ = ~new_new_n379__ & ~new_new_n540__;
  assign new_new_n887__ = ~new_new_n882__ & ~new_new_n885__;
  assign new_new_n888__ = new_new_n886__ & new_new_n887__;
  assign new_new_n889__ = new_new_n859__ & new_new_n888__;
  assign new_new_n890__ = new_new_n881__ & new_new_n889__;
  assign new_new_n891__ = new_new_n869__ & new_new_n876__;
  assign new_new_n892__ = new_new_n890__ & new_new_n891__;
  assign new_new_n893__ = ~new_new_n115__ & new_new_n162__;
  assign new_new_n894__ = ~new_new_n478__ & ~new_new_n893__;
  assign new_new_n895__ = new_new_n87__ & new_new_n218__;
  assign new_new_n896__ = ~new_new_n54__ & ~new_new_n256__;
  assign new_new_n897__ = ~new_new_n116__ & ~new_new_n896__;
  assign new_new_n898__ = ~new_new_n895__ & ~new_new_n897__;
  assign new_new_n899__ = new_new_n894__ & ~new_new_n898__;
  assign new_new_n900__ = new_new_n136__ & new_new_n218__;
  assign new_new_n901__ = ~new_new_n244__ & new_new_n900__;
  assign new_new_n902__ = ~new_new_n364__ & ~new_new_n901__;
  assign new_new_n903__ = new_new_n81__ & new_new_n256__;
  assign new_new_n904__ = ~new_new_n100__ & new_new_n903__;
  assign new_new_n905__ = new_new_n81__ & ~new_new_n116__;
  assign new_new_n906__ = new_new_n347__ & new_new_n905__;
  assign new_new_n907__ = ~new_new_n343__ & ~new_new_n906__;
  assign new_new_n908__ = ~new_new_n904__ & new_new_n907__;
  assign new_new_n909__ = ~new_new_n902__ & ~new_new_n908__;
  assign new_new_n910__ = new_new_n115__ & new_new_n347__;
  assign new_new_n911__ = new_new_n223__ & ~new_new_n910__;
  assign new_new_n912__ = new_new_n227__ & ~new_new_n911__;
  assign new_new_n913__ = ~new_new_n493__ & ~new_new_n912__;
  assign new_new_n914__ = ~new_new_n160__ & new_new_n181__;
  assign new_new_n915__ = ~new_new_n201__ & ~new_new_n914__;
  assign new_new_n916__ = new_new_n244__ & ~new_new_n494__;
  assign new_new_n917__ = ~new_new_n239__ & ~new_new_n916__;
  assign new_new_n918__ = ~new_new_n99__ & new_new_n477__;
  assign new_new_n919__ = ~new_new_n546__ & ~new_new_n918__;
  assign new_new_n920__ = ~new_new_n54__ & new_new_n327__;
  assign new_new_n921__ = ~new_new_n166__ & new_new_n181__;
  assign new_new_n922__ = ~new_new_n250__ & ~new_new_n920__;
  assign new_new_n923__ = ~new_new_n921__ & new_new_n922__;
  assign new_new_n924__ = ~new_new_n662__ & new_new_n923__;
  assign new_new_n925__ = new_new_n100__ & ~new_new_n180__;
  assign new_new_n926__ = new_new_n166__ & ~new_new_n925__;
  assign new_new_n927__ = ~new_new_n100__ & new_new_n190__;
  assign new_new_n928__ = ~new_new_n926__ & ~new_new_n927__;
  assign new_new_n929__ = new_new_n54__ & ~new_new_n195__;
  assign new_new_n930__ = ~new_new_n554__ & ~new_new_n929__;
  assign new_new_n931__ = new_new_n238__ & ~new_new_n244__;
  assign new_new_n932__ = ~new_new_n188__ & new_new_n931__;
  assign new_new_n933__ = new_new_n99__ & new_new_n136__;
  assign new_new_n934__ = new_new_n180__ & new_new_n933__;
  assign new_new_n935__ = ~new_new_n932__ & ~new_new_n934__;
  assign new_new_n936__ = ~new_new_n322__ & ~new_new_n413__;
  assign new_new_n937__ = ~new_new_n709__ & new_new_n936__;
  assign new_new_n938__ = ~new_new_n930__ & new_new_n937__;
  assign new_new_n939__ = new_new_n924__ & ~new_new_n928__;
  assign new_new_n940__ = ~new_new_n935__ & new_new_n939__;
  assign new_new_n941__ = new_new_n938__ & new_new_n940__;
  assign new_new_n942__ = ~new_new_n257__ & ~new_new_n471__;
  assign new_new_n943__ = new_new_n915__ & new_new_n942__;
  assign new_new_n944__ = new_new_n917__ & new_new_n919__;
  assign new_new_n945__ = new_new_n943__ & new_new_n944__;
  assign new_new_n946__ = new_new_n899__ & new_new_n909__;
  assign new_new_n947__ = ~new_new_n913__ & new_new_n946__;
  assign new_new_n948__ = new_new_n945__ & new_new_n947__;
  assign new_new_n949__ = new_new_n892__ & new_new_n948__;
  assign new_new_n950__ = new_new_n941__ & new_new_n949__;
  assign new_new_n951__ = new_new_n223__ & ~new_new_n347__;
  assign new_new_n952__ = new_new_n141__ & new_new_n735__;
  assign new_new_n953__ = new_new_n242__ & ~new_new_n952__;
  assign new_new_n954__ = ~new_new_n248__ & ~new_new_n951__;
  assign new_new_n955__ = ~new_new_n953__ & new_new_n954__;
  assign new_new_n956__ = ~new_new_n54__ & ~new_new_n136__;
  assign new_new_n957__ = new_new_n87__ & new_new_n392__;
  assign new_new_n958__ = ~new_new_n690__ & ~new_new_n925__;
  assign new_new_n959__ = ~new_new_n351__ & ~new_new_n956__;
  assign new_new_n960__ = ~new_new_n446__ & ~new_new_n957__;
  assign new_new_n961__ = new_new_n959__ & new_new_n960__;
  assign new_new_n962__ = ~new_new_n186__ & ~new_new_n451__;
  assign new_new_n963__ = new_new_n958__ & new_new_n962__;
  assign new_new_n964__ = new_new_n961__ & new_new_n963__;
  assign new_new_n965__ = new_new_n213__ & new_new_n663__;
  assign new_new_n966__ = new_new_n125__ & ~new_new_n965__;
  assign new_new_n967__ = ~new_new_n150__ & ~new_new_n966__;
  assign new_new_n968__ = ~new_new_n709__ & new_new_n967__;
  assign new_new_n969__ = ~new_new_n447__ & ~new_new_n475__;
  assign new_new_n970__ = new_new_n256__ & new_new_n347__;
  assign new_new_n971__ = new_new_n125__ & ~new_new_n970__;
  assign new_new_n972__ = new_new_n213__ & new_new_n238__;
  assign new_new_n973__ = new_new_n244__ & ~new_new_n972__;
  assign new_new_n974__ = ~new_new_n457__ & ~new_new_n971__;
  assign new_new_n975__ = ~new_new_n973__ & new_new_n974__;
  assign new_new_n976__ = ~new_new_n124__ & new_new_n249__;
  assign new_new_n977__ = ~new_new_n404__ & ~new_new_n976__;
  assign new_new_n978__ = ~new_new_n506__ & new_new_n977__;
  assign new_new_n979__ = ~new_new_n870__ & new_new_n969__;
  assign new_new_n980__ = new_new_n978__ & new_new_n979__;
  assign new_new_n981__ = new_new_n919__ & new_new_n980__;
  assign new_new_n982__ = new_new_n968__ & new_new_n975__;
  assign new_new_n983__ = new_new_n981__ & new_new_n982__;
  assign new_new_n984__ = ~new_new_n239__ & ~new_new_n730__;
  assign new_new_n985__ = ~new_new_n258__ & new_new_n984__;
  assign new_new_n986__ = ~new_new_n377__ & new_new_n985__;
  assign new_new_n987__ = new_new_n924__ & new_new_n986__;
  assign new_new_n988__ = new_new_n983__ & new_new_n987__;
  assign new_new_n989__ = ~new_new_n124__ & new_new_n273__;
  assign new_new_n990__ = new_new_n180__ & new_new_n347__;
  assign new_new_n991__ = new_new_n162__ & ~new_new_n990__;
  assign new_new_n992__ = new_new_n166__ & new_new_n543__;
  assign new_new_n993__ = ~new_new_n99__ & ~new_new_n110__;
  assign new_new_n994__ = new_new_n141__ & ~new_new_n993__;
  assign new_new_n995__ = new_new_n87__ & ~new_new_n992__;
  assign new_new_n996__ = ~new_new_n994__ & new_new_n995__;
  assign new_new_n997__ = new_new_n326__ & ~new_new_n989__;
  assign new_new_n998__ = ~new_new_n991__ & new_new_n997__;
  assign new_new_n999__ = ~new_new_n996__ & new_new_n998__;
  assign new_new_n1000__ = ~new_new_n222__ & ~new_new_n559__;
  assign new_new_n1001__ = ~new_new_n469__ & new_new_n1000__;
  assign new_new_n1002__ = new_new_n169__ & new_new_n486__;
  assign new_new_n1003__ = new_new_n1001__ & new_new_n1002__;
  assign new_new_n1004__ = new_new_n955__ & new_new_n1003__;
  assign new_new_n1005__ = new_new_n964__ & new_new_n999__;
  assign new_new_n1006__ = new_new_n1004__ & new_new_n1005__;
  assign new_new_n1007__ = new_new_n988__ & new_new_n1006__;
  assign new_new_n1008__ = ~new_new_n950__ & ~new_new_n1007__;
  assign new_new_n1009__ = ~new_new_n430__ & ~new_new_n1008__;
  assign new_new_n1010__ = new_new_n301__ & new_new_n1009__;
  assign new_new_n1011__ = ~new_new_n301__ & ~new_new_n1009__;
  assign new_new_n1012__ = ~new_new_n316__ & ~new_new_n1011__;
  assign new_new_n1013__ = ~new_new_n648__ & ~new_new_n1010__;
  assign new_new_n1014__ = ~new_new_n1012__ & new_new_n1013__;
  assign new_new_n1015__ = ~new_new_n858__ & new_new_n1014__;
  assign new_new_n1016__ = new_new_n858__ & ~new_new_n1014__;
  assign new_new_n1017__ = ~new_new_n1015__ & ~new_new_n1016__;
  assign new_new_n1018__ = ~new_new_n789__ & new_new_n1017__;
  assign new_new_n1019__ = new_new_n308__ & ~new_new_n648__;
  assign new_new_n1020__ = ~new_new_n950__ & ~new_new_n1019__;
  assign new_new_n1021__ = new_new_n115__ & new_new_n270__;
  assign new_new_n1022__ = new_new_n116__ & ~new_new_n1021__;
  assign new_new_n1023__ = ~new_new_n267__ & new_new_n347__;
  assign new_new_n1024__ = ~new_new_n469__ & new_new_n1023__;
  assign new_new_n1025__ = ~new_new_n99__ & ~new_new_n1024__;
  assign new_new_n1026__ = ~new_new_n1022__ & ~new_new_n1025__;
  assign new_new_n1027__ = new_new_n195__ & ~new_new_n797__;
  assign new_new_n1028__ = ~new_new_n81__ & ~new_new_n192__;
  assign new_new_n1029__ = ~new_new_n399__ & ~new_new_n1027__;
  assign new_new_n1030__ = ~new_new_n1028__ & new_new_n1029__;
  assign new_new_n1031__ = new_new_n915__ & new_new_n1030__;
  assign new_new_n1032__ = new_new_n1026__ & new_new_n1031__;
  assign new_new_n1033__ = new_new_n125__ & ~new_new_n174__;
  assign new_new_n1034__ = ~new_new_n447__ & ~new_new_n1033__;
  assign new_new_n1035__ = new_new_n193__ & ~new_new_n227__;
  assign new_new_n1036__ = ~new_new_n181__ & ~new_new_n244__;
  assign new_new_n1037__ = ~new_new_n347__ & ~new_new_n1036__;
  assign new_new_n1038__ = ~new_new_n223__ & ~new_new_n321__;
  assign new_new_n1039__ = new_new_n218__ & new_new_n261__;
  assign new_new_n1040__ = ~new_new_n1038__ & ~new_new_n1039__;
  assign new_new_n1041__ = new_new_n116__ & ~new_new_n719__;
  assign new_new_n1042__ = new_new_n227__ & ~new_new_n1041__;
  assign new_new_n1043__ = ~new_new_n162__ & new_new_n343__;
  assign new_new_n1044__ = ~new_new_n1042__ & ~new_new_n1043__;
  assign new_new_n1045__ = new_new_n148__ & new_new_n160__;
  assign new_new_n1046__ = new_new_n244__ & ~new_new_n1045__;
  assign new_new_n1047__ = ~new_new_n240__ & ~new_new_n1046__;
  assign new_new_n1048__ = ~new_new_n1044__ & new_new_n1047__;
  assign new_new_n1049__ = ~new_new_n99__ & ~new_new_n136__;
  assign new_new_n1050__ = new_new_n141__ & ~new_new_n1049__;
  assign new_new_n1051__ = new_new_n136__ & new_new_n347__;
  assign new_new_n1052__ = ~new_new_n87__ & new_new_n99__;
  assign new_new_n1053__ = ~new_new_n1051__ & ~new_new_n1052__;
  assign new_new_n1054__ = new_new_n115__ & ~new_new_n1053__;
  assign new_new_n1055__ = ~new_new_n1050__ & ~new_new_n1054__;
  assign new_new_n1056__ = ~new_new_n219__ & ~new_new_n1055__;
  assign new_new_n1057__ = ~new_new_n252__ & ~new_new_n730__;
  assign new_new_n1058__ = ~new_new_n870__ & new_new_n1057__;
  assign new_new_n1059__ = new_new_n563__ & new_new_n1058__;
  assign new_new_n1060__ = new_new_n1034__ & ~new_new_n1035__;
  assign new_new_n1061__ = ~new_new_n1037__ & new_new_n1060__;
  assign new_new_n1062__ = ~new_new_n1040__ & new_new_n1059__;
  assign new_new_n1063__ = new_new_n1048__ & new_new_n1056__;
  assign new_new_n1064__ = new_new_n1062__ & new_new_n1063__;
  assign new_new_n1065__ = new_new_n1061__ & new_new_n1064__;
  assign new_new_n1066__ = new_new_n110__ & new_new_n218__;
  assign new_new_n1067__ = new_new_n100__ & ~new_new_n1066__;
  assign new_new_n1068__ = ~new_new_n695__ & ~new_new_n895__;
  assign new_new_n1069__ = new_new_n256__ & ~new_new_n1068__;
  assign new_new_n1070__ = ~new_new_n141__ & ~new_new_n1069__;
  assign new_new_n1071__ = ~new_new_n323__ & ~new_new_n1070__;
  assign new_new_n1072__ = ~new_new_n229__ & ~new_new_n594__;
  assign new_new_n1073__ = ~new_new_n596__ & new_new_n1072__;
  assign new_new_n1074__ = new_new_n958__ & ~new_new_n1067__;
  assign new_new_n1075__ = new_new_n1073__ & new_new_n1074__;
  assign new_new_n1076__ = new_new_n338__ & new_new_n708__;
  assign new_new_n1077__ = new_new_n1075__ & new_new_n1076__;
  assign new_new_n1078__ = new_new_n975__ & new_new_n1077__;
  assign new_new_n1079__ = new_new_n1071__ & new_new_n1078__;
  assign new_new_n1080__ = new_new_n1032__ & new_new_n1065__;
  assign new_new_n1081__ = new_new_n1079__ & new_new_n1080__;
  assign new_new_n1082__ = ~new_new_n1019__ & ~new_new_n1081__;
  assign new_new_n1083__ = ~new_new_n950__ & ~new_new_n1081__;
  assign new_new_n1084__ = new_new_n136__ & new_new_n414__;
  assign new_new_n1085__ = new_new_n181__ & ~new_new_n1084__;
  assign new_new_n1086__ = new_new_n148__ & new_new_n238__;
  assign new_new_n1087__ = ~new_new_n273__ & new_new_n1086__;
  assign new_new_n1088__ = ~new_new_n99__ & ~new_new_n1087__;
  assign new_new_n1089__ = new_new_n270__ & new_new_n910__;
  assign new_new_n1090__ = new_new_n223__ & ~new_new_n1089__;
  assign new_new_n1091__ = ~new_new_n116__ & ~new_new_n1090__;
  assign new_new_n1092__ = new_new_n180__ & new_new_n364__;
  assign new_new_n1093__ = new_new_n910__ & new_new_n1092__;
  assign new_new_n1094__ = ~new_new_n1091__ & ~new_new_n1093__;
  assign new_new_n1095__ = new_new_n81__ & new_new_n180__;
  assign new_new_n1096__ = new_new_n181__ & ~new_new_n1095__;
  assign new_new_n1097__ = new_new_n244__ & ~new_new_n414__;
  assign new_new_n1098__ = ~new_new_n323__ & ~new_new_n373__;
  assign new_new_n1099__ = ~new_new_n1096__ & new_new_n1098__;
  assign new_new_n1100__ = ~new_new_n243__ & ~new_new_n469__;
  assign new_new_n1101__ = ~new_new_n1097__ & new_new_n1100__;
  assign new_new_n1102__ = new_new_n728__ & new_new_n1099__;
  assign new_new_n1103__ = new_new_n1101__ & new_new_n1102__;
  assign new_new_n1104__ = ~new_new_n1085__ & ~new_new_n1088__;
  assign new_new_n1105__ = ~new_new_n1094__ & new_new_n1104__;
  assign new_new_n1106__ = new_new_n1103__ & new_new_n1105__;
  assign new_new_n1107__ = new_new_n160__ & new_new_n180__;
  assign new_new_n1108__ = new_new_n483__ & new_new_n1107__;
  assign new_new_n1109__ = new_new_n162__ & ~new_new_n1108__;
  assign new_new_n1110__ = new_new_n746__ & ~new_new_n1109__;
  assign new_new_n1111__ = new_new_n141__ & ~new_new_n181__;
  assign new_new_n1112__ = ~new_new_n240__ & new_new_n629__;
  assign new_new_n1113__ = ~new_new_n337__ & new_new_n1112__;
  assign new_new_n1114__ = ~new_new_n1111__ & ~new_new_n1113__;
  assign new_new_n1115__ = ~new_new_n201__ & ~new_new_n267__;
  assign new_new_n1116__ = new_new_n81__ & new_new_n174__;
  assign new_new_n1117__ = new_new_n244__ & ~new_new_n1116__;
  assign new_new_n1118__ = ~new_new_n200__ & ~new_new_n422__;
  assign new_new_n1119__ = ~new_new_n54__ & ~new_new_n1118__;
  assign new_new_n1120__ = ~new_new_n277__ & ~new_new_n1119__;
  assign new_new_n1121__ = ~new_new_n478__ & ~new_new_n1117__;
  assign new_new_n1122__ = new_new_n1115__ & new_new_n1121__;
  assign new_new_n1123__ = new_new_n1120__ & new_new_n1122__;
  assign new_new_n1124__ = new_new_n181__ & ~new_new_n270__;
  assign new_new_n1125__ = new_new_n213__ & new_new_n265__;
  assign new_new_n1126__ = new_new_n125__ & ~new_new_n1125__;
  assign new_new_n1127__ = new_new_n100__ & ~new_new_n160__;
  assign new_new_n1128__ = ~new_new_n1124__ & ~new_new_n1127__;
  assign new_new_n1129__ = ~new_new_n137__ & new_new_n1128__;
  assign new_new_n1130__ = ~new_new_n443__ & ~new_new_n451__;
  assign new_new_n1131__ = new_new_n729__ & ~new_new_n1126__;
  assign new_new_n1132__ = new_new_n1130__ & new_new_n1131__;
  assign new_new_n1133__ = new_new_n864__ & new_new_n1129__;
  assign new_new_n1134__ = new_new_n917__ & new_new_n1133__;
  assign new_new_n1135__ = new_new_n1056__ & new_new_n1132__;
  assign new_new_n1136__ = new_new_n1134__ & new_new_n1135__;
  assign new_new_n1137__ = new_new_n162__ & ~new_new_n900__;
  assign new_new_n1138__ = new_new_n125__ & ~new_new_n1089__;
  assign new_new_n1139__ = ~new_new_n222__ & ~new_new_n257__;
  assign new_new_n1140__ = ~new_new_n413__ & ~new_new_n1137__;
  assign new_new_n1141__ = new_new_n1139__ & new_new_n1140__;
  assign new_new_n1142__ = ~new_new_n1138__ & new_new_n1141__;
  assign new_new_n1143__ = new_new_n1110__ & new_new_n1142__;
  assign new_new_n1144__ = ~new_new_n1114__ & new_new_n1123__;
  assign new_new_n1145__ = new_new_n1143__ & new_new_n1144__;
  assign new_new_n1146__ = new_new_n1136__ & new_new_n1145__;
  assign new_new_n1147__ = new_new_n1106__ & new_new_n1146__;
  assign new_new_n1148__ = new_new_n1083__ & new_new_n1147__;
  assign new_new_n1149__ = ~new_new_n1082__ & ~new_new_n1148__;
  assign new_new_n1150__ = ~new_new_n1020__ & new_new_n1149__;
  assign new_new_n1151__ = new_new_n760__ & ~new_new_n842__;
  assign new_new_n1152__ = new_new_n686__ & new_new_n816__;
  assign new_new_n1153__ = ~new_new_n686__ & ~new_new_n816__;
  assign new_new_n1154__ = ~new_new_n1152__ & ~new_new_n1153__;
  assign new_new_n1155__ = new_new_n608__ & new_new_n816__;
  assign new_new_n1156__ = ~new_new_n608__ & ~new_new_n816__;
  assign new_new_n1157__ = ~new_new_n1155__ & ~new_new_n1156__;
  assign new_new_n1158__ = ~new_new_n760__ & new_new_n1154__;
  assign new_new_n1159__ = ~new_new_n1157__ & new_new_n1158__;
  assign new_new_n1160__ = ~new_new_n1151__ & ~new_new_n1159__;
  assign new_new_n1161__ = new_new_n1150__ & ~new_new_n1160__;
  assign new_new_n1162__ = ~new_new_n1150__ & new_new_n1160__;
  assign new_new_n1163__ = ~new_new_n1161__ & ~new_new_n1162__;
  assign new_new_n1164__ = ~new_new_n301__ & ~new_new_n805__;
  assign new_new_n1165__ = new_new_n301__ & new_new_n791__;
  assign new_new_n1166__ = ~new_new_n1164__ & ~new_new_n1165__;
  assign new_new_n1167__ = new_new_n615__ & ~new_new_n805__;
  assign new_new_n1168__ = new_new_n792__ & ~new_new_n1167__;
  assign new_new_n1169__ = ~new_new_n1166__ & ~new_new_n1168__;
  assign new_new_n1170__ = new_new_n1163__ & new_new_n1169__;
  assign new_new_n1171__ = ~new_new_n1161__ & ~new_new_n1170__;
  assign new_new_n1172__ = ~new_new_n437__ & new_new_n950__;
  assign new_new_n1173__ = new_new_n1007__ & new_new_n1172__;
  assign new_new_n1174__ = new_new_n1009__ & ~new_new_n1173__;
  assign new_new_n1175__ = new_new_n430__ & new_new_n1008__;
  assign new_new_n1176__ = ~new_new_n437__ & new_new_n1175__;
  assign new_new_n1177__ = ~new_new_n1174__ & ~new_new_n1176__;
  assign new_new_n1178__ = new_new_n316__ & ~new_new_n648__;
  assign new_new_n1179__ = ~new_new_n1177__ & ~new_new_n1178__;
  assign new_new_n1180__ = new_new_n1177__ & new_new_n1178__;
  assign new_new_n1181__ = new_new_n824__ & new_new_n829__;
  assign new_new_n1182__ = ~new_new_n430__ & ~new_new_n764__;
  assign new_new_n1183__ = new_new_n430__ & new_new_n764__;
  assign new_new_n1184__ = ~new_new_n1182__ & ~new_new_n1183__;
  assign new_new_n1185__ = ~new_new_n767__ & ~new_new_n824__;
  assign new_new_n1186__ = new_new_n1184__ & new_new_n1185__;
  assign new_new_n1187__ = ~new_new_n1181__ & ~new_new_n1186__;
  assign new_new_n1188__ = ~new_new_n1180__ & ~new_new_n1187__;
  assign new_new_n1189__ = ~new_new_n1179__ & ~new_new_n1188__;
  assign new_new_n1190__ = new_new_n1171__ & new_new_n1189__;
  assign new_new_n1191__ = new_new_n301__ & new_new_n316__;
  assign new_new_n1192__ = ~new_new_n301__ & ~new_new_n316__;
  assign new_new_n1193__ = ~new_new_n1191__ & ~new_new_n1192__;
  assign new_new_n1194__ = ~new_new_n648__ & ~new_new_n1193__;
  assign new_new_n1195__ = ~new_new_n1009__ & new_new_n1194__;
  assign new_new_n1196__ = new_new_n1009__ & ~new_new_n1194__;
  assign new_new_n1197__ = ~new_new_n1195__ & ~new_new_n1196__;
  assign new_new_n1198__ = ~new_new_n1190__ & new_new_n1197__;
  assign new_new_n1199__ = new_new_n789__ & ~new_new_n1017__;
  assign new_new_n1200__ = ~new_new_n1171__ & ~new_new_n1189__;
  assign new_new_n1201__ = ~new_new_n1198__ & ~new_new_n1200__;
  assign new_new_n1202__ = ~new_new_n1199__ & new_new_n1201__;
  assign new_new_n1203__ = ~new_new_n1018__ & new_new_n1202__;
  assign new_new_n1204__ = new_new_n1018__ & ~new_new_n1189__;
  assign new_new_n1205__ = new_new_n1197__ & new_new_n1199__;
  assign new_new_n1206__ = ~new_new_n1204__ & ~new_new_n1205__;
  assign new_new_n1207__ = ~new_new_n1171__ & ~new_new_n1206__;
  assign new_new_n1208__ = ~new_new_n1190__ & ~new_new_n1200__;
  assign new_new_n1209__ = ~new_new_n1197__ & new_new_n1208__;
  assign new_new_n1210__ = new_new_n1197__ & ~new_new_n1208__;
  assign new_new_n1211__ = ~new_new_n1209__ & ~new_new_n1210__;
  assign new_new_n1212__ = ~new_new_n1189__ & new_new_n1199__;
  assign new_new_n1213__ = new_new_n1018__ & new_new_n1197__;
  assign new_new_n1214__ = ~new_new_n1212__ & ~new_new_n1213__;
  assign new_new_n1215__ = new_new_n1211__ & ~new_new_n1214__;
  assign new_new_n1216__ = ~new_new_n1203__ & ~new_new_n1207__;
  assign new_new_n1217__ = ~new_new_n1215__ & new_new_n1216__;
  assign new_new_n1218__ = new_new_n1177__ & ~new_new_n1178__;
  assign new_new_n1219__ = ~new_new_n1177__ & new_new_n1178__;
  assign new_new_n1220__ = ~new_new_n1218__ & ~new_new_n1219__;
  assign new_new_n1221__ = new_new_n1187__ & new_new_n1220__;
  assign new_new_n1222__ = ~new_new_n1187__ & ~new_new_n1220__;
  assign new_new_n1223__ = ~new_new_n1221__ & ~new_new_n1222__;
  assign new_new_n1224__ = new_new_n651__ & new_new_n1008__;
  assign new_new_n1225__ = new_new_n950__ & new_new_n1007__;
  assign new_new_n1226__ = ~new_new_n1008__ & ~new_new_n1225__;
  assign new_new_n1227__ = ~new_new_n437__ & new_new_n1226__;
  assign new_new_n1228__ = ~new_new_n1224__ & ~new_new_n1227__;
  assign new_new_n1229__ = new_new_n430__ & ~new_new_n1228__;
  assign new_new_n1230__ = new_new_n651__ & new_new_n1225__;
  assign new_new_n1231__ = ~new_new_n437__ & ~new_new_n1225__;
  assign new_new_n1232__ = new_new_n1009__ & ~new_new_n1230__;
  assign new_new_n1233__ = ~new_new_n1231__ & new_new_n1232__;
  assign new_new_n1234__ = ~new_new_n1229__ & ~new_new_n1233__;
  assign new_new_n1235__ = new_new_n760__ & new_new_n1154__;
  assign new_new_n1236__ = new_new_n615__ & new_new_n686__;
  assign new_new_n1237__ = new_new_n758__ & new_new_n1236__;
  assign new_new_n1238__ = ~new_new_n686__ & new_new_n759__;
  assign new_new_n1239__ = ~new_new_n615__ & new_new_n1238__;
  assign new_new_n1240__ = ~new_new_n1235__ & ~new_new_n1237__;
  assign new_new_n1241__ = ~new_new_n1239__ & new_new_n1240__;
  assign new_new_n1242__ = new_new_n1234__ & new_new_n1241__;
  assign new_new_n1243__ = ~new_new_n1234__ & ~new_new_n1241__;
  assign new_new_n1244__ = ~new_new_n316__ & ~new_new_n791__;
  assign new_new_n1245__ = new_new_n792__ & ~new_new_n1164__;
  assign new_new_n1246__ = new_new_n316__ & new_new_n805__;
  assign new_new_n1247__ = ~new_new_n1244__ & ~new_new_n1246__;
  assign new_new_n1248__ = ~new_new_n1245__ & new_new_n1247__;
  assign new_new_n1249__ = ~new_new_n1243__ & ~new_new_n1248__;
  assign new_new_n1250__ = ~new_new_n1242__ & ~new_new_n1249__;
  assign new_new_n1251__ = ~new_new_n1163__ & ~new_new_n1169__;
  assign new_new_n1252__ = ~new_new_n1170__ & ~new_new_n1251__;
  assign new_new_n1253__ = new_new_n1250__ & new_new_n1252__;
  assign new_new_n1254__ = ~new_new_n1223__ & ~new_new_n1253__;
  assign new_new_n1255__ = ~new_new_n1250__ & ~new_new_n1252__;
  assign new_new_n1256__ = ~new_new_n1254__ & ~new_new_n1255__;
  assign new_new_n1257__ = ~new_new_n615__ & ~new_new_n686__;
  assign new_new_n1258__ = ~new_new_n1236__ & ~new_new_n1257__;
  assign new_new_n1259__ = new_new_n760__ & ~new_new_n1258__;
  assign new_new_n1260__ = new_new_n301__ & new_new_n686__;
  assign new_new_n1261__ = ~new_new_n301__ & ~new_new_n686__;
  assign new_new_n1262__ = ~new_new_n1260__ & ~new_new_n1261__;
  assign new_new_n1263__ = new_new_n301__ & new_new_n608__;
  assign new_new_n1264__ = ~new_new_n301__ & ~new_new_n608__;
  assign new_new_n1265__ = ~new_new_n1263__ & ~new_new_n1264__;
  assign new_new_n1266__ = ~new_new_n760__ & new_new_n1262__;
  assign new_new_n1267__ = ~new_new_n1265__ & new_new_n1266__;
  assign new_new_n1268__ = ~new_new_n1259__ & ~new_new_n1267__;
  assign new_new_n1269__ = new_new_n832__ & new_new_n1226__;
  assign new_new_n1270__ = ~new_new_n764__ & ~new_new_n950__;
  assign new_new_n1271__ = new_new_n764__ & new_new_n950__;
  assign new_new_n1272__ = ~new_new_n1270__ & ~new_new_n1271__;
  assign new_new_n1273__ = ~new_new_n1184__ & ~new_new_n1226__;
  assign new_new_n1274__ = new_new_n1272__ & new_new_n1273__;
  assign new_new_n1275__ = ~new_new_n1269__ & ~new_new_n1274__;
  assign new_new_n1276__ = ~new_new_n1268__ & ~new_new_n1275__;
  assign new_new_n1277__ = new_new_n1268__ & new_new_n1275__;
  assign new_new_n1278__ = new_new_n824__ & ~new_new_n839__;
  assign new_new_n1279__ = new_new_n430__ & new_new_n816__;
  assign new_new_n1280__ = ~new_new_n430__ & ~new_new_n816__;
  assign new_new_n1281__ = ~new_new_n1279__ & ~new_new_n1280__;
  assign new_new_n1282__ = ~new_new_n824__ & new_new_n1157__;
  assign new_new_n1283__ = ~new_new_n1281__ & new_new_n1282__;
  assign new_new_n1284__ = ~new_new_n1278__ & ~new_new_n1283__;
  assign new_new_n1285__ = ~new_new_n1277__ & ~new_new_n1284__;
  assign new_new_n1286__ = ~new_new_n1276__ & ~new_new_n1285__;
  assign new_new_n1287__ = ~new_new_n1184__ & new_new_n1226__;
  assign new_new_n1288__ = new_new_n810__ & new_new_n950__;
  assign new_new_n1289__ = ~new_new_n810__ & ~new_new_n950__;
  assign new_new_n1290__ = ~new_new_n1288__ & ~new_new_n1289__;
  assign new_new_n1291__ = new_new_n430__ & new_new_n810__;
  assign new_new_n1292__ = ~new_new_n430__ & ~new_new_n810__;
  assign new_new_n1293__ = ~new_new_n1291__ & ~new_new_n1292__;
  assign new_new_n1294__ = ~new_new_n1226__ & new_new_n1290__;
  assign new_new_n1295__ = ~new_new_n1293__ & new_new_n1294__;
  assign new_new_n1296__ = ~new_new_n1287__ & ~new_new_n1295__;
  assign new_new_n1297__ = new_new_n760__ & new_new_n1262__;
  assign new_new_n1298__ = new_new_n316__ & new_new_n608__;
  assign new_new_n1299__ = ~new_new_n316__ & ~new_new_n608__;
  assign new_new_n1300__ = ~new_new_n1298__ & ~new_new_n1299__;
  assign new_new_n1301__ = new_new_n316__ & new_new_n686__;
  assign new_new_n1302__ = ~new_new_n316__ & ~new_new_n686__;
  assign new_new_n1303__ = ~new_new_n1301__ & ~new_new_n1302__;
  assign new_new_n1304__ = ~new_new_n760__ & ~new_new_n1303__;
  assign new_new_n1305__ = new_new_n1300__ & new_new_n1304__;
  assign new_new_n1306__ = ~new_new_n1297__ & ~new_new_n1305__;
  assign new_new_n1307__ = ~new_new_n1296__ & ~new_new_n1306__;
  assign new_new_n1308__ = new_new_n1296__ & new_new_n1306__;
  assign new_new_n1309__ = new_new_n824__ & new_new_n1157__;
  assign new_new_n1310__ = ~new_new_n430__ & ~new_new_n615__;
  assign new_new_n1311__ = ~new_new_n608__ & ~new_new_n615__;
  assign new_new_n1312__ = ~new_new_n784__ & ~new_new_n1311__;
  assign new_new_n1313__ = ~new_new_n777__ & ~new_new_n1310__;
  assign new_new_n1314__ = ~new_new_n1312__ & new_new_n1313__;
  assign new_new_n1315__ = ~new_new_n1309__ & ~new_new_n1314__;
  assign new_new_n1316__ = ~new_new_n1308__ & ~new_new_n1315__;
  assign new_new_n1317__ = ~new_new_n1307__ & ~new_new_n1316__;
  assign new_new_n1318__ = ~new_new_n1081__ & ~new_new_n1147__;
  assign new_new_n1319__ = new_new_n950__ & new_new_n1318__;
  assign new_new_n1320__ = new_new_n651__ & new_new_n1319__;
  assign new_new_n1321__ = ~pi22 & ~new_new_n59__;
  assign new_new_n1322__ = pi04 & ~new_new_n1321__;
  assign new_new_n1323__ = ~pi04 & new_new_n1321__;
  assign new_new_n1324__ = ~new_new_n1322__ & ~new_new_n1323__;
  assign new_new_n1325__ = ~new_new_n648__ & ~new_new_n1324__;
  assign new_new_n1326__ = ~new_new_n950__ & new_new_n1147__;
  assign new_new_n1327__ = ~new_new_n651__ & new_new_n1326__;
  assign new_new_n1328__ = new_new_n1081__ & ~new_new_n1327__;
  assign new_new_n1329__ = new_new_n1325__ & ~new_new_n1328__;
  assign new_new_n1330__ = ~new_new_n1147__ & ~new_new_n1325__;
  assign new_new_n1331__ = new_new_n1081__ & new_new_n1147__;
  assign new_new_n1332__ = new_new_n437__ & ~new_new_n950__;
  assign new_new_n1333__ = ~new_new_n1172__ & ~new_new_n1332__;
  assign new_new_n1334__ = ~new_new_n1330__ & ~new_new_n1331__;
  assign new_new_n1335__ = ~new_new_n1333__ & new_new_n1334__;
  assign new_new_n1336__ = ~new_new_n1320__ & ~new_new_n1335__;
  assign new_new_n1337__ = ~new_new_n1329__ & new_new_n1336__;
  assign new_new_n1338__ = ~new_new_n1317__ & ~new_new_n1337__;
  assign new_new_n1339__ = new_new_n1317__ & new_new_n1337__;
  assign new_new_n1340__ = new_new_n791__ & ~new_new_n805__;
  assign new_new_n1341__ = new_new_n316__ & new_new_n1340__;
  assign new_new_n1342__ = ~new_new_n308__ & ~new_new_n648__;
  assign new_new_n1343__ = new_new_n308__ & ~new_new_n791__;
  assign new_new_n1344__ = ~new_new_n1342__ & ~new_new_n1343__;
  assign new_new_n1345__ = ~new_new_n1341__ & new_new_n1344__;
  assign new_new_n1346__ = ~new_new_n1339__ & ~new_new_n1345__;
  assign new_new_n1347__ = ~new_new_n1338__ & ~new_new_n1346__;
  assign new_new_n1348__ = ~new_new_n1286__ & ~new_new_n1347__;
  assign new_new_n1349__ = new_new_n1286__ & new_new_n1347__;
  assign new_new_n1350__ = ~new_new_n1242__ & ~new_new_n1243__;
  assign new_new_n1351__ = ~new_new_n1248__ & new_new_n1350__;
  assign new_new_n1352__ = new_new_n1248__ & ~new_new_n1350__;
  assign new_new_n1353__ = ~new_new_n1351__ & ~new_new_n1352__;
  assign new_new_n1354__ = ~new_new_n1349__ & ~new_new_n1353__;
  assign new_new_n1355__ = ~new_new_n1348__ & ~new_new_n1354__;
  assign new_new_n1356__ = new_new_n310__ & ~new_new_n648__;
  assign new_new_n1357__ = new_new_n1081__ & ~new_new_n1332__;
  assign new_new_n1358__ = new_new_n1356__ & ~new_new_n1357__;
  assign new_new_n1359__ = ~new_new_n950__ & ~new_new_n1356__;
  assign new_new_n1360__ = ~new_new_n437__ & ~new_new_n1081__;
  assign new_new_n1361__ = new_new_n950__ & ~new_new_n1360__;
  assign new_new_n1362__ = ~new_new_n1147__ & ~new_new_n1359__;
  assign new_new_n1363__ = ~new_new_n1361__ & new_new_n1362__;
  assign new_new_n1364__ = ~new_new_n1358__ & ~new_new_n1363__;
  assign new_new_n1365__ = ~new_new_n1019__ & ~new_new_n1364__;
  assign new_new_n1366__ = ~new_new_n1326__ & new_new_n1365__;
  assign new_new_n1367__ = ~new_new_n767__ & new_new_n824__;
  assign new_new_n1368__ = ~new_new_n824__ & ~new_new_n839__;
  assign new_new_n1369__ = new_new_n1293__ & new_new_n1368__;
  assign new_new_n1370__ = ~new_new_n1367__ & ~new_new_n1369__;
  assign new_new_n1371__ = new_new_n1019__ & ~new_new_n1370__;
  assign new_new_n1372__ = new_new_n950__ & new_new_n1371__;
  assign new_new_n1373__ = ~new_new_n1365__ & ~new_new_n1372__;
  assign new_new_n1374__ = new_new_n1081__ & ~new_new_n1373__;
  assign new_new_n1375__ = ~new_new_n1019__ & new_new_n1370__;
  assign new_new_n1376__ = ~new_new_n1149__ & ~new_new_n1375__;
  assign new_new_n1377__ = ~new_new_n1020__ & new_new_n1364__;
  assign new_new_n1378__ = ~new_new_n1370__ & ~new_new_n1377__;
  assign new_new_n1379__ = ~new_new_n1366__ & ~new_new_n1378__;
  assign new_new_n1380__ = ~new_new_n1376__ & new_new_n1379__;
  assign new_new_n1381__ = ~new_new_n1374__ & new_new_n1380__;
  assign new_new_n1382__ = ~new_new_n1355__ & ~new_new_n1381__;
  assign new_new_n1383__ = new_new_n1169__ & new_new_n1223__;
  assign new_new_n1384__ = ~new_new_n1169__ & ~new_new_n1223__;
  assign new_new_n1385__ = ~new_new_n1383__ & ~new_new_n1384__;
  assign new_new_n1386__ = new_new_n1163__ & ~new_new_n1250__;
  assign new_new_n1387__ = ~new_new_n1163__ & new_new_n1250__;
  assign new_new_n1388__ = ~new_new_n1386__ & ~new_new_n1387__;
  assign new_new_n1389__ = new_new_n1385__ & ~new_new_n1388__;
  assign new_new_n1390__ = new_new_n1355__ & new_new_n1381__;
  assign new_new_n1391__ = ~new_new_n1385__ & new_new_n1388__;
  assign new_new_n1392__ = ~new_new_n1389__ & ~new_new_n1391__;
  assign new_new_n1393__ = ~new_new_n1390__ & new_new_n1392__;
  assign new_new_n1394__ = ~new_new_n1382__ & ~new_new_n1393__;
  assign new_new_n1395__ = ~new_new_n1211__ & ~new_new_n1394__;
  assign new_new_n1396__ = new_new_n1226__ & new_new_n1281__;
  assign new_new_n1397__ = new_new_n430__ & new_new_n615__;
  assign new_new_n1398__ = ~new_new_n1225__ & ~new_new_n1397__;
  assign new_new_n1399__ = ~new_new_n1008__ & ~new_new_n1310__;
  assign new_new_n1400__ = ~new_new_n1398__ & ~new_new_n1399__;
  assign new_new_n1401__ = ~new_new_n1396__ & ~new_new_n1400__;
  assign new_new_n1402__ = ~new_new_n308__ & ~new_new_n686__;
  assign new_new_n1403__ = new_new_n308__ & new_new_n686__;
  assign new_new_n1404__ = ~new_new_n1402__ & ~new_new_n1403__;
  assign new_new_n1405__ = new_new_n760__ & ~new_new_n1404__;
  assign new_new_n1406__ = ~new_new_n310__ & ~new_new_n608__;
  assign new_new_n1407__ = new_new_n310__ & new_new_n608__;
  assign new_new_n1408__ = ~new_new_n1406__ & ~new_new_n1407__;
  assign new_new_n1409__ = ~new_new_n310__ & ~new_new_n686__;
  assign new_new_n1410__ = new_new_n310__ & new_new_n686__;
  assign new_new_n1411__ = ~new_new_n1409__ & ~new_new_n1410__;
  assign new_new_n1412__ = ~new_new_n760__ & ~new_new_n1411__;
  assign new_new_n1413__ = new_new_n1408__ & new_new_n1412__;
  assign new_new_n1414__ = ~new_new_n1405__ & ~new_new_n1413__;
  assign new_new_n1415__ = ~new_new_n1401__ & ~new_new_n1414__;
  assign new_new_n1416__ = new_new_n1401__ & new_new_n1414__;
  assign new_new_n1417__ = new_new_n824__ & new_new_n1265__;
  assign new_new_n1418__ = new_new_n316__ & new_new_n430__;
  assign new_new_n1419__ = ~new_new_n316__ & ~new_new_n430__;
  assign new_new_n1420__ = ~new_new_n1418__ & ~new_new_n1419__;
  assign new_new_n1421__ = ~new_new_n824__ & ~new_new_n1300__;
  assign new_new_n1422__ = new_new_n1420__ & new_new_n1421__;
  assign new_new_n1423__ = ~new_new_n1417__ & ~new_new_n1422__;
  assign new_new_n1424__ = ~new_new_n1416__ & ~new_new_n1423__;
  assign new_new_n1425__ = ~new_new_n1415__ & ~new_new_n1424__;
  assign new_new_n1426__ = ~new_new_n805__ & ~new_new_n1324__;
  assign new_new_n1427__ = new_new_n791__ & new_new_n1324__;
  assign new_new_n1428__ = ~new_new_n1426__ & ~new_new_n1427__;
  assign new_new_n1429__ = new_new_n310__ & ~new_new_n805__;
  assign new_new_n1430__ = new_new_n792__ & ~new_new_n1429__;
  assign new_new_n1431__ = ~new_new_n1428__ & ~new_new_n1430__;
  assign new_new_n1432__ = new_new_n1425__ & ~new_new_n1431__;
  assign new_new_n1433__ = ~new_new_n1425__ & new_new_n1431__;
  assign new_new_n1434__ = ~new_new_n87__ & ~new_new_n581__;
  assign new_new_n1435__ = new_new_n54__ & ~new_new_n1434__;
  assign new_new_n1436__ = ~new_new_n87__ & new_new_n124__;
  assign new_new_n1437__ = ~new_new_n581__ & ~new_new_n1436__;
  assign new_new_n1438__ = new_new_n347__ & ~new_new_n1437__;
  assign new_new_n1439__ = ~new_new_n1435__ & ~new_new_n1438__;
  assign new_new_n1440__ = new_new_n181__ & ~new_new_n487__;
  assign new_new_n1441__ = ~new_new_n229__ & ~new_new_n662__;
  assign new_new_n1442__ = ~new_new_n243__ & ~new_new_n730__;
  assign new_new_n1443__ = new_new_n279__ & ~new_new_n337__;
  assign new_new_n1444__ = ~new_new_n863__ & new_new_n1443__;
  assign new_new_n1445__ = new_new_n1115__ & new_new_n1442__;
  assign new_new_n1446__ = new_new_n1441__ & new_new_n1445__;
  assign new_new_n1447__ = new_new_n1444__ & new_new_n1446__;
  assign new_new_n1448__ = ~new_new_n325__ & ~new_new_n451__;
  assign new_new_n1449__ = ~new_new_n546__ & new_new_n1448__;
  assign new_new_n1450__ = ~new_new_n351__ & ~new_new_n377__;
  assign new_new_n1451__ = new_new_n99__ & new_new_n214__;
  assign new_new_n1452__ = new_new_n181__ & ~new_new_n1451__;
  assign new_new_n1453__ = new_new_n100__ & ~new_new_n1045__;
  assign new_new_n1454__ = ~new_new_n244__ & ~new_new_n446__;
  assign new_new_n1455__ = new_new_n218__ & new_new_n414__;
  assign new_new_n1456__ = ~new_new_n1454__ & ~new_new_n1455__;
  assign new_new_n1457__ = ~new_new_n555__ & ~new_new_n1453__;
  assign new_new_n1458__ = new_new_n1450__ & new_new_n1457__;
  assign new_new_n1459__ = ~new_new_n1452__ & ~new_new_n1456__;
  assign new_new_n1460__ = new_new_n1458__ & new_new_n1459__;
  assign new_new_n1461__ = new_new_n584__ & new_new_n1449__;
  assign new_new_n1462__ = new_new_n1460__ & new_new_n1461__;
  assign new_new_n1463__ = new_new_n195__ & ~new_new_n677__;
  assign new_new_n1464__ = new_new_n116__ & ~new_new_n1095__;
  assign new_new_n1465__ = ~new_new_n196__ & new_new_n223__;
  assign new_new_n1466__ = ~new_new_n160__ & ~new_new_n1111__;
  assign new_new_n1467__ = ~new_new_n168__ & ~new_new_n1464__;
  assign new_new_n1468__ = ~new_new_n188__ & ~new_new_n1465__;
  assign new_new_n1469__ = ~new_new_n1466__ & new_new_n1468__;
  assign new_new_n1470__ = new_new_n1467__ & new_new_n1469__;
  assign new_new_n1471__ = ~new_new_n1440__ & ~new_new_n1463__;
  assign new_new_n1472__ = ~new_new_n1439__ & new_new_n1471__;
  assign new_new_n1473__ = new_new_n636__ & new_new_n1472__;
  assign new_new_n1474__ = new_new_n1470__ & new_new_n1473__;
  assign new_new_n1475__ = new_new_n1447__ & new_new_n1462__;
  assign new_new_n1476__ = new_new_n1474__ & new_new_n1475__;
  assign new_new_n1477__ = ~new_new_n1081__ & new_new_n1476__;
  assign new_new_n1478__ = ~new_new_n648__ & ~new_new_n651__;
  assign new_new_n1479__ = new_new_n1477__ & new_new_n1478__;
  assign new_new_n1480__ = new_new_n437__ & new_new_n1081__;
  assign new_new_n1481__ = ~new_new_n651__ & ~new_new_n1081__;
  assign new_new_n1482__ = new_new_n1476__ & ~new_new_n1481__;
  assign new_new_n1483__ = ~new_new_n1480__ & ~new_new_n1482__;
  assign new_new_n1484__ = new_new_n648__ & ~new_new_n1483__;
  assign new_new_n1485__ = new_new_n648__ & ~new_new_n1360__;
  assign new_new_n1486__ = ~new_new_n1360__ & ~new_new_n1480__;
  assign new_new_n1487__ = ~new_new_n648__ & ~new_new_n1486__;
  assign new_new_n1488__ = ~new_new_n1476__ & ~new_new_n1485__;
  assign new_new_n1489__ = ~new_new_n1487__ & new_new_n1488__;
  assign new_new_n1490__ = ~new_new_n1479__ & ~new_new_n1484__;
  assign new_new_n1491__ = ~new_new_n1489__ & new_new_n1490__;
  assign new_new_n1492__ = ~new_new_n648__ & ~new_new_n1491__;
  assign new_new_n1493__ = ~new_new_n1433__ & ~new_new_n1492__;
  assign new_new_n1494__ = ~new_new_n1432__ & ~new_new_n1493__;
  assign new_new_n1495__ = ~new_new_n1318__ & ~new_new_n1331__;
  assign new_new_n1496__ = new_new_n950__ & new_new_n1081__;
  assign new_new_n1497__ = ~new_new_n651__ & ~new_new_n1496__;
  assign new_new_n1498__ = ~new_new_n1495__ & new_new_n1497__;
  assign new_new_n1499__ = new_new_n950__ & ~new_new_n1147__;
  assign new_new_n1500__ = ~new_new_n1326__ & ~new_new_n1499__;
  assign new_new_n1501__ = ~new_new_n1496__ & new_new_n1500__;
  assign new_new_n1502__ = new_new_n437__ & new_new_n1501__;
  assign new_new_n1503__ = ~new_new_n1083__ & ~new_new_n1496__;
  assign new_new_n1504__ = ~new_new_n437__ & ~new_new_n1331__;
  assign new_new_n1505__ = ~new_new_n1503__ & new_new_n1504__;
  assign new_new_n1506__ = ~new_new_n1325__ & ~new_new_n1498__;
  assign new_new_n1507__ = ~new_new_n1505__ & new_new_n1506__;
  assign new_new_n1508__ = ~new_new_n1502__ & new_new_n1507__;
  assign new_new_n1509__ = ~new_new_n1318__ & ~new_new_n1503__;
  assign new_new_n1510__ = new_new_n437__ & new_new_n1509__;
  assign new_new_n1511__ = ~new_new_n437__ & new_new_n1500__;
  assign new_new_n1512__ = new_new_n651__ & ~new_new_n1495__;
  assign new_new_n1513__ = ~new_new_n1511__ & ~new_new_n1512__;
  assign new_new_n1514__ = ~new_new_n1083__ & ~new_new_n1513__;
  assign new_new_n1515__ = new_new_n1325__ & ~new_new_n1510__;
  assign new_new_n1516__ = ~new_new_n1514__ & new_new_n1515__;
  assign new_new_n1517__ = ~new_new_n1508__ & ~new_new_n1516__;
  assign new_new_n1518__ = ~new_new_n1494__ & ~new_new_n1517__;
  assign new_new_n1519__ = new_new_n1494__ & new_new_n1517__;
  assign new_new_n1520__ = ~new_new_n1307__ & ~new_new_n1308__;
  assign new_new_n1521__ = ~new_new_n1315__ & new_new_n1520__;
  assign new_new_n1522__ = new_new_n1315__ & ~new_new_n1520__;
  assign new_new_n1523__ = ~new_new_n1521__ & ~new_new_n1522__;
  assign new_new_n1524__ = ~new_new_n1519__ & ~new_new_n1523__;
  assign new_new_n1525__ = ~new_new_n1518__ & ~new_new_n1524__;
  assign new_new_n1526__ = new_new_n1226__ & ~new_new_n1293__;
  assign new_new_n1527__ = new_new_n816__ & new_new_n950__;
  assign new_new_n1528__ = ~new_new_n816__ & ~new_new_n950__;
  assign new_new_n1529__ = ~new_new_n1527__ & ~new_new_n1528__;
  assign new_new_n1530__ = ~new_new_n1226__ & new_new_n1281__;
  assign new_new_n1531__ = ~new_new_n1529__ & new_new_n1530__;
  assign new_new_n1532__ = ~new_new_n1526__ & ~new_new_n1531__;
  assign new_new_n1533__ = new_new_n760__ & ~new_new_n1303__;
  assign new_new_n1534__ = ~new_new_n308__ & ~new_new_n608__;
  assign new_new_n1535__ = new_new_n308__ & new_new_n608__;
  assign new_new_n1536__ = ~new_new_n1534__ & ~new_new_n1535__;
  assign new_new_n1537__ = ~new_new_n760__ & ~new_new_n1404__;
  assign new_new_n1538__ = new_new_n1536__ & new_new_n1537__;
  assign new_new_n1539__ = ~new_new_n1533__ & ~new_new_n1538__;
  assign new_new_n1540__ = ~new_new_n1532__ & ~new_new_n1539__;
  assign new_new_n1541__ = new_new_n1532__ & new_new_n1539__;
  assign new_new_n1542__ = new_new_n608__ & new_new_n615__;
  assign new_new_n1543__ = ~new_new_n1311__ & ~new_new_n1542__;
  assign new_new_n1544__ = new_new_n824__ & ~new_new_n1543__;
  assign new_new_n1545__ = ~new_new_n301__ & ~new_new_n430__;
  assign new_new_n1546__ = new_new_n301__ & new_new_n430__;
  assign new_new_n1547__ = ~new_new_n1545__ & ~new_new_n1546__;
  assign new_new_n1548__ = ~new_new_n824__ & new_new_n1265__;
  assign new_new_n1549__ = ~new_new_n1547__ & new_new_n1548__;
  assign new_new_n1550__ = ~new_new_n1544__ & ~new_new_n1549__;
  assign new_new_n1551__ = ~new_new_n1541__ & ~new_new_n1550__;
  assign new_new_n1552__ = ~new_new_n1540__ & ~new_new_n1551__;
  assign new_new_n1553__ = new_new_n651__ & new_new_n950__;
  assign new_new_n1554__ = ~new_new_n651__ & ~new_new_n950__;
  assign new_new_n1555__ = ~new_new_n1553__ & ~new_new_n1554__;
  assign new_new_n1556__ = new_new_n1495__ & ~new_new_n1555__;
  assign new_new_n1557__ = ~new_new_n764__ & ~new_new_n1081__;
  assign new_new_n1558__ = new_new_n764__ & new_new_n1081__;
  assign new_new_n1559__ = ~new_new_n1557__ & ~new_new_n1558__;
  assign new_new_n1560__ = ~new_new_n1495__ & ~new_new_n1500__;
  assign new_new_n1561__ = new_new_n1559__ & new_new_n1560__;
  assign new_new_n1562__ = ~new_new_n1556__ & ~new_new_n1561__;
  assign new_new_n1563__ = ~new_new_n1081__ & ~new_new_n1476__;
  assign new_new_n1564__ = new_new_n437__ & ~new_new_n1081__;
  assign new_new_n1565__ = ~new_new_n1563__ & ~new_new_n1564__;
  assign new_new_n1566__ = new_new_n1562__ & new_new_n1565__;
  assign new_new_n1567__ = ~new_new_n1562__ & ~new_new_n1565__;
  assign new_new_n1568__ = ~pi01 & ~pi02;
  assign new_new_n1569__ = ~pi00 & new_new_n1568__;
  assign new_new_n1570__ = ~pi22 & ~new_new_n1569__;
  assign new_new_n1571__ = pi03 & new_new_n1570__;
  assign new_new_n1572__ = ~pi03 & ~new_new_n1570__;
  assign new_new_n1573__ = ~new_new_n1571__ & ~new_new_n1572__;
  assign new_new_n1574__ = ~new_new_n648__ & new_new_n1573__;
  assign new_new_n1575__ = ~new_new_n1567__ & ~new_new_n1574__;
  assign new_new_n1576__ = ~new_new_n1566__ & ~new_new_n1575__;
  assign new_new_n1577__ = ~new_new_n1552__ & new_new_n1576__;
  assign new_new_n1578__ = new_new_n1552__ & ~new_new_n1576__;
  assign new_new_n1579__ = ~new_new_n1577__ & ~new_new_n1578__;
  assign new_new_n1580__ = new_new_n310__ & ~new_new_n791__;
  assign new_new_n1581__ = ~new_new_n310__ & ~new_new_n648__;
  assign new_new_n1582__ = new_new_n308__ & new_new_n1340__;
  assign new_new_n1583__ = ~new_new_n1580__ & ~new_new_n1581__;
  assign new_new_n1584__ = ~new_new_n1582__ & new_new_n1583__;
  assign new_new_n1585__ = new_new_n1579__ & ~new_new_n1584__;
  assign new_new_n1586__ = ~new_new_n1577__ & ~new_new_n1585__;
  assign new_new_n1587__ = new_new_n437__ & new_new_n1503__;
  assign new_new_n1588__ = ~new_new_n1356__ & ~new_new_n1501__;
  assign new_new_n1589__ = ~new_new_n1587__ & new_new_n1588__;
  assign new_new_n1590__ = ~new_new_n437__ & ~new_new_n1500__;
  assign new_new_n1591__ = new_new_n1356__ & ~new_new_n1509__;
  assign new_new_n1592__ = ~new_new_n1590__ & new_new_n1591__;
  assign new_new_n1593__ = ~new_new_n1589__ & ~new_new_n1592__;
  assign new_new_n1594__ = ~new_new_n1586__ & new_new_n1593__;
  assign new_new_n1595__ = new_new_n1586__ & ~new_new_n1593__;
  assign new_new_n1596__ = ~new_new_n1594__ & ~new_new_n1595__;
  assign new_new_n1597__ = ~new_new_n1276__ & ~new_new_n1277__;
  assign new_new_n1598__ = new_new_n1284__ & ~new_new_n1597__;
  assign new_new_n1599__ = ~new_new_n1284__ & new_new_n1597__;
  assign new_new_n1600__ = ~new_new_n1598__ & ~new_new_n1599__;
  assign new_new_n1601__ = new_new_n1596__ & new_new_n1600__;
  assign new_new_n1602__ = ~new_new_n1596__ & ~new_new_n1600__;
  assign new_new_n1603__ = ~new_new_n1601__ & ~new_new_n1602__;
  assign new_new_n1604__ = new_new_n1525__ & new_new_n1603__;
  assign new_new_n1605__ = ~new_new_n1525__ & ~new_new_n1603__;
  assign new_new_n1606__ = ~new_new_n1338__ & ~new_new_n1339__;
  assign new_new_n1607__ = new_new_n1345__ & ~new_new_n1606__;
  assign new_new_n1608__ = ~new_new_n1345__ & new_new_n1606__;
  assign new_new_n1609__ = ~new_new_n1607__ & ~new_new_n1608__;
  assign new_new_n1610__ = ~new_new_n1605__ & new_new_n1609__;
  assign new_new_n1611__ = ~new_new_n1604__ & ~new_new_n1610__;
  assign new_new_n1612__ = ~new_new_n1518__ & ~new_new_n1519__;
  assign new_new_n1613__ = new_new_n1523__ & ~new_new_n1612__;
  assign new_new_n1614__ = ~new_new_n1523__ & new_new_n1612__;
  assign new_new_n1615__ = ~new_new_n1613__ & ~new_new_n1614__;
  assign new_new_n1616__ = ~new_new_n816__ & ~new_new_n1081__;
  assign new_new_n1617__ = new_new_n1499__ & new_new_n1616__;
  assign new_new_n1618__ = ~new_new_n1290__ & new_new_n1495__;
  assign new_new_n1619__ = new_new_n816__ & new_new_n1081__;
  assign new_new_n1620__ = new_new_n1326__ & new_new_n1619__;
  assign new_new_n1621__ = ~new_new_n1617__ & ~new_new_n1620__;
  assign new_new_n1622__ = ~new_new_n1618__ & new_new_n1621__;
  assign new_new_n1623__ = new_new_n760__ & ~new_new_n1411__;
  assign new_new_n1624__ = new_new_n686__ & new_new_n1324__;
  assign new_new_n1625__ = ~new_new_n686__ & ~new_new_n1324__;
  assign new_new_n1626__ = ~new_new_n1624__ & ~new_new_n1625__;
  assign new_new_n1627__ = new_new_n608__ & new_new_n1324__;
  assign new_new_n1628__ = ~new_new_n608__ & ~new_new_n1324__;
  assign new_new_n1629__ = ~new_new_n1627__ & ~new_new_n1628__;
  assign new_new_n1630__ = ~new_new_n760__ & new_new_n1626__;
  assign new_new_n1631__ = ~new_new_n1629__ & new_new_n1630__;
  assign new_new_n1632__ = ~new_new_n1623__ & ~new_new_n1631__;
  assign new_new_n1633__ = new_new_n1622__ & new_new_n1632__;
  assign new_new_n1634__ = ~new_new_n1622__ & ~new_new_n1632__;
  assign new_new_n1635__ = ~new_new_n1633__ & ~new_new_n1634__;
  assign new_new_n1636__ = new_new_n651__ & new_new_n1081__;
  assign new_new_n1637__ = ~new_new_n1481__ & ~new_new_n1636__;
  assign new_new_n1638__ = ~new_new_n1476__ & ~new_new_n1637__;
  assign new_new_n1639__ = new_new_n1476__ & new_new_n1557__;
  assign new_new_n1640__ = ~new_new_n1638__ & ~new_new_n1639__;
  assign new_new_n1641__ = new_new_n1635__ & ~new_new_n1640__;
  assign new_new_n1642__ = ~new_new_n1635__ & new_new_n1640__;
  assign new_new_n1643__ = ~new_new_n1641__ & ~new_new_n1642__;
  assign new_new_n1644__ = new_new_n824__ & ~new_new_n1300__;
  assign new_new_n1645__ = ~new_new_n308__ & ~new_new_n430__;
  assign new_new_n1646__ = new_new_n308__ & new_new_n430__;
  assign new_new_n1647__ = ~new_new_n1645__ & ~new_new_n1646__;
  assign new_new_n1648__ = ~new_new_n824__ & ~new_new_n1536__;
  assign new_new_n1649__ = new_new_n1647__ & new_new_n1648__;
  assign new_new_n1650__ = ~new_new_n1644__ & ~new_new_n1649__;
  assign new_new_n1651__ = ~new_new_n810__ & new_new_n1477__;
  assign new_new_n1652__ = ~new_new_n1476__ & ~new_new_n1559__;
  assign new_new_n1653__ = ~new_new_n1651__ & ~new_new_n1652__;
  assign new_new_n1654__ = ~new_new_n686__ & ~new_new_n758__;
  assign new_new_n1655__ = ~new_new_n759__ & new_new_n1573__;
  assign new_new_n1656__ = new_new_n1654__ & ~new_new_n1655__;
  assign new_new_n1657__ = ~new_new_n1653__ & new_new_n1656__;
  assign new_new_n1658__ = ~new_new_n1310__ & ~new_new_n1397__;
  assign new_new_n1659__ = new_new_n1226__ & ~new_new_n1658__;
  assign new_new_n1660__ = ~new_new_n301__ & new_new_n950__;
  assign new_new_n1661__ = new_new_n301__ & ~new_new_n950__;
  assign new_new_n1662__ = ~new_new_n1660__ & ~new_new_n1661__;
  assign new_new_n1663__ = ~new_new_n1226__ & new_new_n1547__;
  assign new_new_n1664__ = new_new_n1662__ & new_new_n1663__;
  assign new_new_n1665__ = ~new_new_n1659__ & ~new_new_n1664__;
  assign new_new_n1666__ = new_new_n1657__ & ~new_new_n1665__;
  assign new_new_n1667__ = ~new_new_n1657__ & new_new_n1665__;
  assign new_new_n1668__ = ~new_new_n1666__ & ~new_new_n1667__;
  assign new_new_n1669__ = new_new_n1650__ & ~new_new_n1668__;
  assign new_new_n1670__ = ~new_new_n1650__ & new_new_n1668__;
  assign new_new_n1671__ = ~new_new_n1669__ & ~new_new_n1670__;
  assign new_new_n1672__ = new_new_n1340__ & new_new_n1573__;
  assign new_new_n1673__ = new_new_n1495__ & new_new_n1529__;
  assign new_new_n1674__ = new_new_n615__ & ~new_new_n950__;
  assign new_new_n1675__ = ~new_new_n615__ & new_new_n950__;
  assign new_new_n1676__ = ~new_new_n1674__ & ~new_new_n1675__;
  assign new_new_n1677__ = new_new_n1560__ & new_new_n1676__;
  assign new_new_n1678__ = ~new_new_n1673__ & ~new_new_n1677__;
  assign new_new_n1679__ = new_new_n1226__ & new_new_n1547__;
  assign new_new_n1680__ = ~new_new_n1225__ & ~new_new_n1418__;
  assign new_new_n1681__ = ~new_new_n1008__ & ~new_new_n1419__;
  assign new_new_n1682__ = ~new_new_n1680__ & ~new_new_n1681__;
  assign new_new_n1683__ = ~new_new_n1679__ & ~new_new_n1682__;
  assign new_new_n1684__ = ~new_new_n1678__ & ~new_new_n1683__;
  assign new_new_n1685__ = new_new_n1678__ & new_new_n1683__;
  assign new_new_n1686__ = new_new_n824__ & ~new_new_n1536__;
  assign new_new_n1687__ = new_new_n310__ & new_new_n430__;
  assign new_new_n1688__ = ~new_new_n310__ & ~new_new_n430__;
  assign new_new_n1689__ = ~new_new_n1687__ & ~new_new_n1688__;
  assign new_new_n1690__ = ~new_new_n824__ & ~new_new_n1408__;
  assign new_new_n1691__ = new_new_n1689__ & new_new_n1690__;
  assign new_new_n1692__ = ~new_new_n1686__ & ~new_new_n1691__;
  assign new_new_n1693__ = ~new_new_n1685__ & ~new_new_n1692__;
  assign new_new_n1694__ = ~new_new_n1684__ & ~new_new_n1693__;
  assign new_new_n1695__ = ~new_new_n1672__ & new_new_n1694__;
  assign new_new_n1696__ = new_new_n1672__ & ~new_new_n1694__;
  assign new_new_n1697__ = ~new_new_n1695__ & ~new_new_n1696__;
  assign new_new_n1698__ = new_new_n1671__ & ~new_new_n1697__;
  assign new_new_n1699__ = ~new_new_n1671__ & new_new_n1697__;
  assign new_new_n1700__ = ~new_new_n1698__ & ~new_new_n1699__;
  assign new_new_n1701__ = new_new_n1643__ & ~new_new_n1700__;
  assign new_new_n1702__ = ~new_new_n1643__ & new_new_n1700__;
  assign new_new_n1703__ = new_new_n760__ & new_new_n1626__;
  assign new_new_n1704__ = new_new_n608__ & new_new_n1573__;
  assign new_new_n1705__ = new_new_n686__ & new_new_n1573__;
  assign new_new_n1706__ = ~new_new_n757__ & new_new_n1705__;
  assign new_new_n1707__ = ~new_new_n1238__ & ~new_new_n1706__;
  assign new_new_n1708__ = ~new_new_n1704__ & ~new_new_n1707__;
  assign new_new_n1709__ = ~new_new_n1703__ & ~new_new_n1708__;
  assign new_new_n1710__ = new_new_n1318__ & new_new_n1660__;
  assign new_new_n1711__ = new_new_n1495__ & new_new_n1676__;
  assign new_new_n1712__ = new_new_n1331__ & new_new_n1661__;
  assign new_new_n1713__ = ~new_new_n1710__ & ~new_new_n1712__;
  assign new_new_n1714__ = ~new_new_n1711__ & new_new_n1713__;
  assign new_new_n1715__ = new_new_n1226__ & ~new_new_n1420__;
  assign new_new_n1716__ = new_new_n308__ & new_new_n950__;
  assign new_new_n1717__ = ~new_new_n308__ & ~new_new_n950__;
  assign new_new_n1718__ = ~new_new_n1716__ & ~new_new_n1717__;
  assign new_new_n1719__ = ~new_new_n1226__ & ~new_new_n1647__;
  assign new_new_n1720__ = new_new_n1718__ & new_new_n1719__;
  assign new_new_n1721__ = ~new_new_n1715__ & ~new_new_n1720__;
  assign new_new_n1722__ = ~new_new_n1714__ & ~new_new_n1721__;
  assign new_new_n1723__ = new_new_n1714__ & new_new_n1721__;
  assign new_new_n1724__ = new_new_n816__ & ~new_new_n1081__;
  assign new_new_n1725__ = new_new_n1476__ & ~new_new_n1724__;
  assign new_new_n1726__ = new_new_n810__ & ~new_new_n1081__;
  assign new_new_n1727__ = ~new_new_n810__ & new_new_n1081__;
  assign new_new_n1728__ = ~new_new_n1726__ & ~new_new_n1727__;
  assign new_new_n1729__ = ~new_new_n1476__ & ~new_new_n1728__;
  assign new_new_n1730__ = ~new_new_n1725__ & ~new_new_n1729__;
  assign new_new_n1731__ = ~new_new_n1723__ & new_new_n1730__;
  assign new_new_n1732__ = ~new_new_n1722__ & ~new_new_n1731__;
  assign new_new_n1733__ = new_new_n1709__ & new_new_n1732__;
  assign new_new_n1734__ = ~new_new_n1709__ & ~new_new_n1732__;
  assign new_new_n1735__ = new_new_n1653__ & ~new_new_n1656__;
  assign new_new_n1736__ = ~new_new_n1657__ & ~new_new_n1735__;
  assign new_new_n1737__ = ~new_new_n1734__ & ~new_new_n1736__;
  assign new_new_n1738__ = ~new_new_n1733__ & ~new_new_n1737__;
  assign new_new_n1739__ = ~new_new_n1702__ & new_new_n1738__;
  assign new_new_n1740__ = ~new_new_n1701__ & ~new_new_n1739__;
  assign new_new_n1741__ = new_new_n1671__ & ~new_new_n1695__;
  assign new_new_n1742__ = ~new_new_n1696__ & ~new_new_n1741__;
  assign new_new_n1743__ = ~new_new_n1740__ & ~new_new_n1742__;
  assign new_new_n1744__ = new_new_n1740__ & new_new_n1742__;
  assign new_new_n1745__ = ~new_new_n950__ & new_new_n1331__;
  assign new_new_n1746__ = ~new_new_n810__ & new_new_n1745__;
  assign new_new_n1747__ = ~new_new_n1272__ & new_new_n1495__;
  assign new_new_n1748__ = new_new_n1288__ & new_new_n1318__;
  assign new_new_n1749__ = ~new_new_n1746__ & ~new_new_n1748__;
  assign new_new_n1750__ = ~new_new_n1747__ & new_new_n1749__;
  assign new_new_n1751__ = ~new_new_n1491__ & new_new_n1750__;
  assign new_new_n1752__ = new_new_n1491__ & ~new_new_n1750__;
  assign new_new_n1753__ = ~new_new_n1751__ & ~new_new_n1752__;
  assign new_new_n1754__ = new_new_n805__ & new_new_n1573__;
  assign new_new_n1755__ = new_new_n792__ & ~new_new_n1426__;
  assign new_new_n1756__ = ~new_new_n791__ & ~new_new_n1573__;
  assign new_new_n1757__ = ~new_new_n1754__ & ~new_new_n1756__;
  assign new_new_n1758__ = ~new_new_n1755__ & new_new_n1757__;
  assign new_new_n1759__ = new_new_n1753__ & new_new_n1758__;
  assign new_new_n1760__ = ~new_new_n1753__ & ~new_new_n1758__;
  assign new_new_n1761__ = ~new_new_n1759__ & ~new_new_n1760__;
  assign new_new_n1762__ = ~new_new_n1744__ & new_new_n1761__;
  assign new_new_n1763__ = ~new_new_n1633__ & ~new_new_n1640__;
  assign new_new_n1764__ = ~new_new_n1634__ & ~new_new_n1763__;
  assign new_new_n1765__ = new_new_n1650__ & new_new_n1665__;
  assign new_new_n1766__ = ~new_new_n1650__ & ~new_new_n1665__;
  assign new_new_n1767__ = ~new_new_n1657__ & ~new_new_n1766__;
  assign new_new_n1768__ = ~new_new_n1765__ & ~new_new_n1767__;
  assign new_new_n1769__ = ~new_new_n1764__ & new_new_n1768__;
  assign new_new_n1770__ = new_new_n1764__ & ~new_new_n1768__;
  assign new_new_n1771__ = ~new_new_n1769__ & ~new_new_n1770__;
  assign new_new_n1772__ = ~new_new_n1415__ & ~new_new_n1416__;
  assign new_new_n1773__ = ~new_new_n1423__ & new_new_n1772__;
  assign new_new_n1774__ = new_new_n1423__ & ~new_new_n1772__;
  assign new_new_n1775__ = ~new_new_n1773__ & ~new_new_n1774__;
  assign new_new_n1776__ = ~new_new_n1771__ & new_new_n1775__;
  assign new_new_n1777__ = new_new_n1771__ & ~new_new_n1775__;
  assign new_new_n1778__ = ~new_new_n1776__ & ~new_new_n1777__;
  assign new_new_n1779__ = ~new_new_n823__ & new_new_n1573__;
  assign new_new_n1780__ = new_new_n785__ & ~new_new_n1779__;
  assign new_new_n1781__ = ~new_new_n1616__ & ~new_new_n1780__;
  assign new_new_n1782__ = ~new_new_n1616__ & ~new_new_n1619__;
  assign new_new_n1783__ = new_new_n1780__ & ~new_new_n1782__;
  assign new_new_n1784__ = ~new_new_n1476__ & ~new_new_n1781__;
  assign new_new_n1785__ = ~new_new_n1783__ & new_new_n1784__;
  assign new_new_n1786__ = ~new_new_n615__ & ~new_new_n1081__;
  assign new_new_n1787__ = new_new_n1476__ & ~new_new_n1786__;
  assign new_new_n1788__ = ~new_new_n1619__ & ~new_new_n1787__;
  assign new_new_n1789__ = ~new_new_n1780__ & ~new_new_n1788__;
  assign new_new_n1790__ = ~new_new_n615__ & new_new_n1477__;
  assign new_new_n1791__ = new_new_n1780__ & new_new_n1790__;
  assign new_new_n1792__ = ~new_new_n1789__ & ~new_new_n1791__;
  assign new_new_n1793__ = ~new_new_n1785__ & new_new_n1792__;
  assign new_new_n1794__ = new_new_n1780__ & ~new_new_n1793__;
  assign new_new_n1795__ = new_new_n824__ & ~new_new_n1408__;
  assign new_new_n1796__ = new_new_n430__ & new_new_n1324__;
  assign new_new_n1797__ = ~new_new_n430__ & ~new_new_n1324__;
  assign new_new_n1798__ = ~new_new_n1796__ & ~new_new_n1797__;
  assign new_new_n1799__ = ~new_new_n824__ & new_new_n1629__;
  assign new_new_n1800__ = ~new_new_n1798__ & new_new_n1799__;
  assign new_new_n1801__ = ~new_new_n1795__ & ~new_new_n1800__;
  assign new_new_n1802__ = ~new_new_n1794__ & new_new_n1801__;
  assign new_new_n1803__ = new_new_n1226__ & ~new_new_n1647__;
  assign new_new_n1804__ = ~new_new_n1225__ & ~new_new_n1687__;
  assign new_new_n1805__ = ~new_new_n1008__ & ~new_new_n1688__;
  assign new_new_n1806__ = ~new_new_n1804__ & ~new_new_n1805__;
  assign new_new_n1807__ = ~new_new_n1803__ & ~new_new_n1806__;
  assign new_new_n1808__ = new_new_n1495__ & ~new_new_n1662__;
  assign new_new_n1809__ = new_new_n316__ & new_new_n950__;
  assign new_new_n1810__ = ~new_new_n316__ & ~new_new_n950__;
  assign new_new_n1811__ = ~new_new_n1809__ & ~new_new_n1810__;
  assign new_new_n1812__ = ~new_new_n1500__ & new_new_n1503__;
  assign new_new_n1813__ = ~new_new_n1811__ & new_new_n1812__;
  assign new_new_n1814__ = ~new_new_n1808__ & ~new_new_n1813__;
  assign new_new_n1815__ = ~new_new_n1807__ & ~new_new_n1814__;
  assign new_new_n1816__ = new_new_n1807__ & new_new_n1814__;
  assign new_new_n1817__ = new_new_n784__ & new_new_n1704__;
  assign new_new_n1818__ = new_new_n824__ & new_new_n1629__;
  assign new_new_n1819__ = ~new_new_n608__ & ~new_new_n1573__;
  assign new_new_n1820__ = new_new_n823__ & new_new_n1819__;
  assign new_new_n1821__ = ~new_new_n1817__ & ~new_new_n1820__;
  assign new_new_n1822__ = ~new_new_n1818__ & new_new_n1821__;
  assign new_new_n1823__ = ~new_new_n1816__ & ~new_new_n1822__;
  assign new_new_n1824__ = ~new_new_n1815__ & ~new_new_n1823__;
  assign new_new_n1825__ = ~new_new_n1722__ & ~new_new_n1723__;
  assign new_new_n1826__ = new_new_n810__ & new_new_n1563__;
  assign new_new_n1827__ = ~new_new_n1725__ & ~new_new_n1727__;
  assign new_new_n1828__ = ~new_new_n1826__ & new_new_n1827__;
  assign new_new_n1829__ = ~new_new_n1825__ & ~new_new_n1828__;
  assign new_new_n1830__ = new_new_n1730__ & new_new_n1825__;
  assign new_new_n1831__ = ~new_new_n1829__ & ~new_new_n1830__;
  assign new_new_n1832__ = new_new_n1824__ & ~new_new_n1831__;
  assign new_new_n1833__ = new_new_n1802__ & new_new_n1832__;
  assign new_new_n1834__ = new_new_n1794__ & ~new_new_n1801__;
  assign new_new_n1835__ = new_new_n1832__ & ~new_new_n1834__;
  assign new_new_n1836__ = ~new_new_n1824__ & new_new_n1831__;
  assign new_new_n1837__ = new_new_n1802__ & ~new_new_n1836__;
  assign new_new_n1838__ = ~new_new_n1835__ & ~new_new_n1837__;
  assign new_new_n1839__ = ~new_new_n758__ & new_new_n1655__;
  assign new_new_n1840__ = ~new_new_n1838__ & ~new_new_n1839__;
  assign new_new_n1841__ = ~new_new_n1833__ & ~new_new_n1840__;
  assign new_new_n1842__ = ~new_new_n1684__ & ~new_new_n1685__;
  assign new_new_n1843__ = new_new_n1692__ & ~new_new_n1842__;
  assign new_new_n1844__ = ~new_new_n1692__ & new_new_n1842__;
  assign new_new_n1845__ = ~new_new_n1843__ & ~new_new_n1844__;
  assign new_new_n1846__ = new_new_n1841__ & new_new_n1845__;
  assign new_new_n1847__ = ~new_new_n1802__ & new_new_n1839__;
  assign new_new_n1848__ = new_new_n1836__ & new_new_n1847__;
  assign new_new_n1849__ = ~new_new_n1836__ & ~new_new_n1839__;
  assign new_new_n1850__ = ~new_new_n1832__ & new_new_n1834__;
  assign new_new_n1851__ = ~new_new_n1849__ & new_new_n1850__;
  assign new_new_n1852__ = ~new_new_n1848__ & ~new_new_n1851__;
  assign new_new_n1853__ = ~new_new_n1733__ & ~new_new_n1734__;
  assign new_new_n1854__ = ~new_new_n1736__ & new_new_n1853__;
  assign new_new_n1855__ = new_new_n1736__ & ~new_new_n1853__;
  assign new_new_n1856__ = ~new_new_n1854__ & ~new_new_n1855__;
  assign new_new_n1857__ = ~new_new_n1802__ & ~new_new_n1834__;
  assign new_new_n1858__ = ~new_new_n1832__ & ~new_new_n1836__;
  assign new_new_n1859__ = new_new_n1857__ & ~new_new_n1858__;
  assign new_new_n1860__ = ~new_new_n1857__ & new_new_n1858__;
  assign new_new_n1861__ = ~new_new_n1859__ & ~new_new_n1860__;
  assign new_new_n1862__ = new_new_n1839__ & new_new_n1861__;
  assign new_new_n1863__ = ~new_new_n1839__ & ~new_new_n1861__;
  assign new_new_n1864__ = ~new_new_n1862__ & ~new_new_n1863__;
  assign new_new_n1865__ = ~new_new_n1815__ & ~new_new_n1816__;
  assign new_new_n1866__ = new_new_n1822__ & ~new_new_n1865__;
  assign new_new_n1867__ = ~new_new_n1822__ & new_new_n1865__;
  assign new_new_n1868__ = ~new_new_n1866__ & ~new_new_n1867__;
  assign new_new_n1869__ = new_new_n1318__ & new_new_n1716__;
  assign new_new_n1870__ = new_new_n1495__ & ~new_new_n1811__;
  assign new_new_n1871__ = new_new_n1331__ & new_new_n1717__;
  assign new_new_n1872__ = ~new_new_n1869__ & ~new_new_n1871__;
  assign new_new_n1873__ = ~new_new_n1870__ & new_new_n1872__;
  assign new_new_n1874__ = new_new_n1226__ & ~new_new_n1689__;
  assign new_new_n1875__ = new_new_n950__ & ~new_new_n1324__;
  assign new_new_n1876__ = ~new_new_n950__ & new_new_n1324__;
  assign new_new_n1877__ = ~new_new_n1875__ & ~new_new_n1876__;
  assign new_new_n1878__ = ~new_new_n1226__ & new_new_n1798__;
  assign new_new_n1879__ = new_new_n1877__ & new_new_n1878__;
  assign new_new_n1880__ = ~new_new_n1874__ & ~new_new_n1879__;
  assign new_new_n1881__ = ~new_new_n1873__ & ~new_new_n1880__;
  assign new_new_n1882__ = new_new_n1873__ & new_new_n1880__;
  assign new_new_n1883__ = new_new_n301__ & ~new_new_n1081__;
  assign new_new_n1884__ = new_new_n1476__ & ~new_new_n1883__;
  assign new_new_n1885__ = new_new_n615__ & new_new_n1081__;
  assign new_new_n1886__ = ~new_new_n1476__ & ~new_new_n1786__;
  assign new_new_n1887__ = ~new_new_n1885__ & new_new_n1886__;
  assign new_new_n1888__ = ~new_new_n1884__ & ~new_new_n1887__;
  assign new_new_n1889__ = ~new_new_n1882__ & new_new_n1888__;
  assign new_new_n1890__ = ~new_new_n1881__ & ~new_new_n1889__;
  assign new_new_n1891__ = new_new_n1868__ & ~new_new_n1890__;
  assign new_new_n1892__ = ~new_new_n1868__ & new_new_n1890__;
  assign new_new_n1893__ = new_new_n1793__ & ~new_new_n1892__;
  assign new_new_n1894__ = ~new_new_n1891__ & ~new_new_n1893__;
  assign new_new_n1895__ = ~new_new_n1864__ & ~new_new_n1894__;
  assign new_new_n1896__ = ~new_new_n301__ & new_new_n1081__;
  assign new_new_n1897__ = ~new_new_n1883__ & ~new_new_n1896__;
  assign new_new_n1898__ = new_new_n299__ & ~new_new_n1065__;
  assign new_new_n1899__ = ~new_new_n1897__ & ~new_new_n1898__;
  assign new_new_n1900__ = ~new_new_n1476__ & ~new_new_n1899__;
  assign new_new_n1901__ = ~new_new_n316__ & ~new_new_n1081__;
  assign new_new_n1902__ = new_new_n1476__ & ~new_new_n1901__;
  assign new_new_n1903__ = ~new_new_n1900__ & ~new_new_n1902__;
  assign new_new_n1904__ = new_new_n824__ & new_new_n1573__;
  assign new_new_n1905__ = new_new_n1226__ & new_new_n1798__;
  assign new_new_n1906__ = ~new_new_n430__ & ~new_new_n1573__;
  assign new_new_n1907__ = new_new_n1225__ & new_new_n1906__;
  assign new_new_n1908__ = new_new_n1175__ & new_new_n1573__;
  assign new_new_n1909__ = ~new_new_n1905__ & ~new_new_n1907__;
  assign new_new_n1910__ = ~new_new_n1908__ & new_new_n1909__;
  assign new_new_n1911__ = new_new_n1495__ & ~new_new_n1718__;
  assign new_new_n1912__ = ~new_new_n310__ & new_new_n1745__;
  assign new_new_n1913__ = new_new_n310__ & new_new_n1319__;
  assign new_new_n1914__ = ~new_new_n1911__ & ~new_new_n1912__;
  assign new_new_n1915__ = ~new_new_n1913__ & new_new_n1914__;
  assign new_new_n1916__ = new_new_n1910__ & new_new_n1915__;
  assign new_new_n1917__ = new_new_n1226__ & new_new_n1573__;
  assign new_new_n1918__ = new_new_n1009__ & ~new_new_n1917__;
  assign new_new_n1919__ = new_new_n1916__ & ~new_new_n1918__;
  assign new_new_n1920__ = new_new_n1904__ & ~new_new_n1919__;
  assign new_new_n1921__ = ~new_new_n1910__ & ~new_new_n1915__;
  assign new_new_n1922__ = new_new_n1918__ & new_new_n1921__;
  assign new_new_n1923__ = ~new_new_n1920__ & ~new_new_n1922__;
  assign new_new_n1924__ = new_new_n1903__ & ~new_new_n1923__;
  assign new_new_n1925__ = ~new_new_n1915__ & new_new_n1918__;
  assign new_new_n1926__ = ~new_new_n1921__ & ~new_new_n1925__;
  assign new_new_n1927__ = new_new_n1904__ & ~new_new_n1926__;
  assign new_new_n1928__ = ~new_new_n1924__ & ~new_new_n1927__;
  assign new_new_n1929__ = ~new_new_n1916__ & ~new_new_n1921__;
  assign new_new_n1930__ = new_new_n1903__ & new_new_n1918__;
  assign new_new_n1931__ = ~new_new_n1903__ & ~new_new_n1918__;
  assign new_new_n1932__ = ~new_new_n1930__ & ~new_new_n1931__;
  assign new_new_n1933__ = new_new_n1929__ & ~new_new_n1932__;
  assign new_new_n1934__ = ~new_new_n1929__ & new_new_n1932__;
  assign new_new_n1935__ = ~new_new_n1933__ & ~new_new_n1934__;
  assign new_new_n1936__ = pi06 & new_new_n1081__;
  assign new_new_n1937__ = new_new_n304__ & new_new_n1936__;
  assign new_new_n1938__ = ~pi06 & ~new_new_n1081__;
  assign new_new_n1939__ = ~new_new_n1936__ & ~new_new_n1938__;
  assign new_new_n1940__ = new_new_n305__ & new_new_n1939__;
  assign new_new_n1941__ = pi22 & ~new_new_n1939__;
  assign new_new_n1942__ = ~new_new_n1937__ & ~new_new_n1940__;
  assign new_new_n1943__ = ~new_new_n1941__ & new_new_n1942__;
  assign new_new_n1944__ = ~new_new_n1476__ & ~new_new_n1943__;
  assign new_new_n1945__ = ~new_new_n56__ & ~new_new_n1476__;
  assign new_new_n1946__ = ~new_new_n310__ & ~new_new_n1081__;
  assign new_new_n1947__ = ~new_new_n1945__ & new_new_n1946__;
  assign new_new_n1948__ = ~new_new_n1944__ & ~new_new_n1947__;
  assign new_new_n1949__ = ~new_new_n1917__ & new_new_n1948__;
  assign new_new_n1950__ = ~new_new_n308__ & new_new_n1477__;
  assign new_new_n1951__ = new_new_n316__ & new_new_n1081__;
  assign new_new_n1952__ = ~new_new_n1901__ & ~new_new_n1951__;
  assign new_new_n1953__ = ~new_new_n1476__ & ~new_new_n1952__;
  assign new_new_n1954__ = ~new_new_n1950__ & ~new_new_n1953__;
  assign new_new_n1955__ = ~new_new_n1331__ & new_new_n1954__;
  assign new_new_n1956__ = ~new_new_n950__ & ~new_new_n1955__;
  assign new_new_n1957__ = new_new_n1495__ & ~new_new_n1954__;
  assign new_new_n1958__ = new_new_n950__ & ~new_new_n1957__;
  assign new_new_n1959__ = new_new_n310__ & ~new_new_n1956__;
  assign new_new_n1960__ = ~new_new_n1958__ & new_new_n1959__;
  assign new_new_n1961__ = new_new_n310__ & ~new_new_n1331__;
  assign new_new_n1962__ = new_new_n950__ & ~new_new_n1961__;
  assign new_new_n1963__ = ~new_new_n1318__ & ~new_new_n1962__;
  assign new_new_n1964__ = new_new_n1318__ & new_new_n1875__;
  assign new_new_n1965__ = new_new_n1954__ & ~new_new_n1964__;
  assign new_new_n1966__ = ~new_new_n1963__ & new_new_n1965__;
  assign new_new_n1967__ = new_new_n1147__ & new_new_n1324__;
  assign new_new_n1968__ = ~new_new_n1495__ & ~new_new_n1967__;
  assign new_new_n1969__ = ~new_new_n950__ & ~new_new_n1961__;
  assign new_new_n1970__ = ~new_new_n1968__ & new_new_n1969__;
  assign new_new_n1971__ = ~new_new_n1954__ & new_new_n1970__;
  assign new_new_n1972__ = ~new_new_n1319__ & ~new_new_n1954__;
  assign new_new_n1973__ = ~new_new_n1324__ & ~new_new_n1955__;
  assign new_new_n1974__ = ~new_new_n1972__ & new_new_n1973__;
  assign new_new_n1975__ = ~new_new_n1966__ & ~new_new_n1971__;
  assign new_new_n1976__ = ~new_new_n1974__ & new_new_n1975__;
  assign new_new_n1977__ = ~new_new_n1960__ & new_new_n1976__;
  assign new_new_n1978__ = new_new_n1495__ & ~new_new_n1877__;
  assign new_new_n1979__ = ~new_new_n1573__ & new_new_n1745__;
  assign new_new_n1980__ = new_new_n1319__ & new_new_n1573__;
  assign new_new_n1981__ = ~new_new_n1978__ & ~new_new_n1979__;
  assign new_new_n1982__ = ~new_new_n1980__ & new_new_n1981__;
  assign new_new_n1983__ = ~new_new_n1977__ & new_new_n1982__;
  assign new_new_n1984__ = ~new_new_n1949__ & ~new_new_n1983__;
  assign new_new_n1985__ = ~new_new_n1331__ & new_new_n1573__;
  assign new_new_n1986__ = ~new_new_n950__ & ~new_new_n1318__;
  assign new_new_n1987__ = ~new_new_n1985__ & new_new_n1986__;
  assign new_new_n1988__ = ~new_new_n1984__ & ~new_new_n1987__;
  assign new_new_n1989__ = new_new_n1948__ & ~new_new_n1977__;
  assign new_new_n1990__ = new_new_n1977__ & ~new_new_n1982__;
  assign new_new_n1991__ = ~new_new_n1917__ & ~new_new_n1990__;
  assign new_new_n1992__ = ~new_new_n1989__ & ~new_new_n1991__;
  assign new_new_n1993__ = ~new_new_n1988__ & new_new_n1992__;
  assign new_new_n1994__ = ~new_new_n1147__ & new_new_n1573__;
  assign new_new_n1995__ = ~new_new_n1476__ & new_new_n1573__;
  assign new_new_n1996__ = ~new_new_n1324__ & ~new_new_n1995__;
  assign new_new_n1997__ = new_new_n310__ & ~new_new_n1476__;
  assign new_new_n1998__ = ~new_new_n1081__ & ~new_new_n1997__;
  assign new_new_n1999__ = ~new_new_n1994__ & new_new_n1998__;
  assign new_new_n2000__ = ~new_new_n1996__ & new_new_n1999__;
  assign new_new_n2001__ = new_new_n1081__ & new_new_n1997__;
  assign new_new_n2002__ = new_new_n1994__ & new_new_n2001__;
  assign new_new_n2003__ = ~new_new_n2000__ & ~new_new_n2002__;
  assign new_new_n2004__ = ~new_new_n1993__ & new_new_n2003__;
  assign new_new_n2005__ = ~new_new_n1983__ & ~new_new_n1991__;
  assign new_new_n2006__ = new_new_n1948__ & ~new_new_n2005__;
  assign new_new_n2007__ = ~new_new_n1917__ & ~new_new_n1987__;
  assign new_new_n2008__ = ~new_new_n1977__ & new_new_n2007__;
  assign new_new_n2009__ = ~new_new_n2006__ & ~new_new_n2008__;
  assign new_new_n2010__ = ~new_new_n2004__ & new_new_n2009__;
  assign new_new_n2011__ = ~new_new_n1954__ & ~new_new_n1977__;
  assign new_new_n2012__ = ~new_new_n2010__ & new_new_n2011__;
  assign new_new_n2013__ = ~new_new_n1948__ & new_new_n1987__;
  assign new_new_n2014__ = new_new_n1977__ & new_new_n2013__;
  assign new_new_n2015__ = ~new_new_n2012__ & ~new_new_n2014__;
  assign new_new_n2016__ = ~new_new_n1935__ & ~new_new_n2015__;
  assign new_new_n2017__ = new_new_n1935__ & ~new_new_n2011__;
  assign new_new_n2018__ = new_new_n1987__ & new_new_n1989__;
  assign new_new_n2019__ = ~new_new_n2017__ & ~new_new_n2018__;
  assign new_new_n2020__ = new_new_n2010__ & new_new_n2019__;
  assign new_new_n2021__ = ~new_new_n2016__ & ~new_new_n2020__;
  assign new_new_n2022__ = new_new_n1904__ & ~new_new_n1918__;
  assign new_new_n2023__ = new_new_n1903__ & ~new_new_n1915__;
  assign new_new_n2024__ = new_new_n2022__ & ~new_new_n2023__;
  assign new_new_n2025__ = ~new_new_n1925__ & ~new_new_n1930__;
  assign new_new_n2026__ = ~new_new_n2023__ & new_new_n2025__;
  assign new_new_n2027__ = ~new_new_n1904__ & ~new_new_n2026__;
  assign new_new_n2028__ = ~new_new_n2024__ & ~new_new_n2027__;
  assign new_new_n2029__ = new_new_n1910__ & ~new_new_n2028__;
  assign new_new_n2030__ = ~new_new_n1910__ & new_new_n1918__;
  assign new_new_n2031__ = new_new_n1904__ & new_new_n1915__;
  assign new_new_n2032__ = ~new_new_n2030__ & ~new_new_n2031__;
  assign new_new_n2033__ = ~new_new_n1903__ & ~new_new_n2032__;
  assign new_new_n2034__ = new_new_n1915__ & new_new_n1931__;
  assign new_new_n2035__ = ~new_new_n1910__ & ~new_new_n2022__;
  assign new_new_n2036__ = ~new_new_n1925__ & new_new_n2035__;
  assign new_new_n2037__ = ~new_new_n2034__ & new_new_n2036__;
  assign new_new_n2038__ = ~new_new_n2033__ & ~new_new_n2037__;
  assign new_new_n2039__ = ~new_new_n2029__ & new_new_n2038__;
  assign new_new_n2040__ = ~new_new_n1881__ & ~new_new_n1882__;
  assign new_new_n2041__ = ~new_new_n1477__ & ~new_new_n1786__;
  assign new_new_n2042__ = ~new_new_n1885__ & new_new_n2041__;
  assign new_new_n2043__ = ~new_new_n1884__ & ~new_new_n2042__;
  assign new_new_n2044__ = new_new_n2040__ & ~new_new_n2043__;
  assign new_new_n2045__ = new_new_n1888__ & ~new_new_n2040__;
  assign new_new_n2046__ = ~new_new_n2044__ & ~new_new_n2045__;
  assign new_new_n2047__ = new_new_n2039__ & new_new_n2046__;
  assign new_new_n2048__ = ~new_new_n2021__ & ~new_new_n2047__;
  assign new_new_n2049__ = ~new_new_n2039__ & ~new_new_n2046__;
  assign new_new_n2050__ = ~new_new_n2048__ & ~new_new_n2049__;
  assign new_new_n2051__ = new_new_n1928__ & new_new_n2050__;
  assign new_new_n2052__ = new_new_n1864__ & ~new_new_n1891__;
  assign new_new_n2053__ = new_new_n1793__ & ~new_new_n2052__;
  assign new_new_n2054__ = ~new_new_n1864__ & ~new_new_n1892__;
  assign new_new_n2055__ = ~new_new_n2053__ & ~new_new_n2054__;
  assign new_new_n2056__ = ~new_new_n2051__ & ~new_new_n2055__;
  assign new_new_n2057__ = new_new_n1864__ & new_new_n1894__;
  assign new_new_n2058__ = ~new_new_n1928__ & ~new_new_n2057__;
  assign new_new_n2059__ = ~new_new_n2050__ & new_new_n2058__;
  assign new_new_n2060__ = ~new_new_n1895__ & ~new_new_n2059__;
  assign new_new_n2061__ = ~new_new_n2056__ & new_new_n2060__;
  assign new_new_n2062__ = new_new_n1856__ & new_new_n2061__;
  assign new_new_n2063__ = ~new_new_n1701__ & ~new_new_n1702__;
  assign new_new_n2064__ = new_new_n1738__ & ~new_new_n2063__;
  assign new_new_n2065__ = ~new_new_n1738__ & new_new_n2063__;
  assign new_new_n2066__ = ~new_new_n2064__ & ~new_new_n2065__;
  assign new_new_n2067__ = ~new_new_n2062__ & ~new_new_n2066__;
  assign new_new_n2068__ = ~new_new_n1846__ & new_new_n1852__;
  assign new_new_n2069__ = ~new_new_n2067__ & new_new_n2068__;
  assign new_new_n2070__ = ~new_new_n1856__ & ~new_new_n2061__;
  assign new_new_n2071__ = new_new_n1845__ & ~new_new_n1852__;
  assign new_new_n2072__ = new_new_n2066__ & ~new_new_n2071__;
  assign new_new_n2073__ = ~new_new_n1845__ & new_new_n1852__;
  assign new_new_n2074__ = ~new_new_n1841__ & new_new_n2073__;
  assign new_new_n2075__ = ~new_new_n2072__ & ~new_new_n2074__;
  assign new_new_n2076__ = ~new_new_n2070__ & ~new_new_n2075__;
  assign new_new_n2077__ = new_new_n2062__ & new_new_n2066__;
  assign new_new_n2078__ = ~new_new_n2076__ & ~new_new_n2077__;
  assign new_new_n2079__ = ~new_new_n2069__ & new_new_n2078__;
  assign new_new_n2080__ = new_new_n1778__ & ~new_new_n2079__;
  assign new_new_n2081__ = ~new_new_n1769__ & ~new_new_n1775__;
  assign new_new_n2082__ = ~new_new_n1770__ & ~new_new_n2081__;
  assign new_new_n2083__ = ~new_new_n1566__ & ~new_new_n1567__;
  assign new_new_n2084__ = new_new_n1574__ & ~new_new_n2083__;
  assign new_new_n2085__ = ~new_new_n1574__ & new_new_n2083__;
  assign new_new_n2086__ = ~new_new_n2084__ & ~new_new_n2085__;
  assign new_new_n2087__ = ~new_new_n1540__ & ~new_new_n1541__;
  assign new_new_n2088__ = new_new_n1550__ & ~new_new_n2087__;
  assign new_new_n2089__ = ~new_new_n1550__ & new_new_n2087__;
  assign new_new_n2090__ = ~new_new_n2088__ & ~new_new_n2089__;
  assign new_new_n2091__ = new_new_n2086__ & ~new_new_n2090__;
  assign new_new_n2092__ = ~new_new_n2086__ & new_new_n2090__;
  assign new_new_n2093__ = ~new_new_n2091__ & ~new_new_n2092__;
  assign new_new_n2094__ = ~new_new_n1751__ & new_new_n1758__;
  assign new_new_n2095__ = ~new_new_n1752__ & ~new_new_n2094__;
  assign new_new_n2096__ = new_new_n2093__ & new_new_n2095__;
  assign new_new_n2097__ = ~new_new_n2093__ & ~new_new_n2095__;
  assign new_new_n2098__ = ~new_new_n2096__ & ~new_new_n2097__;
  assign new_new_n2099__ = ~new_new_n2082__ & new_new_n2098__;
  assign new_new_n2100__ = new_new_n2082__ & ~new_new_n2098__;
  assign new_new_n2101__ = ~new_new_n2099__ & ~new_new_n2100__;
  assign new_new_n2102__ = ~new_new_n1432__ & ~new_new_n1433__;
  assign new_new_n2103__ = ~new_new_n1492__ & new_new_n2102__;
  assign new_new_n2104__ = new_new_n1492__ & ~new_new_n2102__;
  assign new_new_n2105__ = ~new_new_n2103__ & ~new_new_n2104__;
  assign new_new_n2106__ = new_new_n2101__ & ~new_new_n2105__;
  assign new_new_n2107__ = ~new_new_n2101__ & new_new_n2105__;
  assign new_new_n2108__ = ~new_new_n2106__ & ~new_new_n2107__;
  assign new_new_n2109__ = ~new_new_n2080__ & new_new_n2108__;
  assign new_new_n2110__ = ~new_new_n1743__ & ~new_new_n1762__;
  assign new_new_n2111__ = ~new_new_n2109__ & new_new_n2110__;
  assign new_new_n2112__ = ~new_new_n1778__ & new_new_n2079__;
  assign new_new_n2113__ = new_new_n1744__ & ~new_new_n1761__;
  assign new_new_n2114__ = new_new_n2108__ & ~new_new_n2113__;
  assign new_new_n2115__ = new_new_n1743__ & new_new_n1761__;
  assign new_new_n2116__ = ~new_new_n2114__ & ~new_new_n2115__;
  assign new_new_n2117__ = ~new_new_n2112__ & new_new_n2116__;
  assign new_new_n2118__ = new_new_n2080__ & ~new_new_n2108__;
  assign new_new_n2119__ = ~new_new_n2117__ & ~new_new_n2118__;
  assign new_new_n2120__ = ~new_new_n2111__ & new_new_n2119__;
  assign new_new_n2121__ = ~new_new_n1615__ & new_new_n2120__;
  assign new_new_n2122__ = ~new_new_n2091__ & ~new_new_n2095__;
  assign new_new_n2123__ = ~new_new_n2092__ & ~new_new_n2122__;
  assign new_new_n2124__ = ~new_new_n2099__ & ~new_new_n2105__;
  assign new_new_n2125__ = ~new_new_n2100__ & ~new_new_n2124__;
  assign new_new_n2126__ = ~new_new_n2123__ & ~new_new_n2125__;
  assign new_new_n2127__ = ~new_new_n1604__ & ~new_new_n1605__;
  assign new_new_n2128__ = new_new_n1609__ & new_new_n2127__;
  assign new_new_n2129__ = ~new_new_n1609__ & ~new_new_n2127__;
  assign new_new_n2130__ = ~new_new_n2128__ & ~new_new_n2129__;
  assign new_new_n2131__ = ~new_new_n2126__ & ~new_new_n2130__;
  assign new_new_n2132__ = ~new_new_n1579__ & new_new_n1584__;
  assign new_new_n2133__ = ~new_new_n1585__ & ~new_new_n2132__;
  assign new_new_n2134__ = ~new_new_n2131__ & new_new_n2133__;
  assign new_new_n2135__ = ~new_new_n2121__ & ~new_new_n2134__;
  assign new_new_n2136__ = new_new_n2123__ & new_new_n2125__;
  assign new_new_n2137__ = new_new_n2135__ & new_new_n2136__;
  assign new_new_n2138__ = new_new_n1615__ & ~new_new_n2120__;
  assign new_new_n2139__ = ~new_new_n2135__ & ~new_new_n2138__;
  assign new_new_n2140__ = ~new_new_n2130__ & ~new_new_n2139__;
  assign new_new_n2141__ = new_new_n2133__ & ~new_new_n2136__;
  assign new_new_n2142__ = new_new_n2130__ & ~new_new_n2138__;
  assign new_new_n2143__ = ~new_new_n2126__ & ~new_new_n2141__;
  assign new_new_n2144__ = ~new_new_n2142__ & new_new_n2143__;
  assign new_new_n2145__ = ~new_new_n2137__ & ~new_new_n2144__;
  assign new_new_n2146__ = ~new_new_n2140__ & new_new_n2145__;
  assign new_new_n2147__ = new_new_n1611__ & ~new_new_n2146__;
  assign new_new_n2148__ = ~new_new_n1594__ & ~new_new_n1600__;
  assign new_new_n2149__ = ~new_new_n1595__ & ~new_new_n2148__;
  assign new_new_n2150__ = ~new_new_n1348__ & ~new_new_n1349__;
  assign new_new_n2151__ = ~new_new_n1353__ & new_new_n2150__;
  assign new_new_n2152__ = new_new_n1353__ & ~new_new_n2150__;
  assign new_new_n2153__ = ~new_new_n2151__ & ~new_new_n2152__;
  assign new_new_n2154__ = new_new_n2149__ & new_new_n2153__;
  assign new_new_n2155__ = ~new_new_n2149__ & ~new_new_n2153__;
  assign new_new_n2156__ = ~new_new_n1371__ & ~new_new_n1375__;
  assign new_new_n2157__ = new_new_n1364__ & ~new_new_n1496__;
  assign new_new_n2158__ = ~new_new_n1148__ & ~new_new_n2157__;
  assign new_new_n2159__ = new_new_n2156__ & new_new_n2158__;
  assign new_new_n2160__ = ~new_new_n2156__ & ~new_new_n2158__;
  assign new_new_n2161__ = ~new_new_n2159__ & ~new_new_n2160__;
  assign new_new_n2162__ = ~new_new_n2155__ & ~new_new_n2161__;
  assign new_new_n2163__ = ~new_new_n2154__ & ~new_new_n2162__;
  assign new_new_n2164__ = ~new_new_n2147__ & ~new_new_n2163__;
  assign new_new_n2165__ = ~new_new_n1382__ & ~new_new_n1390__;
  assign new_new_n2166__ = ~new_new_n1385__ & new_new_n2165__;
  assign new_new_n2167__ = new_new_n1385__ & ~new_new_n2165__;
  assign new_new_n2168__ = ~new_new_n2166__ & ~new_new_n2167__;
  assign new_new_n2169__ = new_new_n1388__ & new_new_n2168__;
  assign new_new_n2170__ = ~new_new_n1388__ & ~new_new_n2168__;
  assign new_new_n2171__ = ~new_new_n2169__ & ~new_new_n2170__;
  assign new_new_n2172__ = ~new_new_n2164__ & ~new_new_n2171__;
  assign new_new_n2173__ = ~new_new_n1611__ & new_new_n2146__;
  assign new_new_n2174__ = new_new_n2155__ & new_new_n2161__;
  assign new_new_n2175__ = new_new_n2154__ & ~new_new_n2161__;
  assign new_new_n2176__ = ~new_new_n2171__ & ~new_new_n2175__;
  assign new_new_n2177__ = ~new_new_n2174__ & ~new_new_n2176__;
  assign new_new_n2178__ = ~new_new_n2173__ & ~new_new_n2177__;
  assign new_new_n2179__ = new_new_n2147__ & new_new_n2163__;
  assign new_new_n2180__ = ~new_new_n2178__ & ~new_new_n2179__;
  assign new_new_n2181__ = ~new_new_n2172__ & new_new_n2180__;
  assign new_new_n2182__ = new_new_n1395__ & new_new_n2181__;
  assign new_new_n2183__ = new_new_n1256__ & new_new_n2182__;
  assign new_new_n2184__ = new_new_n1211__ & new_new_n1394__;
  assign new_new_n2185__ = new_new_n2181__ & ~new_new_n2184__;
  assign new_new_n2186__ = ~new_new_n1395__ & ~new_new_n2185__;
  assign new_new_n2187__ = ~new_new_n1256__ & new_new_n2186__;
  assign new_new_n2188__ = ~new_new_n2181__ & new_new_n2184__;
  assign new_new_n2189__ = ~new_new_n2187__ & ~new_new_n2188__;
  assign new_new_n2190__ = ~new_new_n846__ & ~new_new_n847__;
  assign new_new_n2191__ = ~new_new_n853__ & new_new_n2190__;
  assign new_new_n2192__ = new_new_n853__ & ~new_new_n2190__;
  assign new_new_n2193__ = ~new_new_n2191__ & ~new_new_n2192__;
  assign new_new_n2194__ = ~new_new_n2189__ & new_new_n2193__;
  assign new_new_n2195__ = ~new_new_n1256__ & ~new_new_n2182__;
  assign new_new_n2196__ = ~new_new_n2186__ & ~new_new_n2193__;
  assign new_new_n2197__ = ~new_new_n2195__ & new_new_n2196__;
  assign new_new_n2198__ = ~new_new_n1256__ & ~new_new_n2181__;
  assign new_new_n2199__ = new_new_n2184__ & new_new_n2198__;
  assign new_new_n2200__ = ~new_new_n2183__ & ~new_new_n2199__;
  assign new_new_n2201__ = ~new_new_n2197__ & new_new_n2200__;
  assign new_new_n2202__ = ~new_new_n2194__ & new_new_n2201__;
  assign new_new_n2203__ = new_new_n1217__ & ~new_new_n2202__;
  assign new_new_n2204__ = ~new_new_n1217__ & new_new_n2202__;
  assign new_new_n2205__ = ~new_new_n2203__ & ~new_new_n2204__;
  assign new_new_n2206__ = new_new_n2147__ & ~new_new_n2153__;
  assign new_new_n2207__ = ~new_new_n2147__ & new_new_n2153__;
  assign new_new_n2208__ = ~new_new_n2149__ & ~new_new_n2173__;
  assign new_new_n2209__ = ~new_new_n2207__ & new_new_n2208__;
  assign new_new_n2210__ = ~new_new_n2206__ & ~new_new_n2209__;
  assign new_new_n2211__ = new_new_n2161__ & ~new_new_n2210__;
  assign new_new_n2212__ = ~new_new_n2155__ & new_new_n2173__;
  assign new_new_n2213__ = new_new_n2149__ & new_new_n2207__;
  assign new_new_n2214__ = ~new_new_n2212__ & ~new_new_n2213__;
  assign new_new_n2215__ = ~new_new_n2161__ & ~new_new_n2214__;
  assign new_new_n2216__ = new_new_n2154__ & new_new_n2173__;
  assign new_new_n2217__ = ~new_new_n2149__ & new_new_n2206__;
  assign new_new_n2218__ = new_new_n2171__ & ~new_new_n2216__;
  assign new_new_n2219__ = ~new_new_n2217__ & new_new_n2218__;
  assign new_new_n2220__ = ~new_new_n2211__ & new_new_n2219__;
  assign new_new_n2221__ = ~new_new_n2215__ & new_new_n2220__;
  assign new_new_n2222__ = new_new_n2163__ & ~new_new_n2173__;
  assign new_new_n2223__ = ~new_new_n2164__ & ~new_new_n2222__;
  assign new_new_n2224__ = ~new_new_n2147__ & ~new_new_n2173__;
  assign new_new_n2225__ = ~new_new_n2174__ & ~new_new_n2175__;
  assign new_new_n2226__ = new_new_n2224__ & new_new_n2225__;
  assign new_new_n2227__ = ~new_new_n2171__ & ~new_new_n2223__;
  assign new_new_n2228__ = ~new_new_n2226__ & new_new_n2227__;
  assign new_new_n2229__ = ~new_new_n2221__ & ~new_new_n2228__;
  assign new_new_n2230__ = new_new_n244__ & ~new_new_n256__;
  assign new_new_n2231__ = ~new_new_n150__ & ~new_new_n2230__;
  assign new_new_n2232__ = ~new_new_n110__ & ~new_new_n415__;
  assign new_new_n2233__ = new_new_n180__ & new_new_n270__;
  assign new_new_n2234__ = new_new_n100__ & ~new_new_n2233__;
  assign new_new_n2235__ = ~new_new_n323__ & ~new_new_n560__;
  assign new_new_n2236__ = ~new_new_n918__ & ~new_new_n951__;
  assign new_new_n2237__ = new_new_n2235__ & new_new_n2236__;
  assign new_new_n2238__ = ~new_new_n168__ & ~new_new_n2234__;
  assign new_new_n2239__ = new_new_n2237__ & new_new_n2238__;
  assign new_new_n2240__ = new_new_n2231__ & ~new_new_n2232__;
  assign new_new_n2241__ = new_new_n2239__ & new_new_n2240__;
  assign new_new_n2242__ = new_new_n876__ & new_new_n2241__;
  assign new_new_n2243__ = new_new_n213__ & ~new_new_n743__;
  assign new_new_n2244__ = ~new_new_n124__ & ~new_new_n2243__;
  assign new_new_n2245__ = ~new_new_n136__ & ~new_new_n1036__;
  assign new_new_n2246__ = ~new_new_n250__ & ~new_new_n559__;
  assign new_new_n2247__ = ~new_new_n2245__ & new_new_n2246__;
  assign new_new_n2248__ = new_new_n166__ & new_new_n347__;
  assign new_new_n2249__ = new_new_n116__ & ~new_new_n2248__;
  assign new_new_n2250__ = ~new_new_n195__ & ~new_new_n223__;
  assign new_new_n2251__ = ~new_new_n218__ & ~new_new_n2250__;
  assign new_new_n2252__ = ~new_new_n243__ & ~new_new_n383__;
  assign new_new_n2253__ = ~new_new_n2249__ & new_new_n2252__;
  assign new_new_n2254__ = ~new_new_n2251__ & new_new_n2253__;
  assign new_new_n2255__ = new_new_n1110__ & new_new_n2247__;
  assign new_new_n2256__ = new_new_n2254__ & new_new_n2255__;
  assign new_new_n2257__ = new_new_n593__ & new_new_n2256__;
  assign new_new_n2258__ = ~new_new_n325__ & ~new_new_n662__;
  assign new_new_n2259__ = ~new_new_n523__ & new_new_n2258__;
  assign new_new_n2260__ = new_new_n2257__ & new_new_n2259__;
  assign new_new_n2261__ = ~new_new_n115__ & ~new_new_n524__;
  assign new_new_n2262__ = ~new_new_n335__ & ~new_new_n2261__;
  assign new_new_n2263__ = ~new_new_n342__ & new_new_n2262__;
  assign new_new_n2264__ = ~new_new_n2244__ & new_new_n2263__;
  assign new_new_n2265__ = new_new_n234__ & new_new_n2264__;
  assign new_new_n2266__ = new_new_n2242__ & new_new_n2265__;
  assign new_new_n2267__ = new_new_n2260__ & new_new_n2266__;
  assign new_new_n2268__ = ~new_new_n2229__ & ~new_new_n2267__;
  assign new_new_n2269__ = new_new_n2229__ & new_new_n2267__;
  assign new_new_n2270__ = ~new_new_n2154__ & ~new_new_n2155__;
  assign new_new_n2271__ = ~new_new_n2161__ & new_new_n2224__;
  assign new_new_n2272__ = new_new_n2161__ & ~new_new_n2224__;
  assign new_new_n2273__ = ~new_new_n2271__ & ~new_new_n2272__;
  assign new_new_n2274__ = new_new_n2270__ & new_new_n2273__;
  assign new_new_n2275__ = ~new_new_n2270__ & ~new_new_n2273__;
  assign new_new_n2276__ = ~new_new_n2274__ & ~new_new_n2275__;
  assign new_new_n2277__ = new_new_n2120__ & ~new_new_n2125__;
  assign new_new_n2278__ = ~new_new_n1615__ & ~new_new_n2123__;
  assign new_new_n2279__ = new_new_n1615__ & new_new_n2123__;
  assign new_new_n2280__ = new_new_n2133__ & ~new_new_n2279__;
  assign new_new_n2281__ = ~new_new_n2278__ & ~new_new_n2280__;
  assign new_new_n2282__ = new_new_n2277__ & new_new_n2281__;
  assign new_new_n2283__ = ~new_new_n2133__ & new_new_n2279__;
  assign new_new_n2284__ = new_new_n2133__ & new_new_n2278__;
  assign new_new_n2285__ = ~new_new_n2120__ & new_new_n2125__;
  assign new_new_n2286__ = ~new_new_n2277__ & ~new_new_n2285__;
  assign new_new_n2287__ = ~new_new_n2283__ & ~new_new_n2284__;
  assign new_new_n2288__ = new_new_n2286__ & new_new_n2287__;
  assign new_new_n2289__ = ~new_new_n2281__ & new_new_n2285__;
  assign new_new_n2290__ = ~new_new_n2282__ & ~new_new_n2289__;
  assign new_new_n2291__ = ~new_new_n2288__ & new_new_n2290__;
  assign new_new_n2292__ = new_new_n2130__ & ~new_new_n2291__;
  assign new_new_n2293__ = new_new_n2125__ & new_new_n2138__;
  assign new_new_n2294__ = new_new_n2123__ & new_new_n2293__;
  assign new_new_n2295__ = ~new_new_n2125__ & ~new_new_n2138__;
  assign new_new_n2296__ = ~new_new_n2121__ & ~new_new_n2295__;
  assign new_new_n2297__ = new_new_n2123__ & new_new_n2296__;
  assign new_new_n2298__ = ~new_new_n2293__ & ~new_new_n2297__;
  assign new_new_n2299__ = ~new_new_n2133__ & ~new_new_n2298__;
  assign new_new_n2300__ = new_new_n2121__ & ~new_new_n2125__;
  assign new_new_n2301__ = new_new_n2123__ & ~new_new_n2300__;
  assign new_new_n2302__ = new_new_n2133__ & ~new_new_n2296__;
  assign new_new_n2303__ = ~new_new_n2301__ & new_new_n2302__;
  assign new_new_n2304__ = new_new_n2121__ & new_new_n2126__;
  assign new_new_n2305__ = ~new_new_n2294__ & ~new_new_n2304__;
  assign new_new_n2306__ = ~new_new_n2303__ & new_new_n2305__;
  assign new_new_n2307__ = ~new_new_n2299__ & new_new_n2306__;
  assign new_new_n2308__ = ~new_new_n2130__ & ~new_new_n2307__;
  assign new_new_n2309__ = ~new_new_n2292__ & ~new_new_n2308__;
  assign new_new_n2310__ = ~new_new_n595__ & ~new_new_n1124__;
  assign new_new_n2311__ = ~new_new_n594__ & ~new_new_n925__;
  assign new_new_n2312__ = ~new_new_n386__ & new_new_n2311__;
  assign new_new_n2313__ = ~new_new_n443__ & new_new_n2312__;
  assign new_new_n2314__ = ~new_new_n350__ & new_new_n859__;
  assign new_new_n2315__ = new_new_n2310__ & new_new_n2314__;
  assign new_new_n2316__ = new_new_n2313__ & new_new_n2315__;
  assign new_new_n2317__ = new_new_n87__ & new_new_n136__;
  assign new_new_n2318__ = ~new_new_n141__ & ~new_new_n180__;
  assign new_new_n2319__ = ~new_new_n195__ & ~new_new_n2318__;
  assign new_new_n2320__ = ~new_new_n2317__ & ~new_new_n2319__;
  assign new_new_n2321__ = ~new_new_n166__ & new_new_n244__;
  assign new_new_n2322__ = new_new_n166__ & new_new_n658__;
  assign new_new_n2323__ = new_new_n223__ & ~new_new_n2322__;
  assign new_new_n2324__ = ~new_new_n709__ & ~new_new_n744__;
  assign new_new_n2325__ = new_new_n116__ & ~new_new_n174__;
  assign new_new_n2326__ = ~new_new_n250__ & ~new_new_n2325__;
  assign new_new_n2327__ = ~new_new_n619__ & new_new_n2326__;
  assign new_new_n2328__ = new_new_n2324__ & new_new_n2327__;
  assign new_new_n2329__ = new_new_n87__ & new_new_n256__;
  assign new_new_n2330__ = ~new_new_n87__ & new_new_n110__;
  assign new_new_n2331__ = new_new_n141__ & new_new_n2330__;
  assign new_new_n2332__ = ~new_new_n625__ & ~new_new_n2329__;
  assign new_new_n2333__ = ~new_new_n2331__ & new_new_n2332__;
  assign new_new_n2334__ = ~new_new_n54__ & ~new_new_n180__;
  assign new_new_n2335__ = new_new_n115__ & ~new_new_n1033__;
  assign new_new_n2336__ = ~new_new_n124__ & ~new_new_n2335__;
  assign new_new_n2337__ = ~new_new_n259__ & ~new_new_n560__;
  assign new_new_n2338__ = ~new_new_n662__ & new_new_n2337__;
  assign new_new_n2339__ = ~new_new_n2336__ & new_new_n2338__;
  assign new_new_n2340__ = ~new_new_n2333__ & ~new_new_n2334__;
  assign new_new_n2341__ = new_new_n2328__ & new_new_n2340__;
  assign new_new_n2342__ = new_new_n2339__ & new_new_n2341__;
  assign new_new_n2343__ = new_new_n125__ & ~new_new_n270__;
  assign new_new_n2344__ = ~new_new_n163__ & ~new_new_n2343__;
  assign new_new_n2345__ = ~new_new_n117__ & ~new_new_n404__;
  assign new_new_n2346__ = ~new_new_n921__ & new_new_n2345__;
  assign new_new_n2347__ = ~new_new_n150__ & ~new_new_n2321__;
  assign new_new_n2348__ = ~new_new_n2323__ & new_new_n2347__;
  assign new_new_n2349__ = new_new_n378__ & new_new_n2346__;
  assign new_new_n2350__ = ~new_new_n2320__ & new_new_n2344__;
  assign new_new_n2351__ = new_new_n2349__ & new_new_n2350__;
  assign new_new_n2352__ = new_new_n476__ & new_new_n2348__;
  assign new_new_n2353__ = new_new_n2351__ & new_new_n2352__;
  assign new_new_n2354__ = new_new_n2316__ & new_new_n2353__;
  assign new_new_n2355__ = new_new_n2342__ & new_new_n2354__;
  assign new_new_n2356__ = ~new_new_n2281__ & ~new_new_n2284__;
  assign new_new_n2357__ = ~new_new_n2283__ & ~new_new_n2356__;
  assign new_new_n2358__ = new_new_n2286__ & new_new_n2357__;
  assign new_new_n2359__ = ~new_new_n2286__ & ~new_new_n2357__;
  assign new_new_n2360__ = ~new_new_n2358__ & ~new_new_n2359__;
  assign new_new_n2361__ = ~new_new_n2355__ & ~new_new_n2360__;
  assign new_new_n2362__ = new_new_n2355__ & new_new_n2360__;
  assign new_new_n2363__ = ~new_new_n1740__ & new_new_n2079__;
  assign new_new_n2364__ = new_new_n1740__ & ~new_new_n2079__;
  assign new_new_n2365__ = new_new_n1742__ & new_new_n1778__;
  assign new_new_n2366__ = ~new_new_n1761__ & new_new_n2365__;
  assign new_new_n2367__ = ~new_new_n1742__ & ~new_new_n1778__;
  assign new_new_n2368__ = new_new_n1761__ & new_new_n2367__;
  assign new_new_n2369__ = ~new_new_n2366__ & ~new_new_n2368__;
  assign new_new_n2370__ = ~new_new_n2363__ & new_new_n2369__;
  assign new_new_n2371__ = ~new_new_n2364__ & new_new_n2370__;
  assign new_new_n2372__ = ~new_new_n1761__ & ~new_new_n2367__;
  assign new_new_n2373__ = ~new_new_n2365__ & ~new_new_n2372__;
  assign new_new_n2374__ = new_new_n2363__ & ~new_new_n2373__;
  assign new_new_n2375__ = new_new_n2364__ & new_new_n2373__;
  assign new_new_n2376__ = new_new_n2108__ & ~new_new_n2374__;
  assign new_new_n2377__ = ~new_new_n2375__ & new_new_n2376__;
  assign new_new_n2378__ = ~new_new_n2371__ & new_new_n2377__;
  assign new_new_n2379__ = new_new_n1740__ & new_new_n2080__;
  assign new_new_n2380__ = new_new_n1742__ & new_new_n2379__;
  assign new_new_n2381__ = ~new_new_n1740__ & new_new_n2112__;
  assign new_new_n2382__ = new_new_n1742__ & ~new_new_n2381__;
  assign new_new_n2383__ = ~new_new_n1740__ & ~new_new_n2080__;
  assign new_new_n2384__ = ~new_new_n2112__ & ~new_new_n2383__;
  assign new_new_n2385__ = new_new_n1761__ & ~new_new_n2382__;
  assign new_new_n2386__ = ~new_new_n2384__ & new_new_n2385__;
  assign new_new_n2387__ = new_new_n1742__ & new_new_n2384__;
  assign new_new_n2388__ = ~new_new_n2379__ & ~new_new_n2387__;
  assign new_new_n2389__ = ~new_new_n1761__ & ~new_new_n2388__;
  assign new_new_n2390__ = new_new_n1743__ & new_new_n2112__;
  assign new_new_n2391__ = ~new_new_n2108__ & ~new_new_n2390__;
  assign new_new_n2392__ = ~new_new_n2380__ & new_new_n2391__;
  assign new_new_n2393__ = ~new_new_n2386__ & new_new_n2392__;
  assign new_new_n2394__ = ~new_new_n2389__ & new_new_n2393__;
  assign new_new_n2395__ = ~new_new_n2378__ & ~new_new_n2394__;
  assign new_new_n2396__ = ~new_new_n174__ & new_new_n193__;
  assign new_new_n2397__ = new_new_n125__ & ~new_new_n990__;
  assign new_new_n2398__ = ~new_new_n224__ & ~new_new_n447__;
  assign new_new_n2399__ = ~new_new_n921__ & new_new_n2398__;
  assign new_new_n2400__ = ~new_new_n469__ & ~new_new_n2397__;
  assign new_new_n2401__ = new_new_n2399__ & new_new_n2400__;
  assign new_new_n2402__ = ~new_new_n553__ & new_new_n871__;
  assign new_new_n2403__ = new_new_n2310__ & ~new_new_n2396__;
  assign new_new_n2404__ = new_new_n2402__ & new_new_n2403__;
  assign new_new_n2405__ = new_new_n2401__ & new_new_n2404__;
  assign new_new_n2406__ = new_new_n81__ & new_new_n124__;
  assign new_new_n2407__ = ~new_new_n124__ & ~new_new_n160__;
  assign new_new_n2408__ = ~new_new_n195__ & ~new_new_n2407__;
  assign new_new_n2409__ = ~new_new_n2406__ & ~new_new_n2408__;
  assign new_new_n2410__ = new_new_n2344__ & ~new_new_n2409__;
  assign new_new_n2411__ = ~new_new_n560__ & new_new_n967__;
  assign new_new_n2412__ = new_new_n116__ & ~new_new_n368__;
  assign new_new_n2413__ = ~new_new_n141__ & ~new_new_n256__;
  assign new_new_n2414__ = ~new_new_n218__ & ~new_new_n448__;
  assign new_new_n2415__ = ~new_new_n351__ & ~new_new_n744__;
  assign new_new_n2416__ = ~new_new_n2414__ & new_new_n2415__;
  assign new_new_n2417__ = ~new_new_n323__ & ~new_new_n2412__;
  assign new_new_n2418__ = ~new_new_n2413__ & new_new_n2417__;
  assign new_new_n2419__ = ~new_new_n342__ & new_new_n2418__;
  assign new_new_n2420__ = ~new_new_n367__ & new_new_n2419__;
  assign new_new_n2421__ = new_new_n2410__ & new_new_n2411__;
  assign new_new_n2422__ = new_new_n2416__ & new_new_n2421__;
  assign new_new_n2423__ = new_new_n2420__ & new_new_n2422__;
  assign new_new_n2424__ = new_new_n227__ & new_new_n497__;
  assign new_new_n2425__ = ~new_new_n448__ & ~new_new_n2424__;
  assign new_new_n2426__ = new_new_n347__ & ~new_new_n570__;
  assign new_new_n2427__ = ~new_new_n335__ & new_new_n2426__;
  assign new_new_n2428__ = ~new_new_n54__ & ~new_new_n2427__;
  assign new_new_n2429__ = ~new_new_n457__ & ~new_new_n993__;
  assign new_new_n2430__ = new_new_n406__ & new_new_n2429__;
  assign new_new_n2431__ = new_new_n708__ & ~new_new_n2425__;
  assign new_new_n2432__ = ~new_new_n2428__ & new_new_n2431__;
  assign new_new_n2433__ = new_new_n375__ & new_new_n2430__;
  assign new_new_n2434__ = new_new_n881__ & new_new_n2433__;
  assign new_new_n2435__ = new_new_n2432__ & new_new_n2434__;
  assign new_new_n2436__ = new_new_n2405__ & new_new_n2435__;
  assign new_new_n2437__ = new_new_n2423__ & new_new_n2436__;
  assign new_new_n2438__ = ~new_new_n2395__ & new_new_n2437__;
  assign new_new_n2439__ = ~new_new_n2362__ & ~new_new_n2438__;
  assign new_new_n2440__ = ~new_new_n2361__ & ~new_new_n2439__;
  assign new_new_n2441__ = ~new_new_n2309__ & ~new_new_n2440__;
  assign new_new_n2442__ = new_new_n2309__ & new_new_n2440__;
  assign new_new_n2443__ = new_new_n162__ & ~new_new_n483__;
  assign new_new_n2444__ = new_new_n160__ & ~new_new_n373__;
  assign new_new_n2445__ = ~new_new_n343__ & ~new_new_n2444__;
  assign new_new_n2446__ = new_new_n174__ & new_new_n180__;
  assign new_new_n2447__ = new_new_n162__ & ~new_new_n2446__;
  assign new_new_n2448__ = ~new_new_n744__ & ~new_new_n2447__;
  assign new_new_n2449__ = ~new_new_n2445__ & new_new_n2448__;
  assign new_new_n2450__ = new_new_n924__ & new_new_n2449__;
  assign new_new_n2451__ = new_new_n213__ & new_new_n347__;
  assign new_new_n2452__ = new_new_n992__ & new_new_n2451__;
  assign new_new_n2453__ = new_new_n116__ & ~new_new_n2452__;
  assign new_new_n2454__ = ~new_new_n87__ & ~new_new_n483__;
  assign new_new_n2455__ = ~new_new_n54__ & new_new_n2454__;
  assign new_new_n2456__ = new_new_n162__ & ~new_new_n903__;
  assign new_new_n2457__ = ~new_new_n187__ & ~new_new_n2455__;
  assign new_new_n2458__ = ~new_new_n2456__ & new_new_n2457__;
  assign new_new_n2459__ = new_new_n148__ & new_new_n265__;
  assign new_new_n2460__ = new_new_n181__ & ~new_new_n2459__;
  assign new_new_n2461__ = ~new_new_n115__ & new_new_n195__;
  assign new_new_n2462__ = ~new_new_n150__ & ~new_new_n594__;
  assign new_new_n2463__ = ~new_new_n2443__ & ~new_new_n2460__;
  assign new_new_n2464__ = ~new_new_n2461__ & new_new_n2463__;
  assign new_new_n2465__ = new_new_n2462__ & new_new_n2464__;
  assign new_new_n2466__ = ~new_new_n2453__ & new_new_n2458__;
  assign new_new_n2467__ = new_new_n2465__ & new_new_n2466__;
  assign new_new_n2468__ = new_new_n2450__ & new_new_n2467__;
  assign new_new_n2469__ = ~new_new_n213__ & ~new_new_n493__;
  assign new_new_n2470__ = ~new_new_n100__ & new_new_n160__;
  assign new_new_n2471__ = new_new_n347__ & new_new_n492__;
  assign new_new_n2472__ = ~new_new_n2470__ & ~new_new_n2471__;
  assign new_new_n2473__ = new_new_n238__ & new_new_n1051__;
  assign new_new_n2474__ = new_new_n195__ & ~new_new_n2473__;
  assign new_new_n2475__ = ~new_new_n2469__ & ~new_new_n2474__;
  assign new_new_n2476__ = ~new_new_n2472__ & new_new_n2475__;
  assign new_new_n2477__ = ~new_new_n2318__ & ~new_new_n2407__;
  assign new_new_n2478__ = new_new_n87__ & ~new_new_n2477__;
  assign new_new_n2479__ = ~new_new_n239__ & ~new_new_n384__;
  assign new_new_n2480__ = ~new_new_n976__ & new_new_n2479__;
  assign new_new_n2481__ = ~new_new_n243__ & ~new_new_n745__;
  assign new_new_n2482__ = new_new_n2480__ & new_new_n2481__;
  assign new_new_n2483__ = new_new_n470__ & new_new_n915__;
  assign new_new_n2484__ = new_new_n1450__ & ~new_new_n2478__;
  assign new_new_n2485__ = new_new_n2483__ & new_new_n2484__;
  assign new_new_n2486__ = new_new_n975__ & new_new_n2482__;
  assign new_new_n2487__ = new_new_n2485__ & new_new_n2486__;
  assign new_new_n2488__ = new_new_n869__ & new_new_n2476__;
  assign new_new_n2489__ = new_new_n2487__ & new_new_n2488__;
  assign new_new_n2490__ = new_new_n538__ & new_new_n2489__;
  assign new_new_n2491__ = new_new_n2468__ & new_new_n2490__;
  assign new_new_n2492__ = ~new_new_n2442__ & ~new_new_n2491__;
  assign new_new_n2493__ = ~new_new_n2441__ & ~new_new_n2492__;
  assign new_new_n2494__ = ~new_new_n2276__ & ~new_new_n2493__;
  assign new_new_n2495__ = new_new_n2276__ & new_new_n2493__;
  assign new_new_n2496__ = ~new_new_n194__ & ~new_new_n261__;
  assign new_new_n2497__ = new_new_n81__ & new_new_n238__;
  assign new_new_n2498__ = new_new_n110__ & new_new_n2497__;
  assign new_new_n2499__ = new_new_n223__ & ~new_new_n2498__;
  assign new_new_n2500__ = new_new_n81__ & new_new_n115__;
  assign new_new_n2501__ = new_new_n87__ & new_new_n2500__;
  assign new_new_n2502__ = ~new_new_n897__ & ~new_new_n2501__;
  assign new_new_n2503__ = ~new_new_n274__ & ~new_new_n475__;
  assign new_new_n2504__ = ~new_new_n322__ & new_new_n2503__;
  assign new_new_n2505__ = ~new_new_n2499__ & new_new_n2504__;
  assign new_new_n2506__ = ~new_new_n2502__ & new_new_n2505__;
  assign new_new_n2507__ = new_new_n2411__ & ~new_new_n2496__;
  assign new_new_n2508__ = new_new_n2506__ & new_new_n2507__;
  assign new_new_n2509__ = new_new_n2476__ & new_new_n2508__;
  assign new_new_n2510__ = new_new_n2405__ & new_new_n2509__;
  assign new_new_n2511__ = new_new_n391__ & new_new_n2510__;
  assign new_new_n2512__ = ~new_new_n2495__ & ~new_new_n2511__;
  assign new_new_n2513__ = ~new_new_n2494__ & ~new_new_n2512__;
  assign new_new_n2514__ = ~new_new_n2269__ & ~new_new_n2513__;
  assign new_new_n2515__ = ~new_new_n2268__ & ~new_new_n2514__;
  assign new_new_n2516__ = new_new_n1394__ & ~new_new_n2181__;
  assign new_new_n2517__ = ~new_new_n1394__ & new_new_n2181__;
  assign new_new_n2518__ = ~new_new_n2516__ & ~new_new_n2517__;
  assign new_new_n2519__ = ~new_new_n1256__ & new_new_n2518__;
  assign new_new_n2520__ = new_new_n1256__ & ~new_new_n2518__;
  assign new_new_n2521__ = ~new_new_n2519__ & ~new_new_n2520__;
  assign new_new_n2522__ = new_new_n1211__ & ~new_new_n2193__;
  assign new_new_n2523__ = ~new_new_n1211__ & new_new_n2193__;
  assign new_new_n2524__ = ~new_new_n2522__ & ~new_new_n2523__;
  assign new_new_n2525__ = new_new_n2521__ & new_new_n2524__;
  assign new_new_n2526__ = ~new_new_n2521__ & ~new_new_n2524__;
  assign new_new_n2527__ = ~new_new_n2525__ & ~new_new_n2526__;
  assign new_new_n2528__ = ~new_new_n2515__ & ~new_new_n2527__;
  assign new_new_n2529__ = new_new_n2515__ & new_new_n2527__;
  assign new_new_n2530__ = new_new_n54__ & ~new_new_n244__;
  assign new_new_n2531__ = ~new_new_n218__ & ~new_new_n2530__;
  assign new_new_n2532__ = new_new_n115__ & new_new_n180__;
  assign new_new_n2533__ = new_new_n125__ & ~new_new_n2532__;
  assign new_new_n2534__ = new_new_n181__ & ~new_new_n554__;
  assign new_new_n2535__ = new_new_n270__ & new_new_n2317__;
  assign new_new_n2536__ = ~new_new_n99__ & ~new_new_n2535__;
  assign new_new_n2537__ = ~new_new_n2230__ & ~new_new_n2536__;
  assign new_new_n2538__ = ~new_new_n87__ & new_new_n136__;
  assign new_new_n2539__ = new_new_n174__ & new_new_n2538__;
  assign new_new_n2540__ = ~new_new_n2537__ & ~new_new_n2539__;
  assign new_new_n2541__ = new_new_n195__ & ~new_new_n494__;
  assign new_new_n2542__ = new_new_n112__ & ~new_new_n384__;
  assign new_new_n2543__ = ~new_new_n379__ & ~new_new_n2533__;
  assign new_new_n2544__ = ~new_new_n2534__ & ~new_new_n2541__;
  assign new_new_n2545__ = new_new_n2543__ & new_new_n2544__;
  assign new_new_n2546__ = new_new_n864__ & new_new_n2542__;
  assign new_new_n2547__ = ~new_new_n2531__ & new_new_n2546__;
  assign new_new_n2548__ = ~new_new_n935__ & new_new_n2545__;
  assign new_new_n2549__ = ~new_new_n2540__ & new_new_n2548__;
  assign new_new_n2550__ = new_new_n2450__ & new_new_n2547__;
  assign new_new_n2551__ = new_new_n2549__ & new_new_n2550__;
  assign new_new_n2552__ = new_new_n983__ & new_new_n2316__;
  assign new_new_n2553__ = new_new_n2551__ & new_new_n2552__;
  assign new_new_n2554__ = ~new_new_n2529__ & ~new_new_n2553__;
  assign new_new_n2555__ = ~new_new_n2528__ & ~new_new_n2554__;
  assign new_new_n2556__ = ~new_new_n335__ & ~new_new_n1127__;
  assign new_new_n2557__ = ~new_new_n222__ & new_new_n2556__;
  assign new_new_n2558__ = ~new_new_n377__ & ~new_new_n662__;
  assign new_new_n2559__ = ~new_new_n2461__ & new_new_n2558__;
  assign new_new_n2560__ = ~new_new_n2245__ & new_new_n2557__;
  assign new_new_n2561__ = new_new_n2559__ & new_new_n2560__;
  assign new_new_n2562__ = new_new_n909__ & new_new_n1120__;
  assign new_new_n2563__ = new_new_n2561__ & new_new_n2562__;
  assign new_new_n2564__ = new_new_n218__ & new_new_n270__;
  assign new_new_n2565__ = new_new_n181__ & ~new_new_n2564__;
  assign new_new_n2566__ = new_new_n892__ & ~new_new_n2565__;
  assign new_new_n2567__ = ~new_new_n589__ & new_new_n736__;
  assign new_new_n2568__ = ~new_new_n274__ & ~new_new_n328__;
  assign new_new_n2569__ = ~new_new_n2567__ & new_new_n2568__;
  assign new_new_n2570__ = ~new_new_n125__ & new_new_n2497__;
  assign new_new_n2571__ = ~new_new_n365__ & ~new_new_n2570__;
  assign new_new_n2572__ = ~new_new_n921__ & ~new_new_n976__;
  assign new_new_n2573__ = ~new_new_n413__ & new_new_n2572__;
  assign new_new_n2574__ = new_new_n2231__ & new_new_n2573__;
  assign new_new_n2575__ = new_new_n2569__ & ~new_new_n2571__;
  assign new_new_n2576__ = new_new_n2574__ & new_new_n2575__;
  assign new_new_n2577__ = new_new_n203__ & new_new_n2576__;
  assign new_new_n2578__ = new_new_n2563__ & new_new_n2577__;
  assign new_new_n2579__ = new_new_n2566__ & new_new_n2578__;
  assign new_new_n2580__ = new_new_n2555__ & new_new_n2579__;
  assign new_new_n2581__ = ~new_new_n2555__ & ~new_new_n2579__;
  assign new_new_n2582__ = ~new_new_n2580__ & ~new_new_n2581__;
  assign new_new_n2583__ = ~new_new_n2205__ & new_new_n2582__;
  assign new_new_n2584__ = new_new_n2205__ & ~new_new_n2582__;
  assign new_new_n2585__ = ~new_new_n2583__ & ~new_new_n2584__;
  assign new_new_n2586__ = ~new_new_n320__ & new_new_n2585__;
  assign new_new_n2587__ = ~new_new_n2528__ & ~new_new_n2529__;
  assign new_new_n2588__ = new_new_n2553__ & ~new_new_n2587__;
  assign new_new_n2589__ = ~new_new_n2553__ & new_new_n2587__;
  assign new_new_n2590__ = ~new_new_n2588__ & ~new_new_n2589__;
  assign new_new_n2591__ = ~new_new_n318__ & ~new_new_n1191__;
  assign new_new_n2592__ = ~new_new_n311__ & ~new_new_n1192__;
  assign new_new_n2593__ = ~new_new_n2591__ & ~new_new_n2592__;
  assign new_new_n2594__ = new_new_n2590__ & new_new_n2593__;
  assign new_new_n2595__ = ~new_new_n2586__ & ~new_new_n2594__;
  assign new_new_n2596__ = ~new_new_n311__ & ~new_new_n318__;
  assign new_new_n2597__ = ~new_new_n2268__ & ~new_new_n2269__;
  assign new_new_n2598__ = new_new_n2513__ & ~new_new_n2597__;
  assign new_new_n2599__ = ~new_new_n2513__ & new_new_n2597__;
  assign new_new_n2600__ = ~new_new_n2598__ & ~new_new_n2599__;
  assign new_new_n2601__ = ~new_new_n2494__ & ~new_new_n2495__;
  assign new_new_n2602__ = new_new_n2511__ & ~new_new_n2601__;
  assign new_new_n2603__ = ~new_new_n2511__ & new_new_n2601__;
  assign new_new_n2604__ = ~new_new_n2602__ & ~new_new_n2603__;
  assign new_new_n2605__ = ~new_new_n2441__ & ~new_new_n2442__;
  assign new_new_n2606__ = new_new_n2491__ & ~new_new_n2605__;
  assign new_new_n2607__ = ~new_new_n2491__ & new_new_n2605__;
  assign new_new_n2608__ = ~new_new_n2606__ & ~new_new_n2607__;
  assign new_new_n2609__ = ~new_new_n2604__ & new_new_n2608__;
  assign new_new_n2610__ = new_new_n2395__ & ~new_new_n2437__;
  assign new_new_n2611__ = ~new_new_n2438__ & ~new_new_n2610__;
  assign new_new_n2612__ = ~new_new_n2600__ & ~new_new_n2611__;
  assign new_new_n2613__ = ~new_new_n2609__ & ~new_new_n2612__;
  assign new_new_n2614__ = ~new_new_n2600__ & ~new_new_n2604__;
  assign new_new_n2615__ = ~new_new_n2361__ & ~new_new_n2362__;
  assign new_new_n2616__ = new_new_n2438__ & ~new_new_n2615__;
  assign new_new_n2617__ = ~new_new_n2438__ & new_new_n2615__;
  assign new_new_n2618__ = ~new_new_n2616__ & ~new_new_n2617__;
  assign new_new_n2619__ = ~new_new_n2614__ & new_new_n2618__;
  assign new_new_n2620__ = ~new_new_n2613__ & new_new_n2619__;
  assign new_new_n2621__ = new_new_n2604__ & ~new_new_n2608__;
  assign new_new_n2622__ = new_new_n2600__ & new_new_n2621__;
  assign new_new_n2623__ = ~new_new_n2614__ & ~new_new_n2622__;
  assign new_new_n2624__ = ~new_new_n2618__ & ~new_new_n2623__;
  assign new_new_n2625__ = new_new_n2611__ & ~new_new_n2615__;
  assign new_new_n2626__ = new_new_n2604__ & new_new_n2625__;
  assign new_new_n2627__ = new_new_n2600__ & new_new_n2626__;
  assign new_new_n2628__ = ~new_new_n2614__ & ~new_new_n2627__;
  assign new_new_n2629__ = ~new_new_n2608__ & ~new_new_n2628__;
  assign new_new_n2630__ = ~new_new_n2620__ & ~new_new_n2624__;
  assign new_new_n2631__ = ~new_new_n2629__ & new_new_n2630__;
  assign new_new_n2632__ = new_new_n2604__ & new_new_n2608__;
  assign new_new_n2633__ = ~new_new_n2600__ & new_new_n2632__;
  assign new_new_n2634__ = new_new_n2631__ & ~new_new_n2633__;
  assign new_new_n2635__ = ~new_new_n2600__ & new_new_n2634__;
  assign new_new_n2636__ = new_new_n2600__ & ~new_new_n2631__;
  assign new_new_n2637__ = ~new_new_n2635__ & ~new_new_n2636__;
  assign new_new_n2638__ = new_new_n2590__ & ~new_new_n2637__;
  assign new_new_n2639__ = new_new_n2590__ & ~new_new_n2634__;
  assign new_new_n2640__ = ~new_new_n2600__ & ~new_new_n2634__;
  assign new_new_n2641__ = ~new_new_n2590__ & ~new_new_n2640__;
  assign new_new_n2642__ = ~new_new_n2639__ & ~new_new_n2641__;
  assign new_new_n2643__ = new_new_n2511__ & ~new_new_n2642__;
  assign new_new_n2644__ = ~new_new_n2590__ & new_new_n2600__;
  assign new_new_n2645__ = new_new_n2634__ & new_new_n2644__;
  assign new_new_n2646__ = ~new_new_n2639__ & ~new_new_n2645__;
  assign new_new_n2647__ = ~new_new_n2511__ & new_new_n2646__;
  assign new_new_n2648__ = new_new_n2601__ & ~new_new_n2647__;
  assign new_new_n2649__ = ~new_new_n2643__ & new_new_n2648__;
  assign new_new_n2650__ = new_new_n2511__ & new_new_n2646__;
  assign new_new_n2651__ = ~new_new_n2511__ & ~new_new_n2642__;
  assign new_new_n2652__ = ~new_new_n2601__ & ~new_new_n2650__;
  assign new_new_n2653__ = ~new_new_n2651__ & new_new_n2652__;
  assign new_new_n2654__ = ~new_new_n2638__ & ~new_new_n2649__;
  assign new_new_n2655__ = ~new_new_n2653__ & new_new_n2654__;
  assign new_new_n2656__ = ~new_new_n2600__ & ~new_new_n2655__;
  assign new_new_n2657__ = new_new_n2590__ & ~new_new_n2656__;
  assign new_new_n2658__ = ~new_new_n2585__ & ~new_new_n2657__;
  assign new_new_n2659__ = new_new_n2608__ & new_new_n2618__;
  assign new_new_n2660__ = ~new_new_n2604__ & ~new_new_n2659__;
  assign new_new_n2661__ = new_new_n2600__ & ~new_new_n2660__;
  assign new_new_n2662__ = ~new_new_n2590__ & ~new_new_n2661__;
  assign new_new_n2663__ = new_new_n2585__ & ~new_new_n2662__;
  assign new_new_n2664__ = ~new_new_n2658__ & ~new_new_n2663__;
  assign new_new_n2665__ = new_new_n166__ & new_new_n2498__;
  assign new_new_n2666__ = new_new_n88__ & ~new_new_n141__;
  assign new_new_n2667__ = ~new_new_n125__ & ~new_new_n2666__;
  assign new_new_n2668__ = ~new_new_n2665__ & ~new_new_n2667__;
  assign new_new_n2669__ = ~new_new_n54__ & ~new_new_n347__;
  assign new_new_n2670__ = new_new_n141__ & ~new_new_n2669__;
  assign new_new_n2671__ = new_new_n174__ & new_new_n970__;
  assign new_new_n2672__ = ~new_new_n87__ & ~new_new_n2671__;
  assign new_new_n2673__ = new_new_n148__ & ~new_new_n2672__;
  assign new_new_n2674__ = ~new_new_n2670__ & ~new_new_n2673__;
  assign new_new_n2675__ = ~new_new_n392__ & ~new_new_n571__;
  assign new_new_n2676__ = ~new_new_n243__ & new_new_n2675__;
  assign new_new_n2677__ = ~new_new_n2668__ & new_new_n2676__;
  assign new_new_n2678__ = ~new_new_n2674__ & new_new_n2677__;
  assign new_new_n2679__ = new_new_n116__ & ~new_new_n347__;
  assign new_new_n2680__ = new_new_n115__ & ~new_new_n2679__;
  assign new_new_n2681__ = ~new_new_n415__ & ~new_new_n2680__;
  assign new_new_n2682__ = ~new_new_n227__ & ~new_new_n2250__;
  assign new_new_n2683__ = ~new_new_n100__ & ~new_new_n244__;
  assign new_new_n2684__ = ~new_new_n270__ & ~new_new_n2683__;
  assign new_new_n2685__ = ~new_new_n116__ & ~new_new_n2684__;
  assign new_new_n2686__ = ~new_new_n641__ & ~new_new_n2685__;
  assign new_new_n2687__ = ~new_new_n192__ & new_new_n472__;
  assign new_new_n2688__ = ~new_new_n213__ & ~new_new_n245__;
  assign new_new_n2689__ = ~new_new_n219__ & ~new_new_n976__;
  assign new_new_n2690__ = ~new_new_n403__ & new_new_n2689__;
  assign new_new_n2691__ = ~new_new_n2321__ & ~new_new_n2687__;
  assign new_new_n2692__ = new_new_n2690__ & new_new_n2691__;
  assign new_new_n2693__ = new_new_n728__ & ~new_new_n2682__;
  assign new_new_n2694__ = ~new_new_n2688__ & new_new_n2693__;
  assign new_new_n2695__ = new_new_n2416__ & new_new_n2692__;
  assign new_new_n2696__ = new_new_n2694__ & new_new_n2695__;
  assign new_new_n2697__ = new_new_n593__ & ~new_new_n2686__;
  assign new_new_n2698__ = new_new_n2696__ & new_new_n2697__;
  assign new_new_n2699__ = ~new_new_n2681__ & new_new_n2698__;
  assign new_new_n2700__ = new_new_n223__ & ~new_new_n903__;
  assign new_new_n2701__ = new_new_n162__ & ~new_new_n2233__;
  assign new_new_n2702__ = ~new_new_n443__ & ~new_new_n469__;
  assign new_new_n2703__ = ~new_new_n2700__ & ~new_new_n2701__;
  assign new_new_n2704__ = new_new_n2702__ & new_new_n2703__;
  assign new_new_n2705__ = new_new_n1034__ & new_new_n1441__;
  assign new_new_n2706__ = new_new_n2704__ & new_new_n2705__;
  assign new_new_n2707__ = ~new_new_n115__ & ~new_new_n180__;
  assign new_new_n2708__ = new_new_n99__ & ~new_new_n393__;
  assign new_new_n2709__ = new_new_n87__ & ~new_new_n2532__;
  assign new_new_n2710__ = ~new_new_n2708__ & new_new_n2709__;
  assign new_new_n2711__ = ~new_new_n730__ & ~new_new_n993__;
  assign new_new_n2712__ = ~new_new_n2707__ & new_new_n2711__;
  assign new_new_n2713__ = ~new_new_n185__ & ~new_new_n709__;
  assign new_new_n2714__ = ~new_new_n971__ & new_new_n2713__;
  assign new_new_n2715__ = new_new_n915__ & new_new_n2712__;
  assign new_new_n2716__ = ~new_new_n2710__ & new_new_n2715__;
  assign new_new_n2717__ = new_new_n1449__ & new_new_n2714__;
  assign new_new_n2718__ = new_new_n2716__ & new_new_n2717__;
  assign new_new_n2719__ = new_new_n2706__ & new_new_n2718__;
  assign new_new_n2720__ = new_new_n2678__ & new_new_n2719__;
  assign new_new_n2721__ = new_new_n2699__ & new_new_n2720__;
  assign new_new_n2722__ = ~new_new_n2205__ & ~new_new_n2580__;
  assign new_new_n2723__ = ~new_new_n2581__ & ~new_new_n2722__;
  assign new_new_n2724__ = ~new_new_n2721__ & ~new_new_n2723__;
  assign new_new_n2725__ = new_new_n2721__ & new_new_n2723__;
  assign new_new_n2726__ = ~new_new_n2724__ & ~new_new_n2725__;
  assign new_new_n2727__ = ~new_new_n857__ & ~new_new_n1014__;
  assign new_new_n2728__ = ~new_new_n856__ & ~new_new_n2727__;
  assign new_new_n2729__ = ~new_new_n775__ & ~new_new_n787__;
  assign new_new_n2730__ = ~new_new_n774__ & ~new_new_n2729__;
  assign new_new_n2731__ = ~new_new_n437__ & new_new_n686__;
  assign new_new_n2732__ = new_new_n437__ & ~new_new_n686__;
  assign new_new_n2733__ = ~new_new_n2731__ & ~new_new_n2732__;
  assign new_new_n2734__ = new_new_n760__ & ~new_new_n2733__;
  assign new_new_n2735__ = new_new_n689__ & ~new_new_n760__;
  assign new_new_n2736__ = ~new_new_n829__ & new_new_n2735__;
  assign new_new_n2737__ = ~new_new_n2734__ & ~new_new_n2736__;
  assign new_new_n2738__ = new_new_n2730__ & new_new_n2737__;
  assign new_new_n2739__ = ~new_new_n2730__ & ~new_new_n2737__;
  assign new_new_n2740__ = ~new_new_n2738__ & ~new_new_n2739__;
  assign new_new_n2741__ = ~new_new_n791__ & new_new_n810__;
  assign new_new_n2742__ = ~new_new_n648__ & ~new_new_n810__;
  assign new_new_n2743__ = new_new_n764__ & new_new_n1340__;
  assign new_new_n2744__ = ~new_new_n2741__ & ~new_new_n2742__;
  assign new_new_n2745__ = ~new_new_n2743__ & new_new_n2744__;
  assign new_new_n2746__ = ~new_new_n2740__ & new_new_n2745__;
  assign new_new_n2747__ = new_new_n2740__ & ~new_new_n2745__;
  assign new_new_n2748__ = ~new_new_n2746__ & ~new_new_n2747__;
  assign new_new_n2749__ = ~new_new_n2728__ & ~new_new_n2748__;
  assign new_new_n2750__ = new_new_n2728__ & new_new_n2748__;
  assign new_new_n2751__ = ~new_new_n2749__ & ~new_new_n2750__;
  assign new_new_n2752__ = new_new_n615__ & ~new_new_n816__;
  assign new_new_n2753__ = ~new_new_n615__ & new_new_n816__;
  assign new_new_n2754__ = ~new_new_n2752__ & ~new_new_n2753__;
  assign new_new_n2755__ = ~new_new_n648__ & new_new_n2754__;
  assign new_new_n2756__ = ~new_new_n785__ & new_new_n2755__;
  assign new_new_n2757__ = new_new_n785__ & ~new_new_n2755__;
  assign new_new_n2758__ = ~new_new_n2756__ & ~new_new_n2757__;
  assign new_new_n2759__ = ~new_new_n1018__ & ~new_new_n1202__;
  assign new_new_n2760__ = ~new_new_n1217__ & ~new_new_n2184__;
  assign new_new_n2761__ = new_new_n2193__ & ~new_new_n2760__;
  assign new_new_n2762__ = ~new_new_n2198__ & ~new_new_n2761__;
  assign new_new_n2763__ = new_new_n1395__ & new_new_n2762__;
  assign new_new_n2764__ = new_new_n1256__ & new_new_n2181__;
  assign new_new_n2765__ = ~new_new_n2762__ & ~new_new_n2764__;
  assign new_new_n2766__ = ~new_new_n1217__ & ~new_new_n2765__;
  assign new_new_n2767__ = ~new_new_n1395__ & new_new_n2193__;
  assign new_new_n2768__ = new_new_n1217__ & ~new_new_n2764__;
  assign new_new_n2769__ = ~new_new_n2184__ & ~new_new_n2767__;
  assign new_new_n2770__ = ~new_new_n2768__ & new_new_n2769__;
  assign new_new_n2771__ = ~new_new_n2763__ & ~new_new_n2770__;
  assign new_new_n2772__ = ~new_new_n2766__ & new_new_n2771__;
  assign new_new_n2773__ = ~new_new_n2759__ & new_new_n2772__;
  assign new_new_n2774__ = new_new_n2759__ & ~new_new_n2772__;
  assign new_new_n2775__ = ~new_new_n2773__ & ~new_new_n2774__;
  assign new_new_n2776__ = new_new_n2758__ & ~new_new_n2775__;
  assign new_new_n2777__ = ~new_new_n2758__ & new_new_n2775__;
  assign new_new_n2778__ = ~new_new_n2776__ & ~new_new_n2777__;
  assign new_new_n2779__ = new_new_n2751__ & new_new_n2778__;
  assign new_new_n2780__ = ~new_new_n2751__ & ~new_new_n2778__;
  assign new_new_n2781__ = ~new_new_n2779__ & ~new_new_n2780__;
  assign new_new_n2782__ = new_new_n2726__ & ~new_new_n2781__;
  assign new_new_n2783__ = ~new_new_n2726__ & new_new_n2781__;
  assign new_new_n2784__ = ~new_new_n2782__ & ~new_new_n2783__;
  assign new_new_n2785__ = ~new_new_n2664__ & ~new_new_n2784__;
  assign new_new_n2786__ = new_new_n2596__ & new_new_n2785__;
  assign new_new_n2787__ = new_new_n2595__ & ~new_new_n2786__;
  assign new_new_n2788__ = new_new_n301__ & ~new_new_n2787__;
  assign new_new_n2789__ = new_new_n316__ & ~new_new_n2784__;
  assign new_new_n2790__ = ~new_new_n316__ & new_new_n2784__;
  assign new_new_n2791__ = new_new_n2596__ & ~new_new_n2789__;
  assign new_new_n2792__ = ~new_new_n2790__ & new_new_n2791__;
  assign new_new_n2793__ = new_new_n2664__ & new_new_n2792__;
  assign new_new_n2794__ = ~new_new_n2664__ & new_new_n2784__;
  assign new_new_n2795__ = new_new_n2596__ & ~new_new_n2794__;
  assign new_new_n2796__ = ~new_new_n301__ & new_new_n2595__;
  assign new_new_n2797__ = ~new_new_n2795__ & new_new_n2796__;
  assign new_new_n2798__ = ~new_new_n2793__ & ~new_new_n2797__;
  assign new_new_n2799__ = ~new_new_n2788__ & new_new_n2798__;
  assign new_new_n2800__ = ~new_new_n301__ & new_new_n615__;
  assign new_new_n2801__ = ~new_new_n810__ & ~new_new_n816__;
  assign new_new_n2802__ = new_new_n2800__ & new_new_n2801__;
  assign new_new_n2803__ = new_new_n301__ & ~new_new_n615__;
  assign new_new_n2804__ = new_new_n816__ & new_new_n2803__;
  assign new_new_n2805__ = new_new_n810__ & new_new_n2804__;
  assign new_new_n2806__ = ~new_new_n2802__ & ~new_new_n2805__;
  assign new_new_n2807__ = new_new_n2618__ & ~new_new_n2806__;
  assign new_new_n2808__ = ~new_new_n2800__ & ~new_new_n2803__;
  assign new_new_n2809__ = new_new_n2754__ & ~new_new_n2808__;
  assign new_new_n2810__ = new_new_n2608__ & new_new_n2809__;
  assign new_new_n2811__ = ~new_new_n2807__ & ~new_new_n2810__;
  assign new_new_n2812__ = ~new_new_n2438__ & ~new_new_n2609__;
  assign new_new_n2813__ = ~new_new_n2621__ & new_new_n2812__;
  assign new_new_n2814__ = new_new_n2437__ & new_new_n2609__;
  assign new_new_n2815__ = ~new_new_n2621__ & ~new_new_n2814__;
  assign new_new_n2816__ = ~new_new_n2395__ & ~new_new_n2815__;
  assign new_new_n2817__ = new_new_n2615__ & ~new_new_n2813__;
  assign new_new_n2818__ = ~new_new_n2816__ & new_new_n2817__;
  assign new_new_n2819__ = ~new_new_n2608__ & new_new_n2611__;
  assign new_new_n2820__ = new_new_n2615__ & ~new_new_n2819__;
  assign new_new_n2821__ = ~new_new_n2438__ & new_new_n2608__;
  assign new_new_n2822__ = ~new_new_n2608__ & ~new_new_n2610__;
  assign new_new_n2823__ = ~new_new_n2821__ & ~new_new_n2822__;
  assign new_new_n2824__ = ~new_new_n2820__ & ~new_new_n2823__;
  assign new_new_n2825__ = new_new_n2604__ & new_new_n2824__;
  assign new_new_n2826__ = ~new_new_n2615__ & new_new_n2823__;
  assign new_new_n2827__ = ~new_new_n2604__ & new_new_n2826__;
  assign new_new_n2828__ = ~new_new_n2825__ & ~new_new_n2827__;
  assign new_new_n2829__ = ~new_new_n2818__ & new_new_n2828__;
  assign new_new_n2830__ = ~new_new_n2604__ & new_new_n2829__;
  assign new_new_n2831__ = new_new_n2808__ & ~new_new_n2830__;
  assign new_new_n2832__ = new_new_n810__ & ~new_new_n2831__;
  assign new_new_n2833__ = ~new_new_n2604__ & ~new_new_n2829__;
  assign new_new_n2834__ = ~new_new_n816__ & ~new_new_n2833__;
  assign new_new_n2835__ = new_new_n2604__ & new_new_n2829__;
  assign new_new_n2836__ = new_new_n816__ & ~new_new_n2835__;
  assign new_new_n2837__ = new_new_n2808__ & ~new_new_n2834__;
  assign new_new_n2838__ = ~new_new_n2836__ & new_new_n2837__;
  assign new_new_n2839__ = ~new_new_n2832__ & ~new_new_n2838__;
  assign new_new_n2840__ = new_new_n2811__ & ~new_new_n2839__;
  assign new_new_n2841__ = new_new_n2604__ & ~new_new_n2829__;
  assign new_new_n2842__ = new_new_n2808__ & new_new_n2841__;
  assign new_new_n2843__ = new_new_n2811__ & ~new_new_n2842__;
  assign new_new_n2844__ = ~new_new_n810__ & ~new_new_n2843__;
  assign new_new_n2845__ = ~new_new_n2840__ & ~new_new_n2844__;
  assign new_new_n2846__ = ~new_new_n764__ & ~new_new_n810__;
  assign new_new_n2847__ = new_new_n764__ & new_new_n810__;
  assign new_new_n2848__ = ~new_new_n2846__ & ~new_new_n2847__;
  assign new_new_n2849__ = ~new_new_n2611__ & new_new_n2848__;
  assign new_new_n2850__ = new_new_n2618__ & ~new_new_n2803__;
  assign new_new_n2851__ = new_new_n2611__ & ~new_new_n2850__;
  assign new_new_n2852__ = new_new_n816__ & ~new_new_n2611__;
  assign new_new_n2853__ = new_new_n2800__ & ~new_new_n2852__;
  assign new_new_n2854__ = ~new_new_n2804__ & ~new_new_n2853__;
  assign new_new_n2855__ = ~new_new_n2851__ & new_new_n2854__;
  assign new_new_n2856__ = new_new_n2618__ & new_new_n2809__;
  assign new_new_n2857__ = ~new_new_n2611__ & ~new_new_n2806__;
  assign new_new_n2858__ = new_new_n810__ & new_new_n816__;
  assign new_new_n2859__ = ~new_new_n2801__ & ~new_new_n2858__;
  assign new_new_n2860__ = new_new_n2625__ & ~new_new_n2859__;
  assign new_new_n2861__ = new_new_n2608__ & new_new_n2860__;
  assign new_new_n2862__ = ~new_new_n2608__ & ~new_new_n2860__;
  assign new_new_n2863__ = new_new_n2808__ & ~new_new_n2861__;
  assign new_new_n2864__ = ~new_new_n2862__ & new_new_n2863__;
  assign new_new_n2865__ = ~new_new_n2856__ & ~new_new_n2857__;
  assign new_new_n2866__ = ~new_new_n2864__ & new_new_n2865__;
  assign new_new_n2867__ = new_new_n810__ & ~new_new_n2855__;
  assign new_new_n2868__ = new_new_n2866__ & new_new_n2867__;
  assign new_new_n2869__ = ~new_new_n2849__ & ~new_new_n2868__;
  assign new_new_n2870__ = ~new_new_n2845__ & ~new_new_n2869__;
  assign new_new_n2871__ = new_new_n2604__ & new_new_n2809__;
  assign new_new_n2872__ = new_new_n2608__ & ~new_new_n2806__;
  assign new_new_n2873__ = ~new_new_n2871__ & ~new_new_n2872__;
  assign new_new_n2874__ = new_new_n2600__ & new_new_n2808__;
  assign new_new_n2875__ = new_new_n2634__ & new_new_n2874__;
  assign new_new_n2876__ = new_new_n2873__ & ~new_new_n2875__;
  assign new_new_n2877__ = ~new_new_n810__ & ~new_new_n2876__;
  assign new_new_n2878__ = new_new_n816__ & ~new_new_n2636__;
  assign new_new_n2879__ = ~new_new_n816__ & ~new_new_n2635__;
  assign new_new_n2880__ = new_new_n2808__ & ~new_new_n2878__;
  assign new_new_n2881__ = ~new_new_n2879__ & new_new_n2880__;
  assign new_new_n2882__ = ~new_new_n2640__ & new_new_n2808__;
  assign new_new_n2883__ = new_new_n810__ & new_new_n2873__;
  assign new_new_n2884__ = ~new_new_n2882__ & new_new_n2883__;
  assign new_new_n2885__ = ~new_new_n2877__ & ~new_new_n2881__;
  assign new_new_n2886__ = ~new_new_n2884__ & new_new_n2885__;
  assign new_new_n2887__ = new_new_n2870__ & ~new_new_n2886__;
  assign new_new_n2888__ = ~new_new_n2870__ & new_new_n2886__;
  assign new_new_n2889__ = ~new_new_n2887__ & ~new_new_n2888__;
  assign new_new_n2890__ = new_new_n2625__ & new_new_n2848__;
  assign new_new_n2891__ = ~new_new_n2618__ & ~new_new_n2847__;
  assign new_new_n2892__ = ~new_new_n2846__ & ~new_new_n2891__;
  assign new_new_n2893__ = ~new_new_n651__ & ~new_new_n2892__;
  assign new_new_n2894__ = new_new_n651__ & new_new_n2892__;
  assign new_new_n2895__ = ~new_new_n2611__ & ~new_new_n2893__;
  assign new_new_n2896__ = ~new_new_n2894__ & new_new_n2895__;
  assign new_new_n2897__ = ~new_new_n2890__ & ~new_new_n2896__;
  assign new_new_n2898__ = ~new_new_n2889__ & new_new_n2897__;
  assign new_new_n2899__ = new_new_n2889__ & ~new_new_n2897__;
  assign new_new_n2900__ = ~new_new_n2898__ & ~new_new_n2899__;
  assign new_new_n2901__ = new_new_n2799__ & ~new_new_n2900__;
  assign new_new_n2902__ = ~new_new_n2799__ & new_new_n2900__;
  assign new_new_n2903__ = ~new_new_n2901__ & ~new_new_n2902__;
  assign new_new_n2904__ = new_new_n2593__ & new_new_n2604__;
  assign new_new_n2905__ = ~new_new_n320__ & new_new_n2600__;
  assign new_new_n2906__ = ~new_new_n2904__ & ~new_new_n2905__;
  assign new_new_n2907__ = new_new_n2590__ & ~new_new_n2655__;
  assign new_new_n2908__ = new_new_n2596__ & new_new_n2907__;
  assign new_new_n2909__ = new_new_n2906__ & ~new_new_n2908__;
  assign new_new_n2910__ = ~new_new_n301__ & ~new_new_n2909__;
  assign new_new_n2911__ = ~new_new_n2590__ & new_new_n2655__;
  assign new_new_n2912__ = new_new_n2596__ & ~new_new_n2911__;
  assign new_new_n2913__ = new_new_n301__ & new_new_n2906__;
  assign new_new_n2914__ = ~new_new_n2912__ & new_new_n2913__;
  assign new_new_n2915__ = ~new_new_n2590__ & ~new_new_n2655__;
  assign new_new_n2916__ = ~new_new_n316__ & ~new_new_n2915__;
  assign new_new_n2917__ = new_new_n2590__ & new_new_n2655__;
  assign new_new_n2918__ = new_new_n316__ & ~new_new_n2917__;
  assign new_new_n2919__ = new_new_n2596__ & ~new_new_n2916__;
  assign new_new_n2920__ = ~new_new_n2918__ & new_new_n2919__;
  assign new_new_n2921__ = ~new_new_n2910__ & ~new_new_n2914__;
  assign new_new_n2922__ = ~new_new_n2920__ & new_new_n2921__;
  assign new_new_n2923__ = new_new_n810__ & new_new_n2855__;
  assign new_new_n2924__ = ~new_new_n2866__ & new_new_n2923__;
  assign new_new_n2925__ = new_new_n2866__ & ~new_new_n2923__;
  assign new_new_n2926__ = ~new_new_n2924__ & ~new_new_n2925__;
  assign new_new_n2927__ = ~new_new_n2922__ & ~new_new_n2926__;
  assign new_new_n2928__ = new_new_n2922__ & new_new_n2926__;
  assign new_new_n2929__ = ~new_new_n320__ & new_new_n2604__;
  assign new_new_n2930__ = new_new_n2593__ & new_new_n2608__;
  assign new_new_n2931__ = ~new_new_n2929__ & ~new_new_n2930__;
  assign new_new_n2932__ = new_new_n2596__ & ~new_new_n2640__;
  assign new_new_n2933__ = ~new_new_n301__ & ~new_new_n2932__;
  assign new_new_n2934__ = ~new_new_n316__ & ~new_new_n2636__;
  assign new_new_n2935__ = new_new_n316__ & ~new_new_n2635__;
  assign new_new_n2936__ = new_new_n2596__ & ~new_new_n2934__;
  assign new_new_n2937__ = ~new_new_n2935__ & new_new_n2936__;
  assign new_new_n2938__ = ~new_new_n2933__ & ~new_new_n2937__;
  assign new_new_n2939__ = new_new_n2931__ & ~new_new_n2938__;
  assign new_new_n2940__ = new_new_n2596__ & new_new_n2600__;
  assign new_new_n2941__ = new_new_n2634__ & new_new_n2940__;
  assign new_new_n2942__ = new_new_n2931__ & ~new_new_n2941__;
  assign new_new_n2943__ = new_new_n301__ & ~new_new_n2942__;
  assign new_new_n2944__ = ~new_new_n2939__ & ~new_new_n2943__;
  assign new_new_n2945__ = new_new_n2593__ & new_new_n2618__;
  assign new_new_n2946__ = ~new_new_n320__ & new_new_n2608__;
  assign new_new_n2947__ = ~new_new_n2945__ & ~new_new_n2946__;
  assign new_new_n2948__ = new_new_n2596__ & new_new_n2841__;
  assign new_new_n2949__ = new_new_n2947__ & ~new_new_n2948__;
  assign new_new_n2950__ = ~new_new_n301__ & ~new_new_n2949__;
  assign new_new_n2951__ = ~new_new_n316__ & ~new_new_n2833__;
  assign new_new_n2952__ = new_new_n316__ & ~new_new_n2835__;
  assign new_new_n2953__ = new_new_n2596__ & ~new_new_n2951__;
  assign new_new_n2954__ = ~new_new_n2952__ & new_new_n2953__;
  assign new_new_n2955__ = new_new_n2596__ & ~new_new_n2830__;
  assign new_new_n2956__ = new_new_n301__ & new_new_n2947__;
  assign new_new_n2957__ = ~new_new_n2955__ & new_new_n2956__;
  assign new_new_n2958__ = ~new_new_n2950__ & ~new_new_n2957__;
  assign new_new_n2959__ = ~new_new_n2954__ & new_new_n2958__;
  assign new_new_n2960__ = new_new_n2596__ & ~new_new_n2611__;
  assign new_new_n2961__ = new_new_n2596__ & new_new_n2625__;
  assign new_new_n2962__ = ~new_new_n311__ & ~new_new_n2618__;
  assign new_new_n2963__ = ~new_new_n318__ & ~new_new_n2962__;
  assign new_new_n2964__ = ~new_new_n316__ & ~new_new_n2963__;
  assign new_new_n2965__ = new_new_n316__ & new_new_n2963__;
  assign new_new_n2966__ = ~new_new_n2611__ & ~new_new_n2964__;
  assign new_new_n2967__ = ~new_new_n2965__ & new_new_n2966__;
  assign new_new_n2968__ = ~new_new_n2961__ & ~new_new_n2967__;
  assign new_new_n2969__ = ~new_new_n301__ & ~new_new_n2960__;
  assign new_new_n2970__ = new_new_n2968__ & new_new_n2969__;
  assign new_new_n2971__ = ~new_new_n320__ & new_new_n2618__;
  assign new_new_n2972__ = new_new_n2593__ & ~new_new_n2611__;
  assign new_new_n2973__ = ~new_new_n1193__ & new_new_n2625__;
  assign new_new_n2974__ = new_new_n2608__ & new_new_n2973__;
  assign new_new_n2975__ = ~new_new_n2608__ & ~new_new_n2973__;
  assign new_new_n2976__ = new_new_n2596__ & ~new_new_n2974__;
  assign new_new_n2977__ = ~new_new_n2975__ & new_new_n2976__;
  assign new_new_n2978__ = ~new_new_n2971__ & ~new_new_n2972__;
  assign new_new_n2979__ = ~new_new_n2977__ & new_new_n2978__;
  assign new_new_n2980__ = new_new_n2970__ & new_new_n2979__;
  assign new_new_n2981__ = ~new_new_n2611__ & new_new_n2808__;
  assign new_new_n2982__ = ~new_new_n2980__ & ~new_new_n2981__;
  assign new_new_n2983__ = new_new_n2959__ & ~new_new_n2982__;
  assign new_new_n2984__ = new_new_n2944__ & ~new_new_n2983__;
  assign new_new_n2985__ = ~new_new_n2944__ & new_new_n2983__;
  assign new_new_n2986__ = new_new_n2625__ & new_new_n2808__;
  assign new_new_n2987__ = ~new_new_n2800__ & ~new_new_n2850__;
  assign new_new_n2988__ = new_new_n816__ & new_new_n2987__;
  assign new_new_n2989__ = ~new_new_n816__ & ~new_new_n2987__;
  assign new_new_n2990__ = ~new_new_n2611__ & ~new_new_n2988__;
  assign new_new_n2991__ = ~new_new_n2989__ & new_new_n2990__;
  assign new_new_n2992__ = ~new_new_n2986__ & ~new_new_n2991__;
  assign new_new_n2993__ = ~new_new_n2985__ & new_new_n2992__;
  assign new_new_n2994__ = ~new_new_n2984__ & ~new_new_n2993__;
  assign new_new_n2995__ = ~new_new_n2928__ & ~new_new_n2994__;
  assign new_new_n2996__ = ~new_new_n2927__ & ~new_new_n2995__;
  assign new_new_n2997__ = new_new_n2849__ & new_new_n2868__;
  assign new_new_n2998__ = ~new_new_n2845__ & ~new_new_n2997__;
  assign new_new_n2999__ = new_new_n2869__ & ~new_new_n2998__;
  assign new_new_n3000__ = ~new_new_n2869__ & new_new_n2998__;
  assign new_new_n3001__ = ~new_new_n2999__ & ~new_new_n3000__;
  assign new_new_n3002__ = ~new_new_n2996__ & ~new_new_n3001__;
  assign new_new_n3003__ = new_new_n2593__ & new_new_n2600__;
  assign new_new_n3004__ = ~new_new_n320__ & new_new_n2590__;
  assign new_new_n3005__ = ~new_new_n3003__ & ~new_new_n3004__;
  assign new_new_n3006__ = new_new_n2585__ & new_new_n2590__;
  assign new_new_n3007__ = new_new_n2604__ & new_new_n3006__;
  assign new_new_n3008__ = ~new_new_n2585__ & new_new_n2644__;
  assign new_new_n3009__ = new_new_n2829__ & new_new_n3008__;
  assign new_new_n3010__ = ~new_new_n3007__ & ~new_new_n3009__;
  assign new_new_n3011__ = new_new_n2608__ & ~new_new_n3010__;
  assign new_new_n3012__ = new_new_n2829__ & new_new_n3006__;
  assign new_new_n3013__ = ~new_new_n3008__ & ~new_new_n3012__;
  assign new_new_n3014__ = new_new_n2604__ & ~new_new_n3013__;
  assign new_new_n3015__ = new_new_n2585__ & ~new_new_n2590__;
  assign new_new_n3016__ = ~new_new_n2604__ & new_new_n3015__;
  assign new_new_n3017__ = new_new_n2590__ & ~new_new_n2600__;
  assign new_new_n3018__ = ~new_new_n2585__ & new_new_n3017__;
  assign new_new_n3019__ = ~new_new_n2829__ & new_new_n3018__;
  assign new_new_n3020__ = ~new_new_n3016__ & ~new_new_n3019__;
  assign new_new_n3021__ = ~new_new_n2608__ & ~new_new_n3020__;
  assign new_new_n3022__ = ~new_new_n2829__ & new_new_n3015__;
  assign new_new_n3023__ = ~new_new_n3018__ & ~new_new_n3022__;
  assign new_new_n3024__ = ~new_new_n2604__ & ~new_new_n3023__;
  assign new_new_n3025__ = ~new_new_n2644__ & ~new_new_n3017__;
  assign new_new_n3026__ = new_new_n2585__ & new_new_n3025__;
  assign new_new_n3027__ = ~new_new_n3011__ & ~new_new_n3026__;
  assign new_new_n3028__ = ~new_new_n3014__ & ~new_new_n3021__;
  assign new_new_n3029__ = ~new_new_n3024__ & new_new_n3028__;
  assign new_new_n3030__ = new_new_n3027__ & new_new_n3029__;
  assign new_new_n3031__ = new_new_n2585__ & ~new_new_n3030__;
  assign new_new_n3032__ = new_new_n2596__ & new_new_n3031__;
  assign new_new_n3033__ = new_new_n3005__ & ~new_new_n3032__;
  assign new_new_n3034__ = new_new_n301__ & ~new_new_n3033__;
  assign new_new_n3035__ = new_new_n2585__ & new_new_n3030__;
  assign new_new_n3036__ = ~new_new_n316__ & ~new_new_n3035__;
  assign new_new_n3037__ = ~new_new_n2585__ & ~new_new_n3030__;
  assign new_new_n3038__ = new_new_n316__ & ~new_new_n3037__;
  assign new_new_n3039__ = new_new_n2596__ & ~new_new_n3036__;
  assign new_new_n3040__ = ~new_new_n3038__ & new_new_n3039__;
  assign new_new_n3041__ = ~new_new_n2585__ & new_new_n3030__;
  assign new_new_n3042__ = new_new_n2596__ & ~new_new_n3041__;
  assign new_new_n3043__ = ~new_new_n301__ & new_new_n3005__;
  assign new_new_n3044__ = ~new_new_n3042__ & new_new_n3043__;
  assign new_new_n3045__ = ~new_new_n3034__ & ~new_new_n3044__;
  assign new_new_n3046__ = ~new_new_n3040__ & new_new_n3045__;
  assign new_new_n3047__ = new_new_n2996__ & new_new_n3001__;
  assign new_new_n3048__ = ~new_new_n3002__ & ~new_new_n3047__;
  assign new_new_n3049__ = new_new_n3046__ & new_new_n3048__;
  assign new_new_n3050__ = ~new_new_n3002__ & ~new_new_n3049__;
  assign new_new_n3051__ = new_new_n2903__ & ~new_new_n3050__;
  assign new_new_n3052__ = ~new_new_n2901__ & ~new_new_n3051__;
  assign new_new_n3053__ = ~new_new_n437__ & ~new_new_n651__;
  assign new_new_n3054__ = new_new_n2846__ & new_new_n3053__;
  assign new_new_n3055__ = ~new_new_n651__ & ~new_new_n2611__;
  assign new_new_n3056__ = new_new_n2847__ & ~new_new_n3055__;
  assign new_new_n3057__ = ~new_new_n437__ & new_new_n2846__;
  assign new_new_n3058__ = ~new_new_n2615__ & ~new_new_n3057__;
  assign new_new_n3059__ = new_new_n2611__ & ~new_new_n3058__;
  assign new_new_n3060__ = ~new_new_n3054__ & ~new_new_n3056__;
  assign new_new_n3061__ = ~new_new_n3059__ & new_new_n3060__;
  assign new_new_n3062__ = ~new_new_n437__ & new_new_n3061__;
  assign new_new_n3063__ = new_new_n437__ & new_new_n651__;
  assign new_new_n3064__ = new_new_n2847__ & new_new_n3063__;
  assign new_new_n3065__ = ~new_new_n3054__ & ~new_new_n3064__;
  assign new_new_n3066__ = ~new_new_n2611__ & ~new_new_n3065__;
  assign new_new_n3067__ = ~new_new_n651__ & ~new_new_n764__;
  assign new_new_n3068__ = new_new_n651__ & new_new_n764__;
  assign new_new_n3069__ = ~new_new_n3067__ & ~new_new_n3068__;
  assign new_new_n3070__ = ~new_new_n2848__ & new_new_n3069__;
  assign new_new_n3071__ = new_new_n2618__ & new_new_n3070__;
  assign new_new_n3072__ = ~new_new_n3053__ & ~new_new_n3063__;
  assign new_new_n3073__ = new_new_n2625__ & ~new_new_n3072__;
  assign new_new_n3074__ = new_new_n2608__ & new_new_n3073__;
  assign new_new_n3075__ = ~new_new_n2608__ & ~new_new_n3073__;
  assign new_new_n3076__ = new_new_n2848__ & ~new_new_n3074__;
  assign new_new_n3077__ = ~new_new_n3075__ & new_new_n3076__;
  assign new_new_n3078__ = ~new_new_n3066__ & ~new_new_n3071__;
  assign new_new_n3079__ = ~new_new_n3077__ & new_new_n3078__;
  assign new_new_n3080__ = new_new_n3062__ & ~new_new_n3079__;
  assign new_new_n3081__ = ~new_new_n3062__ & new_new_n3079__;
  assign new_new_n3082__ = ~new_new_n3080__ & ~new_new_n3081__;
  assign new_new_n3083__ = new_new_n2600__ & new_new_n2809__;
  assign new_new_n3084__ = new_new_n2604__ & ~new_new_n2806__;
  assign new_new_n3085__ = ~new_new_n3083__ & ~new_new_n3084__;
  assign new_new_n3086__ = new_new_n2808__ & ~new_new_n2911__;
  assign new_new_n3087__ = ~new_new_n810__ & ~new_new_n3086__;
  assign new_new_n3088__ = ~new_new_n816__ & new_new_n2808__;
  assign new_new_n3089__ = new_new_n2917__ & new_new_n3088__;
  assign new_new_n3090__ = ~new_new_n3087__ & ~new_new_n3089__;
  assign new_new_n3091__ = new_new_n3085__ & ~new_new_n3090__;
  assign new_new_n3092__ = new_new_n2808__ & new_new_n2907__;
  assign new_new_n3093__ = new_new_n3085__ & ~new_new_n3092__;
  assign new_new_n3094__ = new_new_n810__ & ~new_new_n3093__;
  assign new_new_n3095__ = new_new_n816__ & new_new_n2808__;
  assign new_new_n3096__ = new_new_n2915__ & new_new_n3095__;
  assign new_new_n3097__ = ~new_new_n3094__ & ~new_new_n3096__;
  assign new_new_n3098__ = ~new_new_n3091__ & new_new_n3097__;
  assign new_new_n3099__ = ~new_new_n2888__ & ~new_new_n2897__;
  assign new_new_n3100__ = ~new_new_n2887__ & ~new_new_n3099__;
  assign new_new_n3101__ = ~new_new_n3098__ & new_new_n3100__;
  assign new_new_n3102__ = new_new_n3098__ & ~new_new_n3100__;
  assign new_new_n3103__ = ~new_new_n3101__ & ~new_new_n3102__;
  assign new_new_n3104__ = new_new_n3082__ & new_new_n3103__;
  assign new_new_n3105__ = ~new_new_n3082__ & ~new_new_n3103__;
  assign new_new_n3106__ = ~new_new_n3104__ & ~new_new_n3105__;
  assign new_new_n3107__ = new_new_n3052__ & new_new_n3106__;
  assign new_new_n3108__ = ~new_new_n3052__ & ~new_new_n3106__;
  assign new_new_n3109__ = ~new_new_n2658__ & ~new_new_n2784__;
  assign new_new_n3110__ = ~new_new_n2663__ & new_new_n2784__;
  assign new_new_n3111__ = ~new_new_n3109__ & ~new_new_n3110__;
  assign new_new_n3112__ = new_new_n301__ & ~new_new_n3111__;
  assign new_new_n3113__ = ~new_new_n316__ & new_new_n3111__;
  assign new_new_n3114__ = ~new_new_n785__ & ~new_new_n2753__;
  assign new_new_n3115__ = ~new_new_n2752__ & ~new_new_n3114__;
  assign new_new_n3116__ = ~new_new_n810__ & new_new_n3115__;
  assign new_new_n3117__ = new_new_n810__ & ~new_new_n3115__;
  assign new_new_n3118__ = ~new_new_n648__ & ~new_new_n3116__;
  assign new_new_n3119__ = ~new_new_n3117__ & new_new_n3118__;
  assign new_new_n3120__ = ~new_new_n437__ & new_new_n759__;
  assign new_new_n3121__ = new_new_n1654__ & ~new_new_n3120__;
  assign new_new_n3122__ = new_new_n758__ & new_new_n2731__;
  assign new_new_n3123__ = ~new_new_n3121__ & ~new_new_n3122__;
  assign new_new_n3124__ = ~new_new_n764__ & ~new_new_n791__;
  assign new_new_n3125__ = ~new_new_n648__ & ~new_new_n764__;
  assign new_new_n3126__ = new_new_n805__ & ~new_new_n3125__;
  assign new_new_n3127__ = ~new_new_n651__ & new_new_n792__;
  assign new_new_n3128__ = ~new_new_n3124__ & ~new_new_n3126__;
  assign new_new_n3129__ = ~new_new_n3127__ & new_new_n3128__;
  assign new_new_n3130__ = new_new_n3123__ & ~new_new_n3129__;
  assign new_new_n3131__ = ~new_new_n3123__ & new_new_n3129__;
  assign new_new_n3132__ = ~new_new_n3130__ & ~new_new_n3131__;
  assign new_new_n3133__ = ~new_new_n2738__ & ~new_new_n2745__;
  assign new_new_n3134__ = ~new_new_n2739__ & ~new_new_n3133__;
  assign new_new_n3135__ = new_new_n3132__ & ~new_new_n3134__;
  assign new_new_n3136__ = ~new_new_n3132__ & new_new_n3134__;
  assign new_new_n3137__ = ~new_new_n3135__ & ~new_new_n3136__;
  assign new_new_n3138__ = new_new_n3119__ & new_new_n3137__;
  assign new_new_n3139__ = ~new_new_n3119__ & ~new_new_n3137__;
  assign new_new_n3140__ = ~new_new_n3138__ & ~new_new_n3139__;
  assign new_new_n3141__ = ~new_new_n2750__ & ~new_new_n2758__;
  assign new_new_n3142__ = ~new_new_n2749__ & ~new_new_n3141__;
  assign new_new_n3143__ = new_new_n2773__ & new_new_n3142__;
  assign new_new_n3144__ = new_new_n2774__ & ~new_new_n3142__;
  assign new_new_n3145__ = new_new_n2749__ & ~new_new_n2758__;
  assign new_new_n3146__ = new_new_n2750__ & new_new_n2758__;
  assign new_new_n3147__ = ~new_new_n3145__ & ~new_new_n3146__;
  assign new_new_n3148__ = new_new_n2775__ & new_new_n3147__;
  assign new_new_n3149__ = ~new_new_n3143__ & ~new_new_n3144__;
  assign new_new_n3150__ = ~new_new_n3148__ & new_new_n3149__;
  assign new_new_n3151__ = ~new_new_n3140__ & ~new_new_n3150__;
  assign new_new_n3152__ = ~new_new_n2748__ & new_new_n2772__;
  assign new_new_n3153__ = ~new_new_n2759__ & new_new_n3152__;
  assign new_new_n3154__ = ~new_new_n2728__ & new_new_n3153__;
  assign new_new_n3155__ = new_new_n2748__ & ~new_new_n2772__;
  assign new_new_n3156__ = ~new_new_n2759__ & ~new_new_n3155__;
  assign new_new_n3157__ = ~new_new_n3152__ & ~new_new_n3156__;
  assign new_new_n3158__ = new_new_n2728__ & new_new_n3157__;
  assign new_new_n3159__ = new_new_n2759__ & new_new_n3155__;
  assign new_new_n3160__ = ~new_new_n3158__ & ~new_new_n3159__;
  assign new_new_n3161__ = new_new_n2758__ & ~new_new_n3160__;
  assign new_new_n3162__ = new_new_n2728__ & ~new_new_n3153__;
  assign new_new_n3163__ = ~new_new_n2758__ & ~new_new_n3157__;
  assign new_new_n3164__ = ~new_new_n3162__ & new_new_n3163__;
  assign new_new_n3165__ = new_new_n2728__ & new_new_n2759__;
  assign new_new_n3166__ = new_new_n3155__ & new_new_n3165__;
  assign new_new_n3167__ = ~new_new_n3154__ & ~new_new_n3166__;
  assign new_new_n3168__ = ~new_new_n3164__ & new_new_n3167__;
  assign new_new_n3169__ = ~new_new_n3161__ & new_new_n3168__;
  assign new_new_n3170__ = new_new_n3140__ & ~new_new_n3169__;
  assign new_new_n3171__ = ~new_new_n3151__ & ~new_new_n3170__;
  assign new_new_n3172__ = ~new_new_n2724__ & ~new_new_n2781__;
  assign new_new_n3173__ = ~new_new_n2725__ & ~new_new_n3172__;
  assign new_new_n3174__ = ~new_new_n3171__ & new_new_n3173__;
  assign new_new_n3175__ = new_new_n3171__ & ~new_new_n3173__;
  assign new_new_n3176__ = ~new_new_n3174__ & ~new_new_n3175__;
  assign new_new_n3177__ = ~new_new_n141__ & new_new_n1434__;
  assign new_new_n3178__ = ~new_new_n384__ & ~new_new_n404__;
  assign new_new_n3179__ = ~new_new_n2461__ & new_new_n3178__;
  assign new_new_n3180__ = new_new_n871__ & new_new_n3179__;
  assign new_new_n3181__ = ~new_new_n3177__ & new_new_n3180__;
  assign new_new_n3182__ = ~new_new_n201__ & ~new_new_n373__;
  assign new_new_n3183__ = ~new_new_n457__ & ~new_new_n617__;
  assign new_new_n3184__ = new_new_n3182__ & new_new_n3183__;
  assign new_new_n3185__ = ~new_new_n700__ & new_new_n3184__;
  assign new_new_n3186__ = new_new_n600__ & new_new_n3185__;
  assign new_new_n3187__ = new_new_n3181__ & new_new_n3186__;
  assign new_new_n3188__ = new_new_n81__ & new_new_n213__;
  assign new_new_n3189__ = new_new_n148__ & new_new_n3188__;
  assign new_new_n3190__ = new_new_n116__ & ~new_new_n3189__;
  assign new_new_n3191__ = ~new_new_n224__ & ~new_new_n359__;
  assign new_new_n3192__ = ~new_new_n921__ & new_new_n3191__;
  assign new_new_n3193__ = ~new_new_n861__ & new_new_n2337__;
  assign new_new_n3194__ = ~new_new_n3190__ & new_new_n3193__;
  assign new_new_n3195__ = ~new_new_n523__ & new_new_n3192__;
  assign new_new_n3196__ = new_new_n3194__ & new_new_n3195__;
  assign new_new_n3197__ = new_new_n727__ & new_new_n3196__;
  assign new_new_n3198__ = new_new_n550__ & new_new_n3197__;
  assign new_new_n3199__ = new_new_n2698__ & new_new_n3198__;
  assign new_new_n3200__ = new_new_n3187__ & new_new_n3199__;
  assign new_new_n3201__ = new_new_n3176__ & new_new_n3200__;
  assign new_new_n3202__ = ~new_new_n3176__ & ~new_new_n3200__;
  assign new_new_n3203__ = ~new_new_n3201__ & ~new_new_n3202__;
  assign new_new_n3204__ = ~new_new_n3113__ & ~new_new_n3203__;
  assign new_new_n3205__ = new_new_n3113__ & new_new_n3203__;
  assign new_new_n3206__ = ~new_new_n3204__ & ~new_new_n3205__;
  assign new_new_n3207__ = new_new_n2596__ & ~new_new_n3112__;
  assign new_new_n3208__ = ~new_new_n3206__ & new_new_n3207__;
  assign new_new_n3209__ = new_new_n2585__ & new_new_n2593__;
  assign new_new_n3210__ = ~new_new_n320__ & ~new_new_n2784__;
  assign new_new_n3211__ = ~new_new_n3209__ & ~new_new_n3210__;
  assign new_new_n3212__ = ~new_new_n301__ & ~new_new_n3211__;
  assign new_new_n3213__ = ~new_new_n3111__ & new_new_n3203__;
  assign new_new_n3214__ = new_new_n2596__ & ~new_new_n3213__;
  assign new_new_n3215__ = new_new_n301__ & new_new_n3211__;
  assign new_new_n3216__ = ~new_new_n3214__ & new_new_n3215__;
  assign new_new_n3217__ = ~new_new_n3212__ & ~new_new_n3216__;
  assign new_new_n3218__ = ~new_new_n3208__ & new_new_n3217__;
  assign new_new_n3219__ = ~new_new_n3107__ & ~new_new_n3218__;
  assign new_new_n3220__ = ~new_new_n3108__ & ~new_new_n3219__;
  assign new_new_n3221__ = ~new_new_n3107__ & new_new_n3220__;
  assign new_new_n3222__ = ~new_new_n3108__ & new_new_n3219__;
  assign new_new_n3223__ = ~new_new_n3218__ & ~new_new_n3222__;
  assign new_new_n3224__ = ~new_new_n3221__ & ~new_new_n3223__;
  assign new_new_n3225__ = ~new_new_n2903__ & new_new_n3050__;
  assign new_new_n3226__ = ~new_new_n3051__ & ~new_new_n3225__;
  assign new_new_n3227__ = ~new_new_n3046__ & ~new_new_n3048__;
  assign new_new_n3228__ = ~new_new_n3049__ & ~new_new_n3227__;
  assign new_new_n3229__ = ~pi22 & ~new_new_n57__;
  assign new_new_n3230__ = pi02 & ~new_new_n3229__;
  assign new_new_n3231__ = ~pi02 & ~pi22;
  assign new_new_n3232__ = ~new_new_n57__ & new_new_n3231__;
  assign new_new_n3233__ = ~new_new_n3230__ & ~new_new_n3232__;
  assign new_new_n3234__ = ~new_new_n1573__ & new_new_n3233__;
  assign new_new_n3235__ = new_new_n1573__ & ~new_new_n3233__;
  assign new_new_n3236__ = ~new_new_n3234__ & ~new_new_n3235__;
  assign new_new_n3237__ = new_new_n1324__ & ~new_new_n1573__;
  assign new_new_n3238__ = ~new_new_n1324__ & new_new_n1573__;
  assign new_new_n3239__ = ~new_new_n3237__ & ~new_new_n3238__;
  assign new_new_n3240__ = ~new_new_n3236__ & new_new_n3239__;
  assign new_new_n3241__ = new_new_n2585__ & new_new_n3240__;
  assign new_new_n3242__ = new_new_n1324__ & new_new_n3234__;
  assign new_new_n3243__ = new_new_n310__ & ~new_new_n3242__;
  assign new_new_n3244__ = ~new_new_n310__ & new_new_n3233__;
  assign new_new_n3245__ = ~new_new_n310__ & ~new_new_n3238__;
  assign new_new_n3246__ = ~new_new_n3244__ & ~new_new_n3245__;
  assign new_new_n3247__ = ~new_new_n3243__ & new_new_n3246__;
  assign new_new_n3248__ = new_new_n2590__ & new_new_n3247__;
  assign new_new_n3249__ = ~new_new_n3241__ & ~new_new_n3248__;
  assign new_new_n3250__ = new_new_n2785__ & new_new_n3236__;
  assign new_new_n3251__ = new_new_n3249__ & ~new_new_n3250__;
  assign new_new_n3252__ = new_new_n310__ & ~new_new_n3251__;
  assign new_new_n3253__ = new_new_n1324__ & ~new_new_n2784__;
  assign new_new_n3254__ = ~new_new_n1324__ & new_new_n2784__;
  assign new_new_n3255__ = new_new_n3236__ & ~new_new_n3253__;
  assign new_new_n3256__ = ~new_new_n3254__ & new_new_n3255__;
  assign new_new_n3257__ = new_new_n2664__ & new_new_n3256__;
  assign new_new_n3258__ = ~new_new_n2794__ & new_new_n3236__;
  assign new_new_n3259__ = ~new_new_n310__ & new_new_n3249__;
  assign new_new_n3260__ = ~new_new_n3258__ & new_new_n3259__;
  assign new_new_n3261__ = ~new_new_n3257__ & ~new_new_n3260__;
  assign new_new_n3262__ = ~new_new_n3252__ & new_new_n3261__;
  assign new_new_n3263__ = ~new_new_n2959__ & new_new_n2982__;
  assign new_new_n3264__ = ~new_new_n2983__ & ~new_new_n3263__;
  assign new_new_n3265__ = new_new_n2980__ & new_new_n2981__;
  assign new_new_n3266__ = ~new_new_n3264__ & ~new_new_n3265__;
  assign new_new_n3267__ = ~new_new_n1324__ & new_new_n3236__;
  assign new_new_n3268__ = new_new_n3037__ & new_new_n3267__;
  assign new_new_n3269__ = new_new_n2600__ & new_new_n3247__;
  assign new_new_n3270__ = new_new_n2590__ & new_new_n3240__;
  assign new_new_n3271__ = ~new_new_n3269__ & ~new_new_n3270__;
  assign new_new_n3272__ = ~new_new_n3041__ & new_new_n3236__;
  assign new_new_n3273__ = new_new_n310__ & ~new_new_n3272__;
  assign new_new_n3274__ = new_new_n1324__ & new_new_n3236__;
  assign new_new_n3275__ = new_new_n3035__ & new_new_n3274__;
  assign new_new_n3276__ = ~new_new_n3273__ & ~new_new_n3275__;
  assign new_new_n3277__ = new_new_n3271__ & ~new_new_n3276__;
  assign new_new_n3278__ = new_new_n3031__ & new_new_n3236__;
  assign new_new_n3279__ = new_new_n3271__ & ~new_new_n3278__;
  assign new_new_n3280__ = ~new_new_n310__ & ~new_new_n3279__;
  assign new_new_n3281__ = ~new_new_n3268__ & ~new_new_n3280__;
  assign new_new_n3282__ = ~new_new_n3277__ & new_new_n3281__;
  assign new_new_n3283__ = new_new_n3266__ & new_new_n3282__;
  assign new_new_n3284__ = ~new_new_n3266__ & ~new_new_n3282__;
  assign new_new_n3285__ = new_new_n2604__ & new_new_n3247__;
  assign new_new_n3286__ = new_new_n2600__ & new_new_n3240__;
  assign new_new_n3287__ = ~new_new_n3285__ & ~new_new_n3286__;
  assign new_new_n3288__ = new_new_n2907__ & new_new_n3236__;
  assign new_new_n3289__ = new_new_n3287__ & ~new_new_n3288__;
  assign new_new_n3290__ = ~new_new_n310__ & ~new_new_n3289__;
  assign new_new_n3291__ = ~new_new_n2911__ & new_new_n3236__;
  assign new_new_n3292__ = new_new_n310__ & new_new_n3287__;
  assign new_new_n3293__ = ~new_new_n3291__ & new_new_n3292__;
  assign new_new_n3294__ = ~new_new_n1324__ & ~new_new_n2915__;
  assign new_new_n3295__ = new_new_n1324__ & ~new_new_n2917__;
  assign new_new_n3296__ = new_new_n3236__ & ~new_new_n3294__;
  assign new_new_n3297__ = ~new_new_n3295__ & new_new_n3296__;
  assign new_new_n3298__ = ~new_new_n3290__ & ~new_new_n3293__;
  assign new_new_n3299__ = ~new_new_n3297__ & new_new_n3298__;
  assign new_new_n3300__ = ~new_new_n301__ & ~new_new_n2970__;
  assign new_new_n3301__ = new_new_n2979__ & ~new_new_n3300__;
  assign new_new_n3302__ = ~new_new_n2979__ & new_new_n3300__;
  assign new_new_n3303__ = ~new_new_n3301__ & ~new_new_n3302__;
  assign new_new_n3304__ = new_new_n3299__ & ~new_new_n3303__;
  assign new_new_n3305__ = ~new_new_n3299__ & new_new_n3303__;
  assign new_new_n3306__ = new_new_n310__ & ~new_new_n1324__;
  assign new_new_n3307__ = ~new_new_n310__ & new_new_n1324__;
  assign new_new_n3308__ = ~new_new_n3306__ & ~new_new_n3307__;
  assign new_new_n3309__ = ~new_new_n3239__ & new_new_n3308__;
  assign new_new_n3310__ = new_new_n2608__ & new_new_n3309__;
  assign new_new_n3311__ = new_new_n2604__ & new_new_n3239__;
  assign new_new_n3312__ = ~new_new_n3236__ & ~new_new_n3310__;
  assign new_new_n3313__ = ~new_new_n3311__ & new_new_n3312__;
  assign new_new_n3314__ = new_new_n2640__ & new_new_n3236__;
  assign new_new_n3315__ = ~new_new_n3313__ & ~new_new_n3314__;
  assign new_new_n3316__ = ~new_new_n310__ & ~new_new_n3315__;
  assign new_new_n3317__ = ~new_new_n1324__ & ~new_new_n2636__;
  assign new_new_n3318__ = new_new_n1324__ & ~new_new_n2635__;
  assign new_new_n3319__ = new_new_n3236__ & ~new_new_n3317__;
  assign new_new_n3320__ = ~new_new_n3318__ & new_new_n3319__;
  assign new_new_n3321__ = ~new_new_n2634__ & new_new_n3236__;
  assign new_new_n3322__ = ~new_new_n2600__ & new_new_n3236__;
  assign new_new_n3323__ = new_new_n310__ & ~new_new_n3313__;
  assign new_new_n3324__ = ~new_new_n3322__ & new_new_n3323__;
  assign new_new_n3325__ = ~new_new_n3321__ & new_new_n3324__;
  assign new_new_n3326__ = ~new_new_n3320__ & ~new_new_n3325__;
  assign new_new_n3327__ = ~new_new_n3316__ & new_new_n3326__;
  assign new_new_n3328__ = new_new_n2618__ & new_new_n3247__;
  assign new_new_n3329__ = new_new_n2608__ & new_new_n3240__;
  assign new_new_n3330__ = new_new_n2829__ & new_new_n3308__;
  assign new_new_n3331__ = ~new_new_n2604__ & ~new_new_n3308__;
  assign new_new_n3332__ = new_new_n3236__ & ~new_new_n3331__;
  assign new_new_n3333__ = ~new_new_n3330__ & new_new_n3332__;
  assign new_new_n3334__ = ~new_new_n3328__ & ~new_new_n3329__;
  assign new_new_n3335__ = ~new_new_n3333__ & new_new_n3334__;
  assign new_new_n3336__ = new_new_n310__ & ~new_new_n3335__;
  assign new_new_n3337__ = ~new_new_n3236__ & ~new_new_n3239__;
  assign new_new_n3338__ = new_new_n2611__ & new_new_n2615__;
  assign new_new_n3339__ = ~new_new_n3337__ & ~new_new_n3338__;
  assign new_new_n3340__ = new_new_n3235__ & new_new_n3306__;
  assign new_new_n3341__ = new_new_n2625__ & new_new_n3308__;
  assign new_new_n3342__ = ~new_new_n2608__ & new_new_n3341__;
  assign new_new_n3343__ = new_new_n2608__ & ~new_new_n3341__;
  assign new_new_n3344__ = new_new_n3236__ & ~new_new_n3342__;
  assign new_new_n3345__ = ~new_new_n3343__ & new_new_n3344__;
  assign new_new_n3346__ = ~new_new_n2618__ & new_new_n3240__;
  assign new_new_n3347__ = new_new_n2611__ & new_new_n3337__;
  assign new_new_n3348__ = ~new_new_n3340__ & ~new_new_n3347__;
  assign new_new_n3349__ = ~new_new_n3346__ & new_new_n3348__;
  assign new_new_n3350__ = ~new_new_n3345__ & new_new_n3349__;
  assign new_new_n3351__ = new_new_n310__ & ~new_new_n3339__;
  assign new_new_n3352__ = ~new_new_n3350__ & new_new_n3351__;
  assign new_new_n3353__ = ~new_new_n2960__ & ~new_new_n3352__;
  assign new_new_n3354__ = ~new_new_n310__ & new_new_n3335__;
  assign new_new_n3355__ = ~new_new_n3336__ & ~new_new_n3353__;
  assign new_new_n3356__ = ~new_new_n3354__ & new_new_n3355__;
  assign new_new_n3357__ = ~new_new_n3327__ & ~new_new_n3356__;
  assign new_new_n3358__ = new_new_n3327__ & new_new_n3356__;
  assign new_new_n3359__ = new_new_n2968__ & ~new_new_n3358__;
  assign new_new_n3360__ = ~new_new_n3357__ & ~new_new_n3359__;
  assign new_new_n3361__ = ~new_new_n3305__ & ~new_new_n3360__;
  assign new_new_n3362__ = ~new_new_n3304__ & ~new_new_n3361__;
  assign new_new_n3363__ = ~new_new_n3284__ & ~new_new_n3362__;
  assign new_new_n3364__ = ~new_new_n3283__ & ~new_new_n3363__;
  assign new_new_n3365__ = ~new_new_n3262__ & ~new_new_n3364__;
  assign new_new_n3366__ = new_new_n3262__ & new_new_n3364__;
  assign new_new_n3367__ = ~new_new_n2984__ & ~new_new_n2985__;
  assign new_new_n3368__ = new_new_n2992__ & new_new_n3367__;
  assign new_new_n3369__ = ~new_new_n2992__ & ~new_new_n3367__;
  assign new_new_n3370__ = ~new_new_n3368__ & ~new_new_n3369__;
  assign new_new_n3371__ = ~new_new_n3366__ & new_new_n3370__;
  assign new_new_n3372__ = ~new_new_n3365__ & ~new_new_n3371__;
  assign new_new_n3373__ = new_new_n310__ & ~new_new_n3111__;
  assign new_new_n3374__ = ~new_new_n1324__ & new_new_n3111__;
  assign new_new_n3375__ = ~new_new_n3203__ & ~new_new_n3374__;
  assign new_new_n3376__ = new_new_n3203__ & new_new_n3374__;
  assign new_new_n3377__ = ~new_new_n3375__ & ~new_new_n3376__;
  assign new_new_n3378__ = new_new_n3236__ & ~new_new_n3373__;
  assign new_new_n3379__ = ~new_new_n3377__ & new_new_n3378__;
  assign new_new_n3380__ = new_new_n2585__ & new_new_n3247__;
  assign new_new_n3381__ = ~new_new_n2784__ & new_new_n3240__;
  assign new_new_n3382__ = ~new_new_n3380__ & ~new_new_n3381__;
  assign new_new_n3383__ = ~new_new_n310__ & ~new_new_n3382__;
  assign new_new_n3384__ = ~new_new_n3213__ & new_new_n3236__;
  assign new_new_n3385__ = new_new_n310__ & new_new_n3382__;
  assign new_new_n3386__ = ~new_new_n3384__ & new_new_n3385__;
  assign new_new_n3387__ = ~new_new_n3383__ & ~new_new_n3386__;
  assign new_new_n3388__ = ~new_new_n3379__ & new_new_n3387__;
  assign new_new_n3389__ = ~new_new_n3372__ & new_new_n3388__;
  assign new_new_n3390__ = new_new_n3372__ & ~new_new_n3388__;
  assign new_new_n3391__ = ~new_new_n2927__ & ~new_new_n2928__;
  assign new_new_n3392__ = new_new_n2994__ & ~new_new_n3391__;
  assign new_new_n3393__ = ~new_new_n2994__ & new_new_n3391__;
  assign new_new_n3394__ = ~new_new_n3392__ & ~new_new_n3393__;
  assign new_new_n3395__ = ~new_new_n3390__ & new_new_n3394__;
  assign new_new_n3396__ = ~new_new_n3389__ & ~new_new_n3395__;
  assign new_new_n3397__ = new_new_n3228__ & ~new_new_n3396__;
  assign new_new_n3398__ = ~new_new_n2784__ & new_new_n3247__;
  assign new_new_n3399__ = ~new_new_n3203__ & new_new_n3240__;
  assign new_new_n3400__ = ~new_new_n3398__ & ~new_new_n3399__;
  assign new_new_n3401__ = ~new_new_n3115__ & ~new_new_n3134__;
  assign new_new_n3402__ = new_new_n3115__ & new_new_n3134__;
  assign new_new_n3403__ = new_new_n810__ & new_new_n3132__;
  assign new_new_n3404__ = ~new_new_n3402__ & new_new_n3403__;
  assign new_new_n3405__ = ~new_new_n3401__ & ~new_new_n3404__;
  assign new_new_n3406__ = ~new_new_n648__ & ~new_new_n3405__;
  assign new_new_n3407__ = ~new_new_n648__ & new_new_n810__;
  assign new_new_n3408__ = ~new_new_n648__ & ~new_new_n3115__;
  assign new_new_n3409__ = new_new_n3134__ & ~new_new_n3408__;
  assign new_new_n3410__ = ~new_new_n3132__ & ~new_new_n3407__;
  assign new_new_n3411__ = ~new_new_n3409__ & new_new_n3410__;
  assign new_new_n3412__ = ~new_new_n3406__ & ~new_new_n3411__;
  assign new_new_n3413__ = ~new_new_n3140__ & ~new_new_n3152__;
  assign new_new_n3414__ = ~new_new_n3165__ & ~new_new_n3413__;
  assign new_new_n3415__ = ~new_new_n2758__ & new_new_n3414__;
  assign new_new_n3416__ = new_new_n3140__ & ~new_new_n3165__;
  assign new_new_n3417__ = new_new_n2758__ & ~new_new_n3416__;
  assign new_new_n3418__ = ~new_new_n3155__ & ~new_new_n3417__;
  assign new_new_n3419__ = ~new_new_n3152__ & ~new_new_n3418__;
  assign new_new_n3420__ = new_new_n3140__ & ~new_new_n3419__;
  assign new_new_n3421__ = ~new_new_n3414__ & ~new_new_n3418__;
  assign new_new_n3422__ = ~new_new_n2728__ & ~new_new_n2759__;
  assign new_new_n3423__ = ~new_new_n3421__ & new_new_n3422__;
  assign new_new_n3424__ = ~new_new_n3415__ & ~new_new_n3420__;
  assign new_new_n3425__ = ~new_new_n3423__ & new_new_n3424__;
  assign new_new_n3426__ = new_new_n3412__ & ~new_new_n3425__;
  assign new_new_n3427__ = ~new_new_n3412__ & new_new_n3425__;
  assign new_new_n3428__ = ~new_new_n3426__ & ~new_new_n3427__;
  assign new_new_n3429__ = ~new_new_n648__ & new_new_n2848__;
  assign new_new_n3430__ = ~new_new_n1654__ & ~new_new_n3429__;
  assign new_new_n3431__ = new_new_n805__ & ~new_new_n1478__;
  assign new_new_n3432__ = ~new_new_n651__ & ~new_new_n791__;
  assign new_new_n3433__ = new_new_n437__ & new_new_n791__;
  assign new_new_n3434__ = ~new_new_n3432__ & ~new_new_n3433__;
  assign new_new_n3435__ = new_new_n648__ & ~new_new_n3434__;
  assign new_new_n3436__ = ~new_new_n3431__ & ~new_new_n3435__;
  assign new_new_n3437__ = ~new_new_n3430__ & ~new_new_n3436__;
  assign new_new_n3438__ = new_new_n3430__ & new_new_n3436__;
  assign new_new_n3439__ = new_new_n3130__ & ~new_new_n3438__;
  assign new_new_n3440__ = ~new_new_n3437__ & new_new_n3439__;
  assign new_new_n3441__ = new_new_n810__ & ~new_new_n3430__;
  assign new_new_n3442__ = new_new_n3123__ & new_new_n3441__;
  assign new_new_n3443__ = new_new_n3436__ & new_new_n3442__;
  assign new_new_n3444__ = ~new_new_n3129__ & ~new_new_n3436__;
  assign new_new_n3445__ = new_new_n3430__ & new_new_n3444__;
  assign new_new_n3446__ = ~new_new_n3443__ & ~new_new_n3445__;
  assign new_new_n3447__ = ~new_new_n648__ & ~new_new_n3446__;
  assign new_new_n3448__ = new_new_n648__ & new_new_n3437__;
  assign new_new_n3449__ = ~new_new_n3407__ & new_new_n3438__;
  assign new_new_n3450__ = ~new_new_n3448__ & ~new_new_n3449__;
  assign new_new_n3451__ = new_new_n3129__ & ~new_new_n3450__;
  assign new_new_n3452__ = new_new_n648__ & new_new_n3438__;
  assign new_new_n3453__ = ~new_new_n3437__ & ~new_new_n3452__;
  assign new_new_n3454__ = ~new_new_n3123__ & ~new_new_n3453__;
  assign new_new_n3455__ = ~new_new_n3440__ & ~new_new_n3451__;
  assign new_new_n3456__ = ~new_new_n3454__ & new_new_n3455__;
  assign new_new_n3457__ = ~new_new_n3447__ & new_new_n3456__;
  assign new_new_n3458__ = ~new_new_n3428__ & new_new_n3457__;
  assign new_new_n3459__ = new_new_n3428__ & ~new_new_n3457__;
  assign new_new_n3460__ = ~new_new_n3458__ & ~new_new_n3459__;
  assign new_new_n3461__ = ~new_new_n181__ & ~new_new_n670__;
  assign new_new_n3462__ = ~new_new_n2500__ & ~new_new_n3461__;
  assign new_new_n3463__ = new_new_n116__ & ~new_new_n1066__;
  assign new_new_n3464__ = ~new_new_n163__ & ~new_new_n277__;
  assign new_new_n3465__ = ~new_new_n507__ & ~new_new_n709__;
  assign new_new_n3466__ = ~new_new_n861__ & new_new_n862__;
  assign new_new_n3467__ = ~new_new_n3463__ & new_new_n3466__;
  assign new_new_n3468__ = new_new_n3464__ & new_new_n3465__;
  assign new_new_n3469__ = new_new_n728__ & new_new_n872__;
  assign new_new_n3470__ = ~new_new_n3462__ & new_new_n3469__;
  assign new_new_n3471__ = new_new_n3467__ & new_new_n3468__;
  assign new_new_n3472__ = new_new_n375__ & new_new_n3471__;
  assign new_new_n3473__ = new_new_n723__ & new_new_n3470__;
  assign new_new_n3474__ = new_new_n999__ & new_new_n3473__;
  assign new_new_n3475__ = new_new_n3472__ & new_new_n3474__;
  assign new_new_n3476__ = new_new_n1079__ & new_new_n3475__;
  assign new_new_n3477__ = ~new_new_n3460__ & ~new_new_n3476__;
  assign new_new_n3478__ = new_new_n3460__ & new_new_n3476__;
  assign new_new_n3479__ = ~new_new_n3477__ & ~new_new_n3478__;
  assign new_new_n3480__ = ~new_new_n3174__ & new_new_n3200__;
  assign new_new_n3481__ = ~new_new_n3175__ & ~new_new_n3480__;
  assign new_new_n3482__ = ~new_new_n3479__ & new_new_n3481__;
  assign new_new_n3483__ = ~new_new_n1071__ & ~new_new_n3460__;
  assign new_new_n3484__ = new_new_n3481__ & ~new_new_n3483__;
  assign new_new_n3485__ = new_new_n3479__ & ~new_new_n3484__;
  assign new_new_n3486__ = ~new_new_n3482__ & ~new_new_n3485__;
  assign new_new_n3487__ = ~new_new_n3109__ & new_new_n3203__;
  assign new_new_n3488__ = ~new_new_n3110__ & ~new_new_n3203__;
  assign new_new_n3489__ = ~new_new_n3487__ & ~new_new_n3488__;
  assign new_new_n3490__ = ~new_new_n3486__ & ~new_new_n3489__;
  assign new_new_n3491__ = new_new_n3236__ & new_new_n3490__;
  assign new_new_n3492__ = new_new_n3400__ & ~new_new_n3491__;
  assign new_new_n3493__ = new_new_n310__ & ~new_new_n3492__;
  assign new_new_n3494__ = ~new_new_n1324__ & new_new_n3486__;
  assign new_new_n3495__ = new_new_n1324__ & ~new_new_n3486__;
  assign new_new_n3496__ = new_new_n3236__ & ~new_new_n3494__;
  assign new_new_n3497__ = ~new_new_n3495__ & new_new_n3496__;
  assign new_new_n3498__ = new_new_n3489__ & new_new_n3497__;
  assign new_new_n3499__ = new_new_n3486__ & ~new_new_n3489__;
  assign new_new_n3500__ = new_new_n3236__ & ~new_new_n3499__;
  assign new_new_n3501__ = ~new_new_n310__ & new_new_n3400__;
  assign new_new_n3502__ = ~new_new_n3500__ & new_new_n3501__;
  assign new_new_n3503__ = ~new_new_n3498__ & ~new_new_n3502__;
  assign new_new_n3504__ = ~new_new_n3493__ & new_new_n3503__;
  assign new_new_n3505__ = ~new_new_n3228__ & new_new_n3396__;
  assign new_new_n3506__ = ~new_new_n3504__ & ~new_new_n3505__;
  assign new_new_n3507__ = ~new_new_n3397__ & ~new_new_n3506__;
  assign new_new_n3508__ = ~new_new_n3226__ & new_new_n3507__;
  assign new_new_n3509__ = new_new_n3226__ & ~new_new_n3507__;
  assign new_new_n3510__ = ~new_new_n3203__ & new_new_n3247__;
  assign new_new_n3511__ = new_new_n3240__ & ~new_new_n3486__;
  assign new_new_n3512__ = ~new_new_n3510__ & ~new_new_n3511__;
  assign new_new_n3513__ = ~new_new_n3486__ & ~new_new_n3487__;
  assign new_new_n3514__ = new_new_n3486__ & ~new_new_n3488__;
  assign new_new_n3515__ = ~new_new_n3513__ & ~new_new_n3514__;
  assign new_new_n3516__ = ~new_new_n115__ & ~new_new_n448__;
  assign new_new_n3517__ = new_new_n256__ & new_new_n270__;
  assign new_new_n3518__ = new_new_n100__ & ~new_new_n3517__;
  assign new_new_n3519__ = ~new_new_n89__ & ~new_new_n1124__;
  assign new_new_n3520__ = ~new_new_n507__ & new_new_n3519__;
  assign new_new_n3521__ = ~new_new_n3518__ & new_new_n3520__;
  assign new_new_n3522__ = new_new_n110__ & new_new_n148__;
  assign new_new_n3523__ = new_new_n181__ & ~new_new_n3522__;
  assign new_new_n3524__ = new_new_n100__ & ~new_new_n663__;
  assign new_new_n3525__ = new_new_n213__ & new_new_n227__;
  assign new_new_n3526__ = new_new_n195__ & ~new_new_n3525__;
  assign new_new_n3527__ = ~new_new_n373__ & ~new_new_n3524__;
  assign new_new_n3528__ = ~new_new_n3523__ & new_new_n3527__;
  assign new_new_n3529__ = ~new_new_n3526__ & new_new_n3528__;
  assign new_new_n3530__ = ~new_new_n3516__ & new_new_n3529__;
  assign new_new_n3531__ = new_new_n3521__ & new_new_n3530__;
  assign new_new_n3532__ = ~new_new_n343__ & ~new_new_n347__;
  assign new_new_n3533__ = ~new_new_n238__ & new_new_n736__;
  assign new_new_n3534__ = ~new_new_n2321__ & ~new_new_n3533__;
  assign new_new_n3535__ = new_new_n731__ & new_new_n3534__;
  assign new_new_n3536__ = ~new_new_n176__ & ~new_new_n559__;
  assign new_new_n3537__ = ~new_new_n328__ & ~new_new_n925__;
  assign new_new_n3538__ = ~new_new_n976__ & new_new_n3537__;
  assign new_new_n3539__ = ~new_new_n240__ & new_new_n3536__;
  assign new_new_n3540__ = ~new_new_n498__ & ~new_new_n3532__;
  assign new_new_n3541__ = new_new_n3539__ & new_new_n3540__;
  assign new_new_n3542__ = new_new_n3538__ & new_new_n3541__;
  assign new_new_n3543__ = new_new_n3535__ & new_new_n3542__;
  assign new_new_n3544__ = new_new_n402__ & new_new_n2706__;
  assign new_new_n3545__ = new_new_n3543__ & new_new_n3544__;
  assign new_new_n3546__ = new_new_n3531__ & new_new_n3545__;
  assign new_new_n3547__ = new_new_n2423__ & new_new_n3546__;
  assign new_new_n3548__ = ~new_new_n3478__ & new_new_n3484__;
  assign new_new_n3549__ = ~new_new_n3477__ & ~new_new_n3548__;
  assign new_new_n3550__ = new_new_n3547__ & new_new_n3549__;
  assign new_new_n3551__ = ~new_new_n3547__ & ~new_new_n3549__;
  assign new_new_n3552__ = ~new_new_n3550__ & ~new_new_n3551__;
  assign new_new_n3553__ = new_new_n651__ & ~new_new_n3433__;
  assign new_new_n3554__ = new_new_n1654__ & ~new_new_n2847__;
  assign new_new_n3555__ = ~new_new_n2846__ & ~new_new_n3554__;
  assign new_new_n3556__ = ~new_new_n3553__ & ~new_new_n3555__;
  assign new_new_n3557__ = ~new_new_n651__ & new_new_n3433__;
  assign new_new_n3558__ = ~new_new_n648__ & ~new_new_n3557__;
  assign new_new_n3559__ = ~new_new_n3556__ & new_new_n3558__;
  assign new_new_n3560__ = new_new_n791__ & new_new_n3559__;
  assign new_new_n3561__ = new_new_n437__ & ~new_new_n648__;
  assign new_new_n3562__ = ~new_new_n3555__ & new_new_n3561__;
  assign new_new_n3563__ = ~new_new_n3560__ & ~new_new_n3562__;
  assign new_new_n3564__ = ~new_new_n651__ & ~new_new_n3563__;
  assign new_new_n3565__ = ~new_new_n437__ & ~new_new_n791__;
  assign new_new_n3566__ = ~new_new_n3559__ & ~new_new_n3565__;
  assign new_new_n3567__ = ~new_new_n437__ & ~new_new_n3555__;
  assign new_new_n3568__ = ~new_new_n648__ & ~new_new_n3433__;
  assign new_new_n3569__ = ~new_new_n3567__ & new_new_n3568__;
  assign new_new_n3570__ = ~new_new_n3566__ & ~new_new_n3569__;
  assign new_new_n3571__ = ~new_new_n3564__ & ~new_new_n3570__;
  assign new_new_n3572__ = ~new_new_n3442__ & ~new_new_n3444__;
  assign new_new_n3573__ = ~new_new_n648__ & ~new_new_n3572__;
  assign new_new_n3574__ = ~new_new_n3437__ & ~new_new_n3439__;
  assign new_new_n3575__ = ~new_new_n3573__ & new_new_n3574__;
  assign new_new_n3576__ = new_new_n3571__ & new_new_n3575__;
  assign new_new_n3577__ = ~new_new_n3571__ & ~new_new_n3575__;
  assign new_new_n3578__ = ~new_new_n3576__ & ~new_new_n3577__;
  assign new_new_n3579__ = ~new_new_n3427__ & new_new_n3457__;
  assign new_new_n3580__ = ~new_new_n3426__ & ~new_new_n3579__;
  assign new_new_n3581__ = new_new_n3578__ & ~new_new_n3580__;
  assign new_new_n3582__ = ~new_new_n3578__ & new_new_n3580__;
  assign new_new_n3583__ = ~new_new_n3581__ & ~new_new_n3582__;
  assign new_new_n3584__ = new_new_n3552__ & ~new_new_n3583__;
  assign new_new_n3585__ = ~new_new_n3552__ & new_new_n3583__;
  assign new_new_n3586__ = ~new_new_n3584__ & ~new_new_n3585__;
  assign new_new_n3587__ = ~new_new_n3515__ & ~new_new_n3586__;
  assign new_new_n3588__ = new_new_n3236__ & new_new_n3587__;
  assign new_new_n3589__ = new_new_n3512__ & ~new_new_n3588__;
  assign new_new_n3590__ = ~new_new_n310__ & ~new_new_n3589__;
  assign new_new_n3591__ = new_new_n1324__ & new_new_n3586__;
  assign new_new_n3592__ = ~new_new_n1324__ & ~new_new_n3586__;
  assign new_new_n3593__ = new_new_n3236__ & new_new_n3515__;
  assign new_new_n3594__ = ~new_new_n3591__ & ~new_new_n3592__;
  assign new_new_n3595__ = new_new_n3593__ & new_new_n3594__;
  assign new_new_n3596__ = ~new_new_n3515__ & new_new_n3586__;
  assign new_new_n3597__ = new_new_n3236__ & ~new_new_n3596__;
  assign new_new_n3598__ = new_new_n310__ & new_new_n3512__;
  assign new_new_n3599__ = ~new_new_n3597__ & new_new_n3598__;
  assign new_new_n3600__ = ~new_new_n3595__ & ~new_new_n3599__;
  assign new_new_n3601__ = ~new_new_n3590__ & new_new_n3600__;
  assign new_new_n3602__ = ~new_new_n3509__ & ~new_new_n3601__;
  assign new_new_n3603__ = ~new_new_n3508__ & ~new_new_n3602__;
  assign new_new_n3604__ = new_new_n310__ & new_new_n3240__;
  assign new_new_n3605__ = ~new_new_n3586__ & new_new_n3604__;
  assign new_new_n3606__ = ~new_new_n3236__ & ~new_new_n3238__;
  assign new_new_n3607__ = new_new_n3586__ & new_new_n3606__;
  assign new_new_n3608__ = new_new_n3235__ & new_new_n3494__;
  assign new_new_n3609__ = ~new_new_n3242__ & ~new_new_n3608__;
  assign new_new_n3610__ = ~new_new_n3607__ & new_new_n3609__;
  assign new_new_n3611__ = ~new_new_n310__ & ~new_new_n3610__;
  assign new_new_n3612__ = ~new_new_n3605__ & ~new_new_n3611__;
  assign new_new_n3613__ = ~new_new_n3236__ & ~new_new_n3612__;
  assign new_new_n3614__ = new_new_n3234__ & new_new_n3495__;
  assign new_new_n3615__ = new_new_n181__ & ~new_new_n256__;
  assign new_new_n3616__ = ~new_new_n351__ & ~new_new_n3615__;
  assign new_new_n3617__ = new_new_n181__ & ~new_new_n1021__;
  assign new_new_n3618__ = ~new_new_n918__ & ~new_new_n976__;
  assign new_new_n3619__ = ~new_new_n2234__ & new_new_n3618__;
  assign new_new_n3620__ = ~new_new_n3617__ & new_new_n3619__;
  assign new_new_n3621__ = new_new_n125__ & ~new_new_n589__;
  assign new_new_n3622__ = ~new_new_n323__ & ~new_new_n877__;
  assign new_new_n3623__ = new_new_n112__ & new_new_n3622__;
  assign new_new_n3624__ = ~new_new_n2321__ & new_new_n3616__;
  assign new_new_n3625__ = ~new_new_n3621__ & new_new_n3624__;
  assign new_new_n3626__ = new_new_n3623__ & new_new_n3625__;
  assign new_new_n3627__ = new_new_n264__ & new_new_n3620__;
  assign new_new_n3628__ = new_new_n3626__ & new_new_n3627__;
  assign new_new_n3629__ = new_new_n869__ & new_new_n3628__;
  assign new_new_n3630__ = new_new_n1032__ & new_new_n3629__;
  assign new_new_n3631__ = new_new_n2260__ & new_new_n3630__;
  assign new_new_n3632__ = ~new_new_n3550__ & new_new_n3583__;
  assign new_new_n3633__ = ~new_new_n3551__ & ~new_new_n3632__;
  assign new_new_n3634__ = new_new_n3631__ & new_new_n3633__;
  assign new_new_n3635__ = ~new_new_n3631__ & ~new_new_n3633__;
  assign new_new_n3636__ = ~new_new_n3634__ & ~new_new_n3635__;
  assign new_new_n3637__ = ~new_new_n3566__ & ~new_new_n3580__;
  assign new_new_n3638__ = ~new_new_n3571__ & new_new_n3637__;
  assign new_new_n3639__ = ~new_new_n3571__ & new_new_n3580__;
  assign new_new_n3640__ = ~new_new_n3637__ & ~new_new_n3639__;
  assign new_new_n3641__ = ~new_new_n3575__ & ~new_new_n3640__;
  assign new_new_n3642__ = ~new_new_n3576__ & ~new_new_n3580__;
  assign new_new_n3643__ = new_new_n3566__ & ~new_new_n3642__;
  assign new_new_n3644__ = ~new_new_n3638__ & ~new_new_n3643__;
  assign new_new_n3645__ = ~new_new_n3641__ & new_new_n3644__;
  assign new_new_n3646__ = new_new_n3636__ & ~new_new_n3645__;
  assign new_new_n3647__ = ~new_new_n3566__ & new_new_n3642__;
  assign new_new_n3648__ = ~new_new_n3577__ & ~new_new_n3643__;
  assign new_new_n3649__ = ~new_new_n3647__ & new_new_n3648__;
  assign new_new_n3650__ = ~new_new_n3636__ & new_new_n3649__;
  assign new_new_n3651__ = ~new_new_n3646__ & ~new_new_n3650__;
  assign new_new_n3652__ = ~new_new_n3513__ & new_new_n3586__;
  assign new_new_n3653__ = ~new_new_n3514__ & ~new_new_n3586__;
  assign new_new_n3654__ = ~new_new_n3652__ & ~new_new_n3653__;
  assign new_new_n3655__ = ~new_new_n1324__ & new_new_n3654__;
  assign new_new_n3656__ = new_new_n310__ & ~new_new_n3654__;
  assign new_new_n3657__ = ~new_new_n3655__ & ~new_new_n3656__;
  assign new_new_n3658__ = ~new_new_n3651__ & ~new_new_n3657__;
  assign new_new_n3659__ = new_new_n3651__ & new_new_n3657__;
  assign new_new_n3660__ = new_new_n3236__ & new_new_n3612__;
  assign new_new_n3661__ = ~new_new_n3658__ & new_new_n3660__;
  assign new_new_n3662__ = ~new_new_n3659__ & new_new_n3661__;
  assign new_new_n3663__ = ~new_new_n3613__ & ~new_new_n3614__;
  assign new_new_n3664__ = ~new_new_n3662__ & new_new_n3663__;
  assign new_new_n3665__ = ~new_new_n3603__ & new_new_n3664__;
  assign new_new_n3666__ = new_new_n3603__ & ~new_new_n3664__;
  assign new_new_n3667__ = ~new_new_n3665__ & ~new_new_n3666__;
  assign new_new_n3668__ = new_new_n3224__ & new_new_n3667__;
  assign new_new_n3669__ = ~new_new_n3224__ & ~new_new_n3667__;
  assign new_new_n3670__ = ~new_new_n3668__ & ~new_new_n3669__;
  assign new_new_n3671__ = ~new_new_n3634__ & ~new_new_n3649__;
  assign new_new_n3672__ = ~new_new_n3635__ & ~new_new_n3671__;
  assign new_new_n3673__ = new_new_n166__ & new_new_n629__;
  assign new_new_n3674__ = ~new_new_n343__ & ~new_new_n3673__;
  assign new_new_n3675__ = new_new_n181__ & ~new_new_n2446__;
  assign new_new_n3676__ = ~new_new_n115__ & ~new_new_n2683__;
  assign new_new_n3677__ = new_new_n110__ & new_new_n347__;
  assign new_new_n3678__ = new_new_n629__ & new_new_n3677__;
  assign new_new_n3679__ = new_new_n125__ & ~new_new_n3678__;
  assign new_new_n3680__ = ~new_new_n337__ & ~new_new_n409__;
  assign new_new_n3681__ = ~new_new_n2321__ & new_new_n3680__;
  assign new_new_n3682__ = ~new_new_n3676__ & ~new_new_n3679__;
  assign new_new_n3683__ = new_new_n3681__ & new_new_n3682__;
  assign new_new_n3684__ = new_new_n894__ & ~new_new_n3675__;
  assign new_new_n3685__ = ~new_new_n3674__ & new_new_n3684__;
  assign new_new_n3686__ = new_new_n740__ & new_new_n3685__;
  assign new_new_n3687__ = new_new_n1071__ & new_new_n3683__;
  assign new_new_n3688__ = new_new_n3686__ & new_new_n3687__;
  assign new_new_n3689__ = new_new_n1462__ & new_new_n2316__;
  assign new_new_n3690__ = new_new_n3688__ & new_new_n3689__;
  assign new_new_n3691__ = new_new_n3672__ & new_new_n3690__;
  assign new_new_n3692__ = ~new_new_n195__ & new_new_n270__;
  assign new_new_n3693__ = ~new_new_n227__ & ~new_new_n3692__;
  assign new_new_n3694__ = ~new_new_n176__ & ~new_new_n2343__;
  assign new_new_n3695__ = ~new_new_n3693__ & new_new_n3694__;
  assign new_new_n3696__ = new_new_n227__ & ~new_new_n595__;
  assign new_new_n3697__ = new_new_n99__ & ~new_new_n162__;
  assign new_new_n3698__ = ~new_new_n3696__ & ~new_new_n3697__;
  assign new_new_n3699__ = new_new_n223__ & ~new_new_n1051__;
  assign new_new_n3700__ = ~new_new_n596__ & ~new_new_n3699__;
  assign new_new_n3701__ = ~new_new_n893__ & ~new_new_n2230__;
  assign new_new_n3702__ = new_new_n3700__ & new_new_n3701__;
  assign new_new_n3703__ = new_new_n160__ & ~new_new_n475__;
  assign new_new_n3704__ = ~new_new_n455__ & ~new_new_n3703__;
  assign new_new_n3705__ = ~new_new_n89__ & ~new_new_n257__;
  assign new_new_n3706__ = ~new_new_n2461__ & ~new_new_n2565__;
  assign new_new_n3707__ = new_new_n3705__ & new_new_n3706__;
  assign new_new_n3708__ = ~new_new_n3704__ & new_new_n3707__;
  assign new_new_n3709__ = new_new_n3535__ & ~new_new_n3698__;
  assign new_new_n3710__ = new_new_n3702__ & new_new_n3709__;
  assign new_new_n3711__ = new_new_n3708__ & new_new_n3710__;
  assign new_new_n3712__ = new_new_n160__ & new_new_n3188__;
  assign new_new_n3713__ = new_new_n223__ & ~new_new_n3712__;
  assign new_new_n3714__ = ~new_new_n187__ & ~new_new_n560__;
  assign new_new_n3715__ = ~new_new_n546__ & new_new_n3714__;
  assign new_new_n3716__ = ~new_new_n617__ & ~new_new_n3713__;
  assign new_new_n3717__ = new_new_n3715__ & new_new_n3716__;
  assign new_new_n3718__ = new_new_n151__ & ~new_new_n523__;
  assign new_new_n3719__ = new_new_n2324__ & new_new_n3718__;
  assign new_new_n3720__ = new_new_n3695__ & new_new_n3717__;
  assign new_new_n3721__ = new_new_n3719__ & new_new_n3720__;
  assign new_new_n3722__ = new_new_n382__ & new_new_n3721__;
  assign new_new_n3723__ = new_new_n358__ & new_new_n3722__;
  assign new_new_n3724__ = new_new_n3711__ & new_new_n3723__;
  assign new_new_n3725__ = ~new_new_n3691__ & ~new_new_n3724__;
  assign new_new_n3726__ = new_new_n3691__ & new_new_n3724__;
  assign new_new_n3727__ = ~new_new_n3725__ & ~new_new_n3726__;
  assign new_new_n3728__ = pi00 & pi01;
  assign new_new_n3729__ = pi02 & new_new_n3728__;
  assign new_new_n3730__ = ~new_new_n1568__ & ~new_new_n3729__;
  assign new_new_n3731__ = ~new_new_n3727__ & ~new_new_n3730__;
  assign new_new_n3732__ = ~new_new_n3672__ & ~new_new_n3690__;
  assign new_new_n3733__ = ~new_new_n3691__ & ~new_new_n3732__;
  assign new_new_n3734__ = pi01 & new_new_n3733__;
  assign new_new_n3735__ = ~pi01 & pi02;
  assign new_new_n3736__ = ~new_new_n3651__ & new_new_n3735__;
  assign new_new_n3737__ = ~pi00 & ~new_new_n3736__;
  assign new_new_n3738__ = ~new_new_n3734__ & new_new_n3737__;
  assign new_new_n3739__ = ~new_new_n3731__ & ~new_new_n3738__;
  assign new_new_n3740__ = new_new_n3651__ & ~new_new_n3652__;
  assign new_new_n3741__ = new_new_n3724__ & ~new_new_n3740__;
  assign new_new_n3742__ = ~new_new_n3652__ & ~new_new_n3724__;
  assign new_new_n3743__ = new_new_n3733__ & ~new_new_n3742__;
  assign new_new_n3744__ = ~new_new_n3741__ & new_new_n3743__;
  assign new_new_n3745__ = ~new_new_n3651__ & ~new_new_n3653__;
  assign new_new_n3746__ = new_new_n3672__ & new_new_n3724__;
  assign new_new_n3747__ = ~new_new_n3672__ & ~new_new_n3724__;
  assign new_new_n3748__ = ~new_new_n3746__ & ~new_new_n3747__;
  assign new_new_n3749__ = ~new_new_n3733__ & ~new_new_n3745__;
  assign new_new_n3750__ = ~new_new_n3748__ & new_new_n3749__;
  assign new_new_n3751__ = ~new_new_n3653__ & ~new_new_n3747__;
  assign new_new_n3752__ = ~new_new_n3733__ & ~new_new_n3751__;
  assign new_new_n3753__ = new_new_n3724__ & ~new_new_n3732__;
  assign new_new_n3754__ = ~new_new_n3651__ & ~new_new_n3753__;
  assign new_new_n3755__ = ~new_new_n3752__ & new_new_n3754__;
  assign new_new_n3756__ = ~new_new_n3744__ & ~new_new_n3750__;
  assign new_new_n3757__ = ~new_new_n3755__ & new_new_n3756__;
  assign new_new_n3758__ = ~new_new_n3231__ & new_new_n3757__;
  assign new_new_n3759__ = ~pi01 & ~pi22;
  assign new_new_n3760__ = pi01 & pi22;
  assign new_new_n3761__ = ~new_new_n3759__ & ~new_new_n3760__;
  assign new_new_n3762__ = ~new_new_n3757__ & new_new_n3761__;
  assign new_new_n3763__ = pi00 & ~new_new_n3758__;
  assign new_new_n3764__ = ~new_new_n3762__ & new_new_n3763__;
  assign new_new_n3765__ = pi02 & pi22;
  assign new_new_n3766__ = ~pi01 & ~new_new_n3757__;
  assign new_new_n3767__ = new_new_n3765__ & ~new_new_n3766__;
  assign new_new_n3768__ = ~pi02 & pi22;
  assign new_new_n3769__ = pi01 & ~pi02;
  assign new_new_n3770__ = ~new_new_n3735__ & ~new_new_n3769__;
  assign new_new_n3771__ = ~pi00 & ~new_new_n3768__;
  assign new_new_n3772__ = ~new_new_n3770__ & new_new_n3771__;
  assign new_new_n3773__ = ~new_new_n3767__ & ~new_new_n3772__;
  assign new_new_n3774__ = ~new_new_n3764__ & new_new_n3773__;
  assign new_new_n3775__ = new_new_n3739__ & ~new_new_n3774__;
  assign new_new_n3776__ = ~new_new_n3231__ & ~new_new_n3765__;
  assign new_new_n3777__ = ~new_new_n3759__ & new_new_n3776__;
  assign new_new_n3778__ = ~new_new_n1569__ & new_new_n3777__;
  assign new_new_n3779__ = ~new_new_n3739__ & new_new_n3778__;
  assign new_new_n3780__ = ~new_new_n3775__ & ~new_new_n3779__;
  assign new_new_n3781__ = pi01 & ~new_new_n3586__;
  assign new_new_n3782__ = ~new_new_n3486__ & new_new_n3735__;
  assign new_new_n3783__ = ~new_new_n3781__ & ~new_new_n3782__;
  assign new_new_n3784__ = ~new_new_n3233__ & ~new_new_n3783__;
  assign new_new_n3785__ = new_new_n3233__ & new_new_n3783__;
  assign new_new_n3786__ = ~pi00 & ~new_new_n3784__;
  assign new_new_n3787__ = ~new_new_n3785__ & new_new_n3786__;
  assign new_new_n3788__ = new_new_n3654__ & ~new_new_n3770__;
  assign new_new_n3789__ = new_new_n3233__ & ~new_new_n3788__;
  assign new_new_n3790__ = ~new_new_n3233__ & new_new_n3788__;
  assign new_new_n3791__ = ~new_new_n3789__ & ~new_new_n3790__;
  assign new_new_n3792__ = new_new_n3651__ & new_new_n3791__;
  assign new_new_n3793__ = ~new_new_n3651__ & ~new_new_n3791__;
  assign new_new_n3794__ = pi00 & ~new_new_n3792__;
  assign new_new_n3795__ = ~new_new_n3793__ & new_new_n3794__;
  assign new_new_n3796__ = ~new_new_n3787__ & ~new_new_n3795__;
  assign new_new_n3797__ = new_new_n3489__ & ~new_new_n3770__;
  assign new_new_n3798__ = new_new_n3486__ & new_new_n3797__;
  assign new_new_n3799__ = ~new_new_n3486__ & ~new_new_n3797__;
  assign new_new_n3800__ = pi00 & ~new_new_n3798__;
  assign new_new_n3801__ = ~new_new_n3799__ & new_new_n3800__;
  assign new_new_n3802__ = ~new_new_n2784__ & new_new_n3735__;
  assign new_new_n3803__ = pi01 & ~new_new_n3203__;
  assign new_new_n3804__ = ~pi00 & ~new_new_n3802__;
  assign new_new_n3805__ = ~new_new_n3803__ & new_new_n3804__;
  assign new_new_n3806__ = ~new_new_n3801__ & ~new_new_n3805__;
  assign new_new_n3807__ = ~new_new_n3283__ & ~new_new_n3284__;
  assign new_new_n3808__ = ~new_new_n3362__ & new_new_n3807__;
  assign new_new_n3809__ = new_new_n3362__ & ~new_new_n3807__;
  assign new_new_n3810__ = ~new_new_n3808__ & ~new_new_n3809__;
  assign new_new_n3811__ = ~new_new_n3233__ & new_new_n3810__;
  assign new_new_n3812__ = pi01 & new_new_n2585__;
  assign new_new_n3813__ = new_new_n2590__ & new_new_n3735__;
  assign new_new_n3814__ = ~new_new_n3812__ & ~new_new_n3813__;
  assign new_new_n3815__ = ~new_new_n3233__ & ~new_new_n3814__;
  assign new_new_n3816__ = new_new_n3233__ & new_new_n3814__;
  assign new_new_n3817__ = ~pi00 & ~new_new_n3815__;
  assign new_new_n3818__ = ~new_new_n3816__ & new_new_n3817__;
  assign new_new_n3819__ = new_new_n2664__ & ~new_new_n3770__;
  assign new_new_n3820__ = ~new_new_n2784__ & new_new_n3233__;
  assign new_new_n3821__ = new_new_n2784__ & ~new_new_n3233__;
  assign new_new_n3822__ = ~new_new_n3820__ & ~new_new_n3821__;
  assign new_new_n3823__ = new_new_n3819__ & ~new_new_n3822__;
  assign new_new_n3824__ = ~new_new_n3819__ & new_new_n3822__;
  assign new_new_n3825__ = pi00 & ~new_new_n3823__;
  assign new_new_n3826__ = ~new_new_n3824__ & new_new_n3825__;
  assign new_new_n3827__ = ~new_new_n3818__ & ~new_new_n3826__;
  assign new_new_n3828__ = new_new_n3335__ & ~new_new_n3352__;
  assign new_new_n3829__ = ~new_new_n308__ & ~new_new_n2611__;
  assign new_new_n3830__ = ~new_new_n3828__ & new_new_n3829__;
  assign new_new_n3831__ = ~new_new_n310__ & new_new_n2611__;
  assign new_new_n3832__ = ~new_new_n3829__ & ~new_new_n3831__;
  assign new_new_n3833__ = new_new_n3828__ & new_new_n3832__;
  assign new_new_n3834__ = new_new_n310__ & ~new_new_n3352__;
  assign new_new_n3835__ = new_new_n2611__ & ~new_new_n3834__;
  assign new_new_n3836__ = ~new_new_n3335__ & new_new_n3835__;
  assign new_new_n3837__ = ~new_new_n3830__ & ~new_new_n3836__;
  assign new_new_n3838__ = ~new_new_n3833__ & new_new_n3837__;
  assign new_new_n3839__ = pi00 & new_new_n3770__;
  assign new_new_n3840__ = new_new_n2585__ & new_new_n3839__;
  assign new_new_n3841__ = new_new_n2600__ & new_new_n3735__;
  assign new_new_n3842__ = pi01 & new_new_n2590__;
  assign new_new_n3843__ = ~new_new_n3841__ & ~new_new_n3842__;
  assign new_new_n3844__ = ~pi00 & ~new_new_n3843__;
  assign new_new_n3845__ = ~new_new_n3840__ & ~new_new_n3844__;
  assign new_new_n3846__ = ~pi01 & ~new_new_n3030__;
  assign new_new_n3847__ = new_new_n3765__ & ~new_new_n3846__;
  assign new_new_n3848__ = ~new_new_n3030__ & new_new_n3761__;
  assign new_new_n3849__ = new_new_n3030__ & ~new_new_n3231__;
  assign new_new_n3850__ = pi00 & ~new_new_n3848__;
  assign new_new_n3851__ = ~new_new_n3849__ & new_new_n3850__;
  assign new_new_n3852__ = ~new_new_n3772__ & ~new_new_n3847__;
  assign new_new_n3853__ = ~new_new_n3851__ & new_new_n3852__;
  assign new_new_n3854__ = new_new_n3845__ & ~new_new_n3853__;
  assign new_new_n3855__ = pi00 & ~new_new_n3030__;
  assign new_new_n3856__ = new_new_n3735__ & ~new_new_n3855__;
  assign new_new_n3857__ = new_new_n3776__ & ~new_new_n3845__;
  assign new_new_n3858__ = ~new_new_n3856__ & new_new_n3857__;
  assign new_new_n3859__ = ~new_new_n3854__ & ~new_new_n3858__;
  assign new_new_n3860__ = new_new_n3838__ & new_new_n3859__;
  assign new_new_n3861__ = new_new_n2625__ & new_new_n3236__;
  assign new_new_n3862__ = new_new_n2618__ & ~new_new_n3234__;
  assign new_new_n3863__ = ~new_new_n3235__ & ~new_new_n3862__;
  assign new_new_n3864__ = new_new_n1324__ & new_new_n3863__;
  assign new_new_n3865__ = ~new_new_n1324__ & ~new_new_n3863__;
  assign new_new_n3866__ = ~new_new_n2611__ & ~new_new_n3864__;
  assign new_new_n3867__ = ~new_new_n3865__ & new_new_n3866__;
  assign new_new_n3868__ = ~new_new_n3861__ & ~new_new_n3867__;
  assign new_new_n3869__ = new_new_n2618__ & new_new_n3735__;
  assign new_new_n3870__ = pi01 & new_new_n2608__;
  assign new_new_n3871__ = ~pi00 & ~new_new_n3869__;
  assign new_new_n3872__ = ~new_new_n3870__ & new_new_n3871__;
  assign new_new_n3873__ = new_new_n2604__ & new_new_n3770__;
  assign new_new_n3874__ = ~new_new_n2829__ & ~new_new_n3770__;
  assign new_new_n3875__ = pi00 & ~new_new_n3873__;
  assign new_new_n3876__ = ~new_new_n3874__ & new_new_n3875__;
  assign new_new_n3877__ = ~new_new_n3872__ & ~new_new_n3876__;
  assign new_new_n3878__ = ~new_new_n3233__ & ~new_new_n3877__;
  assign new_new_n3879__ = new_new_n2615__ & new_new_n2819__;
  assign new_new_n3880__ = new_new_n3878__ & new_new_n3879__;
  assign new_new_n3881__ = new_new_n1573__ & new_new_n3877__;
  assign new_new_n3882__ = ~new_new_n3878__ & ~new_new_n3881__;
  assign new_new_n3883__ = ~new_new_n2611__ & ~new_new_n3235__;
  assign new_new_n3884__ = ~new_new_n3882__ & new_new_n3883__;
  assign new_new_n3885__ = ~new_new_n3880__ & ~new_new_n3884__;
  assign new_new_n3886__ = new_new_n3868__ & new_new_n3885__;
  assign new_new_n3887__ = ~new_new_n3868__ & ~new_new_n3885__;
  assign new_new_n3888__ = new_new_n2600__ & ~new_new_n3730__;
  assign new_new_n3889__ = pi01 & ~new_new_n2604__;
  assign new_new_n3890__ = ~new_new_n2608__ & new_new_n3735__;
  assign new_new_n3891__ = ~pi00 & ~new_new_n3890__;
  assign new_new_n3892__ = ~new_new_n3889__ & new_new_n3891__;
  assign new_new_n3893__ = ~new_new_n3888__ & ~new_new_n3892__;
  assign new_new_n3894__ = ~new_new_n3778__ & ~new_new_n3893__;
  assign new_new_n3895__ = pi00 & new_new_n3231__;
  assign new_new_n3896__ = ~new_new_n3765__ & ~new_new_n3895__;
  assign new_new_n3897__ = ~new_new_n2634__ & ~new_new_n3896__;
  assign new_new_n3898__ = pi00 & ~new_new_n3761__;
  assign new_new_n3899__ = new_new_n2634__ & new_new_n3898__;
  assign new_new_n3900__ = pi01 & new_new_n3765__;
  assign new_new_n3901__ = ~new_new_n3772__ & ~new_new_n3900__;
  assign new_new_n3902__ = new_new_n3893__ & new_new_n3901__;
  assign new_new_n3903__ = ~new_new_n3897__ & new_new_n3902__;
  assign new_new_n3904__ = ~new_new_n3899__ & new_new_n3903__;
  assign new_new_n3905__ = ~new_new_n3894__ & ~new_new_n3904__;
  assign new_new_n3906__ = ~new_new_n3887__ & ~new_new_n3905__;
  assign new_new_n3907__ = ~new_new_n3886__ & ~new_new_n3906__;
  assign new_new_n3908__ = ~new_new_n3838__ & ~new_new_n3859__;
  assign new_new_n3909__ = new_new_n2590__ & new_new_n3839__;
  assign new_new_n3910__ = new_new_n2604__ & new_new_n3735__;
  assign new_new_n3911__ = pi01 & new_new_n2600__;
  assign new_new_n3912__ = ~new_new_n3910__ & ~new_new_n3911__;
  assign new_new_n3913__ = ~pi00 & ~new_new_n3912__;
  assign new_new_n3914__ = ~new_new_n3909__ & ~new_new_n3913__;
  assign new_new_n3915__ = ~pi01 & ~new_new_n2655__;
  assign new_new_n3916__ = new_new_n3765__ & ~new_new_n3915__;
  assign new_new_n3917__ = ~new_new_n2655__ & new_new_n3761__;
  assign new_new_n3918__ = new_new_n2655__ & ~new_new_n3231__;
  assign new_new_n3919__ = pi00 & ~new_new_n3917__;
  assign new_new_n3920__ = ~new_new_n3918__ & new_new_n3919__;
  assign new_new_n3921__ = ~new_new_n3772__ & ~new_new_n3916__;
  assign new_new_n3922__ = ~new_new_n3920__ & new_new_n3921__;
  assign new_new_n3923__ = new_new_n3914__ & ~new_new_n3922__;
  assign new_new_n3924__ = pi00 & ~new_new_n2655__;
  assign new_new_n3925__ = new_new_n3735__ & ~new_new_n3924__;
  assign new_new_n3926__ = new_new_n3776__ & ~new_new_n3914__;
  assign new_new_n3927__ = ~new_new_n3925__ & new_new_n3926__;
  assign new_new_n3928__ = ~new_new_n3923__ & ~new_new_n3927__;
  assign new_new_n3929__ = ~new_new_n3907__ & new_new_n3928__;
  assign new_new_n3930__ = ~new_new_n3908__ & new_new_n3929__;
  assign new_new_n3931__ = new_new_n3907__ & ~new_new_n3928__;
  assign new_new_n3932__ = new_new_n3237__ & new_new_n3244__;
  assign new_new_n3933__ = new_new_n3350__ & ~new_new_n3932__;
  assign new_new_n3934__ = new_new_n1324__ & ~new_new_n2611__;
  assign new_new_n3935__ = new_new_n3235__ & ~new_new_n3934__;
  assign new_new_n3936__ = new_new_n2611__ & ~new_new_n3862__;
  assign new_new_n3937__ = new_new_n3243__ & ~new_new_n3935__;
  assign new_new_n3938__ = ~new_new_n3936__ & new_new_n3937__;
  assign new_new_n3939__ = ~new_new_n3933__ & new_new_n3938__;
  assign new_new_n3940__ = new_new_n3933__ & ~new_new_n3938__;
  assign new_new_n3941__ = ~new_new_n3939__ & ~new_new_n3940__;
  assign new_new_n3942__ = ~new_new_n3931__ & new_new_n3941__;
  assign new_new_n3943__ = ~new_new_n3908__ & new_new_n3942__;
  assign new_new_n3944__ = ~new_new_n3860__ & ~new_new_n3930__;
  assign new_new_n3945__ = ~new_new_n3943__ & new_new_n3944__;
  assign new_new_n3946__ = ~new_new_n3827__ & new_new_n3945__;
  assign new_new_n3947__ = new_new_n3827__ & ~new_new_n3945__;
  assign new_new_n3948__ = ~new_new_n3357__ & ~new_new_n3358__;
  assign new_new_n3949__ = ~new_new_n2968__ & new_new_n3948__;
  assign new_new_n3950__ = new_new_n2968__ & ~new_new_n3948__;
  assign new_new_n3951__ = ~new_new_n3949__ & ~new_new_n3950__;
  assign new_new_n3952__ = ~new_new_n3947__ & new_new_n3951__;
  assign new_new_n3953__ = ~new_new_n3946__ & ~new_new_n3952__;
  assign new_new_n3954__ = new_new_n3111__ & ~new_new_n3770__;
  assign new_new_n3955__ = ~new_new_n3203__ & ~new_new_n3954__;
  assign new_new_n3956__ = new_new_n3203__ & new_new_n3954__;
  assign new_new_n3957__ = pi00 & ~new_new_n3955__;
  assign new_new_n3958__ = ~new_new_n3956__ & new_new_n3957__;
  assign new_new_n3959__ = new_new_n2585__ & new_new_n3735__;
  assign new_new_n3960__ = pi01 & ~new_new_n2784__;
  assign new_new_n3961__ = ~pi00 & ~new_new_n3959__;
  assign new_new_n3962__ = ~new_new_n3960__ & new_new_n3961__;
  assign new_new_n3963__ = ~new_new_n3958__ & ~new_new_n3962__;
  assign new_new_n3964__ = ~new_new_n3810__ & ~new_new_n3963__;
  assign new_new_n3965__ = new_new_n3233__ & new_new_n3963__;
  assign new_new_n3966__ = ~new_new_n3964__ & ~new_new_n3965__;
  assign new_new_n3967__ = new_new_n3953__ & new_new_n3966__;
  assign new_new_n3968__ = ~new_new_n3811__ & ~new_new_n3967__;
  assign new_new_n3969__ = new_new_n3806__ & ~new_new_n3968__;
  assign new_new_n3970__ = new_new_n3233__ & new_new_n3810__;
  assign new_new_n3971__ = ~new_new_n3810__ & new_new_n3963__;
  assign new_new_n3972__ = ~new_new_n3233__ & ~new_new_n3963__;
  assign new_new_n3973__ = ~new_new_n3971__ & ~new_new_n3972__;
  assign new_new_n3974__ = new_new_n3953__ & new_new_n3973__;
  assign new_new_n3975__ = ~new_new_n3970__ & ~new_new_n3974__;
  assign new_new_n3976__ = ~new_new_n3806__ & ~new_new_n3975__;
  assign new_new_n3977__ = ~new_new_n3806__ & new_new_n3973__;
  assign new_new_n3978__ = ~new_new_n3233__ & new_new_n3953__;
  assign new_new_n3979__ = ~new_new_n3966__ & ~new_new_n3978__;
  assign new_new_n3980__ = new_new_n3806__ & ~new_new_n3979__;
  assign new_new_n3981__ = new_new_n3233__ & ~new_new_n3806__;
  assign new_new_n3982__ = ~new_new_n3810__ & ~new_new_n3981__;
  assign new_new_n3983__ = new_new_n3953__ & ~new_new_n3982__;
  assign new_new_n3984__ = ~new_new_n3977__ & ~new_new_n3983__;
  assign new_new_n3985__ = ~new_new_n3980__ & new_new_n3984__;
  assign new_new_n3986__ = ~new_new_n3304__ & ~new_new_n3305__;
  assign new_new_n3987__ = ~new_new_n3360__ & new_new_n3986__;
  assign new_new_n3988__ = new_new_n3360__ & ~new_new_n3986__;
  assign new_new_n3989__ = ~new_new_n3987__ & ~new_new_n3988__;
  assign new_new_n3990__ = ~new_new_n3985__ & new_new_n3989__;
  assign new_new_n3991__ = ~new_new_n3969__ & ~new_new_n3976__;
  assign new_new_n3992__ = ~new_new_n3990__ & new_new_n3991__;
  assign new_new_n3993__ = new_new_n3515__ & ~new_new_n3770__;
  assign new_new_n3994__ = new_new_n3233__ & ~new_new_n3993__;
  assign new_new_n3995__ = ~new_new_n3233__ & new_new_n3993__;
  assign new_new_n3996__ = ~new_new_n3994__ & ~new_new_n3995__;
  assign new_new_n3997__ = new_new_n3586__ & new_new_n3996__;
  assign new_new_n3998__ = ~new_new_n3586__ & ~new_new_n3996__;
  assign new_new_n3999__ = pi00 & ~new_new_n3997__;
  assign new_new_n4000__ = ~new_new_n3998__ & new_new_n3999__;
  assign new_new_n4001__ = pi01 & ~new_new_n3486__;
  assign new_new_n4002__ = ~new_new_n3203__ & new_new_n3735__;
  assign new_new_n4003__ = ~new_new_n4001__ & ~new_new_n4002__;
  assign new_new_n4004__ = ~new_new_n3233__ & new_new_n4003__;
  assign new_new_n4005__ = new_new_n3233__ & ~new_new_n4003__;
  assign new_new_n4006__ = ~pi00 & ~new_new_n4004__;
  assign new_new_n4007__ = ~new_new_n4005__ & new_new_n4006__;
  assign new_new_n4008__ = ~new_new_n4000__ & ~new_new_n4007__;
  assign new_new_n4009__ = ~new_new_n3992__ & ~new_new_n4008__;
  assign new_new_n4010__ = new_new_n3992__ & new_new_n4008__;
  assign new_new_n4011__ = ~new_new_n3365__ & ~new_new_n3366__;
  assign new_new_n4012__ = ~new_new_n3370__ & ~new_new_n4011__;
  assign new_new_n4013__ = new_new_n3370__ & new_new_n4011__;
  assign new_new_n4014__ = ~new_new_n4012__ & ~new_new_n4013__;
  assign new_new_n4015__ = ~new_new_n4010__ & new_new_n4014__;
  assign new_new_n4016__ = ~new_new_n4009__ & ~new_new_n4015__;
  assign new_new_n4017__ = ~new_new_n3796__ & new_new_n4016__;
  assign new_new_n4018__ = new_new_n3796__ & ~new_new_n4016__;
  assign new_new_n4019__ = ~new_new_n3389__ & ~new_new_n3390__;
  assign new_new_n4020__ = new_new_n3394__ & ~new_new_n4019__;
  assign new_new_n4021__ = ~new_new_n3394__ & new_new_n4019__;
  assign new_new_n4022__ = ~new_new_n4020__ & ~new_new_n4021__;
  assign new_new_n4023__ = ~new_new_n4018__ & new_new_n4022__;
  assign new_new_n4024__ = ~new_new_n3740__ & ~new_new_n3745__;
  assign new_new_n4025__ = pi02 & ~new_new_n4024__;
  assign new_new_n4026__ = pi01 & new_new_n4024__;
  assign new_new_n4027__ = ~new_new_n4025__ & ~new_new_n4026__;
  assign new_new_n4028__ = new_new_n3229__ & ~new_new_n3733__;
  assign new_new_n4029__ = ~new_new_n3229__ & new_new_n3733__;
  assign new_new_n4030__ = ~new_new_n4028__ & ~new_new_n4029__;
  assign new_new_n4031__ = new_new_n4027__ & new_new_n4030__;
  assign new_new_n4032__ = ~new_new_n4027__ & ~new_new_n4030__;
  assign new_new_n4033__ = pi00 & ~new_new_n4031__;
  assign new_new_n4034__ = ~new_new_n4032__ & new_new_n4033__;
  assign new_new_n4035__ = new_new_n3586__ & new_new_n3735__;
  assign new_new_n4036__ = ~new_new_n3651__ & new_new_n3776__;
  assign new_new_n4037__ = new_new_n3651__ & ~new_new_n3776__;
  assign new_new_n4038__ = pi01 & ~new_new_n4036__;
  assign new_new_n4039__ = ~new_new_n4037__ & new_new_n4038__;
  assign new_new_n4040__ = ~pi00 & ~new_new_n4035__;
  assign new_new_n4041__ = ~new_new_n4039__ & new_new_n4040__;
  assign new_new_n4042__ = ~new_new_n4034__ & ~new_new_n4041__;
  assign new_new_n4043__ = ~new_new_n3397__ & ~new_new_n3505__;
  assign new_new_n4044__ = ~new_new_n3504__ & new_new_n4043__;
  assign new_new_n4045__ = new_new_n3504__ & ~new_new_n4043__;
  assign new_new_n4046__ = ~new_new_n4044__ & ~new_new_n4045__;
  assign new_new_n4047__ = new_new_n4042__ & ~new_new_n4046__;
  assign new_new_n4048__ = ~new_new_n4017__ & ~new_new_n4047__;
  assign new_new_n4049__ = ~new_new_n4023__ & new_new_n4048__;
  assign new_new_n4050__ = ~new_new_n4042__ & new_new_n4046__;
  assign new_new_n4051__ = ~new_new_n4049__ & ~new_new_n4050__;
  assign new_new_n4052__ = new_new_n3780__ & ~new_new_n4051__;
  assign new_new_n4053__ = ~new_new_n3780__ & new_new_n4051__;
  assign new_new_n4054__ = ~new_new_n3508__ & ~new_new_n3509__;
  assign new_new_n4055__ = new_new_n3601__ & new_new_n4054__;
  assign new_new_n4056__ = ~new_new_n3601__ & ~new_new_n4054__;
  assign new_new_n4057__ = ~new_new_n4055__ & ~new_new_n4056__;
  assign new_new_n4058__ = ~new_new_n4053__ & new_new_n4057__;
  assign new_new_n4059__ = ~new_new_n4052__ & ~new_new_n4058__;
  assign new_new_n4060__ = new_new_n3670__ & new_new_n4059__;
  assign new_new_n4061__ = new_new_n148__ & ~new_new_n570__;
  assign new_new_n4062__ = ~new_new_n200__ & new_new_n4061__;
  assign new_new_n4063__ = ~new_new_n691__ & new_new_n4062__;
  assign new_new_n4064__ = ~new_new_n124__ & ~new_new_n4063__;
  assign new_new_n4065__ = new_new_n256__ & ~new_new_n472__;
  assign new_new_n4066__ = ~new_new_n2454__ & new_new_n4065__;
  assign new_new_n4067__ = ~new_new_n54__ & ~new_new_n4066__;
  assign new_new_n4068__ = new_new_n195__ & ~new_new_n1095__;
  assign new_new_n4069__ = new_new_n160__ & ~new_new_n248__;
  assign new_new_n4070__ = ~new_new_n893__ & ~new_new_n4068__;
  assign new_new_n4071__ = new_new_n1443__ & new_new_n4070__;
  assign new_new_n4072__ = new_new_n2448__ & new_new_n4069__;
  assign new_new_n4073__ = new_new_n4071__ & new_new_n4072__;
  assign new_new_n4074__ = ~new_new_n4064__ & ~new_new_n4067__;
  assign new_new_n4075__ = new_new_n4073__ & new_new_n4074__;
  assign new_new_n4076__ = new_new_n684__ & new_new_n3181__;
  assign new_new_n4077__ = new_new_n4075__ & new_new_n4076__;
  assign new_new_n4078__ = new_new_n638__ & new_new_n4077__;
  assign new_new_n4079__ = ~new_new_n3726__ & new_new_n4078__;
  assign new_new_n4080__ = new_new_n3726__ & ~new_new_n4078__;
  assign new_new_n4081__ = ~new_new_n4079__ & ~new_new_n4080__;
  assign new_new_n4082__ = new_new_n3733__ & new_new_n3740__;
  assign new_new_n4083__ = ~new_new_n3745__ & ~new_new_n3747__;
  assign new_new_n4084__ = ~new_new_n3733__ & ~new_new_n4083__;
  assign new_new_n4085__ = ~new_new_n3753__ & ~new_new_n4082__;
  assign new_new_n4086__ = ~new_new_n4084__ & new_new_n4085__;
  assign new_new_n4087__ = ~new_new_n3770__ & new_new_n4086__;
  assign new_new_n4088__ = ~new_new_n4081__ & new_new_n4087__;
  assign new_new_n4089__ = new_new_n4081__ & ~new_new_n4087__;
  assign new_new_n4090__ = ~new_new_n4088__ & ~new_new_n4089__;
  assign new_new_n4091__ = pi00 & ~new_new_n4090__;
  assign new_new_n4092__ = pi01 & ~new_new_n3727__;
  assign new_new_n4093__ = ~new_new_n3733__ & new_new_n3735__;
  assign new_new_n4094__ = ~new_new_n4092__ & ~new_new_n4093__;
  assign new_new_n4095__ = ~pi00 & ~new_new_n4094__;
  assign new_new_n4096__ = ~new_new_n4091__ & ~new_new_n4095__;
  assign new_new_n4097__ = new_new_n3233__ & ~new_new_n4096__;
  assign new_new_n4098__ = ~new_new_n3233__ & new_new_n4096__;
  assign new_new_n4099__ = ~new_new_n4097__ & ~new_new_n4098__;
  assign new_new_n4100__ = new_new_n4060__ & ~new_new_n4099__;
  assign new_new_n4101__ = new_new_n2593__ & ~new_new_n2784__;
  assign new_new_n4102__ = ~new_new_n320__ & ~new_new_n3203__;
  assign new_new_n4103__ = ~new_new_n4101__ & ~new_new_n4102__;
  assign new_new_n4104__ = new_new_n2596__ & new_new_n3490__;
  assign new_new_n4105__ = new_new_n4103__ & ~new_new_n4104__;
  assign new_new_n4106__ = ~new_new_n301__ & ~new_new_n4105__;
  assign new_new_n4107__ = ~new_new_n316__ & ~new_new_n3486__;
  assign new_new_n4108__ = new_new_n316__ & new_new_n3486__;
  assign new_new_n4109__ = new_new_n2596__ & ~new_new_n4107__;
  assign new_new_n4110__ = ~new_new_n4108__ & new_new_n4109__;
  assign new_new_n4111__ = new_new_n3489__ & new_new_n4110__;
  assign new_new_n4112__ = new_new_n2596__ & ~new_new_n3499__;
  assign new_new_n4113__ = new_new_n301__ & new_new_n4103__;
  assign new_new_n4114__ = ~new_new_n4112__ & new_new_n4113__;
  assign new_new_n4115__ = ~new_new_n4111__ & ~new_new_n4114__;
  assign new_new_n4116__ = ~new_new_n4106__ & new_new_n4115__;
  assign new_new_n4117__ = new_new_n2600__ & ~new_new_n2806__;
  assign new_new_n4118__ = new_new_n2590__ & new_new_n2809__;
  assign new_new_n4119__ = ~new_new_n4117__ & ~new_new_n4118__;
  assign new_new_n4120__ = new_new_n2808__ & new_new_n3031__;
  assign new_new_n4121__ = new_new_n4119__ & ~new_new_n4120__;
  assign new_new_n4122__ = new_new_n810__ & ~new_new_n4121__;
  assign new_new_n4123__ = ~new_new_n816__ & ~new_new_n3035__;
  assign new_new_n4124__ = new_new_n816__ & ~new_new_n3037__;
  assign new_new_n4125__ = new_new_n2808__ & ~new_new_n4123__;
  assign new_new_n4126__ = ~new_new_n4124__ & new_new_n4125__;
  assign new_new_n4127__ = new_new_n2808__ & ~new_new_n3041__;
  assign new_new_n4128__ = ~new_new_n810__ & new_new_n4119__;
  assign new_new_n4129__ = ~new_new_n4127__ & new_new_n4128__;
  assign new_new_n4130__ = ~new_new_n4122__ & ~new_new_n4129__;
  assign new_new_n4131__ = ~new_new_n4126__ & new_new_n4130__;
  assign new_new_n4132__ = ~new_new_n3069__ & ~new_new_n3072__;
  assign new_new_n4133__ = new_new_n2618__ & new_new_n4132__;
  assign new_new_n4134__ = new_new_n2608__ & new_new_n3069__;
  assign new_new_n4135__ = ~new_new_n2848__ & ~new_new_n4133__;
  assign new_new_n4136__ = ~new_new_n4134__ & new_new_n4135__;
  assign new_new_n4137__ = new_new_n2604__ & new_new_n3072__;
  assign new_new_n4138__ = ~new_new_n2829__ & ~new_new_n3072__;
  assign new_new_n4139__ = new_new_n2848__ & ~new_new_n4137__;
  assign new_new_n4140__ = ~new_new_n4138__ & new_new_n4139__;
  assign new_new_n4141__ = ~new_new_n4136__ & ~new_new_n4140__;
  assign new_new_n4142__ = ~new_new_n3061__ & new_new_n3079__;
  assign new_new_n4143__ = ~new_new_n2611__ & new_new_n4142__;
  assign new_new_n4144__ = ~new_new_n437__ & new_new_n2611__;
  assign new_new_n4145__ = ~new_new_n4142__ & new_new_n4144__;
  assign new_new_n4146__ = ~new_new_n4143__ & ~new_new_n4145__;
  assign new_new_n4147__ = ~new_new_n4141__ & new_new_n4146__;
  assign new_new_n4148__ = new_new_n4141__ & new_new_n4145__;
  assign new_new_n4149__ = ~new_new_n4147__ & ~new_new_n4148__;
  assign new_new_n4150__ = new_new_n4131__ & new_new_n4149__;
  assign new_new_n4151__ = ~new_new_n4131__ & ~new_new_n4149__;
  assign new_new_n4152__ = ~new_new_n4150__ & ~new_new_n4151__;
  assign new_new_n4153__ = ~new_new_n3082__ & ~new_new_n3102__;
  assign new_new_n4154__ = ~new_new_n3101__ & ~new_new_n4153__;
  assign new_new_n4155__ = new_new_n4152__ & ~new_new_n4154__;
  assign new_new_n4156__ = ~new_new_n4152__ & new_new_n4154__;
  assign new_new_n4157__ = ~new_new_n4155__ & ~new_new_n4156__;
  assign new_new_n4158__ = ~new_new_n4116__ & new_new_n4157__;
  assign new_new_n4159__ = new_new_n4116__ & ~new_new_n4157__;
  assign new_new_n4160__ = ~new_new_n4158__ & ~new_new_n4159__;
  assign new_new_n4161__ = new_new_n3220__ & new_new_n4160__;
  assign new_new_n4162__ = ~new_new_n3220__ & ~new_new_n4160__;
  assign new_new_n4163__ = ~new_new_n4161__ & ~new_new_n4162__;
  assign new_new_n4164__ = new_new_n3240__ & new_new_n3651__;
  assign new_new_n4165__ = new_new_n3247__ & ~new_new_n3586__;
  assign new_new_n4166__ = ~new_new_n4164__ & ~new_new_n4165__;
  assign new_new_n4167__ = ~new_new_n3733__ & ~new_new_n4024__;
  assign new_new_n4168__ = new_new_n3236__ & new_new_n4167__;
  assign new_new_n4169__ = new_new_n4166__ & ~new_new_n4168__;
  assign new_new_n4170__ = new_new_n310__ & ~new_new_n4169__;
  assign new_new_n4171__ = ~new_new_n1324__ & new_new_n3733__;
  assign new_new_n4172__ = new_new_n1324__ & ~new_new_n3733__;
  assign new_new_n4173__ = new_new_n3236__ & new_new_n4024__;
  assign new_new_n4174__ = ~new_new_n4171__ & ~new_new_n4172__;
  assign new_new_n4175__ = new_new_n4173__ & new_new_n4174__;
  assign new_new_n4176__ = new_new_n3733__ & ~new_new_n4024__;
  assign new_new_n4177__ = new_new_n3236__ & ~new_new_n4176__;
  assign new_new_n4178__ = ~new_new_n310__ & new_new_n4166__;
  assign new_new_n4179__ = ~new_new_n4177__ & new_new_n4178__;
  assign new_new_n4180__ = ~new_new_n4175__ & ~new_new_n4179__;
  assign new_new_n4181__ = ~new_new_n4170__ & new_new_n4180__;
  assign new_new_n4182__ = ~new_new_n3224__ & ~new_new_n3665__;
  assign new_new_n4183__ = ~new_new_n3666__ & ~new_new_n4182__;
  assign new_new_n4184__ = ~new_new_n4181__ & ~new_new_n4183__;
  assign new_new_n4185__ = new_new_n4181__ & new_new_n4183__;
  assign new_new_n4186__ = ~new_new_n4184__ & ~new_new_n4185__;
  assign new_new_n4187__ = ~pi22 & ~new_new_n4078__;
  assign new_new_n4188__ = pi22 & new_new_n4078__;
  assign new_new_n4189__ = ~new_new_n4187__ & ~new_new_n4188__;
  assign new_new_n4190__ = new_new_n3726__ & ~new_new_n4189__;
  assign new_new_n4191__ = ~new_new_n3726__ & new_new_n4189__;
  assign new_new_n4192__ = ~new_new_n4190__ & ~new_new_n4191__;
  assign new_new_n4193__ = new_new_n3769__ & ~new_new_n4192__;
  assign new_new_n4194__ = ~pi01 & ~new_new_n3727__;
  assign new_new_n4195__ = pi01 & new_new_n4191__;
  assign new_new_n4196__ = pi02 & ~new_new_n4190__;
  assign new_new_n4197__ = ~new_new_n4194__ & new_new_n4196__;
  assign new_new_n4198__ = ~new_new_n4195__ & new_new_n4197__;
  assign new_new_n4199__ = ~new_new_n4193__ & ~new_new_n4198__;
  assign new_new_n4200__ = ~pi00 & ~new_new_n4199__;
  assign new_new_n4201__ = new_new_n3726__ & new_new_n4078__;
  assign new_new_n4202__ = new_new_n162__ & ~new_new_n663__;
  assign new_new_n4203__ = ~new_new_n100__ & ~new_new_n4202__;
  assign new_new_n4204__ = new_new_n180__ & new_new_n629__;
  assign new_new_n4205__ = ~new_new_n339__ & new_new_n4204__;
  assign new_new_n4206__ = ~new_new_n4203__ & ~new_new_n4205__;
  assign new_new_n4207__ = new_new_n244__ & ~new_new_n2248__;
  assign new_new_n4208__ = new_new_n174__ & new_new_n677__;
  assign new_new_n4209__ = new_new_n125__ & ~new_new_n4208__;
  assign new_new_n4210__ = ~new_new_n175__ & ~new_new_n662__;
  assign new_new_n4211__ = ~new_new_n4207__ & new_new_n4210__;
  assign new_new_n4212__ = ~new_new_n667__ & new_new_n864__;
  assign new_new_n4213__ = ~new_new_n4209__ & new_new_n4212__;
  assign new_new_n4214__ = ~new_new_n622__ & new_new_n4211__;
  assign new_new_n4215__ = ~new_new_n795__ & ~new_new_n4206__;
  assign new_new_n4216__ = new_new_n4214__ & new_new_n4215__;
  assign new_new_n4217__ = new_new_n636__ & new_new_n4213__;
  assign new_new_n4218__ = new_new_n684__ & new_new_n4217__;
  assign new_new_n4219__ = new_new_n4216__ & new_new_n4218__;
  assign new_new_n4220__ = ~new_new_n4201__ & new_new_n4219__;
  assign new_new_n4221__ = new_new_n4201__ & ~new_new_n4219__;
  assign new_new_n4222__ = ~new_new_n4220__ & ~new_new_n4221__;
  assign new_new_n4223__ = new_new_n3776__ & new_new_n4222__;
  assign new_new_n4224__ = ~new_new_n3740__ & new_new_n4078__;
  assign new_new_n4225__ = ~new_new_n3724__ & ~new_new_n4224__;
  assign new_new_n4226__ = new_new_n3733__ & ~new_new_n4225__;
  assign new_new_n4227__ = ~new_new_n3745__ & ~new_new_n4078__;
  assign new_new_n4228__ = ~new_new_n3725__ & ~new_new_n3746__;
  assign new_new_n4229__ = ~new_new_n4227__ & new_new_n4228__;
  assign new_new_n4230__ = ~new_new_n4226__ & ~new_new_n4229__;
  assign new_new_n4231__ = ~new_new_n4081__ & ~new_new_n4230__;
  assign new_new_n4232__ = new_new_n4081__ & new_new_n4230__;
  assign new_new_n4233__ = ~new_new_n4231__ & ~new_new_n4232__;
  assign new_new_n4234__ = ~new_new_n3776__ & ~new_new_n4222__;
  assign new_new_n4235__ = ~new_new_n4223__ & ~new_new_n4234__;
  assign new_new_n4236__ = ~new_new_n4233__ & new_new_n4235__;
  assign new_new_n4237__ = new_new_n3761__ & new_new_n4222__;
  assign new_new_n4238__ = ~new_new_n3761__ & ~new_new_n4222__;
  assign new_new_n4239__ = ~new_new_n4237__ & ~new_new_n4238__;
  assign new_new_n4240__ = new_new_n4233__ & new_new_n4239__;
  assign new_new_n4241__ = pi00 & ~new_new_n4236__;
  assign new_new_n4242__ = ~new_new_n4240__ & new_new_n4241__;
  assign new_new_n4243__ = ~new_new_n4200__ & ~new_new_n4242__;
  assign new_new_n4244__ = new_new_n4186__ & ~new_new_n4243__;
  assign new_new_n4245__ = ~new_new_n4186__ & new_new_n4243__;
  assign new_new_n4246__ = ~new_new_n4244__ & ~new_new_n4245__;
  assign new_new_n4247__ = new_new_n4163__ & new_new_n4246__;
  assign new_new_n4248__ = ~new_new_n4163__ & ~new_new_n4246__;
  assign new_new_n4249__ = ~new_new_n4247__ & ~new_new_n4248__;
  assign new_new_n4250__ = new_new_n4100__ & ~new_new_n4249__;
  assign new_new_n4251__ = ~new_new_n3670__ & ~new_new_n4059__;
  assign new_new_n4252__ = ~new_new_n4099__ & ~new_new_n4251__;
  assign new_new_n4253__ = ~new_new_n4060__ & ~new_new_n4252__;
  assign new_new_n4254__ = new_new_n4249__ & new_new_n4253__;
  assign new_new_n4255__ = new_new_n4099__ & new_new_n4251__;
  assign new_new_n4256__ = new_new_n4254__ & ~new_new_n4255__;
  assign new_new_n4257__ = ~new_new_n4100__ & new_new_n4249__;
  assign new_new_n4258__ = ~new_new_n162__ & new_new_n493__;
  assign new_new_n4259__ = new_new_n223__ & ~new_new_n1095__;
  assign new_new_n4260__ = ~new_new_n141__ & new_new_n422__;
  assign new_new_n4261__ = new_new_n218__ & ~new_new_n4259__;
  assign new_new_n4262__ = ~new_new_n4260__ & new_new_n4261__;
  assign new_new_n4263__ = ~new_new_n4258__ & ~new_new_n4262__;
  assign new_new_n4264__ = new_new_n162__ & ~new_new_n797__;
  assign new_new_n4265__ = new_new_n256__ & new_new_n2532__;
  assign new_new_n4266__ = new_new_n116__ & ~new_new_n4265__;
  assign new_new_n4267__ = ~new_new_n4264__ & ~new_new_n4266__;
  assign new_new_n4268__ = new_new_n136__ & new_new_n166__;
  assign new_new_n4269__ = new_new_n125__ & ~new_new_n4268__;
  assign new_new_n4270__ = new_new_n470__ & ~new_new_n4269__;
  assign new_new_n4271__ = ~new_new_n4263__ & new_new_n4270__;
  assign new_new_n4272__ = new_new_n4267__ & new_new_n4271__;
  assign new_new_n4273__ = ~new_new_n274__ & ~new_new_n925__;
  assign new_new_n4274__ = new_new_n195__ & ~new_new_n238__;
  assign new_new_n4275__ = ~new_new_n141__ & ~new_new_n2538__;
  assign new_new_n4276__ = ~new_new_n2329__ & new_new_n4275__;
  assign new_new_n4277__ = new_new_n116__ & ~new_new_n2451__;
  assign new_new_n4278__ = ~new_new_n223__ & ~new_new_n4277__;
  assign new_new_n4279__ = ~new_new_n116__ & new_new_n213__;
  assign new_new_n4280__ = new_new_n270__ & new_new_n4279__;
  assign new_new_n4281__ = ~new_new_n4278__ & ~new_new_n4280__;
  assign new_new_n4282__ = ~new_new_n229__ & ~new_new_n921__;
  assign new_new_n4283__ = ~new_new_n240__ & new_new_n4282__;
  assign new_new_n4284__ = ~new_new_n4276__ & new_new_n4283__;
  assign new_new_n4285__ = ~new_new_n4281__ & new_new_n4284__;
  assign new_new_n4286__ = new_new_n2247__ & new_new_n4285__;
  assign new_new_n4287__ = new_new_n1123__ & new_new_n4286__;
  assign new_new_n4288__ = ~new_new_n457__ & ~new_new_n4274__;
  assign new_new_n4289__ = new_new_n476__ & new_new_n4288__;
  assign new_new_n4290__ = new_new_n4287__ & new_new_n4289__;
  assign new_new_n4291__ = ~new_new_n181__ & ~new_new_n195__;
  assign new_new_n4292__ = new_new_n180__ & new_new_n4291__;
  assign new_new_n4293__ = ~new_new_n452__ & ~new_new_n4292__;
  assign new_new_n4294__ = ~new_new_n971__ & ~new_new_n4293__;
  assign new_new_n4295__ = ~new_new_n89__ & ~new_new_n404__;
  assign new_new_n4296__ = ~new_new_n690__ & new_new_n4295__;
  assign new_new_n4297__ = ~new_new_n257__ & new_new_n4273__;
  assign new_new_n4298__ = new_new_n4296__ & new_new_n4297__;
  assign new_new_n4299__ = new_new_n2339__ & new_new_n4298__;
  assign new_new_n4300__ = new_new_n4294__ & new_new_n4299__;
  assign new_new_n4301__ = new_new_n4272__ & new_new_n4300__;
  assign new_new_n4302__ = new_new_n4290__ & new_new_n4301__;
  assign new_new_n4303__ = ~new_new_n4255__ & ~new_new_n4302__;
  assign new_new_n4304__ = ~new_new_n4257__ & new_new_n4303__;
  assign new_new_n4305__ = ~new_new_n4250__ & ~new_new_n4304__;
  assign new_new_n4306__ = ~new_new_n4256__ & new_new_n4305__;
  assign new_new_n4307__ = ~new_new_n297__ & ~new_new_n4306__;
  assign new_new_n4308__ = ~new_new_n4249__ & ~new_new_n4253__;
  assign new_new_n4309__ = ~new_new_n4254__ & ~new_new_n4308__;
  assign new_new_n4310__ = ~new_new_n4302__ & ~new_new_n4309__;
  assign new_new_n4311__ = ~new_new_n4307__ & ~new_new_n4310__;
  assign new_new_n4312__ = new_new_n3247__ & new_new_n3651__;
  assign new_new_n4313__ = new_new_n3240__ & ~new_new_n3733__;
  assign new_new_n4314__ = ~new_new_n4312__ & ~new_new_n4313__;
  assign new_new_n4315__ = ~new_new_n3727__ & ~new_new_n3757__;
  assign new_new_n4316__ = new_new_n3236__ & new_new_n4315__;
  assign new_new_n4317__ = new_new_n4314__ & ~new_new_n4316__;
  assign new_new_n4318__ = new_new_n310__ & ~new_new_n4317__;
  assign new_new_n4319__ = ~new_new_n3727__ & new_new_n3757__;
  assign new_new_n4320__ = ~new_new_n1324__ & ~new_new_n4319__;
  assign new_new_n4321__ = new_new_n3727__ & ~new_new_n3757__;
  assign new_new_n4322__ = new_new_n1324__ & ~new_new_n4321__;
  assign new_new_n4323__ = new_new_n3236__ & ~new_new_n4320__;
  assign new_new_n4324__ = ~new_new_n4322__ & new_new_n4323__;
  assign new_new_n4325__ = new_new_n3727__ & new_new_n3757__;
  assign new_new_n4326__ = new_new_n3236__ & ~new_new_n4325__;
  assign new_new_n4327__ = ~new_new_n310__ & new_new_n4314__;
  assign new_new_n4328__ = ~new_new_n4326__ & new_new_n4327__;
  assign new_new_n4329__ = ~new_new_n4318__ & ~new_new_n4328__;
  assign new_new_n4330__ = ~new_new_n4324__ & new_new_n4329__;
  assign new_new_n4331__ = new_new_n2593__ & ~new_new_n3203__;
  assign new_new_n4332__ = ~new_new_n320__ & ~new_new_n3486__;
  assign new_new_n4333__ = ~new_new_n4331__ & ~new_new_n4332__;
  assign new_new_n4334__ = new_new_n2596__ & new_new_n3587__;
  assign new_new_n4335__ = new_new_n4333__ & ~new_new_n4334__;
  assign new_new_n4336__ = ~new_new_n301__ & ~new_new_n4335__;
  assign new_new_n4337__ = new_new_n316__ & new_new_n3586__;
  assign new_new_n4338__ = ~new_new_n316__ & ~new_new_n3586__;
  assign new_new_n4339__ = new_new_n2596__ & new_new_n3515__;
  assign new_new_n4340__ = ~new_new_n4337__ & ~new_new_n4338__;
  assign new_new_n4341__ = new_new_n4339__ & new_new_n4340__;
  assign new_new_n4342__ = new_new_n2596__ & ~new_new_n3596__;
  assign new_new_n4343__ = new_new_n301__ & new_new_n4333__;
  assign new_new_n4344__ = ~new_new_n4342__ & new_new_n4343__;
  assign new_new_n4345__ = ~new_new_n4341__ & ~new_new_n4344__;
  assign new_new_n4346__ = ~new_new_n4336__ & new_new_n4345__;
  assign new_new_n4347__ = new_new_n2585__ & new_new_n2809__;
  assign new_new_n4348__ = new_new_n2590__ & ~new_new_n2806__;
  assign new_new_n4349__ = ~new_new_n4347__ & ~new_new_n4348__;
  assign new_new_n4350__ = new_new_n2785__ & new_new_n2808__;
  assign new_new_n4351__ = new_new_n4349__ & ~new_new_n4350__;
  assign new_new_n4352__ = ~new_new_n810__ & ~new_new_n4351__;
  assign new_new_n4353__ = new_new_n816__ & new_new_n2784__;
  assign new_new_n4354__ = ~new_new_n816__ & ~new_new_n2784__;
  assign new_new_n4355__ = new_new_n2808__ & ~new_new_n4353__;
  assign new_new_n4356__ = ~new_new_n4354__ & new_new_n4355__;
  assign new_new_n4357__ = new_new_n2664__ & new_new_n4356__;
  assign new_new_n4358__ = ~new_new_n2794__ & new_new_n2808__;
  assign new_new_n4359__ = new_new_n810__ & new_new_n4349__;
  assign new_new_n4360__ = ~new_new_n4358__ & new_new_n4359__;
  assign new_new_n4361__ = ~new_new_n4357__ & ~new_new_n4360__;
  assign new_new_n4362__ = ~new_new_n4352__ & new_new_n4361__;
  assign new_new_n4363__ = ~new_new_n4150__ & ~new_new_n4154__;
  assign new_new_n4364__ = ~new_new_n4151__ & ~new_new_n4363__;
  assign new_new_n4365__ = new_new_n4362__ & ~new_new_n4364__;
  assign new_new_n4366__ = ~new_new_n4362__ & new_new_n4364__;
  assign new_new_n4367__ = ~new_new_n4365__ & ~new_new_n4366__;
  assign new_new_n4368__ = new_new_n2608__ & new_new_n4132__;
  assign new_new_n4369__ = new_new_n2604__ & new_new_n3069__;
  assign new_new_n4370__ = ~new_new_n2848__ & ~new_new_n4368__;
  assign new_new_n4371__ = ~new_new_n4369__ & new_new_n4370__;
  assign new_new_n4372__ = new_new_n2600__ & new_new_n3072__;
  assign new_new_n4373__ = new_new_n2634__ & ~new_new_n3072__;
  assign new_new_n4374__ = new_new_n2848__ & ~new_new_n4372__;
  assign new_new_n4375__ = ~new_new_n4373__ & new_new_n4374__;
  assign new_new_n4376__ = ~new_new_n4371__ & ~new_new_n4375__;
  assign new_new_n4377__ = ~new_new_n437__ & ~new_new_n2611__;
  assign new_new_n4378__ = ~new_new_n4142__ & ~new_new_n4377__;
  assign new_new_n4379__ = ~new_new_n4141__ & ~new_new_n4378__;
  assign new_new_n4380__ = new_new_n2618__ & new_new_n4379__;
  assign new_new_n4381__ = ~new_new_n2618__ & ~new_new_n4379__;
  assign new_new_n4382__ = ~new_new_n4380__ & ~new_new_n4381__;
  assign new_new_n4383__ = ~new_new_n437__ & ~new_new_n4382__;
  assign new_new_n4384__ = new_new_n4376__ & new_new_n4383__;
  assign new_new_n4385__ = ~new_new_n4376__ & ~new_new_n4380__;
  assign new_new_n4386__ = ~new_new_n4383__ & new_new_n4385__;
  assign new_new_n4387__ = ~new_new_n4384__ & ~new_new_n4386__;
  assign new_new_n4388__ = ~new_new_n4367__ & ~new_new_n4387__;
  assign new_new_n4389__ = new_new_n4376__ & ~new_new_n4380__;
  assign new_new_n4390__ = ~new_new_n4383__ & ~new_new_n4389__;
  assign new_new_n4391__ = ~new_new_n4384__ & ~new_new_n4390__;
  assign new_new_n4392__ = new_new_n4367__ & new_new_n4391__;
  assign new_new_n4393__ = ~new_new_n4388__ & ~new_new_n4392__;
  assign new_new_n4394__ = ~new_new_n3220__ & ~new_new_n4159__;
  assign new_new_n4395__ = ~new_new_n4158__ & ~new_new_n4394__;
  assign new_new_n4396__ = ~new_new_n4393__ & ~new_new_n4395__;
  assign new_new_n4397__ = new_new_n4393__ & new_new_n4395__;
  assign new_new_n4398__ = ~new_new_n4396__ & ~new_new_n4397__;
  assign new_new_n4399__ = new_new_n4346__ & ~new_new_n4398__;
  assign new_new_n4400__ = ~new_new_n4346__ & new_new_n4398__;
  assign new_new_n4401__ = ~new_new_n4399__ & ~new_new_n4400__;
  assign new_new_n4402__ = ~new_new_n4163__ & ~new_new_n4185__;
  assign new_new_n4403__ = ~new_new_n4184__ & ~new_new_n4402__;
  assign new_new_n4404__ = new_new_n4401__ & ~new_new_n4403__;
  assign new_new_n4405__ = ~new_new_n4401__ & new_new_n4403__;
  assign new_new_n4406__ = ~new_new_n4404__ & ~new_new_n4405__;
  assign new_new_n4407__ = ~new_new_n4330__ & new_new_n4406__;
  assign new_new_n4408__ = new_new_n4330__ & ~new_new_n4406__;
  assign new_new_n4409__ = ~new_new_n4407__ & ~new_new_n4408__;
  assign new_new_n4410__ = new_new_n4243__ & ~new_new_n4249__;
  assign new_new_n4411__ = ~new_new_n4254__ & ~new_new_n4410__;
  assign new_new_n4412__ = new_new_n4201__ & new_new_n4219__;
  assign new_new_n4413__ = ~new_new_n323__ & ~new_new_n412__;
  assign new_new_n4414__ = ~new_new_n220__ & new_new_n4413__;
  assign new_new_n4415__ = new_new_n628__ & new_new_n4414__;
  assign new_new_n4416__ = new_new_n645__ & new_new_n4415__;
  assign new_new_n4417__ = new_new_n684__ & new_new_n4416__;
  assign new_new_n4418__ = new_new_n804__ & new_new_n4417__;
  assign new_new_n4419__ = ~new_new_n4412__ & new_new_n4418__;
  assign new_new_n4420__ = new_new_n4412__ & ~new_new_n4418__;
  assign new_new_n4421__ = ~new_new_n4419__ & ~new_new_n4420__;
  assign new_new_n4422__ = new_new_n3839__ & new_new_n4421__;
  assign new_new_n4423__ = pi01 & new_new_n4222__;
  assign new_new_n4424__ = new_new_n3735__ & new_new_n4081__;
  assign new_new_n4425__ = ~new_new_n4423__ & ~new_new_n4424__;
  assign new_new_n4426__ = ~pi00 & ~new_new_n4425__;
  assign new_new_n4427__ = ~new_new_n4422__ & ~new_new_n4426__;
  assign new_new_n4428__ = ~new_new_n4078__ & new_new_n4418__;
  assign new_new_n4429__ = ~new_new_n4219__ & new_new_n4428__;
  assign new_new_n4430__ = new_new_n4081__ & new_new_n4418__;
  assign new_new_n4431__ = ~new_new_n3726__ & ~new_new_n4078__;
  assign new_new_n4432__ = ~new_new_n4219__ & new_new_n4431__;
  assign new_new_n4433__ = ~new_new_n4081__ & ~new_new_n4418__;
  assign new_new_n4434__ = ~new_new_n4430__ & ~new_new_n4432__;
  assign new_new_n4435__ = ~new_new_n4433__ & new_new_n4434__;
  assign new_new_n4436__ = ~new_new_n4429__ & ~new_new_n4435__;
  assign new_new_n4437__ = new_new_n4230__ & ~new_new_n4436__;
  assign new_new_n4438__ = new_new_n4222__ & ~new_new_n4431__;
  assign new_new_n4439__ = new_new_n4418__ & ~new_new_n4438__;
  assign new_new_n4440__ = ~new_new_n4219__ & new_new_n4433__;
  assign new_new_n4441__ = ~new_new_n4439__ & ~new_new_n4440__;
  assign new_new_n4442__ = ~new_new_n4230__ & ~new_new_n4441__;
  assign new_new_n4443__ = ~new_new_n4437__ & ~new_new_n4442__;
  assign new_new_n4444__ = ~new_new_n4420__ & new_new_n4443__;
  assign new_new_n4445__ = ~new_new_n3896__ & ~new_new_n4444__;
  assign new_new_n4446__ = new_new_n3898__ & new_new_n4444__;
  assign new_new_n4447__ = new_new_n3901__ & ~new_new_n4445__;
  assign new_new_n4448__ = ~new_new_n4446__ & new_new_n4447__;
  assign new_new_n4449__ = new_new_n4427__ & ~new_new_n4448__;
  assign new_new_n4450__ = new_new_n3777__ & ~new_new_n4427__;
  assign new_new_n4451__ = ~new_new_n4449__ & ~new_new_n4450__;
  assign new_new_n4452__ = ~new_new_n4411__ & new_new_n4451__;
  assign new_new_n4453__ = new_new_n4411__ & ~new_new_n4451__;
  assign new_new_n4454__ = ~new_new_n4452__ & ~new_new_n4453__;
  assign new_new_n4455__ = new_new_n4409__ & new_new_n4454__;
  assign new_new_n4456__ = ~new_new_n4409__ & ~new_new_n4454__;
  assign new_new_n4457__ = ~new_new_n4455__ & ~new_new_n4456__;
  assign new_new_n4458__ = new_new_n4311__ & new_new_n4457__;
  assign new_new_n4459__ = new_new_n223__ & ~new_new_n2500__;
  assign new_new_n4460__ = ~new_new_n321__ & ~new_new_n870__;
  assign new_new_n4461__ = ~new_new_n4459__ & new_new_n4460__;
  assign new_new_n4462__ = new_new_n3702__ & new_new_n4461__;
  assign new_new_n4463__ = new_new_n569__ & new_new_n4462__;
  assign new_new_n4464__ = new_new_n166__ & new_new_n213__;
  assign new_new_n4465__ = new_new_n223__ & ~new_new_n4464__;
  assign new_new_n4466__ = ~new_new_n160__ & ~new_new_n2683__;
  assign new_new_n4467__ = new_new_n115__ & new_new_n238__;
  assign new_new_n4468__ = new_new_n244__ & ~new_new_n4467__;
  assign new_new_n4469__ = ~new_new_n220__ & ~new_new_n403__;
  assign new_new_n4470__ = new_new_n969__ & ~new_new_n4468__;
  assign new_new_n4471__ = new_new_n4469__ & new_new_n4470__;
  assign new_new_n4472__ = ~new_new_n116__ & ~new_new_n413__;
  assign new_new_n4473__ = ~new_new_n793__ & ~new_new_n4472__;
  assign new_new_n4474__ = ~new_new_n245__ & ~new_new_n270__;
  assign new_new_n4475__ = ~new_new_n219__ & ~new_new_n252__;
  assign new_new_n4476__ = ~new_new_n188__ & new_new_n4475__;
  assign new_new_n4477__ = ~new_new_n546__ & ~new_new_n555__;
  assign new_new_n4478__ = ~new_new_n692__ & new_new_n4477__;
  assign new_new_n4479__ = ~new_new_n4474__ & new_new_n4476__;
  assign new_new_n4480__ = new_new_n4478__ & new_new_n4479__;
  assign new_new_n4481__ = new_new_n4471__ & ~new_new_n4473__;
  assign new_new_n4482__ = new_new_n4480__ & new_new_n4481__;
  assign new_new_n4483__ = ~new_new_n337__ & ~new_new_n348__;
  assign new_new_n4484__ = ~new_new_n4466__ & new_new_n4483__;
  assign new_new_n4485__ = new_new_n4482__ & new_new_n4484__;
  assign new_new_n4486__ = ~new_new_n383__ & ~new_new_n404__;
  assign new_new_n4487__ = ~new_new_n571__ & new_new_n4486__;
  assign new_new_n4488__ = ~new_new_n445__ & ~new_new_n471__;
  assign new_new_n4489__ = ~new_new_n595__ & ~new_new_n671__;
  assign new_new_n4490__ = new_new_n3616__ & ~new_new_n4465__;
  assign new_new_n4491__ = new_new_n4489__ & new_new_n4490__;
  assign new_new_n4492__ = new_new_n4487__ & new_new_n4488__;
  assign new_new_n4493__ = new_new_n4491__ & new_new_n4492__;
  assign new_new_n4494__ = new_new_n3695__ & new_new_n4493__;
  assign new_new_n4495__ = new_new_n538__ & new_new_n4494__;
  assign new_new_n4496__ = new_new_n4463__ & new_new_n4495__;
  assign new_new_n4497__ = new_new_n4485__ & new_new_n4496__;
  assign new_new_n4498__ = new_new_n4458__ & new_new_n4497__;
  assign new_new_n4499__ = ~new_new_n4311__ & ~new_new_n4457__;
  assign new_new_n4500__ = ~new_new_n4497__ & new_new_n4499__;
  assign new_new_n4501__ = ~new_new_n4498__ & ~new_new_n4500__;
  assign new_new_n4502__ = pi01 & ~new_new_n4418__;
  assign new_new_n4503__ = ~new_new_n1568__ & ~new_new_n4502__;
  assign new_new_n4504__ = new_new_n4412__ & ~new_new_n4503__;
  assign new_new_n4505__ = ~new_new_n4201__ & ~new_new_n4219__;
  assign new_new_n4506__ = new_new_n3735__ & new_new_n4505__;
  assign new_new_n4507__ = ~new_new_n4412__ & ~new_new_n4502__;
  assign new_new_n4508__ = ~new_new_n4506__ & new_new_n4507__;
  assign new_new_n4509__ = ~pi00 & ~new_new_n4504__;
  assign new_new_n4510__ = ~new_new_n4508__ & new_new_n4509__;
  assign new_new_n4511__ = ~new_new_n181__ & ~new_new_n861__;
  assign new_new_n4512__ = new_new_n227__ & new_new_n238__;
  assign new_new_n4513__ = new_new_n347__ & new_new_n4512__;
  assign new_new_n4514__ = ~new_new_n4511__ & ~new_new_n4513__;
  assign new_new_n4515__ = ~new_new_n136__ & ~new_new_n343__;
  assign new_new_n4516__ = ~new_new_n223__ & ~new_new_n921__;
  assign new_new_n4517__ = new_new_n221__ & new_new_n1095__;
  assign new_new_n4518__ = ~new_new_n4516__ & ~new_new_n4517__;
  assign new_new_n4519__ = ~new_new_n184__ & ~new_new_n384__;
  assign new_new_n4520__ = ~new_new_n4515__ & new_new_n4519__;
  assign new_new_n4521__ = ~new_new_n4518__ & new_new_n4520__;
  assign new_new_n4522__ = new_new_n166__ & new_new_n641__;
  assign new_new_n4523__ = new_new_n116__ & ~new_new_n4522__;
  assign new_new_n4524__ = new_new_n663__ & new_new_n1051__;
  assign new_new_n4525__ = ~new_new_n99__ & ~new_new_n4524__;
  assign new_new_n4526__ = ~new_new_n529__ & ~new_new_n692__;
  assign new_new_n4527__ = ~new_new_n4525__ & new_new_n4526__;
  assign new_new_n4528__ = ~new_new_n4523__ & new_new_n4527__;
  assign new_new_n4529__ = new_new_n3620__ & ~new_new_n4514__;
  assign new_new_n4530__ = new_new_n4521__ & new_new_n4529__;
  assign new_new_n4531__ = new_new_n4528__ & new_new_n4530__;
  assign new_new_n4532__ = new_new_n1106__ & new_new_n4531__;
  assign new_new_n4533__ = new_new_n3770__ & new_new_n4532__;
  assign new_new_n4534__ = new_new_n4078__ & new_new_n4219__;
  assign new_new_n4535__ = ~new_new_n4429__ & ~new_new_n4534__;
  assign new_new_n4536__ = new_new_n4532__ & ~new_new_n4535__;
  assign new_new_n4537__ = ~new_new_n4428__ & ~new_new_n4532__;
  assign new_new_n4538__ = ~new_new_n4534__ & new_new_n4537__;
  assign new_new_n4539__ = new_new_n4230__ & new_new_n4538__;
  assign new_new_n4540__ = ~new_new_n4536__ & ~new_new_n4539__;
  assign new_new_n4541__ = new_new_n4081__ & ~new_new_n4540__;
  assign new_new_n4542__ = ~new_new_n4418__ & new_new_n4532__;
  assign new_new_n4543__ = ~new_new_n4505__ & new_new_n4542__;
  assign new_new_n4544__ = new_new_n4201__ & ~new_new_n4418__;
  assign new_new_n4545__ = ~new_new_n4219__ & ~new_new_n4532__;
  assign new_new_n4546__ = ~new_new_n4431__ & new_new_n4545__;
  assign new_new_n4547__ = ~new_new_n4544__ & new_new_n4546__;
  assign new_new_n4548__ = ~new_new_n4543__ & ~new_new_n4547__;
  assign new_new_n4549__ = ~new_new_n4230__ & ~new_new_n4548__;
  assign new_new_n4550__ = new_new_n4418__ & ~new_new_n4532__;
  assign new_new_n4551__ = ~new_new_n4542__ & ~new_new_n4550__;
  assign new_new_n4552__ = ~new_new_n4430__ & new_new_n4551__;
  assign new_new_n4553__ = new_new_n4230__ & new_new_n4552__;
  assign new_new_n4554__ = ~new_new_n4078__ & ~new_new_n4418__;
  assign new_new_n4555__ = ~new_new_n4532__ & new_new_n4554__;
  assign new_new_n4556__ = ~new_new_n4553__ & ~new_new_n4555__;
  assign new_new_n4557__ = ~new_new_n4219__ & ~new_new_n4556__;
  assign new_new_n4558__ = ~new_new_n4081__ & ~new_new_n4551__;
  assign new_new_n4559__ = ~new_new_n4078__ & new_new_n4550__;
  assign new_new_n4560__ = ~new_new_n4558__ & ~new_new_n4559__;
  assign new_new_n4561__ = new_new_n4219__ & ~new_new_n4560__;
  assign new_new_n4562__ = ~new_new_n4549__ & ~new_new_n4561__;
  assign new_new_n4563__ = ~new_new_n4541__ & new_new_n4562__;
  assign new_new_n4564__ = ~new_new_n4557__ & new_new_n4563__;
  assign new_new_n4565__ = ~new_new_n3770__ & new_new_n4564__;
  assign new_new_n4566__ = pi00 & ~new_new_n4533__;
  assign new_new_n4567__ = ~new_new_n4565__ & new_new_n4566__;
  assign new_new_n4568__ = ~new_new_n4510__ & ~new_new_n4567__;
  assign new_new_n4569__ = new_new_n3233__ & new_new_n4568__;
  assign new_new_n4570__ = ~new_new_n3233__ & ~new_new_n4568__;
  assign new_new_n4571__ = ~new_new_n4569__ & ~new_new_n4570__;
  assign new_new_n4572__ = ~new_new_n4404__ & ~new_new_n4407__;
  assign new_new_n4573__ = new_new_n3604__ & ~new_new_n3727__;
  assign new_new_n4574__ = new_new_n3606__ & new_new_n3727__;
  assign new_new_n4575__ = new_new_n3235__ & new_new_n4171__;
  assign new_new_n4576__ = ~new_new_n3242__ & ~new_new_n4574__;
  assign new_new_n4577__ = ~new_new_n4575__ & new_new_n4576__;
  assign new_new_n4578__ = ~new_new_n310__ & ~new_new_n4577__;
  assign new_new_n4579__ = ~new_new_n4573__ & ~new_new_n4578__;
  assign new_new_n4580__ = ~new_new_n3236__ & ~new_new_n4579__;
  assign new_new_n4581__ = new_new_n3234__ & new_new_n4172__;
  assign new_new_n4582__ = ~new_new_n1324__ & new_new_n4086__;
  assign new_new_n4583__ = new_new_n310__ & ~new_new_n4086__;
  assign new_new_n4584__ = ~new_new_n4582__ & ~new_new_n4583__;
  assign new_new_n4585__ = ~new_new_n4081__ & ~new_new_n4584__;
  assign new_new_n4586__ = new_new_n4081__ & new_new_n4584__;
  assign new_new_n4587__ = new_new_n3236__ & new_new_n4579__;
  assign new_new_n4588__ = ~new_new_n4585__ & ~new_new_n4586__;
  assign new_new_n4589__ = new_new_n4587__ & new_new_n4588__;
  assign new_new_n4590__ = ~new_new_n4580__ & ~new_new_n4581__;
  assign new_new_n4591__ = ~new_new_n4589__ & new_new_n4590__;
  assign new_new_n4592__ = new_new_n4572__ & ~new_new_n4591__;
  assign new_new_n4593__ = ~new_new_n4572__ & new_new_n4591__;
  assign new_new_n4594__ = ~new_new_n4592__ & ~new_new_n4593__;
  assign new_new_n4595__ = ~new_new_n2784__ & new_new_n2809__;
  assign new_new_n4596__ = new_new_n2585__ & ~new_new_n2806__;
  assign new_new_n4597__ = ~new_new_n4595__ & ~new_new_n4596__;
  assign new_new_n4598__ = new_new_n2808__ & ~new_new_n3203__;
  assign new_new_n4599__ = ~new_new_n3111__ & new_new_n4598__;
  assign new_new_n4600__ = new_new_n4597__ & ~new_new_n4599__;
  assign new_new_n4601__ = ~new_new_n810__ & ~new_new_n4600__;
  assign new_new_n4602__ = ~new_new_n816__ & ~new_new_n3203__;
  assign new_new_n4603__ = new_new_n816__ & new_new_n3203__;
  assign new_new_n4604__ = new_new_n2808__ & ~new_new_n4602__;
  assign new_new_n4605__ = ~new_new_n4603__ & new_new_n4604__;
  assign new_new_n4606__ = new_new_n3111__ & new_new_n4605__;
  assign new_new_n4607__ = new_new_n2808__ & ~new_new_n3213__;
  assign new_new_n4608__ = new_new_n810__ & new_new_n4597__;
  assign new_new_n4609__ = ~new_new_n4607__ & new_new_n4608__;
  assign new_new_n4610__ = ~new_new_n4601__ & ~new_new_n4606__;
  assign new_new_n4611__ = ~new_new_n4609__ & new_new_n4610__;
  assign new_new_n4612__ = ~new_new_n4381__ & ~new_new_n4389__;
  assign new_new_n4613__ = ~new_new_n2608__ & ~new_new_n4612__;
  assign new_new_n4614__ = new_new_n2608__ & new_new_n4612__;
  assign new_new_n4615__ = ~new_new_n4613__ & ~new_new_n4614__;
  assign new_new_n4616__ = ~new_new_n437__ & ~new_new_n4615__;
  assign new_new_n4617__ = new_new_n2600__ & new_new_n3070__;
  assign new_new_n4618__ = new_new_n2604__ & ~new_new_n3065__;
  assign new_new_n4619__ = new_new_n2655__ & ~new_new_n3072__;
  assign new_new_n4620__ = ~new_new_n2590__ & new_new_n3072__;
  assign new_new_n4621__ = new_new_n2848__ & ~new_new_n4620__;
  assign new_new_n4622__ = ~new_new_n4619__ & new_new_n4621__;
  assign new_new_n4623__ = ~new_new_n4617__ & ~new_new_n4618__;
  assign new_new_n4624__ = ~new_new_n4622__ & new_new_n4623__;
  assign new_new_n4625__ = new_new_n4616__ & ~new_new_n4624__;
  assign new_new_n4626__ = ~new_new_n4616__ & new_new_n4624__;
  assign new_new_n4627__ = ~new_new_n4625__ & ~new_new_n4626__;
  assign new_new_n4628__ = new_new_n4611__ & new_new_n4627__;
  assign new_new_n4629__ = ~new_new_n4611__ & ~new_new_n4627__;
  assign new_new_n4630__ = ~new_new_n4628__ & ~new_new_n4629__;
  assign new_new_n4631__ = ~new_new_n4366__ & ~new_new_n4387__;
  assign new_new_n4632__ = ~new_new_n4365__ & ~new_new_n4631__;
  assign new_new_n4633__ = ~new_new_n4630__ & new_new_n4632__;
  assign new_new_n4634__ = new_new_n4630__ & ~new_new_n4632__;
  assign new_new_n4635__ = ~new_new_n4633__ & ~new_new_n4634__;
  assign new_new_n4636__ = new_new_n2593__ & ~new_new_n3486__;
  assign new_new_n4637__ = ~new_new_n320__ & ~new_new_n3586__;
  assign new_new_n4638__ = ~new_new_n4636__ & ~new_new_n4637__;
  assign new_new_n4639__ = ~new_new_n301__ & ~new_new_n4638__;
  assign new_new_n4640__ = ~new_new_n3651__ & ~new_new_n3654__;
  assign new_new_n4641__ = new_new_n2596__ & ~new_new_n4640__;
  assign new_new_n4642__ = new_new_n301__ & new_new_n4638__;
  assign new_new_n4643__ = ~new_new_n4641__ & new_new_n4642__;
  assign new_new_n4644__ = new_new_n301__ & ~new_new_n3654__;
  assign new_new_n4645__ = ~new_new_n316__ & new_new_n3654__;
  assign new_new_n4646__ = ~new_new_n3651__ & ~new_new_n4645__;
  assign new_new_n4647__ = new_new_n3651__ & new_new_n4645__;
  assign new_new_n4648__ = new_new_n2596__ & ~new_new_n4644__;
  assign new_new_n4649__ = ~new_new_n4646__ & new_new_n4648__;
  assign new_new_n4650__ = ~new_new_n4647__ & new_new_n4649__;
  assign new_new_n4651__ = ~new_new_n4639__ & ~new_new_n4643__;
  assign new_new_n4652__ = ~new_new_n4650__ & new_new_n4651__;
  assign new_new_n4653__ = ~new_new_n4635__ & ~new_new_n4652__;
  assign new_new_n4654__ = new_new_n4635__ & new_new_n4652__;
  assign new_new_n4655__ = ~new_new_n4653__ & ~new_new_n4654__;
  assign new_new_n4656__ = ~new_new_n4346__ & ~new_new_n4397__;
  assign new_new_n4657__ = ~new_new_n4396__ & ~new_new_n4656__;
  assign new_new_n4658__ = new_new_n4655__ & ~new_new_n4657__;
  assign new_new_n4659__ = ~new_new_n4655__ & new_new_n4657__;
  assign new_new_n4660__ = ~new_new_n4658__ & ~new_new_n4659__;
  assign new_new_n4661__ = new_new_n4594__ & new_new_n4660__;
  assign new_new_n4662__ = ~new_new_n4594__ & ~new_new_n4660__;
  assign new_new_n4663__ = ~new_new_n4661__ & ~new_new_n4662__;
  assign new_new_n4664__ = new_new_n4571__ & new_new_n4663__;
  assign new_new_n4665__ = ~new_new_n4571__ & ~new_new_n4663__;
  assign new_new_n4666__ = ~new_new_n4664__ & ~new_new_n4665__;
  assign new_new_n4667__ = new_new_n4409__ & ~new_new_n4453__;
  assign new_new_n4668__ = ~new_new_n4452__ & ~new_new_n4667__;
  assign new_new_n4669__ = new_new_n4666__ & ~new_new_n4668__;
  assign new_new_n4670__ = ~new_new_n4666__ & new_new_n4668__;
  assign new_new_n4671__ = ~new_new_n4669__ & ~new_new_n4670__;
  assign new_new_n4672__ = new_new_n116__ & ~new_new_n196__;
  assign new_new_n4673__ = ~new_new_n696__ & new_new_n4275__;
  assign new_new_n4674__ = ~new_new_n228__ & ~new_new_n475__;
  assign new_new_n4675__ = ~new_new_n690__ & ~new_new_n918__;
  assign new_new_n4676__ = new_new_n4674__ & new_new_n4675__;
  assign new_new_n4677__ = ~new_new_n322__ & ~new_new_n4672__;
  assign new_new_n4678__ = ~new_new_n4673__ & new_new_n4677__;
  assign new_new_n4679__ = new_new_n470__ & new_new_n4676__;
  assign new_new_n4680__ = new_new_n728__ & new_new_n4679__;
  assign new_new_n4681__ = new_new_n1449__ & new_new_n4678__;
  assign new_new_n4682__ = new_new_n3695__ & new_new_n4681__;
  assign new_new_n4683__ = new_new_n713__ & new_new_n4680__;
  assign new_new_n4684__ = new_new_n4682__ & new_new_n4683__;
  assign new_new_n4685__ = new_new_n502__ & new_new_n2563__;
  assign new_new_n4686__ = new_new_n4684__ & new_new_n4685__;
  assign new_new_n4687__ = ~new_new_n4671__ & ~new_new_n4686__;
  assign new_new_n4688__ = ~new_new_n909__ & ~new_new_n4671__;
  assign new_new_n4689__ = new_new_n4671__ & new_new_n4686__;
  assign new_new_n4690__ = ~new_new_n4688__ & ~new_new_n4689__;
  assign new_new_n4691__ = ~new_new_n4687__ & new_new_n4690__;
  assign new_new_n4692__ = ~new_new_n4501__ & new_new_n4691__;
  assign new_new_n4693__ = new_new_n4501__ & ~new_new_n4691__;
  assign po00 = new_new_n4692__ | new_new_n4693__;
  assign new_new_n4695__ = new_new_n4500__ & new_new_n4687__;
  assign new_new_n4696__ = new_new_n4498__ & new_new_n4689__;
  assign new_new_n4697__ = ~new_new_n4500__ & new_new_n4689__;
  assign new_new_n4698__ = new_new_n4498__ & ~new_new_n4687__;
  assign new_new_n4699__ = ~new_new_n4697__ & ~new_new_n4698__;
  assign new_new_n4700__ = pi22 & ~pi23;
  assign new_new_n4701__ = ~pi22 & pi23;
  assign new_new_n4702__ = ~new_new_n4700__ & ~new_new_n4701__;
  assign new_new_n4703__ = ~new_new_n4699__ & new_new_n4702__;
  assign new_new_n4704__ = ~new_new_n4500__ & ~new_new_n4687__;
  assign new_new_n4705__ = ~new_new_n4498__ & ~new_new_n4702__;
  assign new_new_n4706__ = ~new_new_n4689__ & new_new_n4705__;
  assign new_new_n4707__ = ~new_new_n4704__ & new_new_n4706__;
  assign new_new_n4708__ = ~new_new_n4695__ & ~new_new_n4696__;
  assign new_new_n4709__ = ~new_new_n4707__ & new_new_n4708__;
  assign new_new_n4710__ = ~new_new_n4703__ & new_new_n4709__;
  assign new_new_n4711__ = new_new_n244__ & ~new_new_n663__;
  assign new_new_n4712__ = new_new_n223__ & ~new_new_n4512__;
  assign new_new_n4713__ = ~new_new_n925__ & ~new_new_n1124__;
  assign new_new_n4714__ = ~new_new_n4712__ & new_new_n4713__;
  assign new_new_n4715__ = ~new_new_n186__ & new_new_n4714__;
  assign new_new_n4716__ = ~new_new_n244__ & new_new_n256__;
  assign new_new_n4717__ = ~new_new_n181__ & new_new_n347__;
  assign new_new_n4718__ = ~new_new_n4716__ & ~new_new_n4717__;
  assign new_new_n4719__ = ~new_new_n744__ & ~new_new_n1033__;
  assign new_new_n4720__ = ~new_new_n4718__ & new_new_n4719__;
  assign new_new_n4721__ = ~new_new_n274__ & ~new_new_n921__;
  assign new_new_n4722__ = ~new_new_n951__ & new_new_n4721__;
  assign new_new_n4723__ = ~new_new_n324__ & ~new_new_n471__;
  assign new_new_n4724__ = ~new_new_n4711__ & new_new_n4723__;
  assign new_new_n4725__ = ~new_new_n342__ & new_new_n4722__;
  assign new_new_n4726__ = new_new_n728__ & new_new_n4725__;
  assign new_new_n4727__ = new_new_n3695__ & new_new_n4724__;
  assign new_new_n4728__ = new_new_n4715__ & new_new_n4720__;
  assign new_new_n4729__ = new_new_n4727__ & new_new_n4728__;
  assign new_new_n4730__ = new_new_n4726__ & new_new_n4729__;
  assign new_new_n4731__ = new_new_n2678__ & new_new_n4482__;
  assign new_new_n4732__ = new_new_n4730__ & new_new_n4731__;
  assign new_new_n4733__ = new_new_n1324__ & new_new_n4233__;
  assign new_new_n4734__ = ~new_new_n4222__ & ~new_new_n4733__;
  assign new_new_n4735__ = new_new_n4222__ & new_new_n4733__;
  assign new_new_n4736__ = new_new_n3236__ & ~new_new_n4734__;
  assign new_new_n4737__ = ~new_new_n4735__ & new_new_n4736__;
  assign new_new_n4738__ = new_new_n4233__ & new_new_n4737__;
  assign new_new_n4739__ = new_new_n3247__ & ~new_new_n3727__;
  assign new_new_n4740__ = new_new_n3240__ & new_new_n4081__;
  assign new_new_n4741__ = ~new_new_n4739__ & ~new_new_n4740__;
  assign new_new_n4742__ = ~new_new_n4737__ & new_new_n4741__;
  assign new_new_n4743__ = new_new_n310__ & ~new_new_n4742__;
  assign new_new_n4744__ = ~new_new_n4222__ & ~new_new_n4233__;
  assign new_new_n4745__ = new_new_n3236__ & ~new_new_n4744__;
  assign new_new_n4746__ = ~new_new_n310__ & new_new_n4741__;
  assign new_new_n4747__ = ~new_new_n4745__ & new_new_n4746__;
  assign new_new_n4748__ = ~new_new_n4738__ & ~new_new_n4747__;
  assign new_new_n4749__ = ~new_new_n4743__ & new_new_n4748__;
  assign new_new_n4750__ = ~new_new_n4732__ & ~new_new_n4749__;
  assign new_new_n4751__ = new_new_n4732__ & new_new_n4749__;
  assign new_new_n4752__ = ~new_new_n4750__ & ~new_new_n4751__;
  assign new_new_n4753__ = new_new_n2809__ & ~new_new_n3203__;
  assign new_new_n4754__ = ~new_new_n2784__ & ~new_new_n2806__;
  assign new_new_n4755__ = ~new_new_n4753__ & ~new_new_n4754__;
  assign new_new_n4756__ = new_new_n2808__ & new_new_n3490__;
  assign new_new_n4757__ = new_new_n4755__ & ~new_new_n4756__;
  assign new_new_n4758__ = new_new_n810__ & ~new_new_n4757__;
  assign new_new_n4759__ = ~new_new_n816__ & new_new_n3486__;
  assign new_new_n4760__ = new_new_n816__ & ~new_new_n3486__;
  assign new_new_n4761__ = new_new_n2808__ & ~new_new_n4759__;
  assign new_new_n4762__ = ~new_new_n4760__ & new_new_n4761__;
  assign new_new_n4763__ = new_new_n3489__ & new_new_n4762__;
  assign new_new_n4764__ = new_new_n2808__ & ~new_new_n3499__;
  assign new_new_n4765__ = ~new_new_n810__ & new_new_n4755__;
  assign new_new_n4766__ = ~new_new_n4764__ & new_new_n4765__;
  assign new_new_n4767__ = ~new_new_n4763__ & ~new_new_n4766__;
  assign new_new_n4768__ = ~new_new_n4758__ & new_new_n4767__;
  assign new_new_n4769__ = ~new_new_n4611__ & new_new_n4627__;
  assign new_new_n4770__ = ~new_new_n4633__ & ~new_new_n4769__;
  assign new_new_n4771__ = ~new_new_n4768__ & new_new_n4770__;
  assign new_new_n4772__ = new_new_n4768__ & ~new_new_n4770__;
  assign new_new_n4773__ = ~new_new_n4771__ & ~new_new_n4772__;
  assign new_new_n4774__ = ~new_new_n4614__ & ~new_new_n4624__;
  assign new_new_n4775__ = ~new_new_n437__ & ~new_new_n4613__;
  assign new_new_n4776__ = ~new_new_n4774__ & new_new_n4775__;
  assign new_new_n4777__ = new_new_n2604__ & new_new_n4776__;
  assign new_new_n4778__ = ~new_new_n2604__ & ~new_new_n4776__;
  assign new_new_n4779__ = ~new_new_n4777__ & ~new_new_n4778__;
  assign new_new_n4780__ = ~new_new_n437__ & ~new_new_n4779__;
  assign new_new_n4781__ = ~new_new_n2590__ & new_new_n3070__;
  assign new_new_n4782__ = new_new_n2585__ & new_new_n3072__;
  assign new_new_n4783__ = ~new_new_n3030__ & ~new_new_n3072__;
  assign new_new_n4784__ = new_new_n2848__ & ~new_new_n4782__;
  assign new_new_n4785__ = ~new_new_n4783__ & new_new_n4784__;
  assign new_new_n4786__ = ~new_new_n437__ & new_new_n2600__;
  assign new_new_n4787__ = ~new_new_n651__ & new_new_n2846__;
  assign new_new_n4788__ = ~new_new_n4786__ & new_new_n4787__;
  assign new_new_n4789__ = new_new_n437__ & new_new_n2600__;
  assign new_new_n4790__ = new_new_n810__ & new_new_n3068__;
  assign new_new_n4791__ = ~new_new_n4789__ & new_new_n4790__;
  assign new_new_n4792__ = ~new_new_n4788__ & ~new_new_n4791__;
  assign new_new_n4793__ = ~new_new_n4781__ & new_new_n4792__;
  assign new_new_n4794__ = ~new_new_n4785__ & new_new_n4793__;
  assign new_new_n4795__ = new_new_n4780__ & new_new_n4794__;
  assign new_new_n4796__ = ~new_new_n4777__ & ~new_new_n4794__;
  assign new_new_n4797__ = ~new_new_n4780__ & new_new_n4796__;
  assign new_new_n4798__ = ~new_new_n4795__ & ~new_new_n4797__;
  assign new_new_n4799__ = new_new_n4773__ & ~new_new_n4798__;
  assign new_new_n4800__ = ~new_new_n4777__ & new_new_n4794__;
  assign new_new_n4801__ = ~new_new_n4780__ & ~new_new_n4800__;
  assign new_new_n4802__ = ~new_new_n4795__ & ~new_new_n4801__;
  assign new_new_n4803__ = ~new_new_n4773__ & new_new_n4802__;
  assign new_new_n4804__ = ~new_new_n4799__ & ~new_new_n4803__;
  assign new_new_n4805__ = ~new_new_n316__ & ~new_new_n3733__;
  assign new_new_n4806__ = new_new_n316__ & new_new_n3733__;
  assign new_new_n4807__ = ~new_new_n4805__ & ~new_new_n4806__;
  assign new_new_n4808__ = new_new_n4024__ & ~new_new_n4807__;
  assign new_new_n4809__ = new_new_n301__ & new_new_n4167__;
  assign new_new_n4810__ = ~new_new_n4808__ & ~new_new_n4809__;
  assign new_new_n4811__ = new_new_n2596__ & ~new_new_n4810__;
  assign new_new_n4812__ = ~new_new_n320__ & new_new_n3651__;
  assign new_new_n4813__ = new_new_n2593__ & ~new_new_n3586__;
  assign new_new_n4814__ = ~new_new_n4812__ & ~new_new_n4813__;
  assign new_new_n4815__ = new_new_n301__ & ~new_new_n4814__;
  assign new_new_n4816__ = new_new_n2596__ & ~new_new_n4176__;
  assign new_new_n4817__ = ~new_new_n301__ & new_new_n4814__;
  assign new_new_n4818__ = ~new_new_n4816__ & new_new_n4817__;
  assign new_new_n4819__ = ~new_new_n4815__ & ~new_new_n4818__;
  assign new_new_n4820__ = ~new_new_n4811__ & new_new_n4819__;
  assign new_new_n4821__ = new_new_n4804__ & new_new_n4820__;
  assign new_new_n4822__ = ~new_new_n4804__ & ~new_new_n4820__;
  assign new_new_n4823__ = ~new_new_n4821__ & ~new_new_n4822__;
  assign new_new_n4824__ = ~new_new_n4654__ & ~new_new_n4657__;
  assign new_new_n4825__ = ~new_new_n4653__ & ~new_new_n4824__;
  assign new_new_n4826__ = new_new_n4823__ & ~new_new_n4825__;
  assign new_new_n4827__ = ~new_new_n4823__ & new_new_n4825__;
  assign new_new_n4828__ = ~new_new_n4826__ & ~new_new_n4827__;
  assign new_new_n4829__ = new_new_n4412__ & new_new_n4418__;
  assign new_new_n4830__ = pi01 & ~new_new_n4532__;
  assign new_new_n4831__ = ~new_new_n1568__ & ~new_new_n4830__;
  assign new_new_n4832__ = new_new_n4829__ & ~new_new_n4831__;
  assign new_new_n4833__ = ~new_new_n3735__ & ~new_new_n4418__;
  assign new_new_n4834__ = new_new_n4421__ & ~new_new_n4833__;
  assign new_new_n4835__ = ~new_new_n4830__ & ~new_new_n4834__;
  assign new_new_n4836__ = ~pi00 & ~new_new_n4832__;
  assign new_new_n4837__ = ~new_new_n4835__ & new_new_n4836__;
  assign new_new_n4838__ = new_new_n449__ & new_new_n990__;
  assign new_new_n4839__ = new_new_n195__ & ~new_new_n4838__;
  assign new_new_n4840__ = new_new_n181__ & ~new_new_n4467__;
  assign new_new_n4841__ = ~new_new_n219__ & ~new_new_n870__;
  assign new_new_n4842__ = ~new_new_n4840__ & new_new_n4841__;
  assign new_new_n4843__ = ~new_new_n342__ & ~new_new_n4839__;
  assign new_new_n4844__ = new_new_n4842__ & new_new_n4843__;
  assign new_new_n4845__ = new_new_n661__ & new_new_n4844__;
  assign new_new_n4846__ = new_new_n162__ & ~new_new_n543__;
  assign new_new_n4847__ = ~new_new_n248__ & ~new_new_n4846__;
  assign new_new_n4848__ = ~new_new_n379__ & ~new_new_n410__;
  assign new_new_n4849__ = new_new_n562__ & new_new_n4848__;
  assign new_new_n4850__ = new_new_n2310__ & new_new_n4847__;
  assign new_new_n4851__ = new_new_n4849__ & new_new_n4850__;
  assign new_new_n4852__ = new_new_n1470__ & new_new_n4851__;
  assign new_new_n4853__ = new_new_n440__ & new_new_n4852__;
  assign new_new_n4854__ = new_new_n4845__ & new_new_n4853__;
  assign new_new_n4855__ = new_new_n4412__ & new_new_n4532__;
  assign new_new_n4856__ = new_new_n2468__ & new_new_n4854__;
  assign new_new_n4857__ = ~new_new_n4855__ & new_new_n4856__;
  assign new_new_n4858__ = new_new_n3770__ & new_new_n4857__;
  assign new_new_n4859__ = ~new_new_n4421__ & ~new_new_n4532__;
  assign new_new_n4860__ = new_new_n4421__ & new_new_n4532__;
  assign new_new_n4861__ = ~new_new_n4859__ & ~new_new_n4860__;
  assign new_new_n4862__ = new_new_n4857__ & new_new_n4861__;
  assign new_new_n4863__ = ~new_new_n4421__ & new_new_n4857__;
  assign new_new_n4864__ = new_new_n4222__ & new_new_n4863__;
  assign new_new_n4865__ = ~new_new_n4857__ & new_new_n4860__;
  assign new_new_n4866__ = new_new_n4230__ & new_new_n4865__;
  assign new_new_n4867__ = ~new_new_n4864__ & ~new_new_n4866__;
  assign new_new_n4868__ = new_new_n4081__ & ~new_new_n4867__;
  assign new_new_n4869__ = new_new_n4421__ & new_new_n4857__;
  assign new_new_n4870__ = ~new_new_n4222__ & new_new_n4869__;
  assign new_new_n4871__ = ~new_new_n4857__ & new_new_n4859__;
  assign new_new_n4872__ = ~new_new_n4230__ & new_new_n4871__;
  assign new_new_n4873__ = ~new_new_n4870__ & ~new_new_n4872__;
  assign new_new_n4874__ = ~new_new_n4081__ & ~new_new_n4873__;
  assign new_new_n4875__ = new_new_n4230__ & new_new_n4863__;
  assign new_new_n4876__ = new_new_n4222__ & ~new_new_n4865__;
  assign new_new_n4877__ = ~new_new_n4875__ & new_new_n4876__;
  assign new_new_n4878__ = ~new_new_n4230__ & new_new_n4869__;
  assign new_new_n4879__ = ~new_new_n4222__ & ~new_new_n4871__;
  assign new_new_n4880__ = ~new_new_n4878__ & new_new_n4879__;
  assign new_new_n4881__ = ~new_new_n4877__ & ~new_new_n4880__;
  assign new_new_n4882__ = ~new_new_n4862__ & ~new_new_n4868__;
  assign new_new_n4883__ = ~new_new_n4874__ & ~new_new_n4881__;
  assign new_new_n4884__ = new_new_n4882__ & new_new_n4883__;
  assign new_new_n4885__ = ~new_new_n3770__ & ~new_new_n4884__;
  assign new_new_n4886__ = pi00 & ~new_new_n4858__;
  assign new_new_n4887__ = ~new_new_n4885__ & new_new_n4886__;
  assign new_new_n4888__ = ~new_new_n4837__ & ~new_new_n4887__;
  assign new_new_n4889__ = new_new_n3233__ & new_new_n4888__;
  assign new_new_n4890__ = ~new_new_n3233__ & ~new_new_n4888__;
  assign new_new_n4891__ = ~new_new_n4889__ & ~new_new_n4890__;
  assign new_new_n4892__ = ~new_new_n4664__ & ~new_new_n4668__;
  assign new_new_n4893__ = ~new_new_n4665__ & ~new_new_n4892__;
  assign new_new_n4894__ = new_new_n4572__ & new_new_n4591__;
  assign new_new_n4895__ = ~new_new_n4572__ & ~new_new_n4591__;
  assign new_new_n4896__ = ~new_new_n4660__ & ~new_new_n4895__;
  assign new_new_n4897__ = ~new_new_n4894__ & ~new_new_n4896__;
  assign new_new_n4898__ = ~new_new_n4893__ & new_new_n4897__;
  assign new_new_n4899__ = new_new_n4893__ & ~new_new_n4897__;
  assign new_new_n4900__ = ~new_new_n4898__ & ~new_new_n4899__;
  assign new_new_n4901__ = new_new_n4891__ & ~new_new_n4900__;
  assign new_new_n4902__ = ~new_new_n4891__ & new_new_n4900__;
  assign new_new_n4903__ = ~new_new_n4901__ & ~new_new_n4902__;
  assign new_new_n4904__ = new_new_n4828__ & new_new_n4903__;
  assign new_new_n4905__ = ~new_new_n4828__ & ~new_new_n4903__;
  assign new_new_n4906__ = ~new_new_n4904__ & ~new_new_n4905__;
  assign new_new_n4907__ = new_new_n4752__ & new_new_n4906__;
  assign new_new_n4908__ = ~new_new_n4471__ & new_new_n4732__;
  assign new_new_n4909__ = ~new_new_n4752__ & ~new_new_n4908__;
  assign new_new_n4910__ = ~new_new_n4906__ & new_new_n4909__;
  assign new_new_n4911__ = ~new_new_n4907__ & ~new_new_n4910__;
  assign new_new_n4912__ = new_new_n4710__ & new_new_n4911__;
  assign new_new_n4913__ = ~new_new_n4710__ & ~new_new_n4911__;
  assign po01 = new_new_n4912__ | new_new_n4913__;
  assign new_new_n4915__ = new_new_n4222__ & ~new_new_n4231__;
  assign new_new_n4916__ = ~new_new_n4421__ & ~new_new_n4915__;
  assign new_new_n4917__ = ~new_new_n4532__ & ~new_new_n4916__;
  assign new_new_n4918__ = new_new_n4857__ & ~new_new_n4917__;
  assign new_new_n4919__ = ~new_new_n4222__ & ~new_new_n4232__;
  assign new_new_n4920__ = new_new_n4421__ & ~new_new_n4919__;
  assign new_new_n4921__ = new_new_n4532__ & ~new_new_n4920__;
  assign new_new_n4922__ = ~new_new_n4857__ & ~new_new_n4921__;
  assign new_new_n4923__ = ~new_new_n4918__ & ~new_new_n4922__;
  assign new_new_n4924__ = pi01 & new_new_n4923__;
  assign new_new_n4925__ = pi02 & ~new_new_n4923__;
  assign new_new_n4926__ = ~new_new_n4924__ & ~new_new_n4925__;
  assign new_new_n4927__ = pi22 & ~new_new_n4926__;
  assign new_new_n4928__ = ~pi22 & new_new_n4926__;
  assign new_new_n4929__ = pi00 & ~new_new_n4927__;
  assign new_new_n4930__ = ~new_new_n4928__ & new_new_n4929__;
  assign new_new_n4931__ = new_new_n3735__ & new_new_n4532__;
  assign new_new_n4932__ = new_new_n3765__ & ~new_new_n4854__;
  assign new_new_n4933__ = ~new_new_n3776__ & ~new_new_n4857__;
  assign new_new_n4934__ = new_new_n3776__ & new_new_n4857__;
  assign new_new_n4935__ = pi01 & ~new_new_n4932__;
  assign new_new_n4936__ = ~new_new_n4933__ & new_new_n4935__;
  assign new_new_n4937__ = ~new_new_n4934__ & new_new_n4936__;
  assign new_new_n4938__ = ~pi00 & ~new_new_n4931__;
  assign new_new_n4939__ = ~new_new_n4937__ & new_new_n4938__;
  assign new_new_n4940__ = ~new_new_n4930__ & ~new_new_n4939__;
  assign new_new_n4941__ = new_new_n2593__ & new_new_n3651__;
  assign new_new_n4942__ = ~new_new_n320__ & ~new_new_n3733__;
  assign new_new_n4943__ = ~new_new_n4941__ & ~new_new_n4942__;
  assign new_new_n4944__ = new_new_n2596__ & ~new_new_n4325__;
  assign new_new_n4945__ = ~new_new_n301__ & ~new_new_n4944__;
  assign new_new_n4946__ = ~new_new_n316__ & ~new_new_n4319__;
  assign new_new_n4947__ = new_new_n316__ & ~new_new_n4321__;
  assign new_new_n4948__ = new_new_n2596__ & ~new_new_n4946__;
  assign new_new_n4949__ = ~new_new_n4947__ & new_new_n4948__;
  assign new_new_n4950__ = ~new_new_n4945__ & ~new_new_n4949__;
  assign new_new_n4951__ = new_new_n4943__ & ~new_new_n4950__;
  assign new_new_n4952__ = new_new_n2596__ & new_new_n4315__;
  assign new_new_n4953__ = new_new_n4943__ & ~new_new_n4952__;
  assign new_new_n4954__ = new_new_n301__ & ~new_new_n4953__;
  assign new_new_n4955__ = ~new_new_n4951__ & ~new_new_n4954__;
  assign new_new_n4956__ = new_new_n2809__ & ~new_new_n3486__;
  assign new_new_n4957__ = ~new_new_n2806__ & ~new_new_n3203__;
  assign new_new_n4958__ = ~new_new_n4956__ & ~new_new_n4957__;
  assign new_new_n4959__ = new_new_n2808__ & new_new_n3587__;
  assign new_new_n4960__ = new_new_n4958__ & ~new_new_n4959__;
  assign new_new_n4961__ = new_new_n810__ & ~new_new_n4960__;
  assign new_new_n4962__ = ~new_new_n816__ & new_new_n3586__;
  assign new_new_n4963__ = new_new_n816__ & ~new_new_n3586__;
  assign new_new_n4964__ = new_new_n2808__ & new_new_n3515__;
  assign new_new_n4965__ = ~new_new_n4962__ & ~new_new_n4963__;
  assign new_new_n4966__ = new_new_n4964__ & new_new_n4965__;
  assign new_new_n4967__ = new_new_n2808__ & ~new_new_n3596__;
  assign new_new_n4968__ = ~new_new_n810__ & new_new_n4958__;
  assign new_new_n4969__ = ~new_new_n4967__ & new_new_n4968__;
  assign new_new_n4970__ = ~new_new_n4966__ & ~new_new_n4969__;
  assign new_new_n4971__ = ~new_new_n4961__ & new_new_n4970__;
  assign new_new_n4972__ = ~new_new_n4772__ & ~new_new_n4798__;
  assign new_new_n4973__ = ~new_new_n4771__ & ~new_new_n4972__;
  assign new_new_n4974__ = new_new_n4971__ & new_new_n4973__;
  assign new_new_n4975__ = ~new_new_n4971__ & ~new_new_n4973__;
  assign new_new_n4976__ = ~new_new_n4974__ & ~new_new_n4975__;
  assign new_new_n4977__ = new_new_n2590__ & ~new_new_n3065__;
  assign new_new_n4978__ = new_new_n2585__ & new_new_n3070__;
  assign new_new_n4979__ = new_new_n2664__ & ~new_new_n3072__;
  assign new_new_n4980__ = new_new_n2784__ & ~new_new_n4979__;
  assign new_new_n4981__ = ~new_new_n2784__ & new_new_n4979__;
  assign new_new_n4982__ = new_new_n2848__ & ~new_new_n4980__;
  assign new_new_n4983__ = ~new_new_n4981__ & new_new_n4982__;
  assign new_new_n4984__ = ~new_new_n4977__ & ~new_new_n4978__;
  assign new_new_n4985__ = ~new_new_n4983__ & new_new_n4984__;
  assign new_new_n4986__ = new_new_n437__ & ~new_new_n4985__;
  assign new_new_n4987__ = ~new_new_n2600__ & ~new_new_n4985__;
  assign new_new_n4988__ = new_new_n2600__ & new_new_n4985__;
  assign new_new_n4989__ = ~new_new_n4987__ & ~new_new_n4988__;
  assign new_new_n4990__ = ~new_new_n4789__ & ~new_new_n4794__;
  assign new_new_n4991__ = ~new_new_n4776__ & ~new_new_n4990__;
  assign new_new_n4992__ = new_new_n2604__ & ~new_new_n4991__;
  assign new_new_n4993__ = ~new_new_n4989__ & new_new_n4992__;
  assign new_new_n4994__ = new_new_n4776__ & ~new_new_n4794__;
  assign new_new_n4995__ = ~new_new_n4989__ & new_new_n4994__;
  assign new_new_n4996__ = new_new_n437__ & ~new_new_n2600__;
  assign new_new_n4997__ = ~new_new_n4778__ & ~new_new_n4800__;
  assign new_new_n4998__ = ~new_new_n4996__ & ~new_new_n4997__;
  assign new_new_n4999__ = new_new_n4989__ & new_new_n4998__;
  assign new_new_n5000__ = ~new_new_n4986__ & ~new_new_n4993__;
  assign new_new_n5001__ = ~new_new_n4995__ & ~new_new_n4999__;
  assign new_new_n5002__ = new_new_n5000__ & new_new_n5001__;
  assign new_new_n5003__ = ~new_new_n4976__ & new_new_n5002__;
  assign new_new_n5004__ = new_new_n4976__ & ~new_new_n5002__;
  assign new_new_n5005__ = ~new_new_n5003__ & ~new_new_n5004__;
  assign new_new_n5006__ = ~new_new_n4822__ & ~new_new_n4825__;
  assign new_new_n5007__ = ~new_new_n4821__ & ~new_new_n5006__;
  assign new_new_n5008__ = new_new_n5005__ & new_new_n5007__;
  assign new_new_n5009__ = ~new_new_n5005__ & ~new_new_n5007__;
  assign new_new_n5010__ = ~new_new_n5008__ & ~new_new_n5009__;
  assign new_new_n5011__ = new_new_n4955__ & ~new_new_n5010__;
  assign new_new_n5012__ = ~new_new_n4955__ & new_new_n5010__;
  assign new_new_n5013__ = ~new_new_n5011__ & ~new_new_n5012__;
  assign new_new_n5014__ = new_new_n4940__ & new_new_n5013__;
  assign new_new_n5015__ = ~new_new_n4940__ & ~new_new_n5013__;
  assign new_new_n5016__ = ~new_new_n5014__ & ~new_new_n5015__;
  assign new_new_n5017__ = new_new_n4749__ & ~new_new_n4897__;
  assign new_new_n5018__ = ~new_new_n4749__ & new_new_n4897__;
  assign new_new_n5019__ = ~new_new_n4828__ & ~new_new_n5018__;
  assign new_new_n5020__ = ~new_new_n5017__ & ~new_new_n5019__;
  assign new_new_n5021__ = ~new_new_n4891__ & ~new_new_n4893__;
  assign new_new_n5022__ = new_new_n4891__ & new_new_n4893__;
  assign new_new_n5023__ = ~new_new_n5017__ & ~new_new_n5018__;
  assign new_new_n5024__ = new_new_n4828__ & new_new_n5023__;
  assign new_new_n5025__ = ~new_new_n4828__ & ~new_new_n5023__;
  assign new_new_n5026__ = ~new_new_n5024__ & ~new_new_n5025__;
  assign new_new_n5027__ = ~new_new_n5022__ & new_new_n5026__;
  assign new_new_n5028__ = ~new_new_n5021__ & ~new_new_n5027__;
  assign new_new_n5029__ = ~new_new_n5020__ & new_new_n5028__;
  assign new_new_n5030__ = new_new_n5020__ & ~new_new_n5028__;
  assign new_new_n5031__ = ~new_new_n5029__ & ~new_new_n5030__;
  assign new_new_n5032__ = new_new_n4419__ & new_new_n4443__;
  assign new_new_n5033__ = new_new_n3267__ & new_new_n5032__;
  assign new_new_n5034__ = new_new_n3247__ & new_new_n4081__;
  assign new_new_n5035__ = new_new_n3240__ & new_new_n4222__;
  assign new_new_n5036__ = ~new_new_n5034__ & ~new_new_n5035__;
  assign new_new_n5037__ = ~new_new_n4421__ & ~new_new_n4444__;
  assign new_new_n5038__ = new_new_n3236__ & ~new_new_n5037__;
  assign new_new_n5039__ = new_new_n310__ & ~new_new_n5038__;
  assign new_new_n5040__ = new_new_n4421__ & ~new_new_n4443__;
  assign new_new_n5041__ = new_new_n3274__ & new_new_n5040__;
  assign new_new_n5042__ = ~new_new_n5039__ & ~new_new_n5041__;
  assign new_new_n5043__ = new_new_n5036__ & ~new_new_n5042__;
  assign new_new_n5044__ = new_new_n3236__ & new_new_n4421__;
  assign new_new_n5045__ = new_new_n4444__ & new_new_n5044__;
  assign new_new_n5046__ = new_new_n5036__ & ~new_new_n5045__;
  assign new_new_n5047__ = ~new_new_n310__ & ~new_new_n5046__;
  assign new_new_n5048__ = ~new_new_n5033__ & ~new_new_n5047__;
  assign new_new_n5049__ = ~new_new_n5043__ & new_new_n5048__;
  assign new_new_n5050__ = new_new_n5031__ & ~new_new_n5049__;
  assign new_new_n5051__ = ~new_new_n5031__ & new_new_n5049__;
  assign new_new_n5052__ = ~new_new_n5050__ & ~new_new_n5051__;
  assign new_new_n5053__ = new_new_n5016__ & new_new_n5052__;
  assign new_new_n5054__ = ~new_new_n5016__ & ~new_new_n5052__;
  assign new_new_n5055__ = ~new_new_n5053__ & ~new_new_n5054__;
  assign new_new_n5056__ = new_new_n4732__ & new_new_n4911__;
  assign new_new_n5057__ = ~new_new_n4458__ & ~new_new_n4497__;
  assign new_new_n5058__ = ~new_new_n4499__ & ~new_new_n5057__;
  assign new_new_n5059__ = ~new_new_n4689__ & ~new_new_n5058__;
  assign new_new_n5060__ = ~new_new_n4687__ & ~new_new_n5059__;
  assign new_new_n5061__ = ~new_new_n4911__ & new_new_n5060__;
  assign new_new_n5062__ = ~new_new_n5056__ & ~new_new_n5061__;
  assign new_new_n5063__ = new_new_n5055__ & new_new_n5062__;
  assign new_new_n5064__ = ~new_new_n5055__ & ~new_new_n5062__;
  assign new_new_n5065__ = ~new_new_n5063__ & ~new_new_n5064__;
  assign new_new_n5066__ = ~new_new_n124__ & ~new_new_n1051__;
  assign new_new_n5067__ = new_new_n218__ & ~new_new_n5066__;
  assign new_new_n5068__ = ~new_new_n190__ & ~new_new_n5067__;
  assign new_new_n5069__ = new_new_n160__ & new_new_n174__;
  assign new_new_n5070__ = new_new_n116__ & ~new_new_n5069__;
  assign new_new_n5071__ = ~new_new_n328__ & ~new_new_n5070__;
  assign new_new_n5072__ = ~new_new_n5068__ & new_new_n5071__;
  assign new_new_n5073__ = new_new_n238__ & new_new_n265__;
  assign new_new_n5074__ = ~new_new_n277__ & new_new_n5073__;
  assign new_new_n5075__ = new_new_n180__ & new_new_n256__;
  assign new_new_n5076__ = ~new_new_n195__ & new_new_n5075__;
  assign new_new_n5077__ = ~new_new_n2250__ & ~new_new_n5074__;
  assign new_new_n5078__ = ~new_new_n5076__ & new_new_n5077__;
  assign new_new_n5079__ = new_new_n162__ & ~new_new_n174__;
  assign new_new_n5080__ = ~new_new_n918__ & ~new_new_n1124__;
  assign new_new_n5081__ = ~new_new_n161__ & new_new_n5080__;
  assign new_new_n5082__ = ~new_new_n5079__ & new_new_n5081__;
  assign new_new_n5083__ = ~new_new_n694__ & new_new_n5082__;
  assign new_new_n5084__ = new_new_n5072__ & ~new_new_n5078__;
  assign new_new_n5085__ = new_new_n5083__ & new_new_n5084__;
  assign new_new_n5086__ = new_new_n468__ & new_new_n5085__;
  assign new_new_n5087__ = new_new_n209__ & new_new_n5086__;
  assign new_new_n5088__ = ~new_new_n5065__ & new_new_n5087__;
  assign new_new_n5089__ = new_new_n5065__ & ~new_new_n5087__;
  assign new_new_n5090__ = ~new_new_n5088__ & ~new_new_n5089__;
  assign new_new_n5091__ = new_new_n4498__ & new_new_n4687__;
  assign new_new_n5092__ = new_new_n4690__ & ~new_new_n5058__;
  assign new_new_n5093__ = new_new_n4704__ & new_new_n5092__;
  assign new_new_n5094__ = ~new_new_n5091__ & ~new_new_n5093__;
  assign new_new_n5095__ = ~new_new_n4911__ & ~new_new_n5094__;
  assign new_new_n5096__ = new_new_n4696__ & new_new_n4911__;
  assign new_new_n5097__ = ~new_new_n5095__ & ~new_new_n5096__;
  assign new_new_n5098__ = ~new_new_n4702__ & new_new_n5097__;
  assign new_new_n5099__ = ~new_new_n5090__ & ~new_new_n5098__;
  assign new_new_n5100__ = new_new_n4500__ & new_new_n4689__;
  assign new_new_n5101__ = ~new_new_n4498__ & new_new_n5058__;
  assign new_new_n5102__ = new_new_n4691__ & new_new_n5101__;
  assign new_new_n5103__ = ~new_new_n5100__ & ~new_new_n5102__;
  assign new_new_n5104__ = ~new_new_n4911__ & ~new_new_n5103__;
  assign new_new_n5105__ = new_new_n4695__ & new_new_n4911__;
  assign new_new_n5106__ = ~new_new_n5104__ & ~new_new_n5105__;
  assign new_new_n5107__ = new_new_n5099__ & new_new_n5106__;
  assign new_new_n5108__ = new_new_n4702__ & new_new_n5106__;
  assign new_new_n5109__ = new_new_n5097__ & ~new_new_n5108__;
  assign new_new_n5110__ = new_new_n5090__ & new_new_n5109__;
  assign po02 = ~new_new_n5107__ & ~new_new_n5110__;
  assign new_new_n5112__ = ~new_new_n5099__ & ~new_new_n5108__;
  assign new_new_n5113__ = ~pi01 & ~new_new_n4857__;
  assign new_new_n5114__ = new_new_n3230__ & ~new_new_n5113__;
  assign new_new_n5115__ = ~pi00 & ~pi22;
  assign new_new_n5116__ = new_new_n3769__ & new_new_n5115__;
  assign new_new_n5117__ = new_new_n4219__ & ~new_new_n4431__;
  assign new_new_n5118__ = new_new_n4230__ & ~new_new_n5117__;
  assign new_new_n5119__ = ~new_new_n4505__ & ~new_new_n5118__;
  assign new_new_n5120__ = ~new_new_n4418__ & ~new_new_n5119__;
  assign new_new_n5121__ = new_new_n4532__ & ~new_new_n4829__;
  assign new_new_n5122__ = ~new_new_n5120__ & new_new_n5121__;
  assign new_new_n5123__ = new_new_n3776__ & new_new_n5122__;
  assign new_new_n5124__ = new_new_n3231__ & new_new_n4857__;
  assign new_new_n5125__ = ~new_new_n3761__ & ~new_new_n4857__;
  assign new_new_n5126__ = ~new_new_n5124__ & ~new_new_n5125__;
  assign new_new_n5127__ = ~new_new_n5122__ & new_new_n5126__;
  assign new_new_n5128__ = pi00 & ~new_new_n5123__;
  assign new_new_n5129__ = ~new_new_n5127__ & new_new_n5128__;
  assign new_new_n5130__ = ~new_new_n5114__ & ~new_new_n5116__;
  assign new_new_n5131__ = ~new_new_n5129__ & new_new_n5130__;
  assign new_new_n5132__ = new_new_n318__ & new_new_n4805__;
  assign new_new_n5133__ = ~new_new_n301__ & ~new_new_n4086__;
  assign new_new_n5134__ = new_new_n316__ & new_new_n4086__;
  assign new_new_n5135__ = ~new_new_n5133__ & ~new_new_n5134__;
  assign new_new_n5136__ = new_new_n4081__ & new_new_n5135__;
  assign new_new_n5137__ = ~new_new_n4081__ & ~new_new_n5135__;
  assign new_new_n5138__ = new_new_n2596__ & ~new_new_n5136__;
  assign new_new_n5139__ = ~new_new_n5137__ & new_new_n5138__;
  assign new_new_n5140__ = ~new_new_n317__ & ~new_new_n318__;
  assign new_new_n5141__ = new_new_n3727__ & ~new_new_n5140__;
  assign new_new_n5142__ = ~new_new_n318__ & ~new_new_n4806__;
  assign new_new_n5143__ = ~new_new_n311__ & new_new_n316__;
  assign new_new_n5144__ = ~new_new_n5142__ & ~new_new_n5143__;
  assign new_new_n5145__ = ~new_new_n5141__ & ~new_new_n5144__;
  assign new_new_n5146__ = new_new_n301__ & ~new_new_n5145__;
  assign new_new_n5147__ = ~new_new_n301__ & ~new_new_n320__;
  assign new_new_n5148__ = ~new_new_n3727__ & new_new_n5147__;
  assign new_new_n5149__ = ~new_new_n5132__ & ~new_new_n5148__;
  assign new_new_n5150__ = ~new_new_n5146__ & new_new_n5149__;
  assign new_new_n5151__ = ~new_new_n5139__ & new_new_n5150__;
  assign new_new_n5152__ = ~new_new_n2806__ & ~new_new_n3486__;
  assign new_new_n5153__ = new_new_n2809__ & ~new_new_n3586__;
  assign new_new_n5154__ = ~new_new_n5152__ & ~new_new_n5153__;
  assign new_new_n5155__ = new_new_n2808__ & ~new_new_n3654__;
  assign new_new_n5156__ = new_new_n3651__ & new_new_n5155__;
  assign new_new_n5157__ = new_new_n5154__ & ~new_new_n5156__;
  assign new_new_n5158__ = ~new_new_n810__ & ~new_new_n5157__;
  assign new_new_n5159__ = new_new_n816__ & ~new_new_n3651__;
  assign new_new_n5160__ = ~new_new_n816__ & new_new_n3651__;
  assign new_new_n5161__ = new_new_n2808__ & new_new_n3654__;
  assign new_new_n5162__ = ~new_new_n5159__ & new_new_n5161__;
  assign new_new_n5163__ = ~new_new_n5160__ & new_new_n5162__;
  assign new_new_n5164__ = new_new_n2808__ & ~new_new_n4640__;
  assign new_new_n5165__ = new_new_n810__ & new_new_n5154__;
  assign new_new_n5166__ = ~new_new_n5164__ & new_new_n5165__;
  assign new_new_n5167__ = ~new_new_n5158__ & ~new_new_n5163__;
  assign new_new_n5168__ = ~new_new_n5166__ & new_new_n5167__;
  assign new_new_n5169__ = ~new_new_n4975__ & ~new_new_n5002__;
  assign new_new_n5170__ = ~new_new_n4974__ & ~new_new_n5169__;
  assign new_new_n5171__ = new_new_n5168__ & new_new_n5170__;
  assign new_new_n5172__ = ~new_new_n5168__ & ~new_new_n5170__;
  assign new_new_n5173__ = ~new_new_n5171__ & ~new_new_n5172__;
  assign new_new_n5174__ = ~new_new_n2600__ & ~new_new_n4997__;
  assign new_new_n5175__ = ~new_new_n2604__ & new_new_n4794__;
  assign new_new_n5176__ = new_new_n4776__ & ~new_new_n5175__;
  assign new_new_n5177__ = new_new_n2604__ & ~new_new_n4794__;
  assign new_new_n5178__ = ~new_new_n4985__ & ~new_new_n5177__;
  assign new_new_n5179__ = ~new_new_n437__ & ~new_new_n5178__;
  assign new_new_n5180__ = ~new_new_n5176__ & ~new_new_n5179__;
  assign new_new_n5181__ = ~new_new_n4987__ & ~new_new_n5174__;
  assign new_new_n5182__ = ~new_new_n5180__ & new_new_n5181__;
  assign new_new_n5183__ = new_new_n2590__ & new_new_n5182__;
  assign new_new_n5184__ = ~new_new_n2590__ & ~new_new_n5182__;
  assign new_new_n5185__ = ~new_new_n5183__ & ~new_new_n5184__;
  assign new_new_n5186__ = ~new_new_n437__ & ~new_new_n5185__;
  assign new_new_n5187__ = new_new_n2585__ & ~new_new_n3065__;
  assign new_new_n5188__ = ~new_new_n2784__ & new_new_n3070__;
  assign new_new_n5189__ = ~new_new_n3072__ & new_new_n3111__;
  assign new_new_n5190__ = new_new_n3203__ & ~new_new_n5189__;
  assign new_new_n5191__ = ~new_new_n3203__ & new_new_n5189__;
  assign new_new_n5192__ = new_new_n2848__ & ~new_new_n5190__;
  assign new_new_n5193__ = ~new_new_n5191__ & new_new_n5192__;
  assign new_new_n5194__ = ~new_new_n5187__ & ~new_new_n5188__;
  assign new_new_n5195__ = ~new_new_n5193__ & new_new_n5194__;
  assign new_new_n5196__ = new_new_n5186__ & ~new_new_n5195__;
  assign new_new_n5197__ = ~new_new_n5183__ & new_new_n5195__;
  assign new_new_n5198__ = ~new_new_n5186__ & new_new_n5197__;
  assign new_new_n5199__ = ~new_new_n5196__ & ~new_new_n5198__;
  assign new_new_n5200__ = ~new_new_n5173__ & ~new_new_n5199__;
  assign new_new_n5201__ = ~new_new_n5183__ & ~new_new_n5195__;
  assign new_new_n5202__ = ~new_new_n5186__ & ~new_new_n5201__;
  assign new_new_n5203__ = ~new_new_n5196__ & ~new_new_n5202__;
  assign new_new_n5204__ = new_new_n5173__ & new_new_n5203__;
  assign new_new_n5205__ = ~new_new_n5200__ & ~new_new_n5204__;
  assign new_new_n5206__ = new_new_n5151__ & new_new_n5205__;
  assign new_new_n5207__ = ~new_new_n5151__ & ~new_new_n5205__;
  assign new_new_n5208__ = ~new_new_n5206__ & ~new_new_n5207__;
  assign new_new_n5209__ = new_new_n4955__ & ~new_new_n5008__;
  assign new_new_n5210__ = ~new_new_n5009__ & ~new_new_n5209__;
  assign new_new_n5211__ = new_new_n5208__ & ~new_new_n5210__;
  assign new_new_n5212__ = ~new_new_n5208__ & new_new_n5210__;
  assign new_new_n5213__ = ~new_new_n5211__ & ~new_new_n5212__;
  assign new_new_n5214__ = ~new_new_n4532__ & new_new_n4564__;
  assign new_new_n5215__ = new_new_n3267__ & new_new_n5214__;
  assign new_new_n5216__ = new_new_n3240__ & new_new_n4421__;
  assign new_new_n5217__ = new_new_n3247__ & new_new_n4222__;
  assign new_new_n5218__ = ~new_new_n5216__ & ~new_new_n5217__;
  assign new_new_n5219__ = new_new_n4532__ & new_new_n4564__;
  assign new_new_n5220__ = new_new_n3236__ & ~new_new_n5219__;
  assign new_new_n5221__ = ~new_new_n310__ & ~new_new_n5220__;
  assign new_new_n5222__ = new_new_n4532__ & ~new_new_n4564__;
  assign new_new_n5223__ = new_new_n3274__ & new_new_n5222__;
  assign new_new_n5224__ = ~new_new_n5221__ & ~new_new_n5223__;
  assign new_new_n5225__ = new_new_n5218__ & ~new_new_n5224__;
  assign new_new_n5226__ = ~new_new_n4532__ & ~new_new_n4564__;
  assign new_new_n5227__ = new_new_n3236__ & new_new_n5226__;
  assign new_new_n5228__ = new_new_n5218__ & ~new_new_n5227__;
  assign new_new_n5229__ = new_new_n310__ & ~new_new_n5228__;
  assign new_new_n5230__ = ~new_new_n5215__ & ~new_new_n5229__;
  assign new_new_n5231__ = ~new_new_n5225__ & new_new_n5230__;
  assign new_new_n5232__ = new_new_n5213__ & ~new_new_n5231__;
  assign new_new_n5233__ = ~new_new_n5213__ & new_new_n5231__;
  assign new_new_n5234__ = ~new_new_n5232__ & ~new_new_n5233__;
  assign new_new_n5235__ = new_new_n5131__ & new_new_n5234__;
  assign new_new_n5236__ = ~new_new_n5131__ & ~new_new_n5234__;
  assign new_new_n5237__ = ~new_new_n5235__ & ~new_new_n5236__;
  assign new_new_n5238__ = new_new_n5015__ & new_new_n5049__;
  assign new_new_n5239__ = new_new_n5014__ & ~new_new_n5049__;
  assign new_new_n5240__ = ~new_new_n5238__ & ~new_new_n5239__;
  assign new_new_n5241__ = new_new_n5031__ & new_new_n5240__;
  assign new_new_n5242__ = ~new_new_n5015__ & ~new_new_n5049__;
  assign new_new_n5243__ = ~new_new_n5014__ & ~new_new_n5242__;
  assign new_new_n5244__ = new_new_n5030__ & ~new_new_n5243__;
  assign new_new_n5245__ = new_new_n5029__ & new_new_n5243__;
  assign new_new_n5246__ = ~new_new_n5237__ & ~new_new_n5244__;
  assign new_new_n5247__ = ~new_new_n5245__ & new_new_n5246__;
  assign new_new_n5248__ = ~new_new_n5241__ & new_new_n5247__;
  assign new_new_n5249__ = new_new_n4940__ & ~new_new_n5020__;
  assign new_new_n5250__ = new_new_n5028__ & new_new_n5249__;
  assign new_new_n5251__ = new_new_n5013__ & new_new_n5250__;
  assign new_new_n5252__ = ~new_new_n4940__ & new_new_n5020__;
  assign new_new_n5253__ = ~new_new_n5028__ & ~new_new_n5249__;
  assign new_new_n5254__ = ~new_new_n5252__ & ~new_new_n5253__;
  assign new_new_n5255__ = new_new_n5013__ & new_new_n5254__;
  assign new_new_n5256__ = ~new_new_n5250__ & ~new_new_n5255__;
  assign new_new_n5257__ = ~new_new_n5049__ & ~new_new_n5256__;
  assign new_new_n5258__ = ~new_new_n5028__ & new_new_n5252__;
  assign new_new_n5259__ = new_new_n5013__ & ~new_new_n5258__;
  assign new_new_n5260__ = new_new_n5049__ & ~new_new_n5254__;
  assign new_new_n5261__ = ~new_new_n5259__ & new_new_n5260__;
  assign new_new_n5262__ = ~new_new_n5013__ & ~new_new_n5028__;
  assign new_new_n5263__ = new_new_n5252__ & new_new_n5262__;
  assign new_new_n5264__ = new_new_n5237__ & ~new_new_n5251__;
  assign new_new_n5265__ = ~new_new_n5263__ & new_new_n5264__;
  assign new_new_n5266__ = ~new_new_n5261__ & new_new_n5265__;
  assign new_new_n5267__ = ~new_new_n5257__ & new_new_n5266__;
  assign new_new_n5268__ = ~new_new_n5248__ & ~new_new_n5267__;
  assign new_new_n5269__ = ~new_new_n5112__ & new_new_n5268__;
  assign new_new_n5270__ = new_new_n5112__ & ~new_new_n5268__;
  assign new_new_n5271__ = ~new_new_n5269__ & ~new_new_n5270__;
  assign new_new_n5272__ = ~new_new_n162__ & ~new_new_n244__;
  assign new_new_n5273__ = ~new_new_n81__ & ~new_new_n5272__;
  assign new_new_n5274__ = ~new_new_n244__ & new_new_n343__;
  assign new_new_n5275__ = ~new_new_n227__ & ~new_new_n5274__;
  assign new_new_n5276__ = ~new_new_n176__ & ~new_new_n324__;
  assign new_new_n5277__ = new_new_n4273__ & new_new_n5276__;
  assign new_new_n5278__ = ~new_new_n5273__ & ~new_new_n5275__;
  assign new_new_n5279__ = new_new_n5277__ & new_new_n5278__;
  assign new_new_n5280__ = new_new_n899__ & new_new_n4267__;
  assign new_new_n5281__ = new_new_n5279__ & new_new_n5280__;
  assign new_new_n5282__ = new_new_n421__ & new_new_n593__;
  assign new_new_n5283__ = new_new_n2706__ & new_new_n5282__;
  assign new_new_n5284__ = new_new_n1462__ & new_new_n5281__;
  assign new_new_n5285__ = new_new_n5283__ & new_new_n5284__;
  assign new_new_n5286__ = ~new_new_n5064__ & ~new_new_n5087__;
  assign new_new_n5287__ = ~new_new_n5063__ & ~new_new_n5286__;
  assign new_new_n5288__ = new_new_n5285__ & ~new_new_n5287__;
  assign new_new_n5289__ = ~new_new_n5285__ & new_new_n5287__;
  assign new_new_n5290__ = ~new_new_n5288__ & ~new_new_n5289__;
  assign new_new_n5291__ = new_new_n5271__ & new_new_n5290__;
  assign new_new_n5292__ = ~new_new_n5271__ & ~new_new_n5290__;
  assign po03 = new_new_n5291__ | new_new_n5292__;
  assign new_new_n5294__ = new_new_n5268__ & new_new_n5285__;
  assign new_new_n5295__ = ~new_new_n5268__ & ~new_new_n5285__;
  assign new_new_n5296__ = ~new_new_n5294__ & ~new_new_n5295__;
  assign new_new_n5297__ = ~new_new_n5064__ & ~new_new_n5296__;
  assign new_new_n5298__ = ~new_new_n5063__ & new_new_n5296__;
  assign new_new_n5299__ = new_new_n5087__ & ~new_new_n5297__;
  assign new_new_n5300__ = ~new_new_n5298__ & new_new_n5299__;
  assign new_new_n5301__ = new_new_n5286__ & new_new_n5298__;
  assign new_new_n5302__ = ~new_new_n5300__ & ~new_new_n5301__;
  assign new_new_n5303__ = ~new_new_n5097__ & ~new_new_n5302__;
  assign new_new_n5304__ = new_new_n5286__ & new_new_n5296__;
  assign new_new_n5305__ = ~new_new_n5063__ & ~new_new_n5296__;
  assign new_new_n5306__ = ~new_new_n5088__ & ~new_new_n5106__;
  assign new_new_n5307__ = ~new_new_n5304__ & ~new_new_n5305__;
  assign new_new_n5308__ = new_new_n5306__ & new_new_n5307__;
  assign new_new_n5309__ = new_new_n4702__ & ~new_new_n5308__;
  assign new_new_n5310__ = ~new_new_n5303__ & ~new_new_n5309__;
  assign new_new_n5311__ = new_new_n5237__ & new_new_n5262__;
  assign new_new_n5312__ = new_new_n5013__ & new_new_n5028__;
  assign new_new_n5313__ = new_new_n5237__ & ~new_new_n5249__;
  assign new_new_n5314__ = ~new_new_n5237__ & ~new_new_n5252__;
  assign new_new_n5315__ = new_new_n5049__ & ~new_new_n5314__;
  assign new_new_n5316__ = ~new_new_n5313__ & ~new_new_n5315__;
  assign new_new_n5317__ = ~new_new_n5312__ & ~new_new_n5316__;
  assign new_new_n5318__ = ~new_new_n5049__ & ~new_new_n5252__;
  assign new_new_n5319__ = ~new_new_n5237__ & ~new_new_n5262__;
  assign new_new_n5320__ = ~new_new_n5249__ & ~new_new_n5318__;
  assign new_new_n5321__ = ~new_new_n5319__ & new_new_n5320__;
  assign new_new_n5322__ = ~new_new_n5311__ & ~new_new_n5317__;
  assign new_new_n5323__ = ~new_new_n5321__ & new_new_n5322__;
  assign new_new_n5324__ = new_new_n5131__ & ~new_new_n5233__;
  assign new_new_n5325__ = ~new_new_n5232__ & ~new_new_n5324__;
  assign new_new_n5326__ = ~new_new_n5323__ & ~new_new_n5325__;
  assign new_new_n5327__ = new_new_n5323__ & new_new_n5325__;
  assign new_new_n5328__ = ~new_new_n5326__ & ~new_new_n5327__;
  assign new_new_n5329__ = ~new_new_n5206__ & ~new_new_n5210__;
  assign new_new_n5330__ = ~new_new_n5207__ & ~new_new_n5329__;
  assign new_new_n5331__ = new_new_n3247__ & new_new_n4421__;
  assign new_new_n5332__ = new_new_n3240__ & ~new_new_n4532__;
  assign new_new_n5333__ = ~new_new_n5331__ & ~new_new_n5332__;
  assign new_new_n5334__ = new_new_n3236__ & ~new_new_n4857__;
  assign new_new_n5335__ = new_new_n4884__ & new_new_n5334__;
  assign new_new_n5336__ = new_new_n5333__ & ~new_new_n5335__;
  assign new_new_n5337__ = ~new_new_n310__ & ~new_new_n5336__;
  assign new_new_n5338__ = new_new_n4857__ & ~new_new_n4884__;
  assign new_new_n5339__ = new_new_n3236__ & ~new_new_n5338__;
  assign new_new_n5340__ = new_new_n310__ & new_new_n5333__;
  assign new_new_n5341__ = ~new_new_n5339__ & new_new_n5340__;
  assign new_new_n5342__ = ~new_new_n1324__ & ~new_new_n4857__;
  assign new_new_n5343__ = new_new_n1324__ & new_new_n4884__;
  assign new_new_n5344__ = ~new_new_n5342__ & ~new_new_n5343__;
  assign new_new_n5345__ = new_new_n5339__ & new_new_n5344__;
  assign new_new_n5346__ = ~new_new_n5337__ & ~new_new_n5341__;
  assign new_new_n5347__ = ~new_new_n5345__ & new_new_n5346__;
  assign new_new_n5348__ = ~new_new_n5330__ & new_new_n5347__;
  assign new_new_n5349__ = new_new_n5330__ & ~new_new_n5347__;
  assign new_new_n5350__ = ~new_new_n5348__ & ~new_new_n5349__;
  assign new_new_n5351__ = ~new_new_n5171__ & new_new_n5199__;
  assign new_new_n5352__ = ~new_new_n5172__ & ~new_new_n5351__;
  assign new_new_n5353__ = ~new_new_n316__ & new_new_n4233__;
  assign new_new_n5354__ = ~new_new_n4222__ & ~new_new_n5353__;
  assign new_new_n5355__ = new_new_n4222__ & new_new_n5353__;
  assign new_new_n5356__ = new_new_n2596__ & ~new_new_n5354__;
  assign new_new_n5357__ = ~new_new_n5355__ & new_new_n5356__;
  assign new_new_n5358__ = new_new_n4233__ & new_new_n5357__;
  assign new_new_n5359__ = new_new_n2593__ & ~new_new_n3727__;
  assign new_new_n5360__ = ~new_new_n320__ & new_new_n4081__;
  assign new_new_n5361__ = ~new_new_n5359__ & ~new_new_n5360__;
  assign new_new_n5362__ = ~new_new_n5357__ & new_new_n5361__;
  assign new_new_n5363__ = ~new_new_n301__ & ~new_new_n5362__;
  assign new_new_n5364__ = new_new_n2596__ & ~new_new_n4744__;
  assign new_new_n5365__ = new_new_n301__ & new_new_n5361__;
  assign new_new_n5366__ = ~new_new_n5364__ & new_new_n5365__;
  assign new_new_n5367__ = ~new_new_n5358__ & ~new_new_n5366__;
  assign new_new_n5368__ = ~new_new_n5363__ & new_new_n5367__;
  assign new_new_n5369__ = new_new_n5352__ & ~new_new_n5368__;
  assign new_new_n5370__ = ~new_new_n5352__ & new_new_n5368__;
  assign new_new_n5371__ = ~new_new_n5369__ & ~new_new_n5370__;
  assign new_new_n5372__ = new_new_n2809__ & new_new_n3651__;
  assign new_new_n5373__ = ~new_new_n2806__ & ~new_new_n3586__;
  assign new_new_n5374__ = ~new_new_n5372__ & ~new_new_n5373__;
  assign new_new_n5375__ = new_new_n2808__ & new_new_n4167__;
  assign new_new_n5376__ = new_new_n5374__ & ~new_new_n5375__;
  assign new_new_n5377__ = new_new_n810__ & ~new_new_n5376__;
  assign new_new_n5378__ = new_new_n816__ & ~new_new_n3733__;
  assign new_new_n5379__ = ~new_new_n816__ & new_new_n3733__;
  assign new_new_n5380__ = new_new_n2808__ & new_new_n4024__;
  assign new_new_n5381__ = ~new_new_n5378__ & ~new_new_n5379__;
  assign new_new_n5382__ = new_new_n5380__ & new_new_n5381__;
  assign new_new_n5383__ = new_new_n2808__ & ~new_new_n4176__;
  assign new_new_n5384__ = ~new_new_n810__ & new_new_n5374__;
  assign new_new_n5385__ = ~new_new_n5383__ & new_new_n5384__;
  assign new_new_n5386__ = ~new_new_n5382__ & ~new_new_n5385__;
  assign new_new_n5387__ = ~new_new_n5377__ & new_new_n5386__;
  assign new_new_n5388__ = ~new_new_n5184__ & ~new_new_n5201__;
  assign new_new_n5389__ = ~new_new_n437__ & new_new_n2585__;
  assign new_new_n5390__ = ~new_new_n5388__ & new_new_n5389__;
  assign new_new_n5391__ = ~new_new_n437__ & new_new_n5388__;
  assign new_new_n5392__ = ~new_new_n2585__ & new_new_n5391__;
  assign new_new_n5393__ = ~new_new_n5390__ & ~new_new_n5392__;
  assign new_new_n5394__ = new_new_n3070__ & ~new_new_n3203__;
  assign new_new_n5395__ = ~new_new_n2784__ & ~new_new_n3065__;
  assign new_new_n5396__ = ~new_new_n5394__ & ~new_new_n5395__;
  assign new_new_n5397__ = new_new_n2848__ & new_new_n3490__;
  assign new_new_n5398__ = new_new_n5396__ & ~new_new_n5397__;
  assign new_new_n5399__ = ~new_new_n437__ & ~new_new_n5398__;
  assign new_new_n5400__ = new_new_n651__ & new_new_n3486__;
  assign new_new_n5401__ = ~new_new_n651__ & ~new_new_n3486__;
  assign new_new_n5402__ = new_new_n2848__ & ~new_new_n5400__;
  assign new_new_n5403__ = ~new_new_n5401__ & new_new_n5402__;
  assign new_new_n5404__ = new_new_n3489__ & new_new_n5403__;
  assign new_new_n5405__ = new_new_n2848__ & ~new_new_n3499__;
  assign new_new_n5406__ = new_new_n437__ & new_new_n5396__;
  assign new_new_n5407__ = ~new_new_n5405__ & new_new_n5406__;
  assign new_new_n5408__ = ~new_new_n5404__ & ~new_new_n5407__;
  assign new_new_n5409__ = ~new_new_n5399__ & new_new_n5408__;
  assign new_new_n5410__ = ~new_new_n3233__ & new_new_n5409__;
  assign new_new_n5411__ = new_new_n3233__ & ~new_new_n5409__;
  assign new_new_n5412__ = ~new_new_n5410__ & ~new_new_n5411__;
  assign new_new_n5413__ = new_new_n5393__ & ~new_new_n5412__;
  assign new_new_n5414__ = ~new_new_n5393__ & new_new_n5412__;
  assign new_new_n5415__ = ~new_new_n5413__ & ~new_new_n5414__;
  assign new_new_n5416__ = new_new_n5387__ & new_new_n5415__;
  assign new_new_n5417__ = ~new_new_n5387__ & ~new_new_n5415__;
  assign new_new_n5418__ = ~new_new_n5416__ & ~new_new_n5417__;
  assign new_new_n5419__ = new_new_n5371__ & new_new_n5418__;
  assign new_new_n5420__ = ~new_new_n5371__ & ~new_new_n5418__;
  assign new_new_n5421__ = ~new_new_n5419__ & ~new_new_n5420__;
  assign new_new_n5422__ = new_new_n5350__ & ~new_new_n5421__;
  assign new_new_n5423__ = ~new_new_n5350__ & new_new_n5421__;
  assign new_new_n5424__ = ~new_new_n5422__ & ~new_new_n5423__;
  assign new_new_n5425__ = new_new_n5328__ & new_new_n5424__;
  assign new_new_n5426__ = ~new_new_n5328__ & ~new_new_n5424__;
  assign new_new_n5427__ = ~new_new_n5425__ & ~new_new_n5426__;
  assign new_new_n5428__ = new_new_n160__ & new_new_n270__;
  assign new_new_n5429__ = new_new_n116__ & ~new_new_n5428__;
  assign new_new_n5430__ = ~new_new_n793__ & ~new_new_n4717__;
  assign new_new_n5431__ = ~new_new_n4291__ & new_new_n5430__;
  assign new_new_n5432__ = ~new_new_n137__ & ~new_new_n267__;
  assign new_new_n5433__ = ~new_new_n257__ & ~new_new_n2230__;
  assign new_new_n5434__ = ~new_new_n5429__ & new_new_n5433__;
  assign new_new_n5435__ = new_new_n5432__ & new_new_n5434__;
  assign new_new_n5436__ = new_new_n727__ & ~new_new_n5431__;
  assign new_new_n5437__ = new_new_n5435__ & new_new_n5436__;
  assign new_new_n5438__ = new_new_n964__ & new_new_n5437__;
  assign new_new_n5439__ = new_new_n2342__ & new_new_n5438__;
  assign new_new_n5440__ = new_new_n391__ & new_new_n5439__;
  assign new_new_n5441__ = ~new_new_n5427__ & ~new_new_n5440__;
  assign new_new_n5442__ = new_new_n5427__ & new_new_n5440__;
  assign new_new_n5443__ = ~new_new_n5441__ & ~new_new_n5442__;
  assign new_new_n5444__ = ~new_new_n5287__ & ~new_new_n5294__;
  assign new_new_n5445__ = ~new_new_n5295__ & ~new_new_n5444__;
  assign new_new_n5446__ = new_new_n5443__ & ~new_new_n5445__;
  assign new_new_n5447__ = ~new_new_n5443__ & new_new_n5445__;
  assign new_new_n5448__ = ~new_new_n5446__ & ~new_new_n5447__;
  assign new_new_n5449__ = ~new_new_n5310__ & new_new_n5448__;
  assign new_new_n5450__ = new_new_n5303__ & ~new_new_n5308__;
  assign new_new_n5451__ = ~new_new_n5309__ & ~new_new_n5448__;
  assign new_new_n5452__ = ~new_new_n5450__ & new_new_n5451__;
  assign po04 = new_new_n5449__ | new_new_n5452__;
  assign new_new_n5454__ = ~new_new_n5325__ & new_new_n5347__;
  assign new_new_n5455__ = ~new_new_n5323__ & ~new_new_n5330__;
  assign new_new_n5456__ = new_new_n5454__ & new_new_n5455__;
  assign new_new_n5457__ = new_new_n5325__ & ~new_new_n5347__;
  assign new_new_n5458__ = new_new_n5323__ & ~new_new_n5454__;
  assign new_new_n5459__ = ~new_new_n5457__ & ~new_new_n5458__;
  assign new_new_n5460__ = ~new_new_n5330__ & new_new_n5459__;
  assign new_new_n5461__ = new_new_n5326__ & new_new_n5347__;
  assign new_new_n5462__ = ~new_new_n5460__ & ~new_new_n5461__;
  assign new_new_n5463__ = ~new_new_n5421__ & ~new_new_n5462__;
  assign new_new_n5464__ = new_new_n5330__ & ~new_new_n5459__;
  assign new_new_n5465__ = new_new_n5327__ & ~new_new_n5347__;
  assign new_new_n5466__ = ~new_new_n5464__ & ~new_new_n5465__;
  assign new_new_n5467__ = new_new_n5421__ & ~new_new_n5466__;
  assign new_new_n5468__ = new_new_n5323__ & new_new_n5330__;
  assign new_new_n5469__ = new_new_n5457__ & new_new_n5468__;
  assign new_new_n5470__ = new_new_n3240__ & ~new_new_n4857__;
  assign new_new_n5471__ = new_new_n3247__ & ~new_new_n4532__;
  assign new_new_n5472__ = ~new_new_n5470__ & ~new_new_n5471__;
  assign new_new_n5473__ = ~new_new_n310__ & ~new_new_n5472__;
  assign new_new_n5474__ = new_new_n3267__ & new_new_n4923__;
  assign new_new_n5475__ = new_new_n3236__ & new_new_n4923__;
  assign new_new_n5476__ = new_new_n310__ & new_new_n5472__;
  assign new_new_n5477__ = ~new_new_n5475__ & new_new_n5476__;
  assign new_new_n5478__ = ~new_new_n5473__ & ~new_new_n5474__;
  assign new_new_n5479__ = ~new_new_n5477__ & new_new_n5478__;
  assign new_new_n5480__ = new_new_n2585__ & ~new_new_n5412__;
  assign new_new_n5481__ = ~new_new_n5387__ & ~new_new_n5480__;
  assign new_new_n5482__ = new_new_n5387__ & new_new_n5480__;
  assign new_new_n5483__ = ~new_new_n5388__ & ~new_new_n5482__;
  assign new_new_n5484__ = ~new_new_n437__ & ~new_new_n5481__;
  assign new_new_n5485__ = ~new_new_n5483__ & new_new_n5484__;
  assign new_new_n5486__ = ~new_new_n5387__ & ~new_new_n5391__;
  assign new_new_n5487__ = ~new_new_n5389__ & new_new_n5412__;
  assign new_new_n5488__ = ~new_new_n5486__ & new_new_n5487__;
  assign new_new_n5489__ = ~new_new_n5485__ & ~new_new_n5488__;
  assign new_new_n5490__ = ~new_new_n316__ & new_new_n2596__;
  assign new_new_n5491__ = new_new_n5040__ & new_new_n5490__;
  assign new_new_n5492__ = new_new_n2593__ & new_new_n4081__;
  assign new_new_n5493__ = ~new_new_n320__ & new_new_n4222__;
  assign new_new_n5494__ = ~new_new_n5492__ & ~new_new_n5493__;
  assign new_new_n5495__ = new_new_n2596__ & ~new_new_n5037__;
  assign new_new_n5496__ = ~new_new_n301__ & ~new_new_n5495__;
  assign new_new_n5497__ = ~new_new_n318__ & new_new_n5143__;
  assign new_new_n5498__ = new_new_n5032__ & new_new_n5497__;
  assign new_new_n5499__ = ~new_new_n5496__ & ~new_new_n5498__;
  assign new_new_n5500__ = new_new_n5494__ & ~new_new_n5499__;
  assign new_new_n5501__ = new_new_n2596__ & new_new_n4421__;
  assign new_new_n5502__ = new_new_n4444__ & new_new_n5501__;
  assign new_new_n5503__ = new_new_n5494__ & ~new_new_n5502__;
  assign new_new_n5504__ = new_new_n301__ & ~new_new_n5503__;
  assign new_new_n5505__ = ~new_new_n5491__ & ~new_new_n5504__;
  assign new_new_n5506__ = ~new_new_n5500__ & new_new_n5505__;
  assign new_new_n5507__ = new_new_n5489__ & new_new_n5506__;
  assign new_new_n5508__ = ~new_new_n5489__ & ~new_new_n5506__;
  assign new_new_n5509__ = ~new_new_n5507__ & ~new_new_n5508__;
  assign new_new_n5510__ = new_new_n2848__ & new_new_n3596__;
  assign new_new_n5511__ = ~new_new_n3203__ & new_new_n4132__;
  assign new_new_n5512__ = new_new_n3069__ & ~new_new_n3486__;
  assign new_new_n5513__ = ~new_new_n2848__ & ~new_new_n5511__;
  assign new_new_n5514__ = ~new_new_n5512__ & new_new_n5513__;
  assign new_new_n5515__ = ~new_new_n5510__ & ~new_new_n5514__;
  assign new_new_n5516__ = new_new_n437__ & ~new_new_n5515__;
  assign new_new_n5517__ = new_new_n651__ & new_new_n3586__;
  assign new_new_n5518__ = ~new_new_n651__ & ~new_new_n3586__;
  assign new_new_n5519__ = new_new_n2848__ & new_new_n3515__;
  assign new_new_n5520__ = ~new_new_n5517__ & ~new_new_n5518__;
  assign new_new_n5521__ = new_new_n5519__ & new_new_n5520__;
  assign new_new_n5522__ = new_new_n2848__ & ~new_new_n3587__;
  assign new_new_n5523__ = ~new_new_n437__ & ~new_new_n5514__;
  assign new_new_n5524__ = ~new_new_n5522__ & new_new_n5523__;
  assign new_new_n5525__ = ~new_new_n5521__ & ~new_new_n5524__;
  assign new_new_n5526__ = ~new_new_n5516__ & new_new_n5525__;
  assign new_new_n5527__ = new_new_n2809__ & ~new_new_n3733__;
  assign new_new_n5528__ = ~new_new_n2806__ & new_new_n3651__;
  assign new_new_n5529__ = ~new_new_n5527__ & ~new_new_n5528__;
  assign new_new_n5530__ = new_new_n2808__ & new_new_n4315__;
  assign new_new_n5531__ = new_new_n5529__ & ~new_new_n5530__;
  assign new_new_n5532__ = new_new_n810__ & ~new_new_n5531__;
  assign new_new_n5533__ = new_new_n2808__ & ~new_new_n4325__;
  assign new_new_n5534__ = ~new_new_n810__ & ~new_new_n5533__;
  assign new_new_n5535__ = ~new_new_n816__ & ~new_new_n4319__;
  assign new_new_n5536__ = new_new_n816__ & ~new_new_n4321__;
  assign new_new_n5537__ = new_new_n2808__ & ~new_new_n5535__;
  assign new_new_n5538__ = ~new_new_n5536__ & new_new_n5537__;
  assign new_new_n5539__ = ~new_new_n5534__ & ~new_new_n5538__;
  assign new_new_n5540__ = new_new_n5529__ & ~new_new_n5539__;
  assign new_new_n5541__ = ~new_new_n5532__ & ~new_new_n5540__;
  assign new_new_n5542__ = ~new_new_n437__ & ~new_new_n2784__;
  assign new_new_n5543__ = new_new_n5409__ & ~new_new_n5542__;
  assign new_new_n5544__ = ~new_new_n3821__ & ~new_new_n5409__;
  assign new_new_n5545__ = ~new_new_n2585__ & ~new_new_n5543__;
  assign new_new_n5546__ = ~new_new_n5544__ & new_new_n5545__;
  assign new_new_n5547__ = new_new_n437__ & ~new_new_n3233__;
  assign new_new_n5548__ = ~new_new_n5409__ & new_new_n5547__;
  assign new_new_n5549__ = new_new_n3233__ & new_new_n5409__;
  assign new_new_n5550__ = new_new_n2784__ & ~new_new_n5549__;
  assign new_new_n5551__ = new_new_n2585__ & ~new_new_n3820__;
  assign new_new_n5552__ = new_new_n5412__ & ~new_new_n5551__;
  assign new_new_n5553__ = ~new_new_n437__ & ~new_new_n5550__;
  assign new_new_n5554__ = ~new_new_n5552__ & new_new_n5553__;
  assign new_new_n5555__ = ~new_new_n5546__ & ~new_new_n5548__;
  assign new_new_n5556__ = ~new_new_n5554__ & new_new_n5555__;
  assign new_new_n5557__ = new_new_n5541__ & ~new_new_n5556__;
  assign new_new_n5558__ = ~new_new_n5541__ & new_new_n5556__;
  assign new_new_n5559__ = ~new_new_n5557__ & ~new_new_n5558__;
  assign new_new_n5560__ = ~new_new_n5526__ & new_new_n5559__;
  assign new_new_n5561__ = new_new_n5526__ & ~new_new_n5559__;
  assign new_new_n5562__ = ~new_new_n5560__ & ~new_new_n5561__;
  assign new_new_n5563__ = new_new_n5509__ & ~new_new_n5562__;
  assign new_new_n5564__ = ~new_new_n5509__ & new_new_n5562__;
  assign new_new_n5565__ = ~new_new_n5563__ & ~new_new_n5564__;
  assign new_new_n5566__ = new_new_n5479__ & ~new_new_n5565__;
  assign new_new_n5567__ = ~new_new_n5479__ & new_new_n5565__;
  assign new_new_n5568__ = ~new_new_n5566__ & ~new_new_n5567__;
  assign new_new_n5569__ = ~new_new_n5370__ & ~new_new_n5418__;
  assign new_new_n5570__ = ~new_new_n5369__ & ~new_new_n5569__;
  assign new_new_n5571__ = new_new_n5568__ & ~new_new_n5570__;
  assign new_new_n5572__ = ~new_new_n5568__ & new_new_n5570__;
  assign new_new_n5573__ = ~new_new_n5571__ & ~new_new_n5572__;
  assign new_new_n5574__ = ~new_new_n5456__ & ~new_new_n5573__;
  assign new_new_n5575__ = ~new_new_n5469__ & new_new_n5574__;
  assign new_new_n5576__ = ~new_new_n5463__ & new_new_n5575__;
  assign new_new_n5577__ = ~new_new_n5467__ & new_new_n5576__;
  assign new_new_n5578__ = ~new_new_n5349__ & ~new_new_n5421__;
  assign new_new_n5579__ = ~new_new_n5348__ & ~new_new_n5578__;
  assign new_new_n5580__ = new_new_n5326__ & new_new_n5579__;
  assign new_new_n5581__ = new_new_n5349__ & new_new_n5421__;
  assign new_new_n5582__ = new_new_n5348__ & ~new_new_n5421__;
  assign new_new_n5583__ = ~new_new_n5581__ & ~new_new_n5582__;
  assign new_new_n5584__ = new_new_n5328__ & new_new_n5583__;
  assign new_new_n5585__ = new_new_n5327__ & ~new_new_n5579__;
  assign new_new_n5586__ = new_new_n5573__ & ~new_new_n5580__;
  assign new_new_n5587__ = ~new_new_n5585__ & new_new_n5586__;
  assign new_new_n5588__ = ~new_new_n5584__ & new_new_n5587__;
  assign new_new_n5589__ = ~new_new_n5577__ & ~new_new_n5588__;
  assign new_new_n5590__ = ~new_new_n244__ & new_new_n347__;
  assign new_new_n5591__ = new_new_n227__ & ~new_new_n4260__;
  assign new_new_n5592__ = ~new_new_n5590__ & ~new_new_n5591__;
  assign new_new_n5593__ = ~new_new_n335__ & ~new_new_n5592__;
  assign new_new_n5594__ = ~new_new_n457__ & new_new_n623__;
  assign new_new_n5595__ = ~new_new_n616__ & ~new_new_n5594__;
  assign new_new_n5596__ = ~new_new_n540__ & new_new_n864__;
  assign new_new_n5597__ = ~new_new_n2232__ & ~new_new_n2245__;
  assign new_new_n5598__ = new_new_n2569__ & new_new_n5597__;
  assign new_new_n5599__ = new_new_n4720__ & new_new_n5596__;
  assign new_new_n5600__ = new_new_n5593__ & ~new_new_n5595__;
  assign new_new_n5601__ = new_new_n5599__ & new_new_n5600__;
  assign new_new_n5602__ = new_new_n5598__ & new_new_n5601__;
  assign new_new_n5603__ = new_new_n4845__ & new_new_n5602__;
  assign new_new_n5604__ = new_new_n3711__ & new_new_n5603__;
  assign new_new_n5605__ = new_new_n5589__ & ~new_new_n5604__;
  assign new_new_n5606__ = ~new_new_n5589__ & new_new_n5604__;
  assign new_new_n5607__ = ~new_new_n5605__ & ~new_new_n5606__;
  assign new_new_n5608__ = ~new_new_n5427__ & ~new_new_n5445__;
  assign new_new_n5609__ = new_new_n5607__ & new_new_n5608__;
  assign new_new_n5610__ = new_new_n5303__ & ~new_new_n5448__;
  assign new_new_n5611__ = ~new_new_n4702__ & ~new_new_n5610__;
  assign new_new_n5612__ = new_new_n5445__ & ~new_new_n5607__;
  assign new_new_n5613__ = ~new_new_n5611__ & new_new_n5612__;
  assign new_new_n5614__ = ~new_new_n5609__ & ~new_new_n5613__;
  assign new_new_n5615__ = new_new_n5308__ & ~new_new_n5614__;
  assign new_new_n5616__ = new_new_n5607__ & ~new_new_n5611__;
  assign new_new_n5617__ = ~new_new_n5308__ & ~new_new_n5611__;
  assign new_new_n5618__ = ~new_new_n5607__ & ~new_new_n5617__;
  assign new_new_n5619__ = new_new_n5427__ & new_new_n5445__;
  assign new_new_n5620__ = ~new_new_n5616__ & ~new_new_n5619__;
  assign new_new_n5621__ = ~new_new_n5618__ & new_new_n5620__;
  assign new_new_n5622__ = ~new_new_n5615__ & ~new_new_n5621__;
  assign new_new_n5623__ = ~new_new_n5440__ & ~new_new_n5622__;
  assign new_new_n5624__ = new_new_n5442__ & new_new_n5607__;
  assign new_new_n5625__ = new_new_n5308__ & ~new_new_n5427__;
  assign new_new_n5626__ = ~new_new_n5607__ & new_new_n5625__;
  assign new_new_n5627__ = ~new_new_n5624__ & ~new_new_n5626__;
  assign new_new_n5628__ = new_new_n5445__ & ~new_new_n5627__;
  assign new_new_n5629__ = ~new_new_n5607__ & ~new_new_n5608__;
  assign new_new_n5630__ = ~new_new_n5442__ & new_new_n5607__;
  assign new_new_n5631__ = ~new_new_n5308__ & ~new_new_n5629__;
  assign new_new_n5632__ = ~new_new_n5630__ & new_new_n5631__;
  assign new_new_n5633__ = ~new_new_n5628__ & ~new_new_n5632__;
  assign new_new_n5634__ = ~new_new_n5611__ & ~new_new_n5633__;
  assign new_new_n5635__ = new_new_n5442__ & ~new_new_n5607__;
  assign new_new_n5636__ = ~new_new_n5609__ & ~new_new_n5635__;
  assign new_new_n5637__ = new_new_n5611__ & ~new_new_n5636__;
  assign new_new_n5638__ = new_new_n5308__ & ~new_new_n5611__;
  assign new_new_n5639__ = ~new_new_n5445__ & ~new_new_n5638__;
  assign new_new_n5640__ = new_new_n5607__ & ~new_new_n5617__;
  assign new_new_n5641__ = ~new_new_n5441__ & ~new_new_n5613__;
  assign new_new_n5642__ = ~new_new_n5639__ & new_new_n5641__;
  assign new_new_n5643__ = ~new_new_n5640__ & new_new_n5642__;
  assign new_new_n5644__ = ~new_new_n5634__ & ~new_new_n5637__;
  assign new_new_n5645__ = ~new_new_n5643__ & new_new_n5644__;
  assign po05 = new_new_n5623__ | ~new_new_n5645__;
  assign new_new_n5647__ = new_new_n5468__ & ~new_new_n5573__;
  assign new_new_n5648__ = ~new_new_n5457__ & new_new_n5573__;
  assign new_new_n5649__ = ~new_new_n5454__ & ~new_new_n5573__;
  assign new_new_n5650__ = ~new_new_n5421__ & ~new_new_n5649__;
  assign new_new_n5651__ = ~new_new_n5648__ & ~new_new_n5650__;
  assign new_new_n5652__ = ~new_new_n5455__ & new_new_n5651__;
  assign new_new_n5653__ = ~new_new_n5421__ & ~new_new_n5457__;
  assign new_new_n5654__ = ~new_new_n5468__ & new_new_n5573__;
  assign new_new_n5655__ = ~new_new_n5454__ & ~new_new_n5653__;
  assign new_new_n5656__ = ~new_new_n5654__ & new_new_n5655__;
  assign new_new_n5657__ = ~new_new_n5647__ & ~new_new_n5652__;
  assign new_new_n5658__ = ~new_new_n5656__ & new_new_n5657__;
  assign new_new_n5659__ = ~new_new_n5567__ & ~new_new_n5570__;
  assign new_new_n5660__ = ~new_new_n5566__ & ~new_new_n5659__;
  assign new_new_n5661__ = new_new_n5658__ & ~new_new_n5660__;
  assign new_new_n5662__ = ~new_new_n5658__ & new_new_n5660__;
  assign new_new_n5663__ = ~new_new_n5661__ & ~new_new_n5662__;
  assign new_new_n5664__ = ~new_new_n5507__ & ~new_new_n5562__;
  assign new_new_n5665__ = ~new_new_n5508__ & ~new_new_n5664__;
  assign new_new_n5666__ = ~new_new_n320__ & new_new_n4421__;
  assign new_new_n5667__ = new_new_n2593__ & new_new_n4222__;
  assign new_new_n5668__ = ~new_new_n5666__ & ~new_new_n5667__;
  assign new_new_n5669__ = new_new_n2596__ & new_new_n5226__;
  assign new_new_n5670__ = new_new_n5668__ & ~new_new_n5669__;
  assign new_new_n5671__ = new_new_n301__ & ~new_new_n5670__;
  assign new_new_n5672__ = new_new_n2596__ & ~new_new_n5219__;
  assign new_new_n5673__ = ~new_new_n301__ & new_new_n5668__;
  assign new_new_n5674__ = ~new_new_n5672__ & new_new_n5673__;
  assign new_new_n5675__ = new_new_n316__ & ~new_new_n5222__;
  assign new_new_n5676__ = ~new_new_n316__ & ~new_new_n5214__;
  assign new_new_n5677__ = new_new_n2596__ & ~new_new_n5675__;
  assign new_new_n5678__ = ~new_new_n5676__ & new_new_n5677__;
  assign new_new_n5679__ = ~new_new_n5671__ & ~new_new_n5674__;
  assign new_new_n5680__ = ~new_new_n5678__ & new_new_n5679__;
  assign new_new_n5681__ = new_new_n5526__ & ~new_new_n5558__;
  assign new_new_n5682__ = ~new_new_n5557__ & ~new_new_n5681__;
  assign new_new_n5683__ = new_new_n5680__ & new_new_n5682__;
  assign new_new_n5684__ = ~new_new_n5680__ & ~new_new_n5682__;
  assign new_new_n5685__ = ~new_new_n5683__ & ~new_new_n5684__;
  assign new_new_n5686__ = new_new_n2784__ & ~new_new_n5409__;
  assign new_new_n5687__ = ~new_new_n2585__ & ~new_new_n5686__;
  assign new_new_n5688__ = new_new_n5552__ & ~new_new_n5687__;
  assign new_new_n5689__ = ~new_new_n437__ & ~new_new_n3203__;
  assign new_new_n5690__ = ~new_new_n5688__ & new_new_n5689__;
  assign new_new_n5691__ = ~new_new_n2585__ & new_new_n3821__;
  assign new_new_n5692__ = ~new_new_n5409__ & new_new_n5691__;
  assign new_new_n5693__ = new_new_n3820__ & new_new_n5389__;
  assign new_new_n5694__ = new_new_n5409__ & new_new_n5693__;
  assign new_new_n5695__ = ~new_new_n5692__ & ~new_new_n5694__;
  assign new_new_n5696__ = new_new_n3203__ & ~new_new_n5695__;
  assign new_new_n5697__ = ~new_new_n5548__ & ~new_new_n5696__;
  assign new_new_n5698__ = ~new_new_n5690__ & new_new_n5697__;
  assign new_new_n5699__ = new_new_n2809__ & ~new_new_n3727__;
  assign new_new_n5700__ = ~new_new_n2806__ & ~new_new_n3733__;
  assign new_new_n5701__ = ~new_new_n5699__ & ~new_new_n5700__;
  assign new_new_n5702__ = new_new_n2808__ & new_new_n4081__;
  assign new_new_n5703__ = ~new_new_n4086__ & new_new_n5702__;
  assign new_new_n5704__ = new_new_n5701__ & ~new_new_n5703__;
  assign new_new_n5705__ = ~new_new_n810__ & ~new_new_n5704__;
  assign new_new_n5706__ = ~new_new_n816__ & ~new_new_n4081__;
  assign new_new_n5707__ = new_new_n816__ & new_new_n4081__;
  assign new_new_n5708__ = ~new_new_n5706__ & ~new_new_n5707__;
  assign new_new_n5709__ = new_new_n2808__ & new_new_n4086__;
  assign new_new_n5710__ = ~new_new_n5708__ & new_new_n5709__;
  assign new_new_n5711__ = ~new_new_n4081__ & ~new_new_n4086__;
  assign new_new_n5712__ = new_new_n2808__ & ~new_new_n5711__;
  assign new_new_n5713__ = new_new_n810__ & new_new_n5701__;
  assign new_new_n5714__ = ~new_new_n5712__ & new_new_n5713__;
  assign new_new_n5715__ = ~new_new_n5705__ & ~new_new_n5710__;
  assign new_new_n5716__ = ~new_new_n5714__ & new_new_n5715__;
  assign new_new_n5717__ = ~new_new_n437__ & new_new_n3486__;
  assign new_new_n5718__ = new_new_n4787__ & ~new_new_n5717__;
  assign new_new_n5719__ = ~new_new_n437__ & ~new_new_n3651__;
  assign new_new_n5720__ = new_new_n437__ & new_new_n3651__;
  assign new_new_n5721__ = ~new_new_n5719__ & ~new_new_n5720__;
  assign new_new_n5722__ = ~new_new_n3654__ & ~new_new_n5721__;
  assign new_new_n5723__ = ~new_new_n651__ & ~new_new_n3651__;
  assign new_new_n5724__ = new_new_n651__ & new_new_n3651__;
  assign new_new_n5725__ = new_new_n3654__ & ~new_new_n5723__;
  assign new_new_n5726__ = ~new_new_n5724__ & new_new_n5725__;
  assign new_new_n5727__ = new_new_n2848__ & ~new_new_n5722__;
  assign new_new_n5728__ = ~new_new_n5726__ & new_new_n5727__;
  assign new_new_n5729__ = new_new_n2847__ & new_new_n5400__;
  assign new_new_n5730__ = ~new_new_n2848__ & ~new_new_n3068__;
  assign new_new_n5731__ = new_new_n3586__ & new_new_n5730__;
  assign new_new_n5732__ = ~new_new_n5729__ & ~new_new_n5731__;
  assign new_new_n5733__ = new_new_n437__ & ~new_new_n5732__;
  assign new_new_n5734__ = ~new_new_n437__ & ~new_new_n3586__;
  assign new_new_n5735__ = new_new_n3070__ & new_new_n5734__;
  assign new_new_n5736__ = ~new_new_n5718__ & ~new_new_n5735__;
  assign new_new_n5737__ = ~new_new_n5733__ & new_new_n5736__;
  assign new_new_n5738__ = ~new_new_n5728__ & new_new_n5737__;
  assign new_new_n5739__ = ~new_new_n5716__ & new_new_n5738__;
  assign new_new_n5740__ = new_new_n5716__ & ~new_new_n5738__;
  assign new_new_n5741__ = new_new_n5698__ & ~new_new_n5739__;
  assign new_new_n5742__ = ~new_new_n5740__ & ~new_new_n5741__;
  assign new_new_n5743__ = ~new_new_n5739__ & new_new_n5742__;
  assign new_new_n5744__ = ~new_new_n5698__ & ~new_new_n5743__;
  assign new_new_n5745__ = ~new_new_n5740__ & new_new_n5741__;
  assign new_new_n5746__ = ~new_new_n5744__ & ~new_new_n5745__;
  assign new_new_n5747__ = new_new_n5685__ & ~new_new_n5746__;
  assign new_new_n5748__ = ~new_new_n5685__ & new_new_n5746__;
  assign new_new_n5749__ = ~new_new_n5747__ & ~new_new_n5748__;
  assign new_new_n5750__ = ~new_new_n5665__ & new_new_n5749__;
  assign new_new_n5751__ = new_new_n5665__ & ~new_new_n5749__;
  assign new_new_n5752__ = ~new_new_n5750__ & ~new_new_n5751__;
  assign new_new_n5753__ = ~new_new_n310__ & ~new_new_n5342__;
  assign new_new_n5754__ = ~new_new_n3235__ & ~new_new_n3306__;
  assign new_new_n5755__ = ~new_new_n4857__ & new_new_n5754__;
  assign new_new_n5756__ = ~new_new_n5753__ & ~new_new_n5755__;
  assign new_new_n5757__ = ~new_new_n310__ & new_new_n5122__;
  assign new_new_n5758__ = ~new_new_n5122__ & ~new_new_n5342__;
  assign new_new_n5759__ = ~new_new_n3234__ & ~new_new_n5757__;
  assign new_new_n5760__ = ~new_new_n5758__ & new_new_n5759__;
  assign new_new_n5761__ = ~new_new_n5756__ & ~new_new_n5760__;
  assign new_new_n5762__ = new_new_n5752__ & ~new_new_n5761__;
  assign new_new_n5763__ = ~new_new_n5752__ & new_new_n5761__;
  assign new_new_n5764__ = ~new_new_n5762__ & ~new_new_n5763__;
  assign new_new_n5765__ = new_new_n5663__ & new_new_n5764__;
  assign new_new_n5766__ = ~new_new_n5663__ & ~new_new_n5764__;
  assign new_new_n5767__ = ~new_new_n5765__ & ~new_new_n5766__;
  assign new_new_n5768__ = ~new_new_n5440__ & ~new_new_n5619__;
  assign new_new_n5769__ = new_new_n5607__ & ~new_new_n5608__;
  assign new_new_n5770__ = ~new_new_n5768__ & new_new_n5769__;
  assign new_new_n5771__ = ~new_new_n5606__ & ~new_new_n5770__;
  assign new_new_n5772__ = ~new_new_n5767__ & ~new_new_n5771__;
  assign new_new_n5773__ = new_new_n5767__ & new_new_n5771__;
  assign new_new_n5774__ = ~new_new_n5772__ & ~new_new_n5773__;
  assign new_new_n5775__ = new_new_n125__ & ~new_new_n2446__;
  assign new_new_n5776__ = ~new_new_n87__ & ~new_new_n1107__;
  assign new_new_n5777__ = new_new_n238__ & ~new_new_n5776__;
  assign new_new_n5778__ = ~new_new_n524__ & ~new_new_n5777__;
  assign new_new_n5779__ = ~new_new_n274__ & ~new_new_n662__;
  assign new_new_n5780__ = ~new_new_n5775__ & new_new_n5779__;
  assign new_new_n5781__ = ~new_new_n523__ & ~new_new_n2245__;
  assign new_new_n5782__ = new_new_n4847__ & ~new_new_n5778__;
  assign new_new_n5783__ = new_new_n5781__ & new_new_n5782__;
  assign new_new_n5784__ = new_new_n2458__ & new_new_n5780__;
  assign new_new_n5785__ = new_new_n5783__ & new_new_n5784__;
  assign new_new_n5786__ = new_new_n116__ & ~new_new_n658__;
  assign new_new_n5787__ = new_new_n160__ & new_new_n371__;
  assign new_new_n5788__ = new_new_n195__ & ~new_new_n5787__;
  assign new_new_n5789__ = ~new_new_n137__ & ~new_new_n5786__;
  assign new_new_n5790__ = ~new_new_n322__ & ~new_new_n377__;
  assign new_new_n5791__ = ~new_new_n4207__ & new_new_n5790__;
  assign new_new_n5792__ = ~new_new_n5788__ & new_new_n5789__;
  assign new_new_n5793__ = new_new_n5791__ & new_new_n5792__;
  assign new_new_n5794__ = new_new_n2328__ & new_new_n5793__;
  assign new_new_n5795__ = new_new_n5785__ & new_new_n5794__;
  assign new_new_n5796__ = new_new_n4485__ & new_new_n5795__;
  assign new_new_n5797__ = ~new_new_n5774__ & new_new_n5796__;
  assign new_new_n5798__ = new_new_n5774__ & ~new_new_n5796__;
  assign new_new_n5799__ = ~new_new_n5797__ & ~new_new_n5798__;
  assign new_new_n5800__ = new_new_n5441__ & new_new_n5607__;
  assign new_new_n5801__ = ~new_new_n5635__ & ~new_new_n5800__;
  assign new_new_n5802__ = new_new_n5445__ & ~new_new_n5801__;
  assign new_new_n5803__ = new_new_n5446__ & new_new_n5607__;
  assign new_new_n5804__ = ~new_new_n5802__ & ~new_new_n5803__;
  assign new_new_n5805__ = new_new_n5303__ & ~new_new_n5804__;
  assign new_new_n5806__ = ~new_new_n5441__ & ~new_new_n5607__;
  assign new_new_n5807__ = new_new_n5308__ & ~new_new_n5445__;
  assign new_new_n5808__ = ~new_new_n5630__ & new_new_n5807__;
  assign new_new_n5809__ = ~new_new_n5806__ & new_new_n5808__;
  assign new_new_n5810__ = ~new_new_n5805__ & ~new_new_n5809__;
  assign new_new_n5811__ = new_new_n5308__ & new_new_n5448__;
  assign new_new_n5812__ = ~new_new_n5609__ & new_new_n5811__;
  assign new_new_n5813__ = ~new_new_n5629__ & new_new_n5812__;
  assign new_new_n5814__ = ~new_new_n5810__ & ~new_new_n5813__;
  assign new_new_n5815__ = new_new_n4702__ & ~new_new_n5813__;
  assign new_new_n5816__ = ~new_new_n5814__ & ~new_new_n5815__;
  assign new_new_n5817__ = ~new_new_n5799__ & ~new_new_n5816__;
  assign new_new_n5818__ = new_new_n5799__ & new_new_n5816__;
  assign po06 = ~new_new_n5817__ & ~new_new_n5818__;
  assign new_new_n5820__ = ~new_new_n5662__ & ~new_new_n5749__;
  assign new_new_n5821__ = ~new_new_n5661__ & ~new_new_n5820__;
  assign new_new_n5822__ = new_new_n5665__ & ~new_new_n5821__;
  assign new_new_n5823__ = new_new_n5661__ & ~new_new_n5749__;
  assign new_new_n5824__ = ~new_new_n5822__ & ~new_new_n5823__;
  assign new_new_n5825__ = new_new_n5761__ & ~new_new_n5824__;
  assign new_new_n5826__ = ~new_new_n5665__ & new_new_n5821__;
  assign new_new_n5827__ = new_new_n5662__ & new_new_n5749__;
  assign new_new_n5828__ = ~new_new_n5826__ & ~new_new_n5827__;
  assign new_new_n5829__ = ~new_new_n5761__ & ~new_new_n5828__;
  assign new_new_n5830__ = new_new_n5658__ & ~new_new_n5749__;
  assign new_new_n5831__ = new_new_n5660__ & ~new_new_n5665__;
  assign new_new_n5832__ = ~new_new_n5830__ & ~new_new_n5831__;
  assign new_new_n5833__ = ~new_new_n5660__ & new_new_n5665__;
  assign new_new_n5834__ = ~new_new_n5658__ & new_new_n5749__;
  assign new_new_n5835__ = ~new_new_n5833__ & ~new_new_n5834__;
  assign new_new_n5836__ = ~new_new_n5832__ & ~new_new_n5835__;
  assign new_new_n5837__ = ~new_new_n5683__ & ~new_new_n5746__;
  assign new_new_n5838__ = ~new_new_n5684__ & ~new_new_n5837__;
  assign new_new_n5839__ = new_new_n2593__ & new_new_n4421__;
  assign new_new_n5840__ = ~new_new_n320__ & ~new_new_n4532__;
  assign new_new_n5841__ = ~new_new_n5839__ & ~new_new_n5840__;
  assign new_new_n5842__ = new_new_n2596__ & ~new_new_n4857__;
  assign new_new_n5843__ = new_new_n4884__ & new_new_n5842__;
  assign new_new_n5844__ = new_new_n5841__ & ~new_new_n5843__;
  assign new_new_n5845__ = ~new_new_n301__ & ~new_new_n5844__;
  assign new_new_n5846__ = new_new_n2596__ & ~new_new_n5338__;
  assign new_new_n5847__ = new_new_n301__ & new_new_n5841__;
  assign new_new_n5848__ = ~new_new_n5846__ & new_new_n5847__;
  assign new_new_n5849__ = ~new_new_n316__ & ~new_new_n4857__;
  assign new_new_n5850__ = new_new_n316__ & new_new_n4884__;
  assign new_new_n5851__ = ~new_new_n5849__ & ~new_new_n5850__;
  assign new_new_n5852__ = new_new_n5846__ & new_new_n5851__;
  assign new_new_n5853__ = ~new_new_n5845__ & ~new_new_n5848__;
  assign new_new_n5854__ = ~new_new_n5852__ & new_new_n5853__;
  assign new_new_n5855__ = new_new_n5838__ & ~new_new_n5854__;
  assign new_new_n5856__ = ~new_new_n5838__ & new_new_n5854__;
  assign new_new_n5857__ = ~new_new_n5855__ & ~new_new_n5856__;
  assign new_new_n5858__ = new_new_n2809__ & new_new_n4081__;
  assign new_new_n5859__ = ~new_new_n2806__ & ~new_new_n3727__;
  assign new_new_n5860__ = ~new_new_n5858__ & ~new_new_n5859__;
  assign new_new_n5861__ = new_new_n2808__ & ~new_new_n4744__;
  assign new_new_n5862__ = ~new_new_n810__ & ~new_new_n5861__;
  assign new_new_n5863__ = new_new_n2808__ & new_new_n4233__;
  assign new_new_n5864__ = ~new_new_n816__ & new_new_n4222__;
  assign new_new_n5865__ = new_new_n5863__ & new_new_n5864__;
  assign new_new_n5866__ = ~new_new_n5862__ & ~new_new_n5865__;
  assign new_new_n5867__ = new_new_n5860__ & ~new_new_n5866__;
  assign new_new_n5868__ = new_new_n2808__ & new_new_n4222__;
  assign new_new_n5869__ = ~new_new_n4233__ & new_new_n5868__;
  assign new_new_n5870__ = new_new_n5860__ & ~new_new_n5869__;
  assign new_new_n5871__ = new_new_n810__ & ~new_new_n5870__;
  assign new_new_n5872__ = new_new_n816__ & ~new_new_n4222__;
  assign new_new_n5873__ = new_new_n5863__ & new_new_n5872__;
  assign new_new_n5874__ = ~new_new_n5871__ & ~new_new_n5873__;
  assign new_new_n5875__ = ~new_new_n5867__ & new_new_n5874__;
  assign new_new_n5876__ = new_new_n5742__ & new_new_n5875__;
  assign new_new_n5877__ = ~new_new_n5742__ & ~new_new_n5875__;
  assign new_new_n5878__ = ~new_new_n5876__ & ~new_new_n5877__;
  assign new_new_n5879__ = ~new_new_n2585__ & new_new_n2784__;
  assign new_new_n5880__ = new_new_n3203__ & new_new_n5879__;
  assign new_new_n5881__ = ~new_new_n3233__ & ~new_new_n5880__;
  assign new_new_n5882__ = new_new_n2585__ & ~new_new_n2784__;
  assign new_new_n5883__ = ~new_new_n3203__ & new_new_n5882__;
  assign new_new_n5884__ = new_new_n5409__ & new_new_n5883__;
  assign new_new_n5885__ = ~new_new_n5881__ & ~new_new_n5884__;
  assign new_new_n5886__ = ~new_new_n437__ & ~new_new_n5885__;
  assign new_new_n5887__ = ~new_new_n5410__ & ~new_new_n5886__;
  assign new_new_n5888__ = ~new_new_n437__ & ~new_new_n3486__;
  assign new_new_n5889__ = ~new_new_n3065__ & ~new_new_n3586__;
  assign new_new_n5890__ = new_new_n3070__ & new_new_n3651__;
  assign new_new_n5891__ = ~new_new_n3072__ & new_new_n4024__;
  assign new_new_n5892__ = new_new_n3733__ & ~new_new_n5891__;
  assign new_new_n5893__ = ~new_new_n3733__ & new_new_n5891__;
  assign new_new_n5894__ = new_new_n2848__ & ~new_new_n5892__;
  assign new_new_n5895__ = ~new_new_n5893__ & new_new_n5894__;
  assign new_new_n5896__ = ~new_new_n5889__ & ~new_new_n5890__;
  assign new_new_n5897__ = ~new_new_n5895__ & new_new_n5896__;
  assign new_new_n5898__ = ~new_new_n5888__ & new_new_n5897__;
  assign new_new_n5899__ = new_new_n310__ & new_new_n3233__;
  assign new_new_n5900__ = ~new_new_n5898__ & new_new_n5899__;
  assign new_new_n5901__ = new_new_n3233__ & ~new_new_n3486__;
  assign new_new_n5902__ = ~new_new_n3233__ & new_new_n5717__;
  assign new_new_n5903__ = ~new_new_n310__ & new_new_n5897__;
  assign new_new_n5904__ = ~new_new_n5901__ & ~new_new_n5902__;
  assign new_new_n5905__ = new_new_n5903__ & new_new_n5904__;
  assign new_new_n5906__ = ~new_new_n5900__ & ~new_new_n5905__;
  assign new_new_n5907__ = ~new_new_n5887__ & ~new_new_n5906__;
  assign new_new_n5908__ = ~new_new_n3233__ & new_new_n5887__;
  assign new_new_n5909__ = ~new_new_n5717__ & ~new_new_n5908__;
  assign new_new_n5910__ = new_new_n310__ & ~new_new_n5897__;
  assign new_new_n5911__ = new_new_n5887__ & new_new_n5903__;
  assign new_new_n5912__ = ~new_new_n5910__ & ~new_new_n5911__;
  assign new_new_n5913__ = new_new_n5909__ & ~new_new_n5912__;
  assign new_new_n5914__ = new_new_n3233__ & new_new_n5886__;
  assign new_new_n5915__ = ~new_new_n5903__ & ~new_new_n5914__;
  assign new_new_n5916__ = ~new_new_n5909__ & ~new_new_n5910__;
  assign new_new_n5917__ = new_new_n5915__ & new_new_n5916__;
  assign new_new_n5918__ = ~new_new_n5907__ & ~new_new_n5917__;
  assign new_new_n5919__ = ~new_new_n5913__ & new_new_n5918__;
  assign new_new_n5920__ = ~new_new_n5878__ & new_new_n5919__;
  assign new_new_n5921__ = new_new_n5878__ & ~new_new_n5919__;
  assign new_new_n5922__ = ~new_new_n5920__ & ~new_new_n5921__;
  assign new_new_n5923__ = new_new_n5857__ & ~new_new_n5922__;
  assign new_new_n5924__ = ~new_new_n5857__ & new_new_n5922__;
  assign new_new_n5925__ = ~new_new_n5923__ & ~new_new_n5924__;
  assign new_new_n5926__ = ~new_new_n5836__ & new_new_n5925__;
  assign new_new_n5927__ = ~new_new_n5825__ & new_new_n5926__;
  assign new_new_n5928__ = ~new_new_n5829__ & new_new_n5927__;
  assign new_new_n5929__ = new_new_n5751__ & new_new_n5761__;
  assign new_new_n5930__ = new_new_n5750__ & ~new_new_n5761__;
  assign new_new_n5931__ = ~new_new_n5929__ & ~new_new_n5930__;
  assign new_new_n5932__ = new_new_n5663__ & new_new_n5931__;
  assign new_new_n5933__ = ~new_new_n5750__ & new_new_n5761__;
  assign new_new_n5934__ = ~new_new_n5751__ & ~new_new_n5933__;
  assign new_new_n5935__ = new_new_n5662__ & ~new_new_n5934__;
  assign new_new_n5936__ = new_new_n5661__ & new_new_n5934__;
  assign new_new_n5937__ = ~new_new_n5925__ & ~new_new_n5935__;
  assign new_new_n5938__ = ~new_new_n5936__ & new_new_n5937__;
  assign new_new_n5939__ = ~new_new_n5932__ & new_new_n5938__;
  assign new_new_n5940__ = ~new_new_n5928__ & ~new_new_n5939__;
  assign new_new_n5941__ = ~new_new_n125__ & ~new_new_n181__;
  assign new_new_n5942__ = new_new_n371__ & ~new_new_n571__;
  assign new_new_n5943__ = ~new_new_n5941__ & ~new_new_n5942__;
  assign new_new_n5944__ = ~new_new_n100__ & new_new_n5075__;
  assign new_new_n5945__ = new_new_n174__ & new_new_n1095__;
  assign new_new_n5946__ = ~new_new_n2230__ & new_new_n5945__;
  assign new_new_n5947__ = ~new_new_n2683__ & ~new_new_n5944__;
  assign new_new_n5948__ = ~new_new_n5946__ & new_new_n5947__;
  assign new_new_n5949__ = new_new_n279__ & ~new_new_n379__;
  assign new_new_n5950__ = ~new_new_n5943__ & new_new_n5949__;
  assign new_new_n5951__ = new_new_n5593__ & new_new_n5950__;
  assign new_new_n5952__ = ~new_new_n5948__ & new_new_n5951__;
  assign new_new_n5953__ = new_new_n5785__ & new_new_n5952__;
  assign new_new_n5954__ = new_new_n2699__ & new_new_n5953__;
  assign new_new_n5955__ = new_new_n5940__ & ~new_new_n5954__;
  assign new_new_n5956__ = ~new_new_n5940__ & new_new_n5954__;
  assign new_new_n5957__ = ~new_new_n5955__ & ~new_new_n5956__;
  assign new_new_n5958__ = ~new_new_n5772__ & ~new_new_n5796__;
  assign new_new_n5959__ = ~new_new_n5773__ & ~new_new_n5958__;
  assign new_new_n5960__ = new_new_n5957__ & ~new_new_n5959__;
  assign new_new_n5961__ = ~new_new_n5957__ & new_new_n5959__;
  assign new_new_n5962__ = ~new_new_n5960__ & ~new_new_n5961__;
  assign new_new_n5963__ = new_new_n5799__ & new_new_n5813__;
  assign new_new_n5964__ = new_new_n4702__ & ~new_new_n5963__;
  assign new_new_n5965__ = ~new_new_n5817__ & ~new_new_n5964__;
  assign new_new_n5966__ = new_new_n5962__ & ~new_new_n5965__;
  assign new_new_n5967__ = ~new_new_n5799__ & new_new_n5814__;
  assign new_new_n5968__ = ~new_new_n5962__ & ~new_new_n5967__;
  assign new_new_n5969__ = ~new_new_n5964__ & new_new_n5968__;
  assign po07 = new_new_n5966__ | new_new_n5969__;
  assign new_new_n5971__ = new_new_n5962__ & new_new_n5963__;
  assign new_new_n5972__ = ~new_new_n5962__ & new_new_n5967__;
  assign new_new_n5973__ = ~new_new_n4702__ & ~new_new_n5972__;
  assign new_new_n5974__ = ~new_new_n5971__ & ~new_new_n5973__;
  assign new_new_n5975__ = ~new_new_n5956__ & ~new_new_n5959__;
  assign new_new_n5976__ = ~new_new_n5955__ & ~new_new_n5975__;
  assign new_new_n5977__ = ~new_new_n5833__ & new_new_n5925__;
  assign new_new_n5978__ = new_new_n5761__ & ~new_new_n5834__;
  assign new_new_n5979__ = new_new_n5833__ & ~new_new_n5925__;
  assign new_new_n5980__ = ~new_new_n5830__ & ~new_new_n5979__;
  assign new_new_n5981__ = ~new_new_n5978__ & new_new_n5980__;
  assign new_new_n5982__ = ~new_new_n5977__ & ~new_new_n5981__;
  assign new_new_n5983__ = ~new_new_n5834__ & ~new_new_n5925__;
  assign new_new_n5984__ = ~new_new_n5761__ & ~new_new_n5983__;
  assign new_new_n5985__ = ~new_new_n5830__ & new_new_n5925__;
  assign new_new_n5986__ = ~new_new_n5831__ & ~new_new_n5985__;
  assign new_new_n5987__ = ~new_new_n5984__ & new_new_n5986__;
  assign new_new_n5988__ = ~new_new_n5982__ & ~new_new_n5987__;
  assign new_new_n5989__ = ~new_new_n5856__ & new_new_n5922__;
  assign new_new_n5990__ = ~new_new_n5855__ & ~new_new_n5989__;
  assign new_new_n5991__ = new_new_n5988__ & new_new_n5990__;
  assign new_new_n5992__ = ~new_new_n5988__ & ~new_new_n5990__;
  assign new_new_n5993__ = ~new_new_n5991__ & ~new_new_n5992__;
  assign new_new_n5994__ = ~new_new_n320__ & ~new_new_n4857__;
  assign new_new_n5995__ = new_new_n2593__ & ~new_new_n4532__;
  assign new_new_n5996__ = ~new_new_n5994__ & ~new_new_n5995__;
  assign new_new_n5997__ = ~new_new_n301__ & ~new_new_n5996__;
  assign new_new_n5998__ = new_new_n4923__ & new_new_n5490__;
  assign new_new_n5999__ = new_new_n2596__ & new_new_n4923__;
  assign new_new_n6000__ = new_new_n301__ & new_new_n5996__;
  assign new_new_n6001__ = ~new_new_n5999__ & new_new_n6000__;
  assign new_new_n6002__ = ~new_new_n5997__ & ~new_new_n5998__;
  assign new_new_n6003__ = ~new_new_n6001__ & new_new_n6002__;
  assign new_new_n6004__ = ~new_new_n2806__ & new_new_n4081__;
  assign new_new_n6005__ = new_new_n2809__ & new_new_n4222__;
  assign new_new_n6006__ = ~new_new_n6004__ & ~new_new_n6005__;
  assign new_new_n6007__ = new_new_n2808__ & new_new_n4421__;
  assign new_new_n6008__ = new_new_n4444__ & new_new_n6007__;
  assign new_new_n6009__ = new_new_n6006__ & ~new_new_n6008__;
  assign new_new_n6010__ = new_new_n810__ & ~new_new_n6009__;
  assign new_new_n6011__ = new_new_n2808__ & ~new_new_n5037__;
  assign new_new_n6012__ = ~new_new_n810__ & ~new_new_n6011__;
  assign new_new_n6013__ = new_new_n816__ & ~new_new_n5032__;
  assign new_new_n6014__ = ~new_new_n816__ & ~new_new_n5040__;
  assign new_new_n6015__ = new_new_n2808__ & ~new_new_n6013__;
  assign new_new_n6016__ = ~new_new_n6014__ & new_new_n6015__;
  assign new_new_n6017__ = ~new_new_n6012__ & ~new_new_n6016__;
  assign new_new_n6018__ = new_new_n6006__ & ~new_new_n6017__;
  assign new_new_n6019__ = ~new_new_n6010__ & ~new_new_n6018__;
  assign new_new_n6020__ = new_new_n3069__ & ~new_new_n3733__;
  assign new_new_n6021__ = new_new_n3651__ & new_new_n4132__;
  assign new_new_n6022__ = ~new_new_n6020__ & ~new_new_n6021__;
  assign new_new_n6023__ = ~new_new_n2848__ & ~new_new_n6022__;
  assign new_new_n6024__ = new_new_n2848__ & new_new_n4315__;
  assign new_new_n6025__ = ~new_new_n6023__ & ~new_new_n6024__;
  assign new_new_n6026__ = new_new_n437__ & ~new_new_n6025__;
  assign new_new_n6027__ = ~new_new_n651__ & ~new_new_n4319__;
  assign new_new_n6028__ = new_new_n651__ & ~new_new_n4321__;
  assign new_new_n6029__ = new_new_n2848__ & ~new_new_n6027__;
  assign new_new_n6030__ = ~new_new_n6028__ & new_new_n6029__;
  assign new_new_n6031__ = new_new_n2848__ & ~new_new_n4325__;
  assign new_new_n6032__ = ~new_new_n437__ & ~new_new_n6023__;
  assign new_new_n6033__ = ~new_new_n6031__ & new_new_n6032__;
  assign new_new_n6034__ = ~new_new_n6026__ & ~new_new_n6033__;
  assign new_new_n6035__ = ~new_new_n6030__ & new_new_n6034__;
  assign new_new_n6036__ = new_new_n3586__ & ~new_new_n6035__;
  assign new_new_n6037__ = new_new_n437__ & ~new_new_n6035__;
  assign new_new_n6038__ = ~new_new_n6036__ & ~new_new_n6037__;
  assign new_new_n6039__ = new_new_n3244__ & ~new_new_n6038__;
  assign new_new_n6040__ = ~new_new_n3586__ & new_new_n6035__;
  assign new_new_n6041__ = ~new_new_n6036__ & ~new_new_n6040__;
  assign new_new_n6042__ = new_new_n310__ & ~new_new_n3233__;
  assign new_new_n6043__ = ~new_new_n3486__ & ~new_new_n6042__;
  assign new_new_n6044__ = ~new_new_n6041__ & new_new_n6043__;
  assign new_new_n6045__ = new_new_n3244__ & new_new_n6040__;
  assign new_new_n6046__ = ~new_new_n6044__ & ~new_new_n6045__;
  assign new_new_n6047__ = ~new_new_n437__ & ~new_new_n6046__;
  assign new_new_n6048__ = ~new_new_n437__ & ~new_new_n6041__;
  assign new_new_n6049__ = ~new_new_n3244__ & ~new_new_n5888__;
  assign new_new_n6050__ = ~new_new_n6037__ & new_new_n6049__;
  assign new_new_n6051__ = ~new_new_n6048__ & new_new_n6050__;
  assign new_new_n6052__ = ~new_new_n6037__ & new_new_n6042__;
  assign new_new_n6053__ = new_new_n6041__ & new_new_n6052__;
  assign new_new_n6054__ = ~new_new_n6039__ & ~new_new_n6053__;
  assign new_new_n6055__ = ~new_new_n6051__ & new_new_n6054__;
  assign new_new_n6056__ = ~new_new_n6047__ & new_new_n6055__;
  assign new_new_n6057__ = ~new_new_n6019__ & new_new_n6056__;
  assign new_new_n6058__ = new_new_n6019__ & ~new_new_n6056__;
  assign new_new_n6059__ = ~new_new_n6057__ & ~new_new_n6058__;
  assign new_new_n6060__ = ~new_new_n5887__ & new_new_n5910__;
  assign new_new_n6061__ = ~new_new_n437__ & new_new_n3233__;
  assign new_new_n6062__ = new_new_n5903__ & new_new_n6061__;
  assign new_new_n6063__ = ~new_new_n6060__ & ~new_new_n6062__;
  assign new_new_n6064__ = ~new_new_n3486__ & ~new_new_n6063__;
  assign new_new_n6065__ = new_new_n437__ & ~new_new_n5897__;
  assign new_new_n6066__ = ~new_new_n5899__ & ~new_new_n5903__;
  assign new_new_n6067__ = ~new_new_n6065__ & new_new_n6066__;
  assign new_new_n6068__ = ~new_new_n5887__ & ~new_new_n6067__;
  assign new_new_n6069__ = new_new_n5899__ & new_new_n6065__;
  assign new_new_n6070__ = new_new_n310__ & ~new_new_n437__;
  assign new_new_n6071__ = new_new_n5897__ & new_new_n6070__;
  assign new_new_n6072__ = ~new_new_n310__ & ~new_new_n3233__;
  assign new_new_n6073__ = ~new_new_n5887__ & new_new_n6072__;
  assign new_new_n6074__ = ~new_new_n6071__ & ~new_new_n6073__;
  assign new_new_n6075__ = new_new_n3486__ & ~new_new_n6074__;
  assign new_new_n6076__ = ~new_new_n6065__ & ~new_new_n6070__;
  assign new_new_n6077__ = ~new_new_n3233__ & ~new_new_n5910__;
  assign new_new_n6078__ = ~new_new_n6076__ & new_new_n6077__;
  assign new_new_n6079__ = ~new_new_n6069__ & ~new_new_n6075__;
  assign new_new_n6080__ = ~new_new_n6078__ & new_new_n6079__;
  assign new_new_n6081__ = ~new_new_n6064__ & ~new_new_n6068__;
  assign new_new_n6082__ = new_new_n6080__ & new_new_n6081__;
  assign new_new_n6083__ = ~new_new_n6059__ & new_new_n6082__;
  assign new_new_n6084__ = new_new_n6059__ & ~new_new_n6082__;
  assign new_new_n6085__ = ~new_new_n6083__ & ~new_new_n6084__;
  assign new_new_n6086__ = ~new_new_n6003__ & ~new_new_n6085__;
  assign new_new_n6087__ = new_new_n6003__ & new_new_n6085__;
  assign new_new_n6088__ = ~new_new_n6086__ & ~new_new_n6087__;
  assign new_new_n6089__ = ~new_new_n5876__ & ~new_new_n5919__;
  assign new_new_n6090__ = ~new_new_n5877__ & ~new_new_n6089__;
  assign new_new_n6091__ = new_new_n6088__ & ~new_new_n6090__;
  assign new_new_n6092__ = ~new_new_n6088__ & new_new_n6090__;
  assign new_new_n6093__ = ~new_new_n6091__ & ~new_new_n6092__;
  assign new_new_n6094__ = new_new_n5993__ & new_new_n6093__;
  assign new_new_n6095__ = ~new_new_n5993__ & ~new_new_n6093__;
  assign new_new_n6096__ = ~new_new_n6094__ & ~new_new_n6095__;
  assign new_new_n6097__ = ~new_new_n5976__ & ~new_new_n6096__;
  assign new_new_n6098__ = new_new_n5976__ & new_new_n6096__;
  assign new_new_n6099__ = ~new_new_n6097__ & ~new_new_n6098__;
  assign new_new_n6100__ = new_new_n195__ & ~new_new_n1021__;
  assign new_new_n6101__ = new_new_n141__ & ~new_new_n956__;
  assign new_new_n6102__ = new_new_n87__ & ~new_new_n4268__;
  assign new_new_n6103__ = ~new_new_n6101__ & new_new_n6102__;
  assign new_new_n6104__ = new_new_n115__ & new_new_n1045__;
  assign new_new_n6105__ = new_new_n223__ & ~new_new_n6104__;
  assign new_new_n6106__ = new_new_n246__ & new_new_n677__;
  assign new_new_n6107__ = new_new_n244__ & ~new_new_n6106__;
  assign new_new_n6108__ = ~new_new_n348__ & ~new_new_n671__;
  assign new_new_n6109__ = ~new_new_n6105__ & new_new_n6108__;
  assign new_new_n6110__ = ~new_new_n6107__ & new_new_n6109__;
  assign new_new_n6111__ = new_new_n2410__ & new_new_n6110__;
  assign new_new_n6112__ = new_new_n538__ & new_new_n6111__;
  assign new_new_n6113__ = ~new_new_n175__ & ~new_new_n351__;
  assign new_new_n6114__ = ~new_new_n423__ & ~new_new_n1124__;
  assign new_new_n6115__ = new_new_n6113__ & new_new_n6114__;
  assign new_new_n6116__ = new_new_n385__ & ~new_new_n745__;
  assign new_new_n6117__ = ~new_new_n6100__ & new_new_n6116__;
  assign new_new_n6118__ = ~new_new_n6103__ & new_new_n6115__;
  assign new_new_n6119__ = new_new_n6117__ & new_new_n6118__;
  assign new_new_n6120__ = new_new_n955__ & new_new_n6119__;
  assign new_new_n6121__ = new_new_n6112__ & new_new_n6120__;
  assign new_new_n6122__ = new_new_n4290__ & new_new_n6121__;
  assign new_new_n6123__ = ~new_new_n6099__ & new_new_n6122__;
  assign new_new_n6124__ = new_new_n6099__ & ~new_new_n6122__;
  assign new_new_n6125__ = ~new_new_n6123__ & ~new_new_n6124__;
  assign new_new_n6126__ = new_new_n5974__ & ~new_new_n6125__;
  assign new_new_n6127__ = ~new_new_n5974__ & new_new_n6125__;
  assign po08 = ~new_new_n6126__ & ~new_new_n6127__;
  assign new_new_n6129__ = ~new_new_n301__ & ~new_new_n5849__;
  assign new_new_n6130__ = new_new_n301__ & new_new_n5122__;
  assign new_new_n6131__ = new_new_n316__ & ~new_new_n4857__;
  assign new_new_n6132__ = ~new_new_n5122__ & ~new_new_n6131__;
  assign new_new_n6133__ = ~new_new_n318__ & ~new_new_n6130__;
  assign new_new_n6134__ = ~new_new_n6132__ & new_new_n6133__;
  assign new_new_n6135__ = new_new_n301__ & ~new_new_n6131__;
  assign new_new_n6136__ = new_new_n311__ & ~new_new_n6135__;
  assign new_new_n6137__ = ~new_new_n6129__ & ~new_new_n6136__;
  assign new_new_n6138__ = ~new_new_n6134__ & new_new_n6137__;
  assign new_new_n6139__ = new_new_n2809__ & new_new_n4421__;
  assign new_new_n6140__ = ~new_new_n2806__ & new_new_n4222__;
  assign new_new_n6141__ = ~new_new_n6139__ & ~new_new_n6140__;
  assign new_new_n6142__ = new_new_n2808__ & new_new_n5226__;
  assign new_new_n6143__ = new_new_n6141__ & ~new_new_n6142__;
  assign new_new_n6144__ = ~new_new_n810__ & ~new_new_n6143__;
  assign new_new_n6145__ = new_new_n2808__ & ~new_new_n5219__;
  assign new_new_n6146__ = new_new_n810__ & new_new_n6141__;
  assign new_new_n6147__ = ~new_new_n6145__ & new_new_n6146__;
  assign new_new_n6148__ = ~new_new_n816__ & ~new_new_n5222__;
  assign new_new_n6149__ = new_new_n816__ & ~new_new_n5214__;
  assign new_new_n6150__ = new_new_n2808__ & ~new_new_n6148__;
  assign new_new_n6151__ = ~new_new_n6149__ & new_new_n6150__;
  assign new_new_n6152__ = ~new_new_n6144__ & ~new_new_n6147__;
  assign new_new_n6153__ = ~new_new_n6151__ & new_new_n6152__;
  assign new_new_n6154__ = ~new_new_n6036__ & ~new_new_n6043__;
  assign new_new_n6155__ = ~new_new_n437__ & ~new_new_n6154__;
  assign new_new_n6156__ = ~new_new_n3244__ & ~new_new_n6037__;
  assign new_new_n6157__ = ~new_new_n6155__ & new_new_n6156__;
  assign new_new_n6158__ = new_new_n5734__ & new_new_n6035__;
  assign new_new_n6159__ = ~new_new_n6157__ & ~new_new_n6158__;
  assign new_new_n6160__ = new_new_n6153__ & ~new_new_n6159__;
  assign new_new_n6161__ = ~new_new_n6153__ & new_new_n6159__;
  assign new_new_n6162__ = ~new_new_n6160__ & ~new_new_n6161__;
  assign new_new_n6163__ = ~new_new_n437__ & new_new_n3586__;
  assign new_new_n6164__ = ~new_new_n5720__ & ~new_new_n6163__;
  assign new_new_n6165__ = ~new_new_n3733__ & new_new_n4132__;
  assign new_new_n6166__ = new_new_n3069__ & ~new_new_n3727__;
  assign new_new_n6167__ = ~new_new_n2848__ & ~new_new_n6165__;
  assign new_new_n6168__ = ~new_new_n6166__ & new_new_n6167__;
  assign new_new_n6169__ = ~new_new_n3072__ & new_new_n4086__;
  assign new_new_n6170__ = ~new_new_n4081__ & new_new_n6169__;
  assign new_new_n6171__ = new_new_n4081__ & ~new_new_n6169__;
  assign new_new_n6172__ = new_new_n2848__ & ~new_new_n6170__;
  assign new_new_n6173__ = ~new_new_n6171__ & new_new_n6172__;
  assign new_new_n6174__ = ~new_new_n6168__ & ~new_new_n6173__;
  assign new_new_n6175__ = ~new_new_n3651__ & new_new_n6174__;
  assign new_new_n6176__ = new_new_n3651__ & ~new_new_n6174__;
  assign new_new_n6177__ = ~new_new_n6175__ & ~new_new_n6176__;
  assign new_new_n6178__ = ~new_new_n6164__ & ~new_new_n6177__;
  assign new_new_n6179__ = new_new_n6164__ & new_new_n6177__;
  assign new_new_n6180__ = ~new_new_n6178__ & ~new_new_n6179__;
  assign new_new_n6181__ = new_new_n6162__ & new_new_n6180__;
  assign new_new_n6182__ = ~new_new_n6162__ & ~new_new_n6180__;
  assign new_new_n6183__ = ~new_new_n6181__ & ~new_new_n6182__;
  assign new_new_n6184__ = ~new_new_n6138__ & ~new_new_n6183__;
  assign new_new_n6185__ = new_new_n6138__ & new_new_n6183__;
  assign new_new_n6186__ = ~new_new_n6184__ & ~new_new_n6185__;
  assign new_new_n6187__ = ~new_new_n6057__ & ~new_new_n6082__;
  assign new_new_n6188__ = ~new_new_n6058__ & ~new_new_n6187__;
  assign new_new_n6189__ = new_new_n6186__ & ~new_new_n6188__;
  assign new_new_n6190__ = ~new_new_n6186__ & new_new_n6188__;
  assign new_new_n6191__ = ~new_new_n6189__ & ~new_new_n6190__;
  assign new_new_n6192__ = ~new_new_n6087__ & ~new_new_n6090__;
  assign new_new_n6193__ = ~new_new_n6086__ & ~new_new_n6192__;
  assign new_new_n6194__ = new_new_n5992__ & new_new_n6193__;
  assign new_new_n6195__ = new_new_n6086__ & ~new_new_n6090__;
  assign new_new_n6196__ = new_new_n6087__ & new_new_n6090__;
  assign new_new_n6197__ = ~new_new_n6195__ & ~new_new_n6196__;
  assign new_new_n6198__ = new_new_n5993__ & new_new_n6197__;
  assign new_new_n6199__ = new_new_n5991__ & ~new_new_n6193__;
  assign new_new_n6200__ = new_new_n6191__ & ~new_new_n6194__;
  assign new_new_n6201__ = ~new_new_n6199__ & new_new_n6200__;
  assign new_new_n6202__ = ~new_new_n6198__ & new_new_n6201__;
  assign new_new_n6203__ = new_new_n5992__ & ~new_new_n6085__;
  assign new_new_n6204__ = ~new_new_n6003__ & new_new_n6203__;
  assign new_new_n6205__ = new_new_n5991__ & new_new_n6085__;
  assign new_new_n6206__ = ~new_new_n5991__ & ~new_new_n6085__;
  assign new_new_n6207__ = ~new_new_n5992__ & ~new_new_n6206__;
  assign new_new_n6208__ = new_new_n6003__ & new_new_n6207__;
  assign new_new_n6209__ = ~new_new_n6205__ & ~new_new_n6208__;
  assign new_new_n6210__ = new_new_n6090__ & ~new_new_n6209__;
  assign new_new_n6211__ = new_new_n6003__ & ~new_new_n6203__;
  assign new_new_n6212__ = ~new_new_n6090__ & ~new_new_n6207__;
  assign new_new_n6213__ = ~new_new_n6211__ & new_new_n6212__;
  assign new_new_n6214__ = new_new_n5991__ & new_new_n6087__;
  assign new_new_n6215__ = ~new_new_n6191__ & ~new_new_n6214__;
  assign new_new_n6216__ = ~new_new_n6204__ & new_new_n6215__;
  assign new_new_n6217__ = ~new_new_n6213__ & new_new_n6216__;
  assign new_new_n6218__ = ~new_new_n6210__ & new_new_n6217__;
  assign new_new_n6219__ = ~new_new_n6202__ & ~new_new_n6218__;
  assign new_new_n6220__ = new_new_n136__ & new_new_n160__;
  assign new_new_n6221__ = new_new_n162__ & ~new_new_n6220__;
  assign new_new_n6222__ = new_new_n279__ & ~new_new_n446__;
  assign new_new_n6223__ = ~new_new_n377__ & ~new_new_n403__;
  assign new_new_n6224__ = ~new_new_n555__ & ~new_new_n4207__;
  assign new_new_n6225__ = ~new_new_n6221__ & new_new_n6224__;
  assign new_new_n6226__ = new_new_n6222__ & new_new_n6223__;
  assign new_new_n6227__ = new_new_n6225__ & new_new_n6226__;
  assign new_new_n6228__ = new_new_n332__ & new_new_n4715__;
  assign new_new_n6229__ = new_new_n6227__ & new_new_n6228__;
  assign new_new_n6230__ = new_new_n4463__ & new_new_n6229__;
  assign new_new_n6231__ = new_new_n2468__ & new_new_n6230__;
  assign new_new_n6232__ = new_new_n6219__ & new_new_n6231__;
  assign new_new_n6233__ = ~new_new_n6219__ & ~new_new_n6231__;
  assign new_new_n6234__ = ~new_new_n6232__ & ~new_new_n6233__;
  assign new_new_n6235__ = new_new_n6097__ & new_new_n6234__;
  assign new_new_n6236__ = ~new_new_n4702__ & new_new_n6125__;
  assign new_new_n6237__ = ~new_new_n5973__ & ~new_new_n6236__;
  assign new_new_n6238__ = new_new_n5976__ & ~new_new_n6234__;
  assign new_new_n6239__ = new_new_n6237__ & new_new_n6238__;
  assign new_new_n6240__ = ~new_new_n6235__ & ~new_new_n6239__;
  assign new_new_n6241__ = new_new_n5971__ & ~new_new_n6240__;
  assign new_new_n6242__ = new_new_n6234__ & new_new_n6237__;
  assign new_new_n6243__ = new_new_n5974__ & ~new_new_n6236__;
  assign new_new_n6244__ = ~new_new_n6234__ & ~new_new_n6243__;
  assign new_new_n6245__ = ~new_new_n6098__ & ~new_new_n6242__;
  assign new_new_n6246__ = ~new_new_n6244__ & new_new_n6245__;
  assign new_new_n6247__ = ~new_new_n6241__ & ~new_new_n6246__;
  assign new_new_n6248__ = ~new_new_n6122__ & ~new_new_n6247__;
  assign new_new_n6249__ = new_new_n6234__ & ~new_new_n6243__;
  assign new_new_n6250__ = ~new_new_n6096__ & ~new_new_n6122__;
  assign new_new_n6251__ = new_new_n5971__ & new_new_n6237__;
  assign new_new_n6252__ = ~new_new_n5976__ & ~new_new_n6251__;
  assign new_new_n6253__ = ~new_new_n6239__ & ~new_new_n6250__;
  assign new_new_n6254__ = ~new_new_n6249__ & new_new_n6253__;
  assign new_new_n6255__ = ~new_new_n6252__ & new_new_n6254__;
  assign new_new_n6256__ = new_new_n6096__ & new_new_n6122__;
  assign new_new_n6257__ = ~new_new_n6234__ & new_new_n6256__;
  assign new_new_n6258__ = ~new_new_n6235__ & ~new_new_n6257__;
  assign new_new_n6259__ = ~new_new_n6237__ & new_new_n6258__;
  assign new_new_n6260__ = new_new_n6097__ & ~new_new_n6234__;
  assign new_new_n6261__ = new_new_n6234__ & new_new_n6256__;
  assign new_new_n6262__ = ~new_new_n6260__ & ~new_new_n6261__;
  assign new_new_n6263__ = ~new_new_n5971__ & ~new_new_n6262__;
  assign new_new_n6264__ = new_new_n5971__ & ~new_new_n6096__;
  assign new_new_n6265__ = ~new_new_n6234__ & new_new_n6264__;
  assign new_new_n6266__ = ~new_new_n6261__ & ~new_new_n6265__;
  assign new_new_n6267__ = new_new_n5976__ & ~new_new_n6266__;
  assign new_new_n6268__ = ~new_new_n6263__ & ~new_new_n6267__;
  assign new_new_n6269__ = new_new_n6237__ & new_new_n6268__;
  assign new_new_n6270__ = ~new_new_n6259__ & ~new_new_n6269__;
  assign new_new_n6271__ = ~new_new_n6255__ & ~new_new_n6270__;
  assign po09 = new_new_n6248__ | ~new_new_n6271__;
  assign new_new_n6273__ = ~new_new_n6098__ & ~new_new_n6122__;
  assign new_new_n6274__ = new_new_n6234__ & ~new_new_n6273__;
  assign new_new_n6275__ = ~new_new_n6260__ & ~new_new_n6274__;
  assign new_new_n6276__ = new_new_n5971__ & ~new_new_n6123__;
  assign new_new_n6277__ = ~new_new_n6275__ & new_new_n6276__;
  assign new_new_n6278__ = new_new_n4702__ & ~new_new_n6277__;
  assign new_new_n6279__ = new_new_n5972__ & new_new_n6122__;
  assign new_new_n6280__ = new_new_n6097__ & new_new_n6279__;
  assign new_new_n6281__ = ~new_new_n5971__ & new_new_n6122__;
  assign new_new_n6282__ = ~new_new_n5972__ & ~new_new_n6122__;
  assign new_new_n6283__ = new_new_n6099__ & ~new_new_n6281__;
  assign new_new_n6284__ = ~new_new_n6282__ & new_new_n6283__;
  assign new_new_n6285__ = new_new_n6234__ & ~new_new_n6280__;
  assign new_new_n6286__ = ~new_new_n6284__ & new_new_n6285__;
  assign new_new_n6287__ = new_new_n6098__ & new_new_n6279__;
  assign new_new_n6288__ = ~new_new_n5976__ & new_new_n6250__;
  assign new_new_n6289__ = new_new_n5971__ & new_new_n6288__;
  assign new_new_n6290__ = ~new_new_n6234__ & ~new_new_n6289__;
  assign new_new_n6291__ = ~new_new_n6287__ & new_new_n6290__;
  assign new_new_n6292__ = ~new_new_n6277__ & ~new_new_n6291__;
  assign new_new_n6293__ = ~new_new_n6286__ & new_new_n6292__;
  assign new_new_n6294__ = ~new_new_n6278__ & ~new_new_n6293__;
  assign new_new_n6295__ = ~new_new_n6097__ & ~new_new_n6273__;
  assign new_new_n6296__ = ~new_new_n6232__ & ~new_new_n6295__;
  assign new_new_n6297__ = ~new_new_n6233__ & ~new_new_n6296__;
  assign new_new_n6298__ = ~new_new_n2806__ & new_new_n4421__;
  assign new_new_n6299__ = new_new_n2809__ & ~new_new_n4532__;
  assign new_new_n6300__ = ~new_new_n6298__ & ~new_new_n6299__;
  assign new_new_n6301__ = new_new_n2808__ & ~new_new_n4857__;
  assign new_new_n6302__ = new_new_n4884__ & new_new_n6301__;
  assign new_new_n6303__ = new_new_n6300__ & ~new_new_n6302__;
  assign new_new_n6304__ = new_new_n810__ & ~new_new_n6303__;
  assign new_new_n6305__ = new_new_n2808__ & ~new_new_n5338__;
  assign new_new_n6306__ = ~new_new_n810__ & new_new_n6300__;
  assign new_new_n6307__ = ~new_new_n6305__ & new_new_n6306__;
  assign new_new_n6308__ = new_new_n816__ & ~new_new_n4857__;
  assign new_new_n6309__ = ~new_new_n816__ & new_new_n4884__;
  assign new_new_n6310__ = ~new_new_n6308__ & ~new_new_n6309__;
  assign new_new_n6311__ = new_new_n6305__ & new_new_n6310__;
  assign new_new_n6312__ = ~new_new_n6304__ & ~new_new_n6307__;
  assign new_new_n6313__ = ~new_new_n6311__ & new_new_n6312__;
  assign new_new_n6314__ = new_new_n3067__ & ~new_new_n3726__;
  assign new_new_n6315__ = new_new_n437__ & new_new_n4080__;
  assign new_new_n6316__ = ~new_new_n437__ & new_new_n4081__;
  assign new_new_n6317__ = ~new_new_n6315__ & ~new_new_n6316__;
  assign new_new_n6318__ = ~new_new_n3068__ & ~new_new_n6314__;
  assign new_new_n6319__ = ~new_new_n6317__ & new_new_n6318__;
  assign new_new_n6320__ = ~new_new_n3068__ & ~new_new_n4078__;
  assign new_new_n6321__ = new_new_n3068__ & new_new_n3725__;
  assign new_new_n6322__ = ~new_new_n3726__ & ~new_new_n6320__;
  assign new_new_n6323__ = ~new_new_n6321__ & new_new_n6322__;
  assign new_new_n6324__ = ~new_new_n3067__ & ~new_new_n6323__;
  assign new_new_n6325__ = new_new_n437__ & ~new_new_n6324__;
  assign new_new_n6326__ = new_new_n3067__ & ~new_new_n3727__;
  assign new_new_n6327__ = ~new_new_n2848__ & ~new_new_n6326__;
  assign new_new_n6328__ = ~new_new_n6325__ & new_new_n6327__;
  assign new_new_n6329__ = ~new_new_n6319__ & new_new_n6328__;
  assign new_new_n6330__ = ~new_new_n651__ & new_new_n4233__;
  assign new_new_n6331__ = new_new_n437__ & ~new_new_n4233__;
  assign new_new_n6332__ = ~new_new_n6330__ & ~new_new_n6331__;
  assign new_new_n6333__ = new_new_n4222__ & new_new_n6332__;
  assign new_new_n6334__ = ~new_new_n4222__ & ~new_new_n6332__;
  assign new_new_n6335__ = new_new_n2848__ & ~new_new_n6333__;
  assign new_new_n6336__ = ~new_new_n6334__ & new_new_n6335__;
  assign new_new_n6337__ = ~new_new_n6329__ & ~new_new_n6336__;
  assign new_new_n6338__ = new_new_n437__ & new_new_n6174__;
  assign new_new_n6339__ = ~new_new_n3586__ & ~new_new_n6176__;
  assign new_new_n6340__ = ~new_new_n437__ & ~new_new_n6175__;
  assign new_new_n6341__ = ~new_new_n6339__ & new_new_n6340__;
  assign new_new_n6342__ = ~new_new_n6338__ & ~new_new_n6341__;
  assign new_new_n6343__ = ~new_new_n6337__ & ~new_new_n6342__;
  assign new_new_n6344__ = new_new_n6337__ & new_new_n6342__;
  assign new_new_n6345__ = ~new_new_n6343__ & ~new_new_n6344__;
  assign new_new_n6346__ = ~new_new_n3586__ & ~new_new_n3733__;
  assign new_new_n6347__ = new_new_n3586__ & new_new_n3733__;
  assign new_new_n6348__ = ~new_new_n437__ & ~new_new_n6346__;
  assign new_new_n6349__ = ~new_new_n6347__ & new_new_n6348__;
  assign new_new_n6350__ = new_new_n301__ & new_new_n6349__;
  assign new_new_n6351__ = ~new_new_n301__ & ~new_new_n6349__;
  assign new_new_n6352__ = ~new_new_n6350__ & ~new_new_n6351__;
  assign new_new_n6353__ = new_new_n6345__ & ~new_new_n6352__;
  assign new_new_n6354__ = ~new_new_n6345__ & new_new_n6352__;
  assign new_new_n6355__ = ~new_new_n6353__ & ~new_new_n6354__;
  assign new_new_n6356__ = new_new_n6313__ & ~new_new_n6355__;
  assign new_new_n6357__ = ~new_new_n6313__ & new_new_n6355__;
  assign new_new_n6358__ = ~new_new_n6356__ & ~new_new_n6357__;
  assign new_new_n6359__ = ~new_new_n6185__ & ~new_new_n6188__;
  assign new_new_n6360__ = ~new_new_n6184__ & ~new_new_n6359__;
  assign new_new_n6361__ = new_new_n6191__ & new_new_n6193__;
  assign new_new_n6362__ = new_new_n5992__ & ~new_new_n6361__;
  assign new_new_n6363__ = new_new_n6191__ & ~new_new_n6195__;
  assign new_new_n6364__ = ~new_new_n6196__ & ~new_new_n6363__;
  assign new_new_n6365__ = ~new_new_n5991__ & new_new_n6364__;
  assign new_new_n6366__ = ~new_new_n6191__ & ~new_new_n6193__;
  assign new_new_n6367__ = ~new_new_n6362__ & ~new_new_n6366__;
  assign new_new_n6368__ = ~new_new_n6365__ & new_new_n6367__;
  assign new_new_n6369__ = new_new_n6360__ & ~new_new_n6368__;
  assign new_new_n6370__ = ~new_new_n6360__ & new_new_n6368__;
  assign new_new_n6371__ = ~new_new_n6369__ & ~new_new_n6370__;
  assign new_new_n6372__ = ~new_new_n6160__ & ~new_new_n6180__;
  assign new_new_n6373__ = ~new_new_n6161__ & ~new_new_n6372__;
  assign new_new_n6374__ = new_new_n6371__ & ~new_new_n6373__;
  assign new_new_n6375__ = ~new_new_n6371__ & new_new_n6373__;
  assign new_new_n6376__ = ~new_new_n6374__ & ~new_new_n6375__;
  assign new_new_n6377__ = new_new_n6358__ & new_new_n6376__;
  assign new_new_n6378__ = ~new_new_n6358__ & ~new_new_n6376__;
  assign new_new_n6379__ = ~new_new_n6377__ & ~new_new_n6378__;
  assign new_new_n6380__ = ~new_new_n6297__ & new_new_n6379__;
  assign new_new_n6381__ = new_new_n6297__ & ~new_new_n6379__;
  assign new_new_n6382__ = ~new_new_n6380__ & ~new_new_n6381__;
  assign new_new_n6383__ = ~new_new_n136__ & new_new_n223__;
  assign new_new_n6384__ = ~new_new_n619__ & ~new_new_n6383__;
  assign new_new_n6385__ = ~new_new_n243__ & new_new_n6384__;
  assign new_new_n6386__ = new_new_n3616__ & ~new_new_n4207__;
  assign new_new_n6387__ = ~new_new_n4673__ & new_new_n6386__;
  assign new_new_n6388__ = new_new_n4847__ & new_new_n6385__;
  assign new_new_n6389__ = new_new_n6387__ & new_new_n6388__;
  assign new_new_n6390__ = ~new_new_n367__ & new_new_n3695__;
  assign new_new_n6391__ = new_new_n6389__ & new_new_n6390__;
  assign new_new_n6392__ = new_new_n742__ & new_new_n6391__;
  assign new_new_n6393__ = new_new_n4272__ & new_new_n6392__;
  assign new_new_n6394__ = new_new_n1079__ & new_new_n6393__;
  assign new_new_n6395__ = ~new_new_n6382__ & new_new_n6394__;
  assign new_new_n6396__ = new_new_n6382__ & ~new_new_n6394__;
  assign new_new_n6397__ = ~new_new_n6395__ & ~new_new_n6396__;
  assign new_new_n6398__ = new_new_n6294__ & new_new_n6397__;
  assign new_new_n6399__ = ~new_new_n6294__ & ~new_new_n6397__;
  assign po10 = ~new_new_n6398__ & ~new_new_n6399__;
  assign new_new_n6401__ = new_new_n6277__ & new_new_n6397__;
  assign new_new_n6402__ = new_new_n6293__ & ~new_new_n6397__;
  assign new_new_n6403__ = ~new_new_n4702__ & ~new_new_n6402__;
  assign new_new_n6404__ = ~new_new_n6401__ & ~new_new_n6403__;
  assign new_new_n6405__ = new_new_n6356__ & ~new_new_n6373__;
  assign new_new_n6406__ = ~new_new_n6369__ & new_new_n6405__;
  assign new_new_n6407__ = ~new_new_n6356__ & new_new_n6373__;
  assign new_new_n6408__ = new_new_n6370__ & ~new_new_n6407__;
  assign new_new_n6409__ = ~new_new_n3065__ & new_new_n4081__;
  assign new_new_n6410__ = new_new_n3070__ & new_new_n4222__;
  assign new_new_n6411__ = ~new_new_n6409__ & ~new_new_n6410__;
  assign new_new_n6412__ = new_new_n2848__ & ~new_new_n5037__;
  assign new_new_n6413__ = ~new_new_n437__ & ~new_new_n6412__;
  assign new_new_n6414__ = ~new_new_n651__ & ~new_new_n5040__;
  assign new_new_n6415__ = new_new_n651__ & ~new_new_n5032__;
  assign new_new_n6416__ = new_new_n2848__ & ~new_new_n6414__;
  assign new_new_n6417__ = ~new_new_n6415__ & new_new_n6416__;
  assign new_new_n6418__ = ~new_new_n6413__ & ~new_new_n6417__;
  assign new_new_n6419__ = new_new_n6411__ & ~new_new_n6418__;
  assign new_new_n6420__ = new_new_n2848__ & new_new_n4421__;
  assign new_new_n6421__ = new_new_n4444__ & new_new_n6420__;
  assign new_new_n6422__ = new_new_n6411__ & ~new_new_n6421__;
  assign new_new_n6423__ = new_new_n437__ & ~new_new_n6422__;
  assign new_new_n6424__ = ~new_new_n6419__ & ~new_new_n6423__;
  assign new_new_n6425__ = new_new_n301__ & ~new_new_n6347__;
  assign new_new_n6426__ = ~new_new_n6346__ & ~new_new_n6425__;
  assign new_new_n6427__ = ~new_new_n3727__ & ~new_new_n6426__;
  assign new_new_n6428__ = new_new_n3727__ & new_new_n6426__;
  assign new_new_n6429__ = ~new_new_n437__ & ~new_new_n6427__;
  assign new_new_n6430__ = ~new_new_n6428__ & new_new_n6429__;
  assign new_new_n6431__ = ~new_new_n6424__ & new_new_n6430__;
  assign new_new_n6432__ = new_new_n6424__ & ~new_new_n6430__;
  assign new_new_n6433__ = ~new_new_n6431__ & ~new_new_n6432__;
  assign new_new_n6434__ = ~new_new_n6344__ & new_new_n6352__;
  assign new_new_n6435__ = ~new_new_n6343__ & ~new_new_n6434__;
  assign new_new_n6436__ = new_new_n3088__ & new_new_n4923__;
  assign new_new_n6437__ = new_new_n2809__ & ~new_new_n4857__;
  assign new_new_n6438__ = ~new_new_n2806__ & ~new_new_n4532__;
  assign new_new_n6439__ = ~new_new_n6437__ & ~new_new_n6438__;
  assign new_new_n6440__ = ~new_new_n810__ & ~new_new_n6439__;
  assign new_new_n6441__ = new_new_n2808__ & new_new_n4923__;
  assign new_new_n6442__ = new_new_n810__ & new_new_n6439__;
  assign new_new_n6443__ = ~new_new_n6441__ & new_new_n6442__;
  assign new_new_n6444__ = ~new_new_n6436__ & ~new_new_n6440__;
  assign new_new_n6445__ = ~new_new_n6443__ & new_new_n6444__;
  assign new_new_n6446__ = ~new_new_n6435__ & ~new_new_n6445__;
  assign new_new_n6447__ = new_new_n6435__ & new_new_n6445__;
  assign new_new_n6448__ = ~new_new_n6446__ & ~new_new_n6447__;
  assign new_new_n6449__ = new_new_n6433__ & new_new_n6448__;
  assign new_new_n6450__ = ~new_new_n6433__ & ~new_new_n6448__;
  assign new_new_n6451__ = ~new_new_n6449__ & ~new_new_n6450__;
  assign new_new_n6452__ = ~new_new_n6406__ & ~new_new_n6451__;
  assign new_new_n6453__ = ~new_new_n6408__ & new_new_n6452__;
  assign new_new_n6454__ = new_new_n6369__ & ~new_new_n6407__;
  assign new_new_n6455__ = new_new_n6371__ & new_new_n6373__;
  assign new_new_n6456__ = new_new_n6451__ & ~new_new_n6454__;
  assign new_new_n6457__ = ~new_new_n6455__ & new_new_n6456__;
  assign new_new_n6458__ = ~new_new_n6357__ & ~new_new_n6453__;
  assign new_new_n6459__ = ~new_new_n6457__ & new_new_n6458__;
  assign new_new_n6460__ = ~new_new_n6357__ & ~new_new_n6373__;
  assign new_new_n6461__ = new_new_n6370__ & ~new_new_n6460__;
  assign new_new_n6462__ = new_new_n6451__ & ~new_new_n6461__;
  assign new_new_n6463__ = ~new_new_n6374__ & new_new_n6462__;
  assign new_new_n6464__ = new_new_n6360__ & new_new_n6373__;
  assign new_new_n6465__ = ~new_new_n6357__ & ~new_new_n6464__;
  assign new_new_n6466__ = ~new_new_n6360__ & ~new_new_n6373__;
  assign new_new_n6467__ = ~new_new_n6465__ & ~new_new_n6466__;
  assign new_new_n6468__ = ~new_new_n6368__ & new_new_n6467__;
  assign new_new_n6469__ = ~new_new_n6451__ & ~new_new_n6468__;
  assign new_new_n6470__ = ~new_new_n6356__ & ~new_new_n6469__;
  assign new_new_n6471__ = ~new_new_n6463__ & new_new_n6470__;
  assign new_new_n6472__ = new_new_n6357__ & ~new_new_n6451__;
  assign new_new_n6473__ = new_new_n6464__ & new_new_n6472__;
  assign new_new_n6474__ = new_new_n6368__ & new_new_n6473__;
  assign new_new_n6475__ = ~new_new_n6471__ & ~new_new_n6474__;
  assign new_new_n6476__ = ~new_new_n6459__ & new_new_n6475__;
  assign new_new_n6477__ = ~new_new_n6380__ & new_new_n6394__;
  assign new_new_n6478__ = ~new_new_n6381__ & ~new_new_n6477__;
  assign new_new_n6479__ = ~new_new_n6476__ & new_new_n6478__;
  assign new_new_n6480__ = new_new_n6476__ & ~new_new_n6478__;
  assign new_new_n6481__ = ~new_new_n6479__ & ~new_new_n6480__;
  assign new_new_n6482__ = ~new_new_n99__ & ~new_new_n238__;
  assign new_new_n6483__ = new_new_n162__ & ~new_new_n246__;
  assign new_new_n6484__ = new_new_n411__ & ~new_new_n6482__;
  assign new_new_n6485__ = ~new_new_n446__ & ~new_new_n2413__;
  assign new_new_n6486__ = new_new_n6484__ & new_new_n6485__;
  assign new_new_n6487__ = ~new_new_n243__ & ~new_new_n471__;
  assign new_new_n6488__ = ~new_new_n6483__ & new_new_n6487__;
  assign new_new_n6489__ = ~new_new_n667__ & new_new_n6486__;
  assign new_new_n6490__ = new_new_n6488__ & new_new_n6489__;
  assign new_new_n6491__ = new_new_n4521__ & new_new_n6490__;
  assign new_new_n6492__ = new_new_n723__ & new_new_n6491__;
  assign new_new_n6493__ = new_new_n707__ & new_new_n6492__;
  assign new_new_n6494__ = ~new_new_n6481__ & new_new_n6493__;
  assign new_new_n6495__ = new_new_n6481__ & ~new_new_n6493__;
  assign new_new_n6496__ = ~new_new_n6494__ & ~new_new_n6495__;
  assign new_new_n6497__ = ~new_new_n6404__ & ~new_new_n6496__;
  assign new_new_n6498__ = new_new_n6404__ & new_new_n6496__;
  assign po11 = new_new_n6497__ | new_new_n6498__;
  assign new_new_n6500__ = new_new_n223__ & ~new_new_n1116__;
  assign new_new_n6501__ = ~new_new_n100__ & new_new_n110__;
  assign new_new_n6502__ = ~new_new_n365__ & ~new_new_n6501__;
  assign new_new_n6503__ = ~new_new_n257__ & ~new_new_n6500__;
  assign new_new_n6504__ = ~new_new_n6502__ & new_new_n6503__;
  assign new_new_n6505__ = ~new_new_n348__ & ~new_new_n714__;
  assign new_new_n6506__ = ~new_new_n2230__ & new_new_n6505__;
  assign new_new_n6507__ = ~new_new_n3463__ & new_new_n6506__;
  assign new_new_n6508__ = new_new_n894__ & new_new_n6507__;
  assign new_new_n6509__ = new_new_n5072__ & new_new_n6504__;
  assign new_new_n6510__ = new_new_n6508__ & new_new_n6509__;
  assign new_new_n6511__ = new_new_n2257__ & new_new_n6510__;
  assign new_new_n6512__ = new_new_n3187__ & new_new_n6511__;
  assign new_new_n6513__ = new_new_n3070__ & new_new_n4421__;
  assign new_new_n6514__ = ~new_new_n3065__ & new_new_n4222__;
  assign new_new_n6515__ = ~new_new_n6513__ & ~new_new_n6514__;
  assign new_new_n6516__ = new_new_n2848__ & new_new_n5226__;
  assign new_new_n6517__ = new_new_n6515__ & ~new_new_n6516__;
  assign new_new_n6518__ = new_new_n437__ & ~new_new_n6517__;
  assign new_new_n6519__ = new_new_n2848__ & ~new_new_n5219__;
  assign new_new_n6520__ = ~new_new_n437__ & new_new_n6515__;
  assign new_new_n6521__ = ~new_new_n6519__ & new_new_n6520__;
  assign new_new_n6522__ = ~new_new_n651__ & ~new_new_n5214__;
  assign new_new_n6523__ = new_new_n651__ & ~new_new_n5222__;
  assign new_new_n6524__ = new_new_n2848__ & ~new_new_n6522__;
  assign new_new_n6525__ = ~new_new_n6523__ & new_new_n6524__;
  assign new_new_n6526__ = ~new_new_n6518__ & ~new_new_n6521__;
  assign new_new_n6527__ = ~new_new_n6525__ & new_new_n6526__;
  assign new_new_n6528__ = ~new_new_n6451__ & new_new_n6466__;
  assign new_new_n6529__ = ~new_new_n6356__ & new_new_n6451__;
  assign new_new_n6530__ = new_new_n6368__ & ~new_new_n6529__;
  assign new_new_n6531__ = ~new_new_n6357__ & ~new_new_n6451__;
  assign new_new_n6532__ = ~new_new_n6530__ & ~new_new_n6531__;
  assign new_new_n6533__ = ~new_new_n6464__ & ~new_new_n6532__;
  assign new_new_n6534__ = new_new_n6451__ & ~new_new_n6466__;
  assign new_new_n6535__ = ~new_new_n6357__ & new_new_n6368__;
  assign new_new_n6536__ = ~new_new_n6356__ & ~new_new_n6535__;
  assign new_new_n6537__ = ~new_new_n6534__ & ~new_new_n6536__;
  assign new_new_n6538__ = ~new_new_n6528__ & ~new_new_n6533__;
  assign new_new_n6539__ = ~new_new_n6537__ & new_new_n6538__;
  assign new_new_n6540__ = new_new_n6527__ & new_new_n6539__;
  assign new_new_n6541__ = ~new_new_n6527__ & ~new_new_n6539__;
  assign new_new_n6542__ = ~new_new_n6540__ & ~new_new_n6541__;
  assign new_new_n6543__ = ~new_new_n4081__ & new_new_n6426__;
  assign new_new_n6544__ = new_new_n4081__ & ~new_new_n6426__;
  assign new_new_n6545__ = ~new_new_n3727__ & new_new_n6544__;
  assign new_new_n6546__ = ~new_new_n437__ & ~new_new_n6543__;
  assign new_new_n6547__ = ~new_new_n6545__ & new_new_n6546__;
  assign new_new_n6548__ = ~new_new_n6424__ & ~new_new_n6547__;
  assign new_new_n6549__ = ~new_new_n4081__ & new_new_n6424__;
  assign new_new_n6550__ = ~new_new_n3727__ & ~new_new_n6549__;
  assign new_new_n6551__ = new_new_n4081__ & ~new_new_n6424__;
  assign new_new_n6552__ = ~new_new_n6543__ & ~new_new_n6544__;
  assign new_new_n6553__ = ~new_new_n6551__ & new_new_n6552__;
  assign new_new_n6554__ = new_new_n3727__ & ~new_new_n6553__;
  assign new_new_n6555__ = ~new_new_n437__ & ~new_new_n6550__;
  assign new_new_n6556__ = ~new_new_n6554__ & new_new_n6555__;
  assign new_new_n6557__ = ~new_new_n6433__ & ~new_new_n6447__;
  assign new_new_n6558__ = ~new_new_n6446__ & ~new_new_n6557__;
  assign new_new_n6559__ = ~new_new_n6548__ & ~new_new_n6556__;
  assign new_new_n6560__ = ~new_new_n6558__ & new_new_n6559__;
  assign new_new_n6561__ = ~new_new_n437__ & ~new_new_n6544__;
  assign new_new_n6562__ = new_new_n6424__ & ~new_new_n6561__;
  assign new_new_n6563__ = ~new_new_n6316__ & ~new_new_n6426__;
  assign new_new_n6564__ = new_new_n6426__ & ~new_new_n6549__;
  assign new_new_n6565__ = new_new_n3727__ & ~new_new_n6563__;
  assign new_new_n6566__ = ~new_new_n6564__ & new_new_n6565__;
  assign new_new_n6567__ = new_new_n3727__ & ~new_new_n6551__;
  assign new_new_n6568__ = ~new_new_n6544__ & new_new_n6546__;
  assign new_new_n6569__ = ~new_new_n6549__ & new_new_n6568__;
  assign new_new_n6570__ = ~new_new_n6567__ & new_new_n6569__;
  assign new_new_n6571__ = ~new_new_n6562__ & ~new_new_n6566__;
  assign new_new_n6572__ = ~new_new_n6570__ & new_new_n6571__;
  assign new_new_n6573__ = new_new_n6558__ & new_new_n6572__;
  assign new_new_n6574__ = ~new_new_n6560__ & ~new_new_n6573__;
  assign new_new_n6575__ = new_new_n810__ & ~new_new_n6308__;
  assign new_new_n6576__ = ~new_new_n816__ & ~new_new_n4857__;
  assign new_new_n6577__ = ~new_new_n5122__ & ~new_new_n6576__;
  assign new_new_n6578__ = ~new_new_n810__ & new_new_n5122__;
  assign new_new_n6579__ = ~new_new_n2803__ & ~new_new_n6577__;
  assign new_new_n6580__ = ~new_new_n6578__ & new_new_n6579__;
  assign new_new_n6581__ = ~new_new_n810__ & ~new_new_n6576__;
  assign new_new_n6582__ = new_new_n2800__ & ~new_new_n6581__;
  assign new_new_n6583__ = ~new_new_n6575__ & ~new_new_n6582__;
  assign new_new_n6584__ = ~new_new_n6580__ & new_new_n6583__;
  assign new_new_n6585__ = new_new_n6574__ & ~new_new_n6584__;
  assign new_new_n6586__ = ~new_new_n6574__ & new_new_n6584__;
  assign new_new_n6587__ = ~new_new_n6585__ & ~new_new_n6586__;
  assign new_new_n6588__ = new_new_n6542__ & new_new_n6587__;
  assign new_new_n6589__ = ~new_new_n6542__ & ~new_new_n6587__;
  assign new_new_n6590__ = ~new_new_n6588__ & ~new_new_n6589__;
  assign new_new_n6591__ = ~new_new_n6512__ & new_new_n6590__;
  assign new_new_n6592__ = new_new_n6512__ & ~new_new_n6590__;
  assign new_new_n6593__ = ~new_new_n6591__ & ~new_new_n6592__;
  assign new_new_n6594__ = ~new_new_n6479__ & new_new_n6493__;
  assign new_new_n6595__ = ~new_new_n6480__ & ~new_new_n6594__;
  assign new_new_n6596__ = new_new_n6593__ & ~new_new_n6595__;
  assign new_new_n6597__ = ~new_new_n6593__ & new_new_n6595__;
  assign new_new_n6598__ = ~new_new_n6596__ & ~new_new_n6597__;
  assign new_new_n6599__ = new_new_n6496__ & ~new_new_n6598__;
  assign new_new_n6600__ = new_new_n6401__ & new_new_n6599__;
  assign new_new_n6601__ = ~new_new_n4702__ & ~new_new_n6598__;
  assign new_new_n6602__ = ~new_new_n6496__ & new_new_n6598__;
  assign new_new_n6603__ = new_new_n6402__ & new_new_n6602__;
  assign new_new_n6604__ = new_new_n4702__ & new_new_n6598__;
  assign new_new_n6605__ = ~new_new_n6601__ & ~new_new_n6604__;
  assign new_new_n6606__ = ~new_new_n6600__ & new_new_n6605__;
  assign new_new_n6607__ = ~new_new_n6603__ & new_new_n6606__;
  assign new_new_n6608__ = ~po11 & ~new_new_n6599__;
  assign new_new_n6609__ = ~new_new_n6602__ & new_new_n6608__;
  assign po12 = new_new_n6607__ | new_new_n6609__;
  assign new_new_n6611__ = ~new_new_n3065__ & new_new_n4421__;
  assign new_new_n6612__ = new_new_n3070__ & ~new_new_n4532__;
  assign new_new_n6613__ = ~new_new_n6611__ & ~new_new_n6612__;
  assign new_new_n6614__ = new_new_n2848__ & ~new_new_n4857__;
  assign new_new_n6615__ = new_new_n4884__ & new_new_n6614__;
  assign new_new_n6616__ = new_new_n6613__ & ~new_new_n6615__;
  assign new_new_n6617__ = ~new_new_n437__ & ~new_new_n6616__;
  assign new_new_n6618__ = new_new_n2848__ & ~new_new_n5338__;
  assign new_new_n6619__ = ~new_new_n437__ & ~new_new_n6618__;
  assign new_new_n6620__ = ~new_new_n651__ & new_new_n4857__;
  assign new_new_n6621__ = new_new_n651__ & ~new_new_n4884__;
  assign new_new_n6622__ = new_new_n2848__ & ~new_new_n6620__;
  assign new_new_n6623__ = ~new_new_n6621__ & new_new_n6622__;
  assign new_new_n6624__ = new_new_n6613__ & ~new_new_n6623__;
  assign new_new_n6625__ = ~new_new_n6619__ & new_new_n6624__;
  assign new_new_n6626__ = ~new_new_n6617__ & ~new_new_n6625__;
  assign new_new_n6627__ = ~new_new_n3725__ & ~new_new_n4078__;
  assign new_new_n6628__ = ~new_new_n6426__ & ~new_new_n6627__;
  assign new_new_n6629__ = ~new_new_n437__ & ~new_new_n4079__;
  assign new_new_n6630__ = ~new_new_n6628__ & new_new_n6629__;
  assign new_new_n6631__ = ~new_new_n6424__ & ~new_new_n6630__;
  assign new_new_n6632__ = ~new_new_n437__ & ~new_new_n4081__;
  assign new_new_n6633__ = ~new_new_n6428__ & new_new_n6632__;
  assign new_new_n6634__ = ~new_new_n6631__ & ~new_new_n6633__;
  assign new_new_n6635__ = new_new_n6626__ & ~new_new_n6634__;
  assign new_new_n6636__ = ~new_new_n6626__ & new_new_n6634__;
  assign new_new_n6637__ = ~new_new_n6635__ & ~new_new_n6636__;
  assign new_new_n6638__ = ~new_new_n4081__ & new_new_n4219__;
  assign new_new_n6639__ = new_new_n4081__ & new_new_n4222__;
  assign new_new_n6640__ = ~new_new_n437__ & ~new_new_n6638__;
  assign new_new_n6641__ = ~new_new_n6639__ & new_new_n6640__;
  assign new_new_n6642__ = new_new_n810__ & new_new_n6641__;
  assign new_new_n6643__ = ~new_new_n810__ & ~new_new_n6641__;
  assign new_new_n6644__ = ~new_new_n6642__ & ~new_new_n6643__;
  assign new_new_n6645__ = new_new_n6637__ & ~new_new_n6644__;
  assign new_new_n6646__ = ~new_new_n6637__ & new_new_n6644__;
  assign new_new_n6647__ = ~new_new_n6645__ & ~new_new_n6646__;
  assign new_new_n6648__ = new_new_n6539__ & new_new_n6573__;
  assign new_new_n6649__ = new_new_n6527__ & new_new_n6648__;
  assign new_new_n6650__ = ~new_new_n6539__ & new_new_n6560__;
  assign new_new_n6651__ = new_new_n6539__ & ~new_new_n6560__;
  assign new_new_n6652__ = ~new_new_n6573__ & ~new_new_n6651__;
  assign new_new_n6653__ = ~new_new_n6527__ & new_new_n6652__;
  assign new_new_n6654__ = ~new_new_n6650__ & ~new_new_n6653__;
  assign new_new_n6655__ = ~new_new_n6584__ & ~new_new_n6654__;
  assign new_new_n6656__ = ~new_new_n6527__ & ~new_new_n6648__;
  assign new_new_n6657__ = new_new_n6584__ & ~new_new_n6652__;
  assign new_new_n6658__ = ~new_new_n6656__ & new_new_n6657__;
  assign new_new_n6659__ = new_new_n6541__ & new_new_n6560__;
  assign new_new_n6660__ = new_new_n6647__ & ~new_new_n6649__;
  assign new_new_n6661__ = ~new_new_n6659__ & new_new_n6660__;
  assign new_new_n6662__ = ~new_new_n6658__ & new_new_n6661__;
  assign new_new_n6663__ = ~new_new_n6655__ & new_new_n6662__;
  assign new_new_n6664__ = new_new_n6573__ & ~new_new_n6584__;
  assign new_new_n6665__ = ~new_new_n6527__ & ~new_new_n6584__;
  assign new_new_n6666__ = ~new_new_n6573__ & ~new_new_n6665__;
  assign new_new_n6667__ = ~new_new_n6527__ & new_new_n6573__;
  assign new_new_n6668__ = ~new_new_n6666__ & ~new_new_n6667__;
  assign new_new_n6669__ = ~new_new_n6560__ & ~new_new_n6668__;
  assign new_new_n6670__ = ~new_new_n6664__ & ~new_new_n6669__;
  assign new_new_n6671__ = ~new_new_n6539__ & ~new_new_n6670__;
  assign new_new_n6672__ = new_new_n6527__ & new_new_n6584__;
  assign new_new_n6673__ = new_new_n6560__ & new_new_n6672__;
  assign new_new_n6674__ = ~new_new_n6560__ & new_new_n6665__;
  assign new_new_n6675__ = ~new_new_n6666__ & ~new_new_n6674__;
  assign new_new_n6676__ = ~new_new_n6672__ & ~new_new_n6675__;
  assign new_new_n6677__ = new_new_n6539__ & new_new_n6676__;
  assign new_new_n6678__ = ~new_new_n6647__ & ~new_new_n6673__;
  assign new_new_n6679__ = ~new_new_n6671__ & new_new_n6678__;
  assign new_new_n6680__ = ~new_new_n6677__ & new_new_n6679__;
  assign new_new_n6681__ = ~new_new_n6663__ & ~new_new_n6680__;
  assign new_new_n6682__ = ~new_new_n6591__ & ~new_new_n6595__;
  assign new_new_n6683__ = ~new_new_n6592__ & ~new_new_n6682__;
  assign new_new_n6684__ = new_new_n6681__ & new_new_n6683__;
  assign new_new_n6685__ = ~new_new_n6681__ & ~new_new_n6683__;
  assign new_new_n6686__ = ~new_new_n6684__ & ~new_new_n6685__;
  assign new_new_n6687__ = new_new_n218__ & new_new_n2406__;
  assign new_new_n6688__ = ~new_new_n124__ & ~new_new_n3188__;
  assign new_new_n6689__ = new_new_n141__ & ~new_new_n6688__;
  assign new_new_n6690__ = ~new_new_n87__ & ~new_new_n6687__;
  assign new_new_n6691__ = ~new_new_n6689__ & new_new_n6690__;
  assign new_new_n6692__ = ~new_new_n182__ & ~new_new_n261__;
  assign new_new_n6693__ = new_new_n195__ & ~new_new_n798__;
  assign new_new_n6694__ = new_new_n213__ & new_new_n256__;
  assign new_new_n6695__ = new_new_n244__ & ~new_new_n6694__;
  assign new_new_n6696__ = new_new_n223__ & ~new_new_n554__;
  assign new_new_n6697__ = ~new_new_n471__ & ~new_new_n6695__;
  assign new_new_n6698__ = ~new_new_n6696__ & new_new_n6697__;
  assign new_new_n6699__ = ~new_new_n6692__ & ~new_new_n6693__;
  assign new_new_n6700__ = ~new_new_n523__ & new_new_n6699__;
  assign new_new_n6701__ = new_new_n4720__ & new_new_n6700__;
  assign new_new_n6702__ = ~new_new_n6691__ & new_new_n6698__;
  assign new_new_n6703__ = new_new_n6701__ & new_new_n6702__;
  assign new_new_n6704__ = new_new_n1026__ & new_new_n4294__;
  assign new_new_n6705__ = new_new_n6703__ & new_new_n6704__;
  assign new_new_n6706__ = new_new_n3531__ & new_new_n6705__;
  assign new_new_n6707__ = new_new_n209__ & new_new_n6706__;
  assign new_new_n6708__ = ~new_new_n6686__ & new_new_n6707__;
  assign new_new_n6709__ = new_new_n6686__ & ~new_new_n6707__;
  assign new_new_n6710__ = ~new_new_n6708__ & ~new_new_n6709__;
  assign new_new_n6711__ = new_new_n4702__ & ~new_new_n6600__;
  assign new_new_n6712__ = ~new_new_n6603__ & ~new_new_n6711__;
  assign new_new_n6713__ = new_new_n6710__ & new_new_n6712__;
  assign new_new_n6714__ = ~new_new_n6710__ & ~new_new_n6712__;
  assign po13 = ~new_new_n6713__ & ~new_new_n6714__;
  assign new_new_n6716__ = new_new_n6603__ & ~new_new_n6710__;
  assign new_new_n6717__ = new_new_n6600__ & new_new_n6710__;
  assign new_new_n6718__ = new_new_n4702__ & ~new_new_n6717__;
  assign new_new_n6719__ = ~new_new_n6716__ & ~new_new_n6718__;
  assign new_new_n6720__ = ~new_new_n6684__ & new_new_n6707__;
  assign new_new_n6721__ = ~new_new_n6685__ & ~new_new_n6720__;
  assign new_new_n6722__ = ~new_new_n6636__ & ~new_new_n6644__;
  assign new_new_n6723__ = ~new_new_n6635__ & ~new_new_n6722__;
  assign new_new_n6724__ = ~new_new_n6573__ & ~new_new_n6584__;
  assign new_new_n6725__ = ~new_new_n6560__ & ~new_new_n6724__;
  assign new_new_n6726__ = new_new_n6540__ & new_new_n6725__;
  assign new_new_n6727__ = ~new_new_n6540__ & ~new_new_n6725__;
  assign new_new_n6728__ = ~new_new_n6647__ & ~new_new_n6727__;
  assign new_new_n6729__ = new_new_n6560__ & ~new_new_n6584__;
  assign new_new_n6730__ = new_new_n6573__ & new_new_n6584__;
  assign new_new_n6731__ = new_new_n6647__ & ~new_new_n6730__;
  assign new_new_n6732__ = ~new_new_n6729__ & ~new_new_n6731__;
  assign new_new_n6733__ = ~new_new_n6541__ & new_new_n6732__;
  assign new_new_n6734__ = ~new_new_n6726__ & ~new_new_n6733__;
  assign new_new_n6735__ = ~new_new_n6728__ & new_new_n6734__;
  assign new_new_n6736__ = new_new_n6723__ & ~new_new_n6735__;
  assign new_new_n6737__ = ~new_new_n6723__ & new_new_n6735__;
  assign new_new_n6738__ = ~new_new_n6736__ & ~new_new_n6737__;
  assign new_new_n6739__ = ~new_new_n810__ & ~new_new_n5117__;
  assign new_new_n6740__ = ~new_new_n4432__ & ~new_new_n6739__;
  assign new_new_n6741__ = new_new_n4418__ & ~new_new_n6740__;
  assign new_new_n6742__ = ~new_new_n4418__ & new_new_n6740__;
  assign new_new_n6743__ = ~new_new_n6741__ & ~new_new_n6742__;
  assign new_new_n6744__ = new_new_n3069__ & ~new_new_n4857__;
  assign new_new_n6745__ = new_new_n4132__ & ~new_new_n4532__;
  assign new_new_n6746__ = ~new_new_n6744__ & ~new_new_n6745__;
  assign new_new_n6747__ = ~new_new_n2848__ & ~new_new_n6746__;
  assign new_new_n6748__ = new_new_n2848__ & ~new_new_n3072__;
  assign new_new_n6749__ = new_new_n4923__ & new_new_n6748__;
  assign new_new_n6750__ = ~new_new_n6747__ & ~new_new_n6749__;
  assign new_new_n6751__ = ~new_new_n437__ & new_new_n6750__;
  assign new_new_n6752__ = new_new_n437__ & ~new_new_n6750__;
  assign new_new_n6753__ = ~new_new_n6751__ & ~new_new_n6752__;
  assign new_new_n6754__ = new_new_n6743__ & new_new_n6753__;
  assign new_new_n6755__ = ~new_new_n6743__ & new_new_n6750__;
  assign new_new_n6756__ = ~new_new_n6754__ & ~new_new_n6755__;
  assign new_new_n6757__ = new_new_n6738__ & ~new_new_n6756__;
  assign new_new_n6758__ = ~new_new_n6738__ & new_new_n6756__;
  assign new_new_n6759__ = ~new_new_n6757__ & ~new_new_n6758__;
  assign new_new_n6760__ = ~new_new_n6721__ & ~new_new_n6759__;
  assign new_new_n6761__ = new_new_n6721__ & new_new_n6759__;
  assign new_new_n6762__ = ~new_new_n6760__ & ~new_new_n6761__;
  assign new_new_n6763__ = ~new_new_n445__ & ~new_new_n5079__;
  assign new_new_n6764__ = new_new_n100__ & ~new_new_n6106__;
  assign new_new_n6765__ = ~new_new_n185__ & ~new_new_n259__;
  assign new_new_n6766__ = ~new_new_n324__ & ~new_new_n709__;
  assign new_new_n6767__ = ~new_new_n2230__ & ~new_new_n4207__;
  assign new_new_n6768__ = new_new_n6766__ & new_new_n6767__;
  assign new_new_n6769__ = new_new_n241__ & new_new_n6765__;
  assign new_new_n6770__ = new_new_n6763__ & ~new_new_n6764__;
  assign new_new_n6771__ = new_new_n6769__ & new_new_n6770__;
  assign new_new_n6772__ = new_new_n975__ & new_new_n6768__;
  assign new_new_n6773__ = new_new_n6771__ & new_new_n6772__;
  assign new_new_n6774__ = new_new_n999__ & new_new_n6773__;
  assign new_new_n6775__ = new_new_n1447__ & new_new_n6774__;
  assign new_new_n6776__ = new_new_n2423__ & new_new_n6775__;
  assign new_new_n6777__ = ~new_new_n6762__ & new_new_n6776__;
  assign new_new_n6778__ = new_new_n6762__ & ~new_new_n6776__;
  assign new_new_n6779__ = ~new_new_n6777__ & ~new_new_n6778__;
  assign new_new_n6780__ = new_new_n6719__ & new_new_n6779__;
  assign new_new_n6781__ = ~new_new_n6719__ & ~new_new_n6779__;
  assign po14 = ~new_new_n6780__ & ~new_new_n6781__;
  assign new_new_n6783__ = new_new_n125__ & ~new_new_n4512__;
  assign new_new_n6784__ = ~new_new_n404__ & ~new_new_n6783__;
  assign new_new_n6785__ = new_new_n1123__ & new_new_n6784__;
  assign new_new_n6786__ = new_new_n1136__ & new_new_n6785__;
  assign new_new_n6787__ = new_new_n116__ & ~new_new_n275__;
  assign new_new_n6788__ = new_new_n110__ & new_new_n270__;
  assign new_new_n6789__ = new_new_n223__ & ~new_new_n6788__;
  assign new_new_n6790__ = ~new_new_n252__ & ~new_new_n475__;
  assign new_new_n6791__ = ~new_new_n957__ & new_new_n6790__;
  assign new_new_n6792__ = new_new_n112__ & ~new_new_n163__;
  assign new_new_n6793__ = ~new_new_n6787__ & ~new_new_n6789__;
  assign new_new_n6794__ = new_new_n6792__ & new_new_n6793__;
  assign new_new_n6795__ = new_new_n6763__ & new_new_n6791__;
  assign new_new_n6796__ = new_new_n6794__ & new_new_n6795__;
  assign new_new_n6797__ = new_new_n1048__ & new_new_n6504__;
  assign new_new_n6798__ = new_new_n6796__ & new_new_n6797__;
  assign new_new_n6799__ = new_new_n2242__ & new_new_n6798__;
  assign new_new_n6800__ = new_new_n6786__ & new_new_n6799__;
  assign new_new_n6801__ = ~new_new_n2846__ & new_new_n5122__;
  assign new_new_n6802__ = ~new_new_n2847__ & new_new_n3053__;
  assign new_new_n6803__ = ~new_new_n6801__ & new_new_n6802__;
  assign new_new_n6804__ = ~new_new_n2847__ & new_new_n5122__;
  assign new_new_n6805__ = ~new_new_n2846__ & new_new_n3063__;
  assign new_new_n6806__ = ~new_new_n6804__ & new_new_n6805__;
  assign new_new_n6807__ = ~new_new_n6803__ & ~new_new_n6806__;
  assign new_new_n6808__ = ~new_new_n4857__ & ~new_new_n6807__;
  assign new_new_n6809__ = ~new_new_n6736__ & ~new_new_n6756__;
  assign new_new_n6810__ = ~new_new_n6737__ & ~new_new_n6809__;
  assign new_new_n6811__ = new_new_n6808__ & ~new_new_n6810__;
  assign new_new_n6812__ = ~new_new_n437__ & ~new_new_n4532__;
  assign new_new_n6813__ = new_new_n4421__ & new_new_n6812__;
  assign new_new_n6814__ = new_new_n6811__ & new_new_n6813__;
  assign new_new_n6815__ = ~new_new_n4421__ & ~new_new_n6750__;
  assign new_new_n6816__ = ~new_new_n6751__ & ~new_new_n6815__;
  assign new_new_n6817__ = ~new_new_n810__ & ~new_new_n6638__;
  assign new_new_n6818__ = ~new_new_n6639__ & ~new_new_n6817__;
  assign new_new_n6819__ = ~new_new_n6816__ & ~new_new_n6818__;
  assign new_new_n6820__ = ~new_new_n437__ & new_new_n4421__;
  assign new_new_n6821__ = ~new_new_n6753__ & ~new_new_n6820__;
  assign new_new_n6822__ = ~new_new_n6819__ & ~new_new_n6821__;
  assign new_new_n6823__ = ~new_new_n4421__ & new_new_n4532__;
  assign new_new_n6824__ = new_new_n6811__ & ~new_new_n6823__;
  assign new_new_n6825__ = ~new_new_n6808__ & new_new_n6810__;
  assign new_new_n6826__ = ~new_new_n6820__ & ~new_new_n6825__;
  assign new_new_n6827__ = new_new_n4421__ & new_new_n6825__;
  assign new_new_n6828__ = ~new_new_n4532__ & ~new_new_n6827__;
  assign new_new_n6829__ = ~new_new_n437__ & ~new_new_n6828__;
  assign new_new_n6830__ = ~new_new_n6826__ & ~new_new_n6829__;
  assign new_new_n6831__ = ~new_new_n6824__ & ~new_new_n6830__;
  assign new_new_n6832__ = ~new_new_n6822__ & ~new_new_n6831__;
  assign new_new_n6833__ = new_new_n6810__ & ~new_new_n6813__;
  assign new_new_n6834__ = new_new_n4861__ & ~new_new_n6810__;
  assign new_new_n6835__ = ~new_new_n6808__ & ~new_new_n6833__;
  assign new_new_n6836__ = ~new_new_n6834__ & new_new_n6835__;
  assign new_new_n6837__ = new_new_n437__ & ~new_new_n6811__;
  assign new_new_n6838__ = ~new_new_n6825__ & new_new_n6837__;
  assign new_new_n6839__ = ~new_new_n6836__ & ~new_new_n6838__;
  assign new_new_n6840__ = new_new_n6822__ & ~new_new_n6839__;
  assign new_new_n6841__ = ~new_new_n6822__ & new_new_n6827__;
  assign new_new_n6842__ = ~new_new_n437__ & ~new_new_n6808__;
  assign new_new_n6843__ = ~new_new_n6822__ & new_new_n6842__;
  assign new_new_n6844__ = ~new_new_n6810__ & ~new_new_n6843__;
  assign new_new_n6845__ = ~new_new_n4421__ & ~new_new_n6825__;
  assign new_new_n6846__ = ~new_new_n6844__ & new_new_n6845__;
  assign new_new_n6847__ = ~new_new_n6841__ & ~new_new_n6846__;
  assign new_new_n6848__ = new_new_n4532__ & ~new_new_n6847__;
  assign new_new_n6849__ = ~new_new_n6814__ & ~new_new_n6840__;
  assign new_new_n6850__ = ~new_new_n6848__ & new_new_n6849__;
  assign new_new_n6851__ = ~new_new_n6832__ & new_new_n6850__;
  assign new_new_n6852__ = new_new_n6800__ & ~new_new_n6851__;
  assign new_new_n6853__ = ~new_new_n6800__ & new_new_n6851__;
  assign new_new_n6854__ = ~new_new_n6852__ & ~new_new_n6853__;
  assign new_new_n6855__ = ~new_new_n6761__ & new_new_n6776__;
  assign new_new_n6856__ = ~new_new_n6760__ & ~new_new_n6855__;
  assign new_new_n6857__ = new_new_n6854__ & new_new_n6856__;
  assign new_new_n6858__ = ~new_new_n6854__ & ~new_new_n6856__;
  assign new_new_n6859__ = ~new_new_n6857__ & ~new_new_n6858__;
  assign new_new_n6860__ = ~new_new_n4702__ & ~new_new_n6716__;
  assign new_new_n6861__ = ~new_new_n6718__ & new_new_n6779__;
  assign new_new_n6862__ = ~new_new_n6860__ & ~new_new_n6861__;
  assign new_new_n6863__ = ~new_new_n6859__ & new_new_n6862__;
  assign new_new_n6864__ = new_new_n6859__ & ~new_new_n6862__;
  assign po15 = ~new_new_n6863__ & ~new_new_n6864__;
  assign new_new_n6866__ = new_new_n6717__ & new_new_n6779__;
  assign new_new_n6867__ = new_new_n6859__ & new_new_n6866__;
  assign new_new_n6868__ = ~new_new_n4702__ & ~new_new_n6863__;
  assign new_new_n6869__ = ~new_new_n6867__ & ~new_new_n6868__;
  assign new_new_n6870__ = new_new_n6808__ & new_new_n6823__;
  assign new_new_n6871__ = ~new_new_n4532__ & ~new_new_n4829__;
  assign new_new_n6872__ = new_new_n4857__ & ~new_new_n6871__;
  assign new_new_n6873__ = ~new_new_n6870__ & ~new_new_n6872__;
  assign new_new_n6874__ = ~new_new_n437__ & ~new_new_n6873__;
  assign new_new_n6875__ = ~new_new_n4412__ & new_new_n4532__;
  assign new_new_n6876__ = ~new_new_n4420__ & ~new_new_n4550__;
  assign new_new_n6877__ = ~new_new_n6875__ & new_new_n6876__;
  assign new_new_n6878__ = ~new_new_n4857__ & new_new_n6877__;
  assign new_new_n6879__ = ~new_new_n437__ & ~new_new_n4863__;
  assign new_new_n6880__ = ~new_new_n6878__ & new_new_n6879__;
  assign new_new_n6881__ = ~new_new_n6808__ & ~new_new_n6880__;
  assign new_new_n6882__ = ~new_new_n6874__ & ~new_new_n6881__;
  assign new_new_n6883__ = new_new_n6810__ & new_new_n6822__;
  assign new_new_n6884__ = ~new_new_n4532__ & ~new_new_n6808__;
  assign new_new_n6885__ = new_new_n4421__ & ~new_new_n6884__;
  assign new_new_n6886__ = new_new_n6812__ & new_new_n6885__;
  assign new_new_n6887__ = new_new_n6810__ & ~new_new_n6870__;
  assign new_new_n6888__ = ~new_new_n6822__ & ~new_new_n6887__;
  assign new_new_n6889__ = ~new_new_n437__ & ~new_new_n4859__;
  assign new_new_n6890__ = ~new_new_n6885__ & new_new_n6889__;
  assign new_new_n6891__ = ~new_new_n6808__ & ~new_new_n6890__;
  assign new_new_n6892__ = ~new_new_n6886__ & ~new_new_n6891__;
  assign new_new_n6893__ = ~new_new_n6888__ & new_new_n6892__;
  assign new_new_n6894__ = ~new_new_n6883__ & ~new_new_n6893__;
  assign new_new_n6895__ = ~new_new_n6882__ & ~new_new_n6894__;
  assign new_new_n6896__ = new_new_n6882__ & new_new_n6894__;
  assign new_new_n6897__ = ~new_new_n6895__ & ~new_new_n6896__;
  assign new_new_n6898__ = new_new_n54__ & new_new_n124__;
  assign new_new_n6899__ = new_new_n149__ & ~new_new_n6898__;
  assign new_new_n6900__ = new_new_n223__ & ~new_new_n2471__;
  assign new_new_n6901__ = new_new_n125__ & ~new_new_n581__;
  assign new_new_n6902__ = ~new_new_n376__ & ~new_new_n957__;
  assign new_new_n6903__ = ~new_new_n2461__ & ~new_new_n6899__;
  assign new_new_n6904__ = ~new_new_n6901__ & new_new_n6903__;
  assign new_new_n6905__ = new_new_n6902__ & new_new_n6904__;
  assign new_new_n6906__ = new_new_n4471__ & new_new_n6698__;
  assign new_new_n6907__ = ~new_new_n6900__ & new_new_n6906__;
  assign new_new_n6908__ = new_new_n6905__ & new_new_n6907__;
  assign new_new_n6909__ = new_new_n285__ & new_new_n6908__;
  assign new_new_n6910__ = new_new_n2566__ & new_new_n6909__;
  assign new_new_n6911__ = ~new_new_n6897__ & ~new_new_n6910__;
  assign new_new_n6912__ = new_new_n6897__ & new_new_n6910__;
  assign new_new_n6913__ = ~new_new_n6911__ & ~new_new_n6912__;
  assign new_new_n6914__ = ~new_new_n6853__ & ~new_new_n6856__;
  assign new_new_n6915__ = ~new_new_n6852__ & ~new_new_n6914__;
  assign new_new_n6916__ = new_new_n6913__ & ~new_new_n6915__;
  assign new_new_n6917__ = ~new_new_n6913__ & new_new_n6915__;
  assign new_new_n6918__ = ~new_new_n6916__ & ~new_new_n6917__;
  assign new_new_n6919__ = ~new_new_n6869__ & ~new_new_n6918__;
  assign new_new_n6920__ = new_new_n6869__ & new_new_n6918__;
  assign po16 = ~new_new_n6919__ & ~new_new_n6920__;
  assign new_new_n6922__ = ~new_new_n6911__ & ~new_new_n6915__;
  assign new_new_n6923__ = ~new_new_n6912__ & ~new_new_n6922__;
  assign new_new_n6924__ = new_new_n81__ & new_new_n522__;
  assign new_new_n6925__ = ~new_new_n365__ & ~new_new_n6924__;
  assign new_new_n6926__ = ~new_new_n176__ & ~new_new_n409__;
  assign new_new_n6927__ = ~new_new_n386__ & new_new_n6926__;
  assign new_new_n6928__ = ~new_new_n971__ & new_new_n3616__;
  assign new_new_n6929__ = new_new_n6927__ & new_new_n6928__;
  assign new_new_n6930__ = ~new_new_n363__ & ~new_new_n523__;
  assign new_new_n6931__ = new_new_n526__ & new_new_n871__;
  assign new_new_n6932__ = ~new_new_n6925__ & new_new_n6931__;
  assign new_new_n6933__ = new_new_n6929__ & new_new_n6930__;
  assign new_new_n6934__ = new_new_n6932__ & new_new_n6933__;
  assign new_new_n6935__ = new_new_n580__ & new_new_n6934__;
  assign new_new_n6936__ = new_new_n3711__ & new_new_n6935__;
  assign new_new_n6937__ = ~new_new_n6923__ & new_new_n6936__;
  assign new_new_n6938__ = new_new_n6923__ & ~new_new_n6936__;
  assign new_new_n6939__ = ~new_new_n6937__ & ~new_new_n6938__;
  assign new_new_n6940__ = new_new_n6867__ & ~new_new_n6918__;
  assign new_new_n6941__ = new_new_n6716__ & ~new_new_n6779__;
  assign new_new_n6942__ = ~new_new_n6859__ & new_new_n6941__;
  assign new_new_n6943__ = new_new_n6918__ & new_new_n6942__;
  assign new_new_n6944__ = ~new_new_n4702__ & ~new_new_n6943__;
  assign new_new_n6945__ = ~new_new_n6940__ & ~new_new_n6944__;
  assign new_new_n6946__ = new_new_n6939__ & new_new_n6945__;
  assign new_new_n6947__ = ~new_new_n6939__ & ~new_new_n6945__;
  assign po17 = new_new_n6946__ | new_new_n6947__;
  assign new_new_n6949__ = ~new_new_n6923__ & new_new_n6940__;
  assign new_new_n6950__ = ~new_new_n6937__ & new_new_n6943__;
  assign new_new_n6951__ = ~new_new_n6949__ & ~new_new_n6950__;
  assign new_new_n6952__ = ~new_new_n176__ & ~new_new_n328__;
  assign new_new_n6953__ = ~new_new_n384__ & new_new_n6952__;
  assign new_new_n6954__ = ~new_new_n617__ & ~new_new_n991__;
  assign new_new_n6955__ = new_new_n6953__ & new_new_n6954__;
  assign new_new_n6956__ = ~new_new_n694__ & new_new_n6955__;
  assign new_new_n6957__ = new_new_n968__ & new_new_n1056__;
  assign new_new_n6958__ = new_new_n3521__ & new_new_n6957__;
  assign new_new_n6959__ = new_new_n1103__ & new_new_n6956__;
  assign new_new_n6960__ = new_new_n6958__ & new_new_n6959__;
  assign new_new_n6961__ = new_new_n538__ & new_new_n6960__;
  assign new_new_n6962__ = new_new_n4287__ & new_new_n6961__;
  assign new_new_n6963__ = ~new_new_n6951__ & new_new_n6962__;
  assign new_new_n6964__ = new_new_n6938__ & ~new_new_n6962__;
  assign new_new_n6965__ = ~new_new_n6943__ & new_new_n6964__;
  assign new_new_n6966__ = ~new_new_n6963__ & ~new_new_n6965__;
  assign new_new_n6967__ = ~new_new_n4702__ & ~new_new_n6966__;
  assign new_new_n6968__ = ~new_new_n6944__ & new_new_n6962__;
  assign new_new_n6969__ = ~new_new_n6938__ & ~new_new_n6940__;
  assign new_new_n6970__ = ~new_new_n4702__ & ~new_new_n6962__;
  assign new_new_n6971__ = new_new_n6969__ & ~new_new_n6970__;
  assign new_new_n6972__ = ~new_new_n6968__ & new_new_n6971__;
  assign new_new_n6973__ = new_new_n6923__ & new_new_n6962__;
  assign new_new_n6974__ = new_new_n6940__ & new_new_n6973__;
  assign new_new_n6975__ = ~new_new_n6923__ & ~new_new_n6962__;
  assign new_new_n6976__ = new_new_n6943__ & new_new_n6975__;
  assign new_new_n6977__ = ~new_new_n6974__ & ~new_new_n6976__;
  assign new_new_n6978__ = new_new_n6936__ & ~new_new_n6977__;
  assign new_new_n6979__ = ~new_new_n6936__ & new_new_n6962__;
  assign new_new_n6980__ = new_new_n6949__ & new_new_n6979__;
  assign new_new_n6981__ = ~new_new_n6973__ & ~new_new_n6975__;
  assign new_new_n6982__ = new_new_n4702__ & ~new_new_n6939__;
  assign new_new_n6983__ = ~new_new_n6981__ & new_new_n6982__;
  assign new_new_n6984__ = ~new_new_n6972__ & ~new_new_n6980__;
  assign new_new_n6985__ = ~new_new_n6978__ & ~new_new_n6983__;
  assign new_new_n6986__ = new_new_n6984__ & new_new_n6985__;
  assign po18 = new_new_n6967__ | ~new_new_n6986__;
  assign new_new_n6988__ = new_new_n6940__ & ~new_new_n6962__;
  assign new_new_n6989__ = new_new_n6939__ & new_new_n6988__;
  assign new_new_n6990__ = ~new_new_n6939__ & new_new_n6943__;
  assign new_new_n6991__ = new_new_n6981__ & new_new_n6990__;
  assign new_new_n6992__ = ~new_new_n6989__ & ~new_new_n6991__;
  assign new_new_n6993__ = ~new_new_n4702__ & new_new_n6992__;
  assign new_new_n6994__ = new_new_n174__ & new_new_n1021__;
  assign new_new_n6995__ = new_new_n125__ & ~new_new_n6994__;
  assign new_new_n6996__ = new_new_n195__ & ~new_new_n4512__;
  assign new_new_n6997__ = ~new_new_n383__ & ~new_new_n2679__;
  assign new_new_n6998__ = ~new_new_n690__ & new_new_n6997__;
  assign new_new_n6999__ = ~new_new_n6996__ & new_new_n6998__;
  assign new_new_n7000__ = ~new_new_n6995__ & new_new_n6999__;
  assign new_new_n7001__ = new_new_n5593__ & new_new_n7000__;
  assign new_new_n7002__ = new_new_n3683__ & new_new_n7001__;
  assign new_new_n7003__ = new_new_n941__ & new_new_n7002__;
  assign new_new_n7004__ = new_new_n6786__ & new_new_n7003__;
  assign new_new_n7005__ = ~new_new_n6937__ & ~new_new_n6962__;
  assign new_new_n7006__ = ~new_new_n6969__ & new_new_n7005__;
  assign new_new_n7007__ = ~new_new_n7004__ & new_new_n7006__;
  assign new_new_n7008__ = new_new_n7004__ & ~new_new_n7006__;
  assign new_new_n7009__ = ~new_new_n7007__ & ~new_new_n7008__;
  assign new_new_n7010__ = ~new_new_n6993__ & new_new_n7009__;
  assign new_new_n7011__ = new_new_n6993__ & ~new_new_n7009__;
  assign po19 = new_new_n7010__ | new_new_n7011__;
  assign new_new_n7013__ = ~new_new_n100__ & ~new_new_n195__;
  assign new_new_n7014__ = ~new_new_n3712__ & ~new_new_n7013__;
  assign new_new_n7015__ = ~new_new_n267__ & ~new_new_n560__;
  assign new_new_n7016__ = ~new_new_n321__ & new_new_n7015__;
  assign new_new_n7017__ = ~new_new_n617__ & ~new_new_n2230__;
  assign new_new_n7018__ = ~new_new_n2700__ & new_new_n7017__;
  assign new_new_n7019__ = ~new_new_n2245__ & new_new_n7016__;
  assign new_new_n7020__ = ~new_new_n7014__ & new_new_n7019__;
  assign new_new_n7021__ = ~new_new_n795__ & new_new_n7018__;
  assign new_new_n7022__ = new_new_n7020__ & new_new_n7021__;
  assign new_new_n7023__ = new_new_n988__ & new_new_n7022__;
  assign new_new_n7024__ = new_new_n6112__ & new_new_n7023__;
  assign new_new_n7025__ = ~new_new_n7006__ & new_new_n7024__;
  assign new_new_n7026__ = new_new_n7007__ & ~new_new_n7024__;
  assign new_new_n7027__ = ~new_new_n7025__ & ~new_new_n7026__;
  assign new_new_n7028__ = new_new_n6992__ & ~new_new_n7027__;
  assign new_new_n7029__ = new_new_n7009__ & new_new_n7024__;
  assign new_new_n7030__ = ~new_new_n7028__ & ~new_new_n7029__;
  assign new_new_n7031__ = ~new_new_n4702__ & ~new_new_n7030__;
  assign new_new_n7032__ = ~new_new_n7007__ & new_new_n7024__;
  assign new_new_n7033__ = new_new_n4702__ & ~new_new_n7026__;
  assign new_new_n7034__ = ~new_new_n7032__ & new_new_n7033__;
  assign new_new_n7035__ = ~new_new_n7008__ & ~new_new_n7024__;
  assign new_new_n7036__ = ~new_new_n6992__ & ~new_new_n7032__;
  assign new_new_n7037__ = ~new_new_n7035__ & new_new_n7036__;
  assign new_new_n7038__ = ~new_new_n7034__ & ~new_new_n7037__;
  assign po20 = new_new_n7031__ | ~new_new_n7038__;
  assign new_new_n7040__ = ~new_new_n323__ & new_new_n396__;
  assign new_new_n7041__ = new_new_n99__ & new_new_n115__;
  assign new_new_n7042__ = ~new_new_n410__ & new_new_n7041__;
  assign new_new_n7043__ = ~new_new_n7040__ & ~new_new_n7042__;
  assign new_new_n7044__ = ~new_new_n594__ & ~new_new_n7043__;
  assign new_new_n7045__ = new_new_n684__ & new_new_n7044__;
  assign new_new_n7046__ = new_new_n796__ & new_new_n7045__;
  assign new_new_n7047__ = new_new_n648__ & new_new_n7046__;
  assign new_new_n7048__ = new_new_n7026__ & ~new_new_n7047__;
  assign new_new_n7049__ = ~new_new_n7006__ & new_new_n7047__;
  assign new_new_n7050__ = ~new_new_n7048__ & ~new_new_n7049__;
  assign new_new_n7051__ = new_new_n6992__ & ~new_new_n7050__;
  assign new_new_n7052__ = ~new_new_n7026__ & new_new_n7047__;
  assign new_new_n7053__ = new_new_n7008__ & new_new_n7024__;
  assign new_new_n7054__ = new_new_n7052__ & ~new_new_n7053__;
  assign new_new_n7055__ = ~new_new_n7051__ & ~new_new_n7054__;
  assign new_new_n7056__ = ~new_new_n4702__ & ~new_new_n7055__;
  assign new_new_n7057__ = new_new_n4702__ & ~new_new_n7048__;
  assign new_new_n7058__ = ~new_new_n7047__ & ~new_new_n7053__;
  assign new_new_n7059__ = ~new_new_n6992__ & ~new_new_n7058__;
  assign new_new_n7060__ = ~new_new_n7057__ & ~new_new_n7059__;
  assign new_new_n7061__ = ~new_new_n7052__ & ~new_new_n7060__;
  assign po21 = new_new_n7056__ | new_new_n7061__;
  assign new_new_n7063__ = new_new_n792__ & ~new_new_n803__;
  assign new_new_n7064__ = ~new_new_n7048__ & ~new_new_n7063__;
  assign new_new_n7065__ = new_new_n7048__ & new_new_n7063__;
  assign new_new_n7066__ = ~new_new_n7064__ & ~new_new_n7065__;
  assign new_new_n7067__ = ~new_new_n6992__ & new_new_n7047__;
  assign new_new_n7068__ = new_new_n7053__ & new_new_n7067__;
  assign new_new_n7069__ = ~new_new_n4702__ & ~new_new_n7068__;
  assign new_new_n7070__ = ~new_new_n6992__ & new_new_n7048__;
  assign new_new_n7071__ = new_new_n7069__ & ~new_new_n7070__;
  assign new_new_n7072__ = new_new_n7066__ & new_new_n7071__;
  assign new_new_n7073__ = new_new_n7006__ & new_new_n7063__;
  assign new_new_n7074__ = ~new_new_n7064__ & ~new_new_n7073__;
  assign new_new_n7075__ = ~new_new_n7068__ & ~new_new_n7070__;
  assign new_new_n7076__ = ~new_new_n7074__ & ~new_new_n7075__;
  assign new_new_n7077__ = new_new_n4702__ & ~new_new_n7066__;
  assign new_new_n7078__ = ~new_new_n7076__ & ~new_new_n7077__;
  assign po22 = new_new_n7072__ | ~new_new_n7078__;
  assign new_new_n7080__ = new_new_n118__ & new_new_n120__;
  assign new_new_n7081__ = new_new_n7057__ & ~new_new_n7080__;
  assign new_new_n7082__ = new_new_n7063__ & ~new_new_n7080__;
  assign new_new_n7083__ = ~new_new_n7069__ & new_new_n7082__;
  assign new_new_n7084__ = ~pi21 & pi23;
  assign new_new_n7085__ = new_new_n120__ & new_new_n7084__;
  assign new_new_n7086__ = ~new_new_n7063__ & ~new_new_n7085__;
  assign new_new_n7087__ = new_new_n7048__ & new_new_n7086__;
  assign new_new_n7088__ = new_new_n7071__ & new_new_n7087__;
  assign new_new_n7089__ = ~new_new_n7081__ & ~new_new_n7083__;
  assign po23 = ~new_new_n7088__ & new_new_n7089__;
  assign new_new_n7091__ = new_new_n7063__ & ~new_new_n7085__;
  assign new_new_n7092__ = new_new_n7068__ & new_new_n7091__;
  assign po24 = ~new_new_n4702__ & ~new_new_n7092__;
endmodule


