// Benchmark "log2" written by ABC on Wed Jul 13 18:49:08 2022

module log2 ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31;
  wire new_new_n65__, new_new_n66__, new_new_n67__, new_new_n68__,
    new_new_n69__, new_new_n70__, new_new_n71__, new_new_n72__,
    new_new_n73__, new_new_n74__, new_new_n75__, new_new_n76__,
    new_new_n77__, new_new_n78__, new_new_n79__, new_new_n80__,
    new_new_n81__, new_new_n82__, new_new_n83__, new_new_n84__,
    new_new_n85__, new_new_n86__, new_new_n87__, new_new_n88__,
    new_new_n89__, new_new_n90__, new_new_n91__, new_new_n92__,
    new_new_n93__, new_new_n94__, new_new_n95__, new_new_n96__,
    new_new_n97__, new_new_n98__, new_new_n99__, new_new_n100__,
    new_new_n101__, new_new_n102__, new_new_n103__, new_new_n104__,
    new_new_n105__, new_new_n106__, new_new_n107__, new_new_n108__,
    new_new_n109__, new_new_n110__, new_new_n111__, new_new_n112__,
    new_new_n113__, new_new_n114__, new_new_n115__, new_new_n116__,
    new_new_n117__, new_new_n118__, new_new_n119__, new_new_n120__,
    new_new_n121__, new_new_n122__, new_new_n123__, new_new_n124__,
    new_new_n125__, new_new_n126__, new_new_n127__, new_new_n128__,
    new_new_n129__, new_new_n130__, new_new_n131__, new_new_n132__,
    new_new_n133__, new_new_n134__, new_new_n135__, new_new_n136__,
    new_new_n137__, new_new_n138__, new_new_n139__, new_new_n140__,
    new_new_n141__, new_new_n142__, new_new_n143__, new_new_n144__,
    new_new_n145__, new_new_n146__, new_new_n147__, new_new_n148__,
    new_new_n149__, new_new_n150__, new_new_n151__, new_new_n152__,
    new_new_n153__, new_new_n154__, new_new_n155__, new_new_n156__,
    new_new_n157__, new_new_n158__, new_new_n159__, new_new_n160__,
    new_new_n161__, new_new_n162__, new_new_n163__, new_new_n164__,
    new_new_n165__, new_new_n166__, new_new_n167__, new_new_n168__,
    new_new_n169__, new_new_n170__, new_new_n171__, new_new_n172__,
    new_new_n173__, new_new_n174__, new_new_n175__, new_new_n176__,
    new_new_n177__, new_new_n178__, new_new_n179__, new_new_n180__,
    new_new_n181__, new_new_n182__, new_new_n183__, new_new_n184__,
    new_new_n185__, new_new_n186__, new_new_n187__, new_new_n188__,
    new_new_n189__, new_new_n190__, new_new_n191__, new_new_n192__,
    new_new_n193__, new_new_n194__, new_new_n195__, new_new_n196__,
    new_new_n197__, new_new_n198__, new_new_n199__, new_new_n200__,
    new_new_n201__, new_new_n202__, new_new_n203__, new_new_n204__,
    new_new_n205__, new_new_n206__, new_new_n207__, new_new_n208__,
    new_new_n209__, new_new_n210__, new_new_n211__, new_new_n212__,
    new_new_n213__, new_new_n214__, new_new_n215__, new_new_n216__,
    new_new_n217__, new_new_n218__, new_new_n219__, new_new_n220__,
    new_new_n221__, new_new_n222__, new_new_n223__, new_new_n224__,
    new_new_n225__, new_new_n226__, new_new_n227__, new_new_n228__,
    new_new_n229__, new_new_n230__, new_new_n231__, new_new_n232__,
    new_new_n233__, new_new_n234__, new_new_n235__, new_new_n236__,
    new_new_n237__, new_new_n238__, new_new_n239__, new_new_n240__,
    new_new_n241__, new_new_n242__, new_new_n243__, new_new_n244__,
    new_new_n245__, new_new_n246__, new_new_n247__, new_new_n248__,
    new_new_n249__, new_new_n250__, new_new_n251__, new_new_n252__,
    new_new_n253__, new_new_n254__, new_new_n255__, new_new_n256__,
    new_new_n257__, new_new_n258__, new_new_n259__, new_new_n260__,
    new_new_n261__, new_new_n262__, new_new_n263__, new_new_n264__,
    new_new_n265__, new_new_n266__, new_new_n267__, new_new_n268__,
    new_new_n269__, new_new_n270__, new_new_n271__, new_new_n272__,
    new_new_n273__, new_new_n274__, new_new_n275__, new_new_n276__,
    new_new_n277__, new_new_n278__, new_new_n279__, new_new_n280__,
    new_new_n281__, new_new_n282__, new_new_n283__, new_new_n284__,
    new_new_n285__, new_new_n286__, new_new_n287__, new_new_n288__,
    new_new_n289__, new_new_n290__, new_new_n291__, new_new_n292__,
    new_new_n293__, new_new_n294__, new_new_n295__, new_new_n296__,
    new_new_n297__, new_new_n298__, new_new_n299__, new_new_n300__,
    new_new_n301__, new_new_n302__, new_new_n303__, new_new_n304__,
    new_new_n305__, new_new_n306__, new_new_n307__, new_new_n308__,
    new_new_n309__, new_new_n310__, new_new_n311__, new_new_n312__,
    new_new_n313__, new_new_n314__, new_new_n315__, new_new_n316__,
    new_new_n317__, new_new_n318__, new_new_n319__, new_new_n320__,
    new_new_n321__, new_new_n322__, new_new_n323__, new_new_n324__,
    new_new_n325__, new_new_n326__, new_new_n327__, new_new_n328__,
    new_new_n329__, new_new_n330__, new_new_n331__, new_new_n332__,
    new_new_n333__, new_new_n334__, new_new_n335__, new_new_n336__,
    new_new_n337__, new_new_n338__, new_new_n339__, new_new_n340__,
    new_new_n341__, new_new_n342__, new_new_n343__, new_new_n344__,
    new_new_n345__, new_new_n346__, new_new_n347__, new_new_n348__,
    new_new_n349__, new_new_n350__, new_new_n351__, new_new_n352__,
    new_new_n353__, new_new_n354__, new_new_n355__, new_new_n356__,
    new_new_n357__, new_new_n358__, new_new_n359__, new_new_n360__,
    new_new_n361__, new_new_n362__, new_new_n363__, new_new_n364__,
    new_new_n365__, new_new_n366__, new_new_n367__, new_new_n368__,
    new_new_n369__, new_new_n370__, new_new_n371__, new_new_n372__,
    new_new_n373__, new_new_n374__, new_new_n375__, new_new_n376__,
    new_new_n377__, new_new_n378__, new_new_n379__, new_new_n380__,
    new_new_n381__, new_new_n382__, new_new_n383__, new_new_n384__,
    new_new_n385__, new_new_n386__, new_new_n387__, new_new_n388__,
    new_new_n389__, new_new_n390__, new_new_n391__, new_new_n392__,
    new_new_n393__, new_new_n394__, new_new_n395__, new_new_n396__,
    new_new_n397__, new_new_n398__, new_new_n399__, new_new_n400__,
    new_new_n401__, new_new_n402__, new_new_n403__, new_new_n404__,
    new_new_n405__, new_new_n406__, new_new_n407__, new_new_n408__,
    new_new_n409__, new_new_n410__, new_new_n411__, new_new_n412__,
    new_new_n413__, new_new_n414__, new_new_n415__, new_new_n416__,
    new_new_n417__, new_new_n418__, new_new_n419__, new_new_n420__,
    new_new_n421__, new_new_n422__, new_new_n423__, new_new_n424__,
    new_new_n425__, new_new_n426__, new_new_n427__, new_new_n428__,
    new_new_n429__, new_new_n430__, new_new_n431__, new_new_n432__,
    new_new_n433__, new_new_n434__, new_new_n435__, new_new_n436__,
    new_new_n437__, new_new_n438__, new_new_n439__, new_new_n440__,
    new_new_n441__, new_new_n442__, new_new_n443__, new_new_n444__,
    new_new_n445__, new_new_n446__, new_new_n447__, new_new_n448__,
    new_new_n449__, new_new_n450__, new_new_n451__, new_new_n452__,
    new_new_n453__, new_new_n454__, new_new_n455__, new_new_n456__,
    new_new_n457__, new_new_n458__, new_new_n459__, new_new_n460__,
    new_new_n461__, new_new_n462__, new_new_n463__, new_new_n464__,
    new_new_n465__, new_new_n466__, new_new_n467__, new_new_n468__,
    new_new_n469__, new_new_n470__, new_new_n471__, new_new_n472__,
    new_new_n473__, new_new_n474__, new_new_n475__, new_new_n476__,
    new_new_n477__, new_new_n478__, new_new_n479__, new_new_n480__,
    new_new_n481__, new_new_n482__, new_new_n483__, new_new_n484__,
    new_new_n485__, new_new_n486__, new_new_n487__, new_new_n488__,
    new_new_n489__, new_new_n490__, new_new_n491__, new_new_n492__,
    new_new_n493__, new_new_n494__, new_new_n495__, new_new_n496__,
    new_new_n497__, new_new_n498__, new_new_n499__, new_new_n500__,
    new_new_n501__, new_new_n502__, new_new_n503__, new_new_n504__,
    new_new_n505__, new_new_n506__, new_new_n507__, new_new_n508__,
    new_new_n509__, new_new_n510__, new_new_n511__, new_new_n512__,
    new_new_n513__, new_new_n514__, new_new_n515__, new_new_n516__,
    new_new_n517__, new_new_n518__, new_new_n519__, new_new_n520__,
    new_new_n521__, new_new_n522__, new_new_n523__, new_new_n524__,
    new_new_n525__, new_new_n526__, new_new_n527__, new_new_n528__,
    new_new_n529__, new_new_n530__, new_new_n531__, new_new_n532__,
    new_new_n533__, new_new_n534__, new_new_n535__, new_new_n536__,
    new_new_n537__, new_new_n538__, new_new_n539__, new_new_n540__,
    new_new_n541__, new_new_n542__, new_new_n543__, new_new_n544__,
    new_new_n545__, new_new_n546__, new_new_n547__, new_new_n548__,
    new_new_n549__, new_new_n550__, new_new_n551__, new_new_n552__,
    new_new_n553__, new_new_n554__, new_new_n555__, new_new_n556__,
    new_new_n557__, new_new_n558__, new_new_n559__, new_new_n560__,
    new_new_n561__, new_new_n562__, new_new_n563__, new_new_n564__,
    new_new_n565__, new_new_n566__, new_new_n567__, new_new_n568__,
    new_new_n569__, new_new_n570__, new_new_n571__, new_new_n572__,
    new_new_n573__, new_new_n574__, new_new_n575__, new_new_n576__,
    new_new_n577__, new_new_n578__, new_new_n579__, new_new_n580__,
    new_new_n581__, new_new_n582__, new_new_n583__, new_new_n584__,
    new_new_n585__, new_new_n586__, new_new_n587__, new_new_n588__,
    new_new_n589__, new_new_n590__, new_new_n591__, new_new_n592__,
    new_new_n593__, new_new_n594__, new_new_n595__, new_new_n596__,
    new_new_n597__, new_new_n598__, new_new_n599__, new_new_n600__,
    new_new_n601__, new_new_n602__, new_new_n603__, new_new_n604__,
    new_new_n605__, new_new_n606__, new_new_n607__, new_new_n608__,
    new_new_n609__, new_new_n610__, new_new_n611__, new_new_n612__,
    new_new_n613__, new_new_n614__, new_new_n615__, new_new_n616__,
    new_new_n617__, new_new_n618__, new_new_n619__, new_new_n620__,
    new_new_n621__, new_new_n622__, new_new_n623__, new_new_n624__,
    new_new_n625__, new_new_n626__, new_new_n627__, new_new_n628__,
    new_new_n629__, new_new_n630__, new_new_n631__, new_new_n632__,
    new_new_n633__, new_new_n634__, new_new_n635__, new_new_n636__,
    new_new_n637__, new_new_n638__, new_new_n639__, new_new_n640__,
    new_new_n641__, new_new_n642__, new_new_n643__, new_new_n644__,
    new_new_n645__, new_new_n646__, new_new_n647__, new_new_n648__,
    new_new_n649__, new_new_n650__, new_new_n651__, new_new_n652__,
    new_new_n653__, new_new_n654__, new_new_n655__, new_new_n656__,
    new_new_n657__, new_new_n658__, new_new_n659__, new_new_n660__,
    new_new_n661__, new_new_n662__, new_new_n663__, new_new_n664__,
    new_new_n665__, new_new_n666__, new_new_n667__, new_new_n668__,
    new_new_n669__, new_new_n670__, new_new_n671__, new_new_n672__,
    new_new_n673__, new_new_n674__, new_new_n675__, new_new_n676__,
    new_new_n677__, new_new_n678__, new_new_n679__, new_new_n680__,
    new_new_n681__, new_new_n682__, new_new_n683__, new_new_n684__,
    new_new_n685__, new_new_n686__, new_new_n687__, new_new_n688__,
    new_new_n689__, new_new_n690__, new_new_n691__, new_new_n692__,
    new_new_n693__, new_new_n694__, new_new_n695__, new_new_n696__,
    new_new_n697__, new_new_n698__, new_new_n699__, new_new_n700__,
    new_new_n701__, new_new_n702__, new_new_n703__, new_new_n704__,
    new_new_n705__, new_new_n706__, new_new_n707__, new_new_n708__,
    new_new_n709__, new_new_n710__, new_new_n711__, new_new_n712__,
    new_new_n713__, new_new_n714__, new_new_n715__, new_new_n716__,
    new_new_n717__, new_new_n718__, new_new_n719__, new_new_n720__,
    new_new_n721__, new_new_n722__, new_new_n723__, new_new_n724__,
    new_new_n725__, new_new_n726__, new_new_n727__, new_new_n728__,
    new_new_n729__, new_new_n730__, new_new_n731__, new_new_n732__,
    new_new_n733__, new_new_n734__, new_new_n735__, new_new_n736__,
    new_new_n737__, new_new_n738__, new_new_n739__, new_new_n740__,
    new_new_n741__, new_new_n742__, new_new_n743__, new_new_n744__,
    new_new_n745__, new_new_n746__, new_new_n747__, new_new_n748__,
    new_new_n749__, new_new_n750__, new_new_n751__, new_new_n752__,
    new_new_n753__, new_new_n754__, new_new_n755__, new_new_n756__,
    new_new_n757__, new_new_n758__, new_new_n759__, new_new_n760__,
    new_new_n761__, new_new_n762__, new_new_n763__, new_new_n764__,
    new_new_n765__, new_new_n766__, new_new_n767__, new_new_n768__,
    new_new_n769__, new_new_n770__, new_new_n771__, new_new_n772__,
    new_new_n773__, new_new_n774__, new_new_n775__, new_new_n776__,
    new_new_n777__, new_new_n778__, new_new_n779__, new_new_n780__,
    new_new_n781__, new_new_n782__, new_new_n783__, new_new_n784__,
    new_new_n785__, new_new_n786__, new_new_n787__, new_new_n788__,
    new_new_n789__, new_new_n790__, new_new_n791__, new_new_n792__,
    new_new_n793__, new_new_n794__, new_new_n795__, new_new_n796__,
    new_new_n797__, new_new_n798__, new_new_n799__, new_new_n800__,
    new_new_n801__, new_new_n802__, new_new_n803__, new_new_n804__,
    new_new_n805__, new_new_n806__, new_new_n807__, new_new_n808__,
    new_new_n809__, new_new_n810__, new_new_n811__, new_new_n812__,
    new_new_n813__, new_new_n814__, new_new_n815__, new_new_n816__,
    new_new_n817__, new_new_n818__, new_new_n819__, new_new_n820__,
    new_new_n821__, new_new_n822__, new_new_n823__, new_new_n824__,
    new_new_n825__, new_new_n826__, new_new_n827__, new_new_n828__,
    new_new_n829__, new_new_n830__, new_new_n831__, new_new_n832__,
    new_new_n833__, new_new_n834__, new_new_n835__, new_new_n836__,
    new_new_n837__, new_new_n838__, new_new_n839__, new_new_n840__,
    new_new_n841__, new_new_n842__, new_new_n843__, new_new_n844__,
    new_new_n845__, new_new_n846__, new_new_n847__, new_new_n848__,
    new_new_n849__, new_new_n850__, new_new_n851__, new_new_n852__,
    new_new_n853__, new_new_n854__, new_new_n855__, new_new_n856__,
    new_new_n857__, new_new_n858__, new_new_n859__, new_new_n860__,
    new_new_n861__, new_new_n862__, new_new_n863__, new_new_n864__,
    new_new_n865__, new_new_n866__, new_new_n867__, new_new_n868__,
    new_new_n869__, new_new_n870__, new_new_n871__, new_new_n872__,
    new_new_n873__, new_new_n874__, new_new_n875__, new_new_n876__,
    new_new_n877__, new_new_n878__, new_new_n879__, new_new_n880__,
    new_new_n881__, new_new_n882__, new_new_n883__, new_new_n884__,
    new_new_n885__, new_new_n886__, new_new_n887__, new_new_n888__,
    new_new_n889__, new_new_n890__, new_new_n891__, new_new_n892__,
    new_new_n893__, new_new_n894__, new_new_n895__, new_new_n896__,
    new_new_n897__, new_new_n898__, new_new_n899__, new_new_n900__,
    new_new_n901__, new_new_n902__, new_new_n903__, new_new_n904__,
    new_new_n905__, new_new_n906__, new_new_n907__, new_new_n908__,
    new_new_n909__, new_new_n910__, new_new_n911__, new_new_n912__,
    new_new_n913__, new_new_n914__, new_new_n915__, new_new_n916__,
    new_new_n917__, new_new_n918__, new_new_n919__, new_new_n920__,
    new_new_n921__, new_new_n922__, new_new_n923__, new_new_n924__,
    new_new_n925__, new_new_n926__, new_new_n927__, new_new_n928__,
    new_new_n929__, new_new_n930__, new_new_n931__, new_new_n932__,
    new_new_n933__, new_new_n934__, new_new_n935__, new_new_n936__,
    new_new_n937__, new_new_n938__, new_new_n939__, new_new_n940__,
    new_new_n941__, new_new_n942__, new_new_n943__, new_new_n944__,
    new_new_n945__, new_new_n946__, new_new_n947__, new_new_n948__,
    new_new_n949__, new_new_n950__, new_new_n951__, new_new_n952__,
    new_new_n953__, new_new_n954__, new_new_n955__, new_new_n956__,
    new_new_n957__, new_new_n958__, new_new_n959__, new_new_n960__,
    new_new_n961__, new_new_n962__, new_new_n963__, new_new_n964__,
    new_new_n965__, new_new_n966__, new_new_n967__, new_new_n968__,
    new_new_n969__, new_new_n970__, new_new_n971__, new_new_n972__,
    new_new_n973__, new_new_n974__, new_new_n975__, new_new_n976__,
    new_new_n977__, new_new_n978__, new_new_n979__, new_new_n980__,
    new_new_n981__, new_new_n982__, new_new_n983__, new_new_n984__,
    new_new_n985__, new_new_n986__, new_new_n987__, new_new_n988__,
    new_new_n989__, new_new_n990__, new_new_n991__, new_new_n992__,
    new_new_n993__, new_new_n994__, new_new_n995__, new_new_n996__,
    new_new_n997__, new_new_n998__, new_new_n999__, new_new_n1000__,
    new_new_n1001__, new_new_n1002__, new_new_n1003__, new_new_n1004__,
    new_new_n1005__, new_new_n1006__, new_new_n1007__, new_new_n1008__,
    new_new_n1009__, new_new_n1010__, new_new_n1011__, new_new_n1012__,
    new_new_n1013__, new_new_n1014__, new_new_n1015__, new_new_n1016__,
    new_new_n1017__, new_new_n1018__, new_new_n1019__, new_new_n1020__,
    new_new_n1021__, new_new_n1022__, new_new_n1023__, new_new_n1024__,
    new_new_n1025__, new_new_n1026__, new_new_n1027__, new_new_n1028__,
    new_new_n1029__, new_new_n1030__, new_new_n1031__, new_new_n1032__,
    new_new_n1033__, new_new_n1034__, new_new_n1035__, new_new_n1036__,
    new_new_n1037__, new_new_n1038__, new_new_n1039__, new_new_n1040__,
    new_new_n1041__, new_new_n1042__, new_new_n1043__, new_new_n1044__,
    new_new_n1045__, new_new_n1046__, new_new_n1047__, new_new_n1048__,
    new_new_n1049__, new_new_n1050__, new_new_n1051__, new_new_n1052__,
    new_new_n1053__, new_new_n1054__, new_new_n1055__, new_new_n1056__,
    new_new_n1057__, new_new_n1058__, new_new_n1059__, new_new_n1060__,
    new_new_n1061__, new_new_n1062__, new_new_n1063__, new_new_n1064__,
    new_new_n1065__, new_new_n1066__, new_new_n1067__, new_new_n1068__,
    new_new_n1069__, new_new_n1070__, new_new_n1071__, new_new_n1072__,
    new_new_n1073__, new_new_n1074__, new_new_n1075__, new_new_n1076__,
    new_new_n1077__, new_new_n1078__, new_new_n1079__, new_new_n1080__,
    new_new_n1081__, new_new_n1082__, new_new_n1083__, new_new_n1084__,
    new_new_n1085__, new_new_n1086__, new_new_n1087__, new_new_n1088__,
    new_new_n1089__, new_new_n1090__, new_new_n1091__, new_new_n1092__,
    new_new_n1093__, new_new_n1094__, new_new_n1095__, new_new_n1096__,
    new_new_n1097__, new_new_n1098__, new_new_n1099__, new_new_n1100__,
    new_new_n1101__, new_new_n1102__, new_new_n1103__, new_new_n1104__,
    new_new_n1105__, new_new_n1106__, new_new_n1107__, new_new_n1108__,
    new_new_n1109__, new_new_n1110__, new_new_n1111__, new_new_n1112__,
    new_new_n1113__, new_new_n1114__, new_new_n1115__, new_new_n1116__,
    new_new_n1117__, new_new_n1118__, new_new_n1119__, new_new_n1120__,
    new_new_n1121__, new_new_n1122__, new_new_n1123__, new_new_n1124__,
    new_new_n1125__, new_new_n1126__, new_new_n1127__, new_new_n1128__,
    new_new_n1129__, new_new_n1130__, new_new_n1131__, new_new_n1132__,
    new_new_n1133__, new_new_n1134__, new_new_n1135__, new_new_n1136__,
    new_new_n1137__, new_new_n1138__, new_new_n1139__, new_new_n1140__,
    new_new_n1141__, new_new_n1142__, new_new_n1143__, new_new_n1144__,
    new_new_n1145__, new_new_n1146__, new_new_n1147__, new_new_n1148__,
    new_new_n1149__, new_new_n1150__, new_new_n1151__, new_new_n1152__,
    new_new_n1153__, new_new_n1154__, new_new_n1155__, new_new_n1156__,
    new_new_n1157__, new_new_n1158__, new_new_n1159__, new_new_n1160__,
    new_new_n1161__, new_new_n1162__, new_new_n1163__, new_new_n1164__,
    new_new_n1165__, new_new_n1166__, new_new_n1167__, new_new_n1168__,
    new_new_n1169__, new_new_n1170__, new_new_n1171__, new_new_n1172__,
    new_new_n1173__, new_new_n1174__, new_new_n1175__, new_new_n1176__,
    new_new_n1177__, new_new_n1178__, new_new_n1179__, new_new_n1180__,
    new_new_n1181__, new_new_n1182__, new_new_n1183__, new_new_n1184__,
    new_new_n1185__, new_new_n1186__, new_new_n1187__, new_new_n1188__,
    new_new_n1189__, new_new_n1190__, new_new_n1191__, new_new_n1192__,
    new_new_n1193__, new_new_n1194__, new_new_n1195__, new_new_n1196__,
    new_new_n1197__, new_new_n1198__, new_new_n1199__, new_new_n1200__,
    new_new_n1201__, new_new_n1202__, new_new_n1203__, new_new_n1204__,
    new_new_n1205__, new_new_n1206__, new_new_n1207__, new_new_n1208__,
    new_new_n1209__, new_new_n1210__, new_new_n1211__, new_new_n1212__,
    new_new_n1213__, new_new_n1214__, new_new_n1215__, new_new_n1216__,
    new_new_n1217__, new_new_n1218__, new_new_n1219__, new_new_n1220__,
    new_new_n1221__, new_new_n1222__, new_new_n1223__, new_new_n1224__,
    new_new_n1225__, new_new_n1226__, new_new_n1227__, new_new_n1228__,
    new_new_n1229__, new_new_n1230__, new_new_n1231__, new_new_n1232__,
    new_new_n1233__, new_new_n1234__, new_new_n1235__, new_new_n1236__,
    new_new_n1237__, new_new_n1238__, new_new_n1239__, new_new_n1240__,
    new_new_n1241__, new_new_n1242__, new_new_n1243__, new_new_n1244__,
    new_new_n1245__, new_new_n1246__, new_new_n1247__, new_new_n1248__,
    new_new_n1249__, new_new_n1250__, new_new_n1251__, new_new_n1252__,
    new_new_n1253__, new_new_n1254__, new_new_n1255__, new_new_n1256__,
    new_new_n1257__, new_new_n1258__, new_new_n1259__, new_new_n1260__,
    new_new_n1261__, new_new_n1262__, new_new_n1263__, new_new_n1264__,
    new_new_n1265__, new_new_n1266__, new_new_n1267__, new_new_n1268__,
    new_new_n1269__, new_new_n1270__, new_new_n1271__, new_new_n1272__,
    new_new_n1273__, new_new_n1274__, new_new_n1275__, new_new_n1276__,
    new_new_n1277__, new_new_n1278__, new_new_n1279__, new_new_n1280__,
    new_new_n1281__, new_new_n1282__, new_new_n1283__, new_new_n1284__,
    new_new_n1285__, new_new_n1286__, new_new_n1287__, new_new_n1288__,
    new_new_n1289__, new_new_n1290__, new_new_n1291__, new_new_n1292__,
    new_new_n1293__, new_new_n1294__, new_new_n1295__, new_new_n1296__,
    new_new_n1297__, new_new_n1298__, new_new_n1299__, new_new_n1300__,
    new_new_n1301__, new_new_n1302__, new_new_n1303__, new_new_n1304__,
    new_new_n1305__, new_new_n1306__, new_new_n1307__, new_new_n1308__,
    new_new_n1309__, new_new_n1310__, new_new_n1311__, new_new_n1312__,
    new_new_n1313__, new_new_n1314__, new_new_n1315__, new_new_n1316__,
    new_new_n1317__, new_new_n1318__, new_new_n1319__, new_new_n1320__,
    new_new_n1321__, new_new_n1322__, new_new_n1323__, new_new_n1324__,
    new_new_n1325__, new_new_n1326__, new_new_n1327__, new_new_n1328__,
    new_new_n1329__, new_new_n1330__, new_new_n1331__, new_new_n1332__,
    new_new_n1333__, new_new_n1334__, new_new_n1335__, new_new_n1336__,
    new_new_n1337__, new_new_n1338__, new_new_n1339__, new_new_n1340__,
    new_new_n1341__, new_new_n1342__, new_new_n1343__, new_new_n1344__,
    new_new_n1345__, new_new_n1346__, new_new_n1347__, new_new_n1348__,
    new_new_n1349__, new_new_n1350__, new_new_n1351__, new_new_n1352__,
    new_new_n1353__, new_new_n1354__, new_new_n1355__, new_new_n1356__,
    new_new_n1357__, new_new_n1358__, new_new_n1359__, new_new_n1360__,
    new_new_n1361__, new_new_n1362__, new_new_n1363__, new_new_n1364__,
    new_new_n1365__, new_new_n1366__, new_new_n1367__, new_new_n1368__,
    new_new_n1369__, new_new_n1370__, new_new_n1371__, new_new_n1372__,
    new_new_n1373__, new_new_n1374__, new_new_n1375__, new_new_n1376__,
    new_new_n1377__, new_new_n1378__, new_new_n1379__, new_new_n1380__,
    new_new_n1381__, new_new_n1382__, new_new_n1383__, new_new_n1384__,
    new_new_n1385__, new_new_n1386__, new_new_n1387__, new_new_n1388__,
    new_new_n1389__, new_new_n1390__, new_new_n1391__, new_new_n1392__,
    new_new_n1393__, new_new_n1394__, new_new_n1395__, new_new_n1396__,
    new_new_n1397__, new_new_n1398__, new_new_n1399__, new_new_n1400__,
    new_new_n1401__, new_new_n1402__, new_new_n1403__, new_new_n1404__,
    new_new_n1405__, new_new_n1406__, new_new_n1407__, new_new_n1408__,
    new_new_n1409__, new_new_n1410__, new_new_n1411__, new_new_n1412__,
    new_new_n1413__, new_new_n1414__, new_new_n1415__, new_new_n1416__,
    new_new_n1417__, new_new_n1418__, new_new_n1419__, new_new_n1420__,
    new_new_n1421__, new_new_n1422__, new_new_n1423__, new_new_n1424__,
    new_new_n1425__, new_new_n1426__, new_new_n1427__, new_new_n1428__,
    new_new_n1429__, new_new_n1430__, new_new_n1431__, new_new_n1432__,
    new_new_n1433__, new_new_n1434__, new_new_n1435__, new_new_n1436__,
    new_new_n1437__, new_new_n1438__, new_new_n1439__, new_new_n1440__,
    new_new_n1441__, new_new_n1442__, new_new_n1443__, new_new_n1444__,
    new_new_n1445__, new_new_n1446__, new_new_n1447__, new_new_n1448__,
    new_new_n1449__, new_new_n1450__, new_new_n1451__, new_new_n1452__,
    new_new_n1453__, new_new_n1454__, new_new_n1455__, new_new_n1456__,
    new_new_n1457__, new_new_n1458__, new_new_n1459__, new_new_n1460__,
    new_new_n1461__, new_new_n1462__, new_new_n1463__, new_new_n1464__,
    new_new_n1465__, new_new_n1466__, new_new_n1467__, new_new_n1468__,
    new_new_n1469__, new_new_n1470__, new_new_n1471__, new_new_n1472__,
    new_new_n1473__, new_new_n1474__, new_new_n1475__, new_new_n1476__,
    new_new_n1477__, new_new_n1478__, new_new_n1479__, new_new_n1480__,
    new_new_n1481__, new_new_n1482__, new_new_n1483__, new_new_n1484__,
    new_new_n1485__, new_new_n1486__, new_new_n1487__, new_new_n1488__,
    new_new_n1489__, new_new_n1490__, new_new_n1491__, new_new_n1492__,
    new_new_n1493__, new_new_n1494__, new_new_n1495__, new_new_n1496__,
    new_new_n1497__, new_new_n1498__, new_new_n1499__, new_new_n1500__,
    new_new_n1501__, new_new_n1502__, new_new_n1503__, new_new_n1504__,
    new_new_n1505__, new_new_n1506__, new_new_n1507__, new_new_n1508__,
    new_new_n1509__, new_new_n1510__, new_new_n1511__, new_new_n1512__,
    new_new_n1513__, new_new_n1514__, new_new_n1515__, new_new_n1516__,
    new_new_n1517__, new_new_n1518__, new_new_n1519__, new_new_n1520__,
    new_new_n1521__, new_new_n1522__, new_new_n1523__, new_new_n1524__,
    new_new_n1525__, new_new_n1526__, new_new_n1527__, new_new_n1528__,
    new_new_n1529__, new_new_n1530__, new_new_n1531__, new_new_n1532__,
    new_new_n1533__, new_new_n1534__, new_new_n1535__, new_new_n1536__,
    new_new_n1537__, new_new_n1538__, new_new_n1539__, new_new_n1540__,
    new_new_n1541__, new_new_n1542__, new_new_n1543__, new_new_n1544__,
    new_new_n1545__, new_new_n1546__, new_new_n1547__, new_new_n1548__,
    new_new_n1549__, new_new_n1550__, new_new_n1551__, new_new_n1552__,
    new_new_n1553__, new_new_n1554__, new_new_n1555__, new_new_n1556__,
    new_new_n1557__, new_new_n1558__, new_new_n1559__, new_new_n1560__,
    new_new_n1561__, new_new_n1562__, new_new_n1563__, new_new_n1564__,
    new_new_n1565__, new_new_n1566__, new_new_n1567__, new_new_n1568__,
    new_new_n1569__, new_new_n1570__, new_new_n1571__, new_new_n1572__,
    new_new_n1573__, new_new_n1574__, new_new_n1575__, new_new_n1576__,
    new_new_n1577__, new_new_n1578__, new_new_n1579__, new_new_n1580__,
    new_new_n1581__, new_new_n1582__, new_new_n1583__, new_new_n1584__,
    new_new_n1585__, new_new_n1586__, new_new_n1587__, new_new_n1588__,
    new_new_n1589__, new_new_n1590__, new_new_n1591__, new_new_n1592__,
    new_new_n1593__, new_new_n1594__, new_new_n1595__, new_new_n1596__,
    new_new_n1597__, new_new_n1598__, new_new_n1599__, new_new_n1600__,
    new_new_n1601__, new_new_n1602__, new_new_n1603__, new_new_n1604__,
    new_new_n1605__, new_new_n1606__, new_new_n1607__, new_new_n1608__,
    new_new_n1609__, new_new_n1610__, new_new_n1611__, new_new_n1612__,
    new_new_n1613__, new_new_n1614__, new_new_n1615__, new_new_n1616__,
    new_new_n1617__, new_new_n1618__, new_new_n1619__, new_new_n1620__,
    new_new_n1621__, new_new_n1622__, new_new_n1623__, new_new_n1624__,
    new_new_n1625__, new_new_n1626__, new_new_n1627__, new_new_n1628__,
    new_new_n1629__, new_new_n1630__, new_new_n1631__, new_new_n1632__,
    new_new_n1633__, new_new_n1634__, new_new_n1635__, new_new_n1636__,
    new_new_n1637__, new_new_n1638__, new_new_n1639__, new_new_n1640__,
    new_new_n1641__, new_new_n1642__, new_new_n1643__, new_new_n1644__,
    new_new_n1645__, new_new_n1646__, new_new_n1647__, new_new_n1648__,
    new_new_n1649__, new_new_n1650__, new_new_n1651__, new_new_n1652__,
    new_new_n1653__, new_new_n1654__, new_new_n1655__, new_new_n1656__,
    new_new_n1657__, new_new_n1658__, new_new_n1659__, new_new_n1660__,
    new_new_n1661__, new_new_n1662__, new_new_n1663__, new_new_n1664__,
    new_new_n1665__, new_new_n1666__, new_new_n1667__, new_new_n1668__,
    new_new_n1669__, new_new_n1670__, new_new_n1671__, new_new_n1672__,
    new_new_n1673__, new_new_n1674__, new_new_n1675__, new_new_n1676__,
    new_new_n1677__, new_new_n1678__, new_new_n1679__, new_new_n1680__,
    new_new_n1681__, new_new_n1682__, new_new_n1683__, new_new_n1684__,
    new_new_n1685__, new_new_n1686__, new_new_n1687__, new_new_n1688__,
    new_new_n1689__, new_new_n1690__, new_new_n1691__, new_new_n1692__,
    new_new_n1693__, new_new_n1694__, new_new_n1695__, new_new_n1696__,
    new_new_n1697__, new_new_n1698__, new_new_n1699__, new_new_n1700__,
    new_new_n1701__, new_new_n1702__, new_new_n1703__, new_new_n1704__,
    new_new_n1705__, new_new_n1706__, new_new_n1707__, new_new_n1708__,
    new_new_n1709__, new_new_n1710__, new_new_n1711__, new_new_n1712__,
    new_new_n1713__, new_new_n1714__, new_new_n1715__, new_new_n1716__,
    new_new_n1717__, new_new_n1718__, new_new_n1719__, new_new_n1720__,
    new_new_n1721__, new_new_n1722__, new_new_n1723__, new_new_n1724__,
    new_new_n1725__, new_new_n1726__, new_new_n1727__, new_new_n1728__,
    new_new_n1729__, new_new_n1730__, new_new_n1731__, new_new_n1732__,
    new_new_n1733__, new_new_n1734__, new_new_n1735__, new_new_n1736__,
    new_new_n1737__, new_new_n1738__, new_new_n1739__, new_new_n1740__,
    new_new_n1741__, new_new_n1742__, new_new_n1743__, new_new_n1744__,
    new_new_n1745__, new_new_n1746__, new_new_n1747__, new_new_n1748__,
    new_new_n1749__, new_new_n1750__, new_new_n1751__, new_new_n1752__,
    new_new_n1753__, new_new_n1754__, new_new_n1755__, new_new_n1756__,
    new_new_n1757__, new_new_n1758__, new_new_n1759__, new_new_n1760__,
    new_new_n1761__, new_new_n1762__, new_new_n1763__, new_new_n1764__,
    new_new_n1765__, new_new_n1766__, new_new_n1767__, new_new_n1768__,
    new_new_n1769__, new_new_n1770__, new_new_n1771__, new_new_n1772__,
    new_new_n1773__, new_new_n1774__, new_new_n1775__, new_new_n1776__,
    new_new_n1777__, new_new_n1778__, new_new_n1779__, new_new_n1780__,
    new_new_n1781__, new_new_n1782__, new_new_n1783__, new_new_n1784__,
    new_new_n1785__, new_new_n1786__, new_new_n1787__, new_new_n1788__,
    new_new_n1789__, new_new_n1790__, new_new_n1791__, new_new_n1792__,
    new_new_n1793__, new_new_n1794__, new_new_n1795__, new_new_n1796__,
    new_new_n1797__, new_new_n1798__, new_new_n1799__, new_new_n1800__,
    new_new_n1801__, new_new_n1802__, new_new_n1803__, new_new_n1804__,
    new_new_n1805__, new_new_n1806__, new_new_n1807__, new_new_n1808__,
    new_new_n1809__, new_new_n1810__, new_new_n1811__, new_new_n1812__,
    new_new_n1813__, new_new_n1814__, new_new_n1815__, new_new_n1816__,
    new_new_n1817__, new_new_n1818__, new_new_n1819__, new_new_n1820__,
    new_new_n1821__, new_new_n1822__, new_new_n1823__, new_new_n1824__,
    new_new_n1825__, new_new_n1826__, new_new_n1827__, new_new_n1828__,
    new_new_n1829__, new_new_n1830__, new_new_n1831__, new_new_n1832__,
    new_new_n1833__, new_new_n1834__, new_new_n1835__, new_new_n1836__,
    new_new_n1837__, new_new_n1838__, new_new_n1839__, new_new_n1840__,
    new_new_n1841__, new_new_n1842__, new_new_n1843__, new_new_n1844__,
    new_new_n1845__, new_new_n1846__, new_new_n1847__, new_new_n1848__,
    new_new_n1849__, new_new_n1850__, new_new_n1851__, new_new_n1852__,
    new_new_n1853__, new_new_n1854__, new_new_n1855__, new_new_n1856__,
    new_new_n1857__, new_new_n1858__, new_new_n1859__, new_new_n1860__,
    new_new_n1861__, new_new_n1862__, new_new_n1863__, new_new_n1864__,
    new_new_n1865__, new_new_n1866__, new_new_n1867__, new_new_n1868__,
    new_new_n1869__, new_new_n1870__, new_new_n1871__, new_new_n1872__,
    new_new_n1873__, new_new_n1874__, new_new_n1875__, new_new_n1876__,
    new_new_n1877__, new_new_n1878__, new_new_n1879__, new_new_n1880__,
    new_new_n1881__, new_new_n1882__, new_new_n1883__, new_new_n1884__,
    new_new_n1885__, new_new_n1886__, new_new_n1887__, new_new_n1888__,
    new_new_n1889__, new_new_n1890__, new_new_n1891__, new_new_n1892__,
    new_new_n1893__, new_new_n1894__, new_new_n1895__, new_new_n1896__,
    new_new_n1897__, new_new_n1898__, new_new_n1899__, new_new_n1900__,
    new_new_n1901__, new_new_n1902__, new_new_n1903__, new_new_n1904__,
    new_new_n1905__, new_new_n1906__, new_new_n1907__, new_new_n1908__,
    new_new_n1909__, new_new_n1910__, new_new_n1911__, new_new_n1912__,
    new_new_n1913__, new_new_n1914__, new_new_n1915__, new_new_n1916__,
    new_new_n1917__, new_new_n1918__, new_new_n1919__, new_new_n1920__,
    new_new_n1921__, new_new_n1922__, new_new_n1923__, new_new_n1924__,
    new_new_n1925__, new_new_n1926__, new_new_n1927__, new_new_n1928__,
    new_new_n1929__, new_new_n1930__, new_new_n1931__, new_new_n1932__,
    new_new_n1933__, new_new_n1934__, new_new_n1935__, new_new_n1936__,
    new_new_n1937__, new_new_n1938__, new_new_n1939__, new_new_n1940__,
    new_new_n1941__, new_new_n1942__, new_new_n1943__, new_new_n1944__,
    new_new_n1945__, new_new_n1946__, new_new_n1947__, new_new_n1948__,
    new_new_n1949__, new_new_n1950__, new_new_n1951__, new_new_n1952__,
    new_new_n1953__, new_new_n1954__, new_new_n1955__, new_new_n1956__,
    new_new_n1957__, new_new_n1958__, new_new_n1959__, new_new_n1960__,
    new_new_n1961__, new_new_n1962__, new_new_n1963__, new_new_n1964__,
    new_new_n1965__, new_new_n1966__, new_new_n1967__, new_new_n1968__,
    new_new_n1969__, new_new_n1970__, new_new_n1971__, new_new_n1972__,
    new_new_n1973__, new_new_n1974__, new_new_n1975__, new_new_n1976__,
    new_new_n1977__, new_new_n1978__, new_new_n1979__, new_new_n1980__,
    new_new_n1981__, new_new_n1982__, new_new_n1983__, new_new_n1984__,
    new_new_n1985__, new_new_n1986__, new_new_n1987__, new_new_n1988__,
    new_new_n1989__, new_new_n1990__, new_new_n1991__, new_new_n1992__,
    new_new_n1993__, new_new_n1994__, new_new_n1995__, new_new_n1996__,
    new_new_n1997__, new_new_n1998__, new_new_n1999__, new_new_n2000__,
    new_new_n2001__, new_new_n2002__, new_new_n2003__, new_new_n2004__,
    new_new_n2005__, new_new_n2006__, new_new_n2007__, new_new_n2008__,
    new_new_n2009__, new_new_n2010__, new_new_n2011__, new_new_n2012__,
    new_new_n2013__, new_new_n2014__, new_new_n2015__, new_new_n2016__,
    new_new_n2017__, new_new_n2018__, new_new_n2019__, new_new_n2020__,
    new_new_n2021__, new_new_n2022__, new_new_n2023__, new_new_n2024__,
    new_new_n2025__, new_new_n2026__, new_new_n2027__, new_new_n2028__,
    new_new_n2029__, new_new_n2030__, new_new_n2031__, new_new_n2032__,
    new_new_n2033__, new_new_n2034__, new_new_n2035__, new_new_n2036__,
    new_new_n2037__, new_new_n2038__, new_new_n2039__, new_new_n2040__,
    new_new_n2041__, new_new_n2042__, new_new_n2043__, new_new_n2044__,
    new_new_n2045__, new_new_n2046__, new_new_n2047__, new_new_n2048__,
    new_new_n2049__, new_new_n2050__, new_new_n2051__, new_new_n2052__,
    new_new_n2053__, new_new_n2054__, new_new_n2055__, new_new_n2056__,
    new_new_n2057__, new_new_n2058__, new_new_n2059__, new_new_n2060__,
    new_new_n2061__, new_new_n2062__, new_new_n2063__, new_new_n2064__,
    new_new_n2065__, new_new_n2066__, new_new_n2067__, new_new_n2068__,
    new_new_n2069__, new_new_n2070__, new_new_n2071__, new_new_n2072__,
    new_new_n2073__, new_new_n2074__, new_new_n2075__, new_new_n2076__,
    new_new_n2077__, new_new_n2078__, new_new_n2079__, new_new_n2080__,
    new_new_n2081__, new_new_n2082__, new_new_n2083__, new_new_n2084__,
    new_new_n2085__, new_new_n2086__, new_new_n2087__, new_new_n2088__,
    new_new_n2089__, new_new_n2090__, new_new_n2091__, new_new_n2092__,
    new_new_n2093__, new_new_n2094__, new_new_n2095__, new_new_n2096__,
    new_new_n2097__, new_new_n2098__, new_new_n2099__, new_new_n2100__,
    new_new_n2101__, new_new_n2102__, new_new_n2103__, new_new_n2104__,
    new_new_n2105__, new_new_n2106__, new_new_n2107__, new_new_n2108__,
    new_new_n2109__, new_new_n2110__, new_new_n2111__, new_new_n2112__,
    new_new_n2113__, new_new_n2114__, new_new_n2115__, new_new_n2116__,
    new_new_n2117__, new_new_n2118__, new_new_n2119__, new_new_n2120__,
    new_new_n2121__, new_new_n2122__, new_new_n2123__, new_new_n2124__,
    new_new_n2125__, new_new_n2126__, new_new_n2127__, new_new_n2128__,
    new_new_n2129__, new_new_n2130__, new_new_n2131__, new_new_n2132__,
    new_new_n2133__, new_new_n2134__, new_new_n2135__, new_new_n2136__,
    new_new_n2137__, new_new_n2138__, new_new_n2139__, new_new_n2140__,
    new_new_n2141__, new_new_n2142__, new_new_n2143__, new_new_n2144__,
    new_new_n2145__, new_new_n2146__, new_new_n2147__, new_new_n2148__,
    new_new_n2149__, new_new_n2150__, new_new_n2151__, new_new_n2152__,
    new_new_n2153__, new_new_n2154__, new_new_n2155__, new_new_n2156__,
    new_new_n2157__, new_new_n2158__, new_new_n2159__, new_new_n2160__,
    new_new_n2161__, new_new_n2162__, new_new_n2163__, new_new_n2164__,
    new_new_n2165__, new_new_n2166__, new_new_n2167__, new_new_n2168__,
    new_new_n2169__, new_new_n2170__, new_new_n2171__, new_new_n2172__,
    new_new_n2173__, new_new_n2174__, new_new_n2175__, new_new_n2176__,
    new_new_n2177__, new_new_n2178__, new_new_n2179__, new_new_n2180__,
    new_new_n2181__, new_new_n2182__, new_new_n2183__, new_new_n2184__,
    new_new_n2185__, new_new_n2186__, new_new_n2187__, new_new_n2188__,
    new_new_n2189__, new_new_n2190__, new_new_n2191__, new_new_n2192__,
    new_new_n2193__, new_new_n2194__, new_new_n2195__, new_new_n2196__,
    new_new_n2197__, new_new_n2198__, new_new_n2199__, new_new_n2200__,
    new_new_n2201__, new_new_n2202__, new_new_n2203__, new_new_n2204__,
    new_new_n2205__, new_new_n2206__, new_new_n2207__, new_new_n2208__,
    new_new_n2209__, new_new_n2210__, new_new_n2211__, new_new_n2212__,
    new_new_n2213__, new_new_n2214__, new_new_n2215__, new_new_n2216__,
    new_new_n2217__, new_new_n2218__, new_new_n2219__, new_new_n2220__,
    new_new_n2221__, new_new_n2222__, new_new_n2223__, new_new_n2224__,
    new_new_n2225__, new_new_n2226__, new_new_n2227__, new_new_n2228__,
    new_new_n2229__, new_new_n2230__, new_new_n2231__, new_new_n2232__,
    new_new_n2233__, new_new_n2234__, new_new_n2235__, new_new_n2236__,
    new_new_n2237__, new_new_n2238__, new_new_n2239__, new_new_n2240__,
    new_new_n2241__, new_new_n2242__, new_new_n2243__, new_new_n2244__,
    new_new_n2245__, new_new_n2246__, new_new_n2247__, new_new_n2248__,
    new_new_n2249__, new_new_n2250__, new_new_n2251__, new_new_n2252__,
    new_new_n2253__, new_new_n2254__, new_new_n2255__, new_new_n2256__,
    new_new_n2257__, new_new_n2258__, new_new_n2259__, new_new_n2260__,
    new_new_n2261__, new_new_n2262__, new_new_n2263__, new_new_n2264__,
    new_new_n2265__, new_new_n2266__, new_new_n2267__, new_new_n2268__,
    new_new_n2269__, new_new_n2270__, new_new_n2271__, new_new_n2272__,
    new_new_n2273__, new_new_n2274__, new_new_n2275__, new_new_n2276__,
    new_new_n2277__, new_new_n2278__, new_new_n2279__, new_new_n2280__,
    new_new_n2281__, new_new_n2282__, new_new_n2283__, new_new_n2284__,
    new_new_n2285__, new_new_n2286__, new_new_n2287__, new_new_n2288__,
    new_new_n2289__, new_new_n2290__, new_new_n2291__, new_new_n2292__,
    new_new_n2293__, new_new_n2294__, new_new_n2295__, new_new_n2296__,
    new_new_n2297__, new_new_n2298__, new_new_n2299__, new_new_n2300__,
    new_new_n2301__, new_new_n2302__, new_new_n2303__, new_new_n2304__,
    new_new_n2305__, new_new_n2306__, new_new_n2307__, new_new_n2308__,
    new_new_n2309__, new_new_n2310__, new_new_n2311__, new_new_n2312__,
    new_new_n2313__, new_new_n2314__, new_new_n2315__, new_new_n2316__,
    new_new_n2317__, new_new_n2318__, new_new_n2319__, new_new_n2320__,
    new_new_n2321__, new_new_n2322__, new_new_n2323__, new_new_n2324__,
    new_new_n2325__, new_new_n2326__, new_new_n2327__, new_new_n2328__,
    new_new_n2329__, new_new_n2330__, new_new_n2331__, new_new_n2332__,
    new_new_n2333__, new_new_n2334__, new_new_n2335__, new_new_n2336__,
    new_new_n2337__, new_new_n2338__, new_new_n2339__, new_new_n2340__,
    new_new_n2341__, new_new_n2342__, new_new_n2343__, new_new_n2344__,
    new_new_n2345__, new_new_n2346__, new_new_n2347__, new_new_n2348__,
    new_new_n2349__, new_new_n2350__, new_new_n2351__, new_new_n2352__,
    new_new_n2353__, new_new_n2354__, new_new_n2355__, new_new_n2356__,
    new_new_n2357__, new_new_n2358__, new_new_n2359__, new_new_n2360__,
    new_new_n2361__, new_new_n2362__, new_new_n2363__, new_new_n2364__,
    new_new_n2365__, new_new_n2366__, new_new_n2367__, new_new_n2368__,
    new_new_n2369__, new_new_n2370__, new_new_n2371__, new_new_n2372__,
    new_new_n2373__, new_new_n2374__, new_new_n2375__, new_new_n2376__,
    new_new_n2377__, new_new_n2378__, new_new_n2379__, new_new_n2380__,
    new_new_n2381__, new_new_n2382__, new_new_n2383__, new_new_n2384__,
    new_new_n2385__, new_new_n2386__, new_new_n2387__, new_new_n2388__,
    new_new_n2389__, new_new_n2390__, new_new_n2391__, new_new_n2392__,
    new_new_n2393__, new_new_n2394__, new_new_n2395__, new_new_n2396__,
    new_new_n2397__, new_new_n2398__, new_new_n2399__, new_new_n2400__,
    new_new_n2401__, new_new_n2402__, new_new_n2403__, new_new_n2404__,
    new_new_n2405__, new_new_n2406__, new_new_n2407__, new_new_n2408__,
    new_new_n2409__, new_new_n2410__, new_new_n2411__, new_new_n2412__,
    new_new_n2413__, new_new_n2414__, new_new_n2415__, new_new_n2416__,
    new_new_n2417__, new_new_n2418__, new_new_n2419__, new_new_n2420__,
    new_new_n2421__, new_new_n2422__, new_new_n2423__, new_new_n2424__,
    new_new_n2425__, new_new_n2426__, new_new_n2427__, new_new_n2428__,
    new_new_n2429__, new_new_n2430__, new_new_n2431__, new_new_n2432__,
    new_new_n2433__, new_new_n2434__, new_new_n2435__, new_new_n2436__,
    new_new_n2437__, new_new_n2438__, new_new_n2439__, new_new_n2440__,
    new_new_n2441__, new_new_n2442__, new_new_n2443__, new_new_n2444__,
    new_new_n2445__, new_new_n2446__, new_new_n2447__, new_new_n2448__,
    new_new_n2449__, new_new_n2450__, new_new_n2451__, new_new_n2452__,
    new_new_n2453__, new_new_n2454__, new_new_n2455__, new_new_n2456__,
    new_new_n2457__, new_new_n2458__, new_new_n2459__, new_new_n2460__,
    new_new_n2461__, new_new_n2462__, new_new_n2463__, new_new_n2464__,
    new_new_n2465__, new_new_n2466__, new_new_n2467__, new_new_n2468__,
    new_new_n2469__, new_new_n2470__, new_new_n2471__, new_new_n2472__,
    new_new_n2473__, new_new_n2474__, new_new_n2475__, new_new_n2476__,
    new_new_n2477__, new_new_n2478__, new_new_n2479__, new_new_n2480__,
    new_new_n2481__, new_new_n2482__, new_new_n2483__, new_new_n2484__,
    new_new_n2485__, new_new_n2486__, new_new_n2487__, new_new_n2488__,
    new_new_n2489__, new_new_n2490__, new_new_n2491__, new_new_n2492__,
    new_new_n2493__, new_new_n2494__, new_new_n2495__, new_new_n2496__,
    new_new_n2497__, new_new_n2498__, new_new_n2499__, new_new_n2500__,
    new_new_n2501__, new_new_n2502__, new_new_n2503__, new_new_n2504__,
    new_new_n2505__, new_new_n2506__, new_new_n2507__, new_new_n2508__,
    new_new_n2509__, new_new_n2510__, new_new_n2511__, new_new_n2512__,
    new_new_n2513__, new_new_n2514__, new_new_n2515__, new_new_n2516__,
    new_new_n2517__, new_new_n2518__, new_new_n2519__, new_new_n2520__,
    new_new_n2521__, new_new_n2522__, new_new_n2523__, new_new_n2524__,
    new_new_n2525__, new_new_n2526__, new_new_n2527__, new_new_n2528__,
    new_new_n2529__, new_new_n2530__, new_new_n2531__, new_new_n2532__,
    new_new_n2533__, new_new_n2534__, new_new_n2535__, new_new_n2536__,
    new_new_n2537__, new_new_n2538__, new_new_n2539__, new_new_n2540__,
    new_new_n2541__, new_new_n2542__, new_new_n2543__, new_new_n2544__,
    new_new_n2545__, new_new_n2546__, new_new_n2547__, new_new_n2548__,
    new_new_n2549__, new_new_n2550__, new_new_n2551__, new_new_n2552__,
    new_new_n2553__, new_new_n2554__, new_new_n2555__, new_new_n2556__,
    new_new_n2557__, new_new_n2558__, new_new_n2559__, new_new_n2560__,
    new_new_n2561__, new_new_n2562__, new_new_n2563__, new_new_n2564__,
    new_new_n2565__, new_new_n2566__, new_new_n2567__, new_new_n2568__,
    new_new_n2569__, new_new_n2570__, new_new_n2571__, new_new_n2572__,
    new_new_n2573__, new_new_n2574__, new_new_n2575__, new_new_n2576__,
    new_new_n2577__, new_new_n2578__, new_new_n2579__, new_new_n2580__,
    new_new_n2581__, new_new_n2582__, new_new_n2583__, new_new_n2584__,
    new_new_n2585__, new_new_n2586__, new_new_n2587__, new_new_n2588__,
    new_new_n2589__, new_new_n2590__, new_new_n2591__, new_new_n2592__,
    new_new_n2593__, new_new_n2594__, new_new_n2595__, new_new_n2596__,
    new_new_n2597__, new_new_n2598__, new_new_n2599__, new_new_n2600__,
    new_new_n2601__, new_new_n2602__, new_new_n2603__, new_new_n2604__,
    new_new_n2605__, new_new_n2606__, new_new_n2607__, new_new_n2608__,
    new_new_n2609__, new_new_n2610__, new_new_n2611__, new_new_n2612__,
    new_new_n2613__, new_new_n2614__, new_new_n2615__, new_new_n2616__,
    new_new_n2617__, new_new_n2618__, new_new_n2619__, new_new_n2620__,
    new_new_n2621__, new_new_n2622__, new_new_n2623__, new_new_n2624__,
    new_new_n2625__, new_new_n2626__, new_new_n2627__, new_new_n2628__,
    new_new_n2629__, new_new_n2630__, new_new_n2631__, new_new_n2632__,
    new_new_n2633__, new_new_n2634__, new_new_n2635__, new_new_n2636__,
    new_new_n2637__, new_new_n2638__, new_new_n2639__, new_new_n2640__,
    new_new_n2641__, new_new_n2642__, new_new_n2643__, new_new_n2644__,
    new_new_n2645__, new_new_n2646__, new_new_n2647__, new_new_n2648__,
    new_new_n2649__, new_new_n2650__, new_new_n2651__, new_new_n2652__,
    new_new_n2653__, new_new_n2654__, new_new_n2655__, new_new_n2656__,
    new_new_n2657__, new_new_n2658__, new_new_n2659__, new_new_n2660__,
    new_new_n2661__, new_new_n2662__, new_new_n2663__, new_new_n2664__,
    new_new_n2665__, new_new_n2666__, new_new_n2667__, new_new_n2668__,
    new_new_n2669__, new_new_n2670__, new_new_n2671__, new_new_n2672__,
    new_new_n2673__, new_new_n2674__, new_new_n2675__, new_new_n2676__,
    new_new_n2677__, new_new_n2678__, new_new_n2679__, new_new_n2680__,
    new_new_n2681__, new_new_n2682__, new_new_n2683__, new_new_n2684__,
    new_new_n2685__, new_new_n2686__, new_new_n2687__, new_new_n2688__,
    new_new_n2689__, new_new_n2690__, new_new_n2691__, new_new_n2692__,
    new_new_n2693__, new_new_n2694__, new_new_n2695__, new_new_n2696__,
    new_new_n2697__, new_new_n2698__, new_new_n2699__, new_new_n2700__,
    new_new_n2701__, new_new_n2702__, new_new_n2703__, new_new_n2704__,
    new_new_n2705__, new_new_n2706__, new_new_n2707__, new_new_n2708__,
    new_new_n2709__, new_new_n2710__, new_new_n2711__, new_new_n2712__,
    new_new_n2713__, new_new_n2714__, new_new_n2715__, new_new_n2716__,
    new_new_n2717__, new_new_n2718__, new_new_n2719__, new_new_n2720__,
    new_new_n2721__, new_new_n2722__, new_new_n2723__, new_new_n2724__,
    new_new_n2725__, new_new_n2726__, new_new_n2727__, new_new_n2728__,
    new_new_n2729__, new_new_n2730__, new_new_n2731__, new_new_n2732__,
    new_new_n2733__, new_new_n2734__, new_new_n2735__, new_new_n2736__,
    new_new_n2737__, new_new_n2738__, new_new_n2739__, new_new_n2740__,
    new_new_n2741__, new_new_n2742__, new_new_n2743__, new_new_n2744__,
    new_new_n2745__, new_new_n2746__, new_new_n2747__, new_new_n2748__,
    new_new_n2749__, new_new_n2750__, new_new_n2751__, new_new_n2752__,
    new_new_n2753__, new_new_n2754__, new_new_n2755__, new_new_n2756__,
    new_new_n2757__, new_new_n2758__, new_new_n2759__, new_new_n2760__,
    new_new_n2761__, new_new_n2762__, new_new_n2763__, new_new_n2764__,
    new_new_n2765__, new_new_n2766__, new_new_n2767__, new_new_n2768__,
    new_new_n2769__, new_new_n2770__, new_new_n2771__, new_new_n2772__,
    new_new_n2773__, new_new_n2774__, new_new_n2775__, new_new_n2776__,
    new_new_n2777__, new_new_n2778__, new_new_n2779__, new_new_n2780__,
    new_new_n2781__, new_new_n2782__, new_new_n2783__, new_new_n2784__,
    new_new_n2785__, new_new_n2786__, new_new_n2787__, new_new_n2788__,
    new_new_n2789__, new_new_n2790__, new_new_n2791__, new_new_n2792__,
    new_new_n2793__, new_new_n2794__, new_new_n2795__, new_new_n2796__,
    new_new_n2797__, new_new_n2798__, new_new_n2799__, new_new_n2800__,
    new_new_n2801__, new_new_n2802__, new_new_n2803__, new_new_n2804__,
    new_new_n2805__, new_new_n2806__, new_new_n2807__, new_new_n2808__,
    new_new_n2809__, new_new_n2810__, new_new_n2811__, new_new_n2812__,
    new_new_n2813__, new_new_n2814__, new_new_n2815__, new_new_n2816__,
    new_new_n2817__, new_new_n2818__, new_new_n2819__, new_new_n2820__,
    new_new_n2821__, new_new_n2822__, new_new_n2823__, new_new_n2824__,
    new_new_n2825__, new_new_n2826__, new_new_n2827__, new_new_n2828__,
    new_new_n2829__, new_new_n2830__, new_new_n2831__, new_new_n2832__,
    new_new_n2833__, new_new_n2834__, new_new_n2835__, new_new_n2836__,
    new_new_n2837__, new_new_n2838__, new_new_n2839__, new_new_n2840__,
    new_new_n2841__, new_new_n2842__, new_new_n2843__, new_new_n2844__,
    new_new_n2845__, new_new_n2846__, new_new_n2847__, new_new_n2848__,
    new_new_n2849__, new_new_n2850__, new_new_n2851__, new_new_n2852__,
    new_new_n2853__, new_new_n2854__, new_new_n2855__, new_new_n2856__,
    new_new_n2857__, new_new_n2858__, new_new_n2859__, new_new_n2860__,
    new_new_n2861__, new_new_n2862__, new_new_n2863__, new_new_n2864__,
    new_new_n2865__, new_new_n2866__, new_new_n2867__, new_new_n2868__,
    new_new_n2869__, new_new_n2870__, new_new_n2871__, new_new_n2872__,
    new_new_n2873__, new_new_n2874__, new_new_n2875__, new_new_n2876__,
    new_new_n2877__, new_new_n2878__, new_new_n2879__, new_new_n2880__,
    new_new_n2881__, new_new_n2882__, new_new_n2883__, new_new_n2884__,
    new_new_n2885__, new_new_n2886__, new_new_n2887__, new_new_n2888__,
    new_new_n2889__, new_new_n2890__, new_new_n2891__, new_new_n2892__,
    new_new_n2893__, new_new_n2894__, new_new_n2895__, new_new_n2896__,
    new_new_n2897__, new_new_n2898__, new_new_n2899__, new_new_n2900__,
    new_new_n2901__, new_new_n2902__, new_new_n2903__, new_new_n2904__,
    new_new_n2905__, new_new_n2906__, new_new_n2907__, new_new_n2908__,
    new_new_n2909__, new_new_n2910__, new_new_n2911__, new_new_n2912__,
    new_new_n2913__, new_new_n2914__, new_new_n2915__, new_new_n2916__,
    new_new_n2917__, new_new_n2918__, new_new_n2919__, new_new_n2920__,
    new_new_n2921__, new_new_n2922__, new_new_n2923__, new_new_n2924__,
    new_new_n2925__, new_new_n2926__, new_new_n2927__, new_new_n2928__,
    new_new_n2929__, new_new_n2930__, new_new_n2931__, new_new_n2932__,
    new_new_n2933__, new_new_n2934__, new_new_n2935__, new_new_n2936__,
    new_new_n2937__, new_new_n2938__, new_new_n2939__, new_new_n2940__,
    new_new_n2941__, new_new_n2942__, new_new_n2943__, new_new_n2944__,
    new_new_n2945__, new_new_n2946__, new_new_n2947__, new_new_n2948__,
    new_new_n2949__, new_new_n2950__, new_new_n2951__, new_new_n2952__,
    new_new_n2953__, new_new_n2954__, new_new_n2955__, new_new_n2956__,
    new_new_n2957__, new_new_n2958__, new_new_n2959__, new_new_n2960__,
    new_new_n2961__, new_new_n2962__, new_new_n2963__, new_new_n2964__,
    new_new_n2965__, new_new_n2966__, new_new_n2967__, new_new_n2968__,
    new_new_n2969__, new_new_n2970__, new_new_n2971__, new_new_n2972__,
    new_new_n2973__, new_new_n2974__, new_new_n2975__, new_new_n2976__,
    new_new_n2977__, new_new_n2978__, new_new_n2979__, new_new_n2980__,
    new_new_n2981__, new_new_n2982__, new_new_n2983__, new_new_n2984__,
    new_new_n2985__, new_new_n2986__, new_new_n2987__, new_new_n2988__,
    new_new_n2989__, new_new_n2990__, new_new_n2991__, new_new_n2992__,
    new_new_n2993__, new_new_n2994__, new_new_n2995__, new_new_n2996__,
    new_new_n2997__, new_new_n2998__, new_new_n2999__, new_new_n3000__,
    new_new_n3001__, new_new_n3002__, new_new_n3003__, new_new_n3004__,
    new_new_n3005__, new_new_n3006__, new_new_n3007__, new_new_n3008__,
    new_new_n3009__, new_new_n3010__, new_new_n3011__, new_new_n3012__,
    new_new_n3013__, new_new_n3014__, new_new_n3015__, new_new_n3016__,
    new_new_n3017__, new_new_n3018__, new_new_n3019__, new_new_n3020__,
    new_new_n3021__, new_new_n3022__, new_new_n3023__, new_new_n3024__,
    new_new_n3025__, new_new_n3026__, new_new_n3027__, new_new_n3028__,
    new_new_n3029__, new_new_n3030__, new_new_n3031__, new_new_n3032__,
    new_new_n3033__, new_new_n3034__, new_new_n3035__, new_new_n3036__,
    new_new_n3037__, new_new_n3038__, new_new_n3039__, new_new_n3040__,
    new_new_n3041__, new_new_n3042__, new_new_n3043__, new_new_n3044__,
    new_new_n3045__, new_new_n3046__, new_new_n3047__, new_new_n3048__,
    new_new_n3049__, new_new_n3050__, new_new_n3051__, new_new_n3052__,
    new_new_n3053__, new_new_n3054__, new_new_n3055__, new_new_n3056__,
    new_new_n3057__, new_new_n3058__, new_new_n3059__, new_new_n3060__,
    new_new_n3061__, new_new_n3062__, new_new_n3063__, new_new_n3064__,
    new_new_n3065__, new_new_n3066__, new_new_n3067__, new_new_n3068__,
    new_new_n3069__, new_new_n3070__, new_new_n3071__, new_new_n3072__,
    new_new_n3073__, new_new_n3074__, new_new_n3075__, new_new_n3076__,
    new_new_n3077__, new_new_n3078__, new_new_n3079__, new_new_n3080__,
    new_new_n3081__, new_new_n3082__, new_new_n3083__, new_new_n3084__,
    new_new_n3085__, new_new_n3086__, new_new_n3087__, new_new_n3088__,
    new_new_n3089__, new_new_n3090__, new_new_n3091__, new_new_n3092__,
    new_new_n3093__, new_new_n3094__, new_new_n3095__, new_new_n3096__,
    new_new_n3097__, new_new_n3098__, new_new_n3099__, new_new_n3100__,
    new_new_n3101__, new_new_n3102__, new_new_n3103__, new_new_n3104__,
    new_new_n3105__, new_new_n3106__, new_new_n3107__, new_new_n3108__,
    new_new_n3109__, new_new_n3110__, new_new_n3111__, new_new_n3112__,
    new_new_n3113__, new_new_n3114__, new_new_n3115__, new_new_n3116__,
    new_new_n3117__, new_new_n3118__, new_new_n3119__, new_new_n3120__,
    new_new_n3121__, new_new_n3122__, new_new_n3123__, new_new_n3124__,
    new_new_n3125__, new_new_n3126__, new_new_n3127__, new_new_n3128__,
    new_new_n3129__, new_new_n3130__, new_new_n3131__, new_new_n3132__,
    new_new_n3133__, new_new_n3134__, new_new_n3135__, new_new_n3136__,
    new_new_n3137__, new_new_n3138__, new_new_n3139__, new_new_n3140__,
    new_new_n3141__, new_new_n3142__, new_new_n3143__, new_new_n3144__,
    new_new_n3145__, new_new_n3146__, new_new_n3147__, new_new_n3148__,
    new_new_n3149__, new_new_n3150__, new_new_n3151__, new_new_n3152__,
    new_new_n3153__, new_new_n3154__, new_new_n3155__, new_new_n3156__,
    new_new_n3157__, new_new_n3158__, new_new_n3159__, new_new_n3160__,
    new_new_n3161__, new_new_n3162__, new_new_n3163__, new_new_n3164__,
    new_new_n3165__, new_new_n3166__, new_new_n3167__, new_new_n3168__,
    new_new_n3169__, new_new_n3170__, new_new_n3171__, new_new_n3172__,
    new_new_n3173__, new_new_n3174__, new_new_n3175__, new_new_n3176__,
    new_new_n3177__, new_new_n3178__, new_new_n3179__, new_new_n3180__,
    new_new_n3181__, new_new_n3182__, new_new_n3183__, new_new_n3184__,
    new_new_n3185__, new_new_n3186__, new_new_n3187__, new_new_n3188__,
    new_new_n3189__, new_new_n3190__, new_new_n3191__, new_new_n3192__,
    new_new_n3193__, new_new_n3194__, new_new_n3195__, new_new_n3196__,
    new_new_n3197__, new_new_n3198__, new_new_n3199__, new_new_n3200__,
    new_new_n3201__, new_new_n3202__, new_new_n3203__, new_new_n3204__,
    new_new_n3205__, new_new_n3206__, new_new_n3207__, new_new_n3208__,
    new_new_n3209__, new_new_n3210__, new_new_n3211__, new_new_n3212__,
    new_new_n3213__, new_new_n3214__, new_new_n3215__, new_new_n3216__,
    new_new_n3217__, new_new_n3218__, new_new_n3219__, new_new_n3220__,
    new_new_n3221__, new_new_n3222__, new_new_n3223__, new_new_n3224__,
    new_new_n3225__, new_new_n3226__, new_new_n3227__, new_new_n3228__,
    new_new_n3229__, new_new_n3230__, new_new_n3231__, new_new_n3232__,
    new_new_n3233__, new_new_n3234__, new_new_n3235__, new_new_n3236__,
    new_new_n3237__, new_new_n3238__, new_new_n3239__, new_new_n3240__,
    new_new_n3241__, new_new_n3242__, new_new_n3243__, new_new_n3244__,
    new_new_n3245__, new_new_n3246__, new_new_n3247__, new_new_n3248__,
    new_new_n3249__, new_new_n3250__, new_new_n3251__, new_new_n3252__,
    new_new_n3253__, new_new_n3254__, new_new_n3255__, new_new_n3256__,
    new_new_n3257__, new_new_n3258__, new_new_n3259__, new_new_n3260__,
    new_new_n3261__, new_new_n3262__, new_new_n3263__, new_new_n3264__,
    new_new_n3265__, new_new_n3266__, new_new_n3267__, new_new_n3268__,
    new_new_n3269__, new_new_n3270__, new_new_n3271__, new_new_n3272__,
    new_new_n3273__, new_new_n3274__, new_new_n3275__, new_new_n3276__,
    new_new_n3277__, new_new_n3278__, new_new_n3279__, new_new_n3280__,
    new_new_n3281__, new_new_n3282__, new_new_n3283__, new_new_n3284__,
    new_new_n3285__, new_new_n3286__, new_new_n3287__, new_new_n3288__,
    new_new_n3289__, new_new_n3290__, new_new_n3291__, new_new_n3292__,
    new_new_n3293__, new_new_n3294__, new_new_n3295__, new_new_n3296__,
    new_new_n3297__, new_new_n3298__, new_new_n3299__, new_new_n3300__,
    new_new_n3301__, new_new_n3302__, new_new_n3303__, new_new_n3304__,
    new_new_n3305__, new_new_n3306__, new_new_n3307__, new_new_n3308__,
    new_new_n3309__, new_new_n3310__, new_new_n3311__, new_new_n3312__,
    new_new_n3313__, new_new_n3314__, new_new_n3315__, new_new_n3316__,
    new_new_n3317__, new_new_n3318__, new_new_n3319__, new_new_n3320__,
    new_new_n3321__, new_new_n3322__, new_new_n3323__, new_new_n3324__,
    new_new_n3325__, new_new_n3326__, new_new_n3327__, new_new_n3328__,
    new_new_n3329__, new_new_n3330__, new_new_n3331__, new_new_n3332__,
    new_new_n3333__, new_new_n3334__, new_new_n3335__, new_new_n3336__,
    new_new_n3337__, new_new_n3338__, new_new_n3339__, new_new_n3340__,
    new_new_n3341__, new_new_n3342__, new_new_n3343__, new_new_n3344__,
    new_new_n3345__, new_new_n3346__, new_new_n3347__, new_new_n3348__,
    new_new_n3349__, new_new_n3350__, new_new_n3351__, new_new_n3352__,
    new_new_n3353__, new_new_n3354__, new_new_n3355__, new_new_n3356__,
    new_new_n3357__, new_new_n3358__, new_new_n3359__, new_new_n3360__,
    new_new_n3361__, new_new_n3362__, new_new_n3363__, new_new_n3364__,
    new_new_n3365__, new_new_n3366__, new_new_n3367__, new_new_n3368__,
    new_new_n3369__, new_new_n3370__, new_new_n3371__, new_new_n3372__,
    new_new_n3373__, new_new_n3374__, new_new_n3375__, new_new_n3376__,
    new_new_n3377__, new_new_n3378__, new_new_n3379__, new_new_n3380__,
    new_new_n3381__, new_new_n3382__, new_new_n3383__, new_new_n3384__,
    new_new_n3385__, new_new_n3386__, new_new_n3387__, new_new_n3388__,
    new_new_n3389__, new_new_n3390__, new_new_n3391__, new_new_n3392__,
    new_new_n3393__, new_new_n3394__, new_new_n3395__, new_new_n3396__,
    new_new_n3397__, new_new_n3398__, new_new_n3399__, new_new_n3400__,
    new_new_n3401__, new_new_n3402__, new_new_n3403__, new_new_n3404__,
    new_new_n3405__, new_new_n3406__, new_new_n3407__, new_new_n3408__,
    new_new_n3409__, new_new_n3410__, new_new_n3411__, new_new_n3412__,
    new_new_n3413__, new_new_n3414__, new_new_n3415__, new_new_n3416__,
    new_new_n3417__, new_new_n3418__, new_new_n3419__, new_new_n3420__,
    new_new_n3421__, new_new_n3422__, new_new_n3423__, new_new_n3424__,
    new_new_n3425__, new_new_n3426__, new_new_n3427__, new_new_n3428__,
    new_new_n3429__, new_new_n3430__, new_new_n3431__, new_new_n3432__,
    new_new_n3433__, new_new_n3434__, new_new_n3435__, new_new_n3436__,
    new_new_n3437__, new_new_n3438__, new_new_n3439__, new_new_n3440__,
    new_new_n3441__, new_new_n3442__, new_new_n3443__, new_new_n3444__,
    new_new_n3445__, new_new_n3446__, new_new_n3447__, new_new_n3448__,
    new_new_n3449__, new_new_n3450__, new_new_n3451__, new_new_n3452__,
    new_new_n3453__, new_new_n3454__, new_new_n3455__, new_new_n3456__,
    new_new_n3457__, new_new_n3458__, new_new_n3459__, new_new_n3460__,
    new_new_n3461__, new_new_n3462__, new_new_n3463__, new_new_n3464__,
    new_new_n3465__, new_new_n3466__, new_new_n3467__, new_new_n3468__,
    new_new_n3469__, new_new_n3470__, new_new_n3471__, new_new_n3472__,
    new_new_n3473__, new_new_n3474__, new_new_n3475__, new_new_n3476__,
    new_new_n3477__, new_new_n3478__, new_new_n3479__, new_new_n3480__,
    new_new_n3481__, new_new_n3482__, new_new_n3483__, new_new_n3484__,
    new_new_n3485__, new_new_n3486__, new_new_n3487__, new_new_n3488__,
    new_new_n3489__, new_new_n3490__, new_new_n3491__, new_new_n3492__,
    new_new_n3493__, new_new_n3494__, new_new_n3495__, new_new_n3496__,
    new_new_n3497__, new_new_n3498__, new_new_n3499__, new_new_n3500__,
    new_new_n3501__, new_new_n3502__, new_new_n3503__, new_new_n3504__,
    new_new_n3505__, new_new_n3506__, new_new_n3507__, new_new_n3508__,
    new_new_n3509__, new_new_n3510__, new_new_n3511__, new_new_n3512__,
    new_new_n3513__, new_new_n3514__, new_new_n3515__, new_new_n3516__,
    new_new_n3517__, new_new_n3518__, new_new_n3519__, new_new_n3520__,
    new_new_n3521__, new_new_n3522__, new_new_n3523__, new_new_n3524__,
    new_new_n3525__, new_new_n3526__, new_new_n3527__, new_new_n3528__,
    new_new_n3529__, new_new_n3530__, new_new_n3531__, new_new_n3532__,
    new_new_n3533__, new_new_n3534__, new_new_n3535__, new_new_n3536__,
    new_new_n3537__, new_new_n3538__, new_new_n3539__, new_new_n3540__,
    new_new_n3541__, new_new_n3542__, new_new_n3543__, new_new_n3544__,
    new_new_n3545__, new_new_n3546__, new_new_n3547__, new_new_n3548__,
    new_new_n3549__, new_new_n3550__, new_new_n3551__, new_new_n3552__,
    new_new_n3553__, new_new_n3554__, new_new_n3555__, new_new_n3556__,
    new_new_n3557__, new_new_n3558__, new_new_n3559__, new_new_n3560__,
    new_new_n3561__, new_new_n3562__, new_new_n3563__, new_new_n3564__,
    new_new_n3565__, new_new_n3566__, new_new_n3567__, new_new_n3568__,
    new_new_n3569__, new_new_n3570__, new_new_n3571__, new_new_n3572__,
    new_new_n3573__, new_new_n3574__, new_new_n3575__, new_new_n3576__,
    new_new_n3577__, new_new_n3578__, new_new_n3579__, new_new_n3580__,
    new_new_n3581__, new_new_n3582__, new_new_n3583__, new_new_n3584__,
    new_new_n3585__, new_new_n3586__, new_new_n3587__, new_new_n3588__,
    new_new_n3589__, new_new_n3590__, new_new_n3591__, new_new_n3592__,
    new_new_n3593__, new_new_n3594__, new_new_n3595__, new_new_n3596__,
    new_new_n3597__, new_new_n3598__, new_new_n3599__, new_new_n3600__,
    new_new_n3601__, new_new_n3602__, new_new_n3603__, new_new_n3604__,
    new_new_n3605__, new_new_n3606__, new_new_n3607__, new_new_n3608__,
    new_new_n3609__, new_new_n3610__, new_new_n3611__, new_new_n3612__,
    new_new_n3613__, new_new_n3614__, new_new_n3615__, new_new_n3616__,
    new_new_n3617__, new_new_n3618__, new_new_n3619__, new_new_n3620__,
    new_new_n3621__, new_new_n3622__, new_new_n3623__, new_new_n3624__,
    new_new_n3625__, new_new_n3626__, new_new_n3627__, new_new_n3628__,
    new_new_n3629__, new_new_n3630__, new_new_n3631__, new_new_n3632__,
    new_new_n3633__, new_new_n3634__, new_new_n3635__, new_new_n3636__,
    new_new_n3637__, new_new_n3638__, new_new_n3639__, new_new_n3640__,
    new_new_n3641__, new_new_n3642__, new_new_n3643__, new_new_n3644__,
    new_new_n3645__, new_new_n3646__, new_new_n3647__, new_new_n3648__,
    new_new_n3649__, new_new_n3650__, new_new_n3651__, new_new_n3652__,
    new_new_n3653__, new_new_n3654__, new_new_n3655__, new_new_n3656__,
    new_new_n3657__, new_new_n3658__, new_new_n3659__, new_new_n3660__,
    new_new_n3661__, new_new_n3662__, new_new_n3663__, new_new_n3664__,
    new_new_n3665__, new_new_n3666__, new_new_n3667__, new_new_n3668__,
    new_new_n3669__, new_new_n3670__, new_new_n3671__, new_new_n3672__,
    new_new_n3673__, new_new_n3674__, new_new_n3675__, new_new_n3676__,
    new_new_n3677__, new_new_n3678__, new_new_n3679__, new_new_n3680__,
    new_new_n3681__, new_new_n3682__, new_new_n3683__, new_new_n3684__,
    new_new_n3685__, new_new_n3686__, new_new_n3687__, new_new_n3688__,
    new_new_n3689__, new_new_n3690__, new_new_n3691__, new_new_n3692__,
    new_new_n3693__, new_new_n3694__, new_new_n3695__, new_new_n3696__,
    new_new_n3697__, new_new_n3698__, new_new_n3699__, new_new_n3700__,
    new_new_n3701__, new_new_n3702__, new_new_n3703__, new_new_n3704__,
    new_new_n3705__, new_new_n3706__, new_new_n3707__, new_new_n3708__,
    new_new_n3709__, new_new_n3710__, new_new_n3711__, new_new_n3712__,
    new_new_n3713__, new_new_n3714__, new_new_n3715__, new_new_n3716__,
    new_new_n3717__, new_new_n3718__, new_new_n3719__, new_new_n3720__,
    new_new_n3721__, new_new_n3722__, new_new_n3723__, new_new_n3724__,
    new_new_n3725__, new_new_n3726__, new_new_n3727__, new_new_n3728__,
    new_new_n3729__, new_new_n3730__, new_new_n3731__, new_new_n3732__,
    new_new_n3733__, new_new_n3734__, new_new_n3735__, new_new_n3736__,
    new_new_n3737__, new_new_n3738__, new_new_n3739__, new_new_n3740__,
    new_new_n3741__, new_new_n3742__, new_new_n3743__, new_new_n3744__,
    new_new_n3745__, new_new_n3746__, new_new_n3747__, new_new_n3748__,
    new_new_n3749__, new_new_n3750__, new_new_n3751__, new_new_n3752__,
    new_new_n3753__, new_new_n3754__, new_new_n3755__, new_new_n3756__,
    new_new_n3757__, new_new_n3758__, new_new_n3759__, new_new_n3760__,
    new_new_n3761__, new_new_n3762__, new_new_n3763__, new_new_n3764__,
    new_new_n3765__, new_new_n3766__, new_new_n3767__, new_new_n3768__,
    new_new_n3769__, new_new_n3770__, new_new_n3771__, new_new_n3772__,
    new_new_n3773__, new_new_n3774__, new_new_n3775__, new_new_n3776__,
    new_new_n3777__, new_new_n3778__, new_new_n3779__, new_new_n3780__,
    new_new_n3781__, new_new_n3782__, new_new_n3783__, new_new_n3784__,
    new_new_n3785__, new_new_n3786__, new_new_n3787__, new_new_n3788__,
    new_new_n3789__, new_new_n3790__, new_new_n3791__, new_new_n3792__,
    new_new_n3793__, new_new_n3794__, new_new_n3795__, new_new_n3796__,
    new_new_n3797__, new_new_n3798__, new_new_n3799__, new_new_n3800__,
    new_new_n3801__, new_new_n3802__, new_new_n3803__, new_new_n3804__,
    new_new_n3805__, new_new_n3806__, new_new_n3807__, new_new_n3808__,
    new_new_n3809__, new_new_n3810__, new_new_n3811__, new_new_n3812__,
    new_new_n3813__, new_new_n3814__, new_new_n3815__, new_new_n3816__,
    new_new_n3817__, new_new_n3818__, new_new_n3819__, new_new_n3820__,
    new_new_n3821__, new_new_n3822__, new_new_n3823__, new_new_n3824__,
    new_new_n3825__, new_new_n3826__, new_new_n3827__, new_new_n3828__,
    new_new_n3829__, new_new_n3830__, new_new_n3831__, new_new_n3832__,
    new_new_n3833__, new_new_n3834__, new_new_n3835__, new_new_n3836__,
    new_new_n3837__, new_new_n3838__, new_new_n3839__, new_new_n3840__,
    new_new_n3841__, new_new_n3842__, new_new_n3843__, new_new_n3844__,
    new_new_n3845__, new_new_n3846__, new_new_n3847__, new_new_n3848__,
    new_new_n3849__, new_new_n3850__, new_new_n3851__, new_new_n3852__,
    new_new_n3853__, new_new_n3854__, new_new_n3855__, new_new_n3856__,
    new_new_n3857__, new_new_n3858__, new_new_n3859__, new_new_n3860__,
    new_new_n3861__, new_new_n3862__, new_new_n3863__, new_new_n3864__,
    new_new_n3865__, new_new_n3866__, new_new_n3867__, new_new_n3868__,
    new_new_n3869__, new_new_n3870__, new_new_n3871__, new_new_n3872__,
    new_new_n3873__, new_new_n3874__, new_new_n3875__, new_new_n3876__,
    new_new_n3877__, new_new_n3878__, new_new_n3879__, new_new_n3880__,
    new_new_n3881__, new_new_n3882__, new_new_n3883__, new_new_n3884__,
    new_new_n3885__, new_new_n3886__, new_new_n3887__, new_new_n3888__,
    new_new_n3889__, new_new_n3890__, new_new_n3891__, new_new_n3892__,
    new_new_n3893__, new_new_n3894__, new_new_n3895__, new_new_n3896__,
    new_new_n3897__, new_new_n3898__, new_new_n3899__, new_new_n3900__,
    new_new_n3901__, new_new_n3902__, new_new_n3903__, new_new_n3904__,
    new_new_n3905__, new_new_n3906__, new_new_n3907__, new_new_n3908__,
    new_new_n3909__, new_new_n3910__, new_new_n3911__, new_new_n3912__,
    new_new_n3913__, new_new_n3914__, new_new_n3915__, new_new_n3916__,
    new_new_n3917__, new_new_n3918__, new_new_n3919__, new_new_n3920__,
    new_new_n3921__, new_new_n3922__, new_new_n3923__, new_new_n3924__,
    new_new_n3925__, new_new_n3926__, new_new_n3927__, new_new_n3928__,
    new_new_n3929__, new_new_n3930__, new_new_n3931__, new_new_n3932__,
    new_new_n3933__, new_new_n3934__, new_new_n3935__, new_new_n3936__,
    new_new_n3937__, new_new_n3938__, new_new_n3939__, new_new_n3940__,
    new_new_n3941__, new_new_n3942__, new_new_n3943__, new_new_n3944__,
    new_new_n3945__, new_new_n3946__, new_new_n3947__, new_new_n3948__,
    new_new_n3949__, new_new_n3950__, new_new_n3951__, new_new_n3952__,
    new_new_n3953__, new_new_n3954__, new_new_n3955__, new_new_n3956__,
    new_new_n3957__, new_new_n3958__, new_new_n3959__, new_new_n3960__,
    new_new_n3961__, new_new_n3962__, new_new_n3963__, new_new_n3964__,
    new_new_n3965__, new_new_n3966__, new_new_n3967__, new_new_n3968__,
    new_new_n3969__, new_new_n3970__, new_new_n3971__, new_new_n3972__,
    new_new_n3973__, new_new_n3974__, new_new_n3975__, new_new_n3976__,
    new_new_n3977__, new_new_n3978__, new_new_n3979__, new_new_n3980__,
    new_new_n3981__, new_new_n3982__, new_new_n3983__, new_new_n3984__,
    new_new_n3985__, new_new_n3986__, new_new_n3987__, new_new_n3988__,
    new_new_n3989__, new_new_n3990__, new_new_n3991__, new_new_n3992__,
    new_new_n3993__, new_new_n3994__, new_new_n3995__, new_new_n3996__,
    new_new_n3997__, new_new_n3998__, new_new_n3999__, new_new_n4000__,
    new_new_n4001__, new_new_n4002__, new_new_n4003__, new_new_n4004__,
    new_new_n4005__, new_new_n4006__, new_new_n4007__, new_new_n4008__,
    new_new_n4009__, new_new_n4010__, new_new_n4011__, new_new_n4012__,
    new_new_n4013__, new_new_n4014__, new_new_n4015__, new_new_n4016__,
    new_new_n4017__, new_new_n4018__, new_new_n4019__, new_new_n4020__,
    new_new_n4021__, new_new_n4022__, new_new_n4023__, new_new_n4024__,
    new_new_n4025__, new_new_n4026__, new_new_n4027__, new_new_n4028__,
    new_new_n4029__, new_new_n4030__, new_new_n4031__, new_new_n4032__,
    new_new_n4033__, new_new_n4034__, new_new_n4035__, new_new_n4036__,
    new_new_n4037__, new_new_n4038__, new_new_n4039__, new_new_n4040__,
    new_new_n4041__, new_new_n4042__, new_new_n4043__, new_new_n4044__,
    new_new_n4045__, new_new_n4046__, new_new_n4047__, new_new_n4048__,
    new_new_n4049__, new_new_n4050__, new_new_n4051__, new_new_n4052__,
    new_new_n4053__, new_new_n4054__, new_new_n4055__, new_new_n4056__,
    new_new_n4057__, new_new_n4058__, new_new_n4059__, new_new_n4060__,
    new_new_n4061__, new_new_n4062__, new_new_n4063__, new_new_n4064__,
    new_new_n4065__, new_new_n4066__, new_new_n4067__, new_new_n4068__,
    new_new_n4069__, new_new_n4070__, new_new_n4071__, new_new_n4072__,
    new_new_n4073__, new_new_n4074__, new_new_n4075__, new_new_n4076__,
    new_new_n4077__, new_new_n4078__, new_new_n4079__, new_new_n4080__,
    new_new_n4081__, new_new_n4082__, new_new_n4083__, new_new_n4084__,
    new_new_n4085__, new_new_n4086__, new_new_n4087__, new_new_n4088__,
    new_new_n4089__, new_new_n4090__, new_new_n4091__, new_new_n4092__,
    new_new_n4093__, new_new_n4094__, new_new_n4095__, new_new_n4096__,
    new_new_n4097__, new_new_n4098__, new_new_n4099__, new_new_n4100__,
    new_new_n4101__, new_new_n4102__, new_new_n4103__, new_new_n4104__,
    new_new_n4105__, new_new_n4106__, new_new_n4107__, new_new_n4108__,
    new_new_n4109__, new_new_n4110__, new_new_n4111__, new_new_n4112__,
    new_new_n4113__, new_new_n4114__, new_new_n4115__, new_new_n4116__,
    new_new_n4117__, new_new_n4118__, new_new_n4119__, new_new_n4120__,
    new_new_n4121__, new_new_n4122__, new_new_n4123__, new_new_n4124__,
    new_new_n4125__, new_new_n4126__, new_new_n4127__, new_new_n4128__,
    new_new_n4129__, new_new_n4130__, new_new_n4131__, new_new_n4132__,
    new_new_n4133__, new_new_n4134__, new_new_n4135__, new_new_n4136__,
    new_new_n4137__, new_new_n4138__, new_new_n4139__, new_new_n4140__,
    new_new_n4141__, new_new_n4142__, new_new_n4143__, new_new_n4144__,
    new_new_n4145__, new_new_n4146__, new_new_n4147__, new_new_n4148__,
    new_new_n4149__, new_new_n4150__, new_new_n4151__, new_new_n4152__,
    new_new_n4153__, new_new_n4154__, new_new_n4155__, new_new_n4156__,
    new_new_n4157__, new_new_n4158__, new_new_n4159__, new_new_n4160__,
    new_new_n4161__, new_new_n4162__, new_new_n4163__, new_new_n4164__,
    new_new_n4165__, new_new_n4166__, new_new_n4167__, new_new_n4168__,
    new_new_n4169__, new_new_n4170__, new_new_n4171__, new_new_n4172__,
    new_new_n4173__, new_new_n4174__, new_new_n4175__, new_new_n4176__,
    new_new_n4177__, new_new_n4178__, new_new_n4179__, new_new_n4180__,
    new_new_n4181__, new_new_n4182__, new_new_n4183__, new_new_n4184__,
    new_new_n4185__, new_new_n4186__, new_new_n4187__, new_new_n4188__,
    new_new_n4189__, new_new_n4190__, new_new_n4191__, new_new_n4192__,
    new_new_n4193__, new_new_n4194__, new_new_n4195__, new_new_n4196__,
    new_new_n4197__, new_new_n4198__, new_new_n4199__, new_new_n4200__,
    new_new_n4201__, new_new_n4202__, new_new_n4203__, new_new_n4204__,
    new_new_n4205__, new_new_n4206__, new_new_n4207__, new_new_n4208__,
    new_new_n4209__, new_new_n4210__, new_new_n4211__, new_new_n4212__,
    new_new_n4213__, new_new_n4214__, new_new_n4215__, new_new_n4216__,
    new_new_n4217__, new_new_n4218__, new_new_n4219__, new_new_n4220__,
    new_new_n4221__, new_new_n4222__, new_new_n4223__, new_new_n4224__,
    new_new_n4225__, new_new_n4226__, new_new_n4227__, new_new_n4228__,
    new_new_n4229__, new_new_n4230__, new_new_n4231__, new_new_n4232__,
    new_new_n4233__, new_new_n4234__, new_new_n4235__, new_new_n4236__,
    new_new_n4237__, new_new_n4238__, new_new_n4239__, new_new_n4240__,
    new_new_n4241__, new_new_n4242__, new_new_n4243__, new_new_n4244__,
    new_new_n4245__, new_new_n4246__, new_new_n4247__, new_new_n4248__,
    new_new_n4249__, new_new_n4250__, new_new_n4251__, new_new_n4252__,
    new_new_n4253__, new_new_n4254__, new_new_n4255__, new_new_n4256__,
    new_new_n4257__, new_new_n4258__, new_new_n4259__, new_new_n4260__,
    new_new_n4261__, new_new_n4262__, new_new_n4263__, new_new_n4264__,
    new_new_n4265__, new_new_n4266__, new_new_n4267__, new_new_n4268__,
    new_new_n4269__, new_new_n4270__, new_new_n4271__, new_new_n4272__,
    new_new_n4273__, new_new_n4274__, new_new_n4275__, new_new_n4276__,
    new_new_n4277__, new_new_n4278__, new_new_n4279__, new_new_n4280__,
    new_new_n4281__, new_new_n4282__, new_new_n4283__, new_new_n4284__,
    new_new_n4285__, new_new_n4286__, new_new_n4287__, new_new_n4288__,
    new_new_n4289__, new_new_n4290__, new_new_n4291__, new_new_n4292__,
    new_new_n4293__, new_new_n4294__, new_new_n4295__, new_new_n4296__,
    new_new_n4297__, new_new_n4298__, new_new_n4299__, new_new_n4300__,
    new_new_n4301__, new_new_n4302__, new_new_n4303__, new_new_n4304__,
    new_new_n4305__, new_new_n4306__, new_new_n4307__, new_new_n4308__,
    new_new_n4309__, new_new_n4310__, new_new_n4311__, new_new_n4312__,
    new_new_n4313__, new_new_n4314__, new_new_n4315__, new_new_n4316__,
    new_new_n4317__, new_new_n4318__, new_new_n4319__, new_new_n4320__,
    new_new_n4321__, new_new_n4322__, new_new_n4323__, new_new_n4324__,
    new_new_n4325__, new_new_n4326__, new_new_n4327__, new_new_n4328__,
    new_new_n4329__, new_new_n4330__, new_new_n4331__, new_new_n4332__,
    new_new_n4333__, new_new_n4334__, new_new_n4335__, new_new_n4336__,
    new_new_n4337__, new_new_n4338__, new_new_n4339__, new_new_n4340__,
    new_new_n4341__, new_new_n4342__, new_new_n4343__, new_new_n4344__,
    new_new_n4345__, new_new_n4346__, new_new_n4347__, new_new_n4348__,
    new_new_n4349__, new_new_n4350__, new_new_n4351__, new_new_n4352__,
    new_new_n4353__, new_new_n4354__, new_new_n4355__, new_new_n4356__,
    new_new_n4357__, new_new_n4358__, new_new_n4359__, new_new_n4360__,
    new_new_n4361__, new_new_n4362__, new_new_n4363__, new_new_n4364__,
    new_new_n4365__, new_new_n4366__, new_new_n4367__, new_new_n4368__,
    new_new_n4369__, new_new_n4370__, new_new_n4371__, new_new_n4372__,
    new_new_n4373__, new_new_n4374__, new_new_n4375__, new_new_n4376__,
    new_new_n4377__, new_new_n4378__, new_new_n4379__, new_new_n4380__,
    new_new_n4381__, new_new_n4382__, new_new_n4383__, new_new_n4384__,
    new_new_n4385__, new_new_n4386__, new_new_n4387__, new_new_n4388__,
    new_new_n4389__, new_new_n4390__, new_new_n4391__, new_new_n4392__,
    new_new_n4393__, new_new_n4394__, new_new_n4395__, new_new_n4396__,
    new_new_n4397__, new_new_n4398__, new_new_n4399__, new_new_n4400__,
    new_new_n4401__, new_new_n4402__, new_new_n4403__, new_new_n4404__,
    new_new_n4405__, new_new_n4406__, new_new_n4407__, new_new_n4408__,
    new_new_n4409__, new_new_n4410__, new_new_n4411__, new_new_n4412__,
    new_new_n4413__, new_new_n4414__, new_new_n4415__, new_new_n4416__,
    new_new_n4417__, new_new_n4418__, new_new_n4419__, new_new_n4420__,
    new_new_n4421__, new_new_n4422__, new_new_n4423__, new_new_n4424__,
    new_new_n4425__, new_new_n4426__, new_new_n4427__, new_new_n4428__,
    new_new_n4429__, new_new_n4430__, new_new_n4431__, new_new_n4432__,
    new_new_n4433__, new_new_n4434__, new_new_n4435__, new_new_n4436__,
    new_new_n4437__, new_new_n4438__, new_new_n4439__, new_new_n4440__,
    new_new_n4441__, new_new_n4442__, new_new_n4443__, new_new_n4444__,
    new_new_n4445__, new_new_n4446__, new_new_n4447__, new_new_n4448__,
    new_new_n4449__, new_new_n4450__, new_new_n4451__, new_new_n4452__,
    new_new_n4453__, new_new_n4454__, new_new_n4455__, new_new_n4456__,
    new_new_n4457__, new_new_n4458__, new_new_n4459__, new_new_n4460__,
    new_new_n4461__, new_new_n4462__, new_new_n4463__, new_new_n4464__,
    new_new_n4465__, new_new_n4466__, new_new_n4467__, new_new_n4468__,
    new_new_n4469__, new_new_n4470__, new_new_n4471__, new_new_n4472__,
    new_new_n4473__, new_new_n4474__, new_new_n4475__, new_new_n4476__,
    new_new_n4477__, new_new_n4478__, new_new_n4479__, new_new_n4480__,
    new_new_n4481__, new_new_n4482__, new_new_n4483__, new_new_n4484__,
    new_new_n4485__, new_new_n4486__, new_new_n4487__, new_new_n4488__,
    new_new_n4489__, new_new_n4490__, new_new_n4491__, new_new_n4492__,
    new_new_n4493__, new_new_n4494__, new_new_n4495__, new_new_n4496__,
    new_new_n4497__, new_new_n4498__, new_new_n4499__, new_new_n4500__,
    new_new_n4501__, new_new_n4502__, new_new_n4503__, new_new_n4504__,
    new_new_n4505__, new_new_n4506__, new_new_n4507__, new_new_n4508__,
    new_new_n4509__, new_new_n4510__, new_new_n4511__, new_new_n4512__,
    new_new_n4513__, new_new_n4514__, new_new_n4515__, new_new_n4516__,
    new_new_n4517__, new_new_n4518__, new_new_n4519__, new_new_n4520__,
    new_new_n4521__, new_new_n4522__, new_new_n4523__, new_new_n4524__,
    new_new_n4525__, new_new_n4526__, new_new_n4527__, new_new_n4528__,
    new_new_n4529__, new_new_n4530__, new_new_n4531__, new_new_n4532__,
    new_new_n4533__, new_new_n4534__, new_new_n4535__, new_new_n4536__,
    new_new_n4537__, new_new_n4538__, new_new_n4539__, new_new_n4540__,
    new_new_n4541__, new_new_n4542__, new_new_n4543__, new_new_n4544__,
    new_new_n4545__, new_new_n4546__, new_new_n4547__, new_new_n4548__,
    new_new_n4549__, new_new_n4550__, new_new_n4551__, new_new_n4552__,
    new_new_n4553__, new_new_n4554__, new_new_n4555__, new_new_n4556__,
    new_new_n4557__, new_new_n4558__, new_new_n4559__, new_new_n4560__,
    new_new_n4561__, new_new_n4562__, new_new_n4563__, new_new_n4564__,
    new_new_n4565__, new_new_n4566__, new_new_n4567__, new_new_n4568__,
    new_new_n4569__, new_new_n4570__, new_new_n4571__, new_new_n4572__,
    new_new_n4573__, new_new_n4574__, new_new_n4575__, new_new_n4576__,
    new_new_n4577__, new_new_n4578__, new_new_n4579__, new_new_n4580__,
    new_new_n4581__, new_new_n4582__, new_new_n4583__, new_new_n4584__,
    new_new_n4585__, new_new_n4586__, new_new_n4587__, new_new_n4588__,
    new_new_n4589__, new_new_n4590__, new_new_n4591__, new_new_n4592__,
    new_new_n4593__, new_new_n4594__, new_new_n4595__, new_new_n4596__,
    new_new_n4597__, new_new_n4598__, new_new_n4599__, new_new_n4600__,
    new_new_n4601__, new_new_n4602__, new_new_n4603__, new_new_n4604__,
    new_new_n4605__, new_new_n4606__, new_new_n4607__, new_new_n4608__,
    new_new_n4609__, new_new_n4610__, new_new_n4611__, new_new_n4612__,
    new_new_n4613__, new_new_n4614__, new_new_n4615__, new_new_n4616__,
    new_new_n4617__, new_new_n4618__, new_new_n4619__, new_new_n4620__,
    new_new_n4621__, new_new_n4622__, new_new_n4623__, new_new_n4624__,
    new_new_n4625__, new_new_n4626__, new_new_n4627__, new_new_n4628__,
    new_new_n4629__, new_new_n4630__, new_new_n4631__, new_new_n4632__,
    new_new_n4633__, new_new_n4634__, new_new_n4635__, new_new_n4636__,
    new_new_n4637__, new_new_n4638__, new_new_n4639__, new_new_n4640__,
    new_new_n4641__, new_new_n4642__, new_new_n4643__, new_new_n4644__,
    new_new_n4645__, new_new_n4646__, new_new_n4647__, new_new_n4648__,
    new_new_n4649__, new_new_n4650__, new_new_n4651__, new_new_n4652__,
    new_new_n4653__, new_new_n4654__, new_new_n4655__, new_new_n4656__,
    new_new_n4657__, new_new_n4658__, new_new_n4659__, new_new_n4660__,
    new_new_n4661__, new_new_n4662__, new_new_n4663__, new_new_n4664__,
    new_new_n4665__, new_new_n4666__, new_new_n4667__, new_new_n4668__,
    new_new_n4669__, new_new_n4670__, new_new_n4671__, new_new_n4672__,
    new_new_n4673__, new_new_n4674__, new_new_n4675__, new_new_n4676__,
    new_new_n4677__, new_new_n4678__, new_new_n4679__, new_new_n4680__,
    new_new_n4681__, new_new_n4682__, new_new_n4683__, new_new_n4684__,
    new_new_n4685__, new_new_n4686__, new_new_n4687__, new_new_n4688__,
    new_new_n4689__, new_new_n4690__, new_new_n4691__, new_new_n4692__,
    new_new_n4693__, new_new_n4694__, new_new_n4695__, new_new_n4696__,
    new_new_n4697__, new_new_n4698__, new_new_n4699__, new_new_n4700__,
    new_new_n4701__, new_new_n4702__, new_new_n4703__, new_new_n4704__,
    new_new_n4705__, new_new_n4706__, new_new_n4707__, new_new_n4708__,
    new_new_n4709__, new_new_n4710__, new_new_n4711__, new_new_n4712__,
    new_new_n4713__, new_new_n4714__, new_new_n4715__, new_new_n4716__,
    new_new_n4717__, new_new_n4718__, new_new_n4719__, new_new_n4720__,
    new_new_n4721__, new_new_n4722__, new_new_n4723__, new_new_n4724__,
    new_new_n4725__, new_new_n4726__, new_new_n4727__, new_new_n4728__,
    new_new_n4729__, new_new_n4730__, new_new_n4731__, new_new_n4732__,
    new_new_n4733__, new_new_n4734__, new_new_n4735__, new_new_n4736__,
    new_new_n4737__, new_new_n4738__, new_new_n4739__, new_new_n4740__,
    new_new_n4741__, new_new_n4742__, new_new_n4743__, new_new_n4744__,
    new_new_n4745__, new_new_n4746__, new_new_n4747__, new_new_n4748__,
    new_new_n4749__, new_new_n4750__, new_new_n4751__, new_new_n4752__,
    new_new_n4753__, new_new_n4754__, new_new_n4755__, new_new_n4756__,
    new_new_n4757__, new_new_n4758__, new_new_n4759__, new_new_n4760__,
    new_new_n4761__, new_new_n4762__, new_new_n4763__, new_new_n4764__,
    new_new_n4765__, new_new_n4766__, new_new_n4767__, new_new_n4768__,
    new_new_n4769__, new_new_n4770__, new_new_n4771__, new_new_n4772__,
    new_new_n4773__, new_new_n4774__, new_new_n4775__, new_new_n4776__,
    new_new_n4777__, new_new_n4778__, new_new_n4779__, new_new_n4780__,
    new_new_n4781__, new_new_n4782__, new_new_n4783__, new_new_n4784__,
    new_new_n4785__, new_new_n4786__, new_new_n4787__, new_new_n4788__,
    new_new_n4789__, new_new_n4790__, new_new_n4791__, new_new_n4792__,
    new_new_n4793__, new_new_n4794__, new_new_n4795__, new_new_n4796__,
    new_new_n4797__, new_new_n4798__, new_new_n4799__, new_new_n4800__,
    new_new_n4801__, new_new_n4802__, new_new_n4803__, new_new_n4804__,
    new_new_n4805__, new_new_n4806__, new_new_n4807__, new_new_n4808__,
    new_new_n4809__, new_new_n4810__, new_new_n4811__, new_new_n4812__,
    new_new_n4813__, new_new_n4814__, new_new_n4815__, new_new_n4816__,
    new_new_n4817__, new_new_n4818__, new_new_n4819__, new_new_n4820__,
    new_new_n4821__, new_new_n4822__, new_new_n4823__, new_new_n4824__,
    new_new_n4825__, new_new_n4826__, new_new_n4827__, new_new_n4828__,
    new_new_n4829__, new_new_n4830__, new_new_n4831__, new_new_n4832__,
    new_new_n4833__, new_new_n4834__, new_new_n4835__, new_new_n4836__,
    new_new_n4837__, new_new_n4838__, new_new_n4839__, new_new_n4840__,
    new_new_n4841__, new_new_n4842__, new_new_n4843__, new_new_n4844__,
    new_new_n4845__, new_new_n4846__, new_new_n4847__, new_new_n4848__,
    new_new_n4849__, new_new_n4850__, new_new_n4851__, new_new_n4852__,
    new_new_n4853__, new_new_n4854__, new_new_n4855__, new_new_n4856__,
    new_new_n4857__, new_new_n4858__, new_new_n4859__, new_new_n4860__,
    new_new_n4861__, new_new_n4862__, new_new_n4863__, new_new_n4864__,
    new_new_n4865__, new_new_n4866__, new_new_n4867__, new_new_n4868__,
    new_new_n4869__, new_new_n4870__, new_new_n4871__, new_new_n4872__,
    new_new_n4873__, new_new_n4874__, new_new_n4875__, new_new_n4876__,
    new_new_n4877__, new_new_n4878__, new_new_n4879__, new_new_n4880__,
    new_new_n4881__, new_new_n4882__, new_new_n4883__, new_new_n4884__,
    new_new_n4885__, new_new_n4886__, new_new_n4887__, new_new_n4888__,
    new_new_n4889__, new_new_n4890__, new_new_n4891__, new_new_n4892__,
    new_new_n4893__, new_new_n4894__, new_new_n4895__, new_new_n4896__,
    new_new_n4897__, new_new_n4898__, new_new_n4899__, new_new_n4900__,
    new_new_n4901__, new_new_n4902__, new_new_n4903__, new_new_n4904__,
    new_new_n4905__, new_new_n4906__, new_new_n4907__, new_new_n4908__,
    new_new_n4909__, new_new_n4910__, new_new_n4911__, new_new_n4912__,
    new_new_n4913__, new_new_n4914__, new_new_n4915__, new_new_n4916__,
    new_new_n4917__, new_new_n4918__, new_new_n4919__, new_new_n4920__,
    new_new_n4921__, new_new_n4922__, new_new_n4923__, new_new_n4924__,
    new_new_n4925__, new_new_n4926__, new_new_n4927__, new_new_n4928__,
    new_new_n4929__, new_new_n4930__, new_new_n4931__, new_new_n4932__,
    new_new_n4933__, new_new_n4934__, new_new_n4935__, new_new_n4936__,
    new_new_n4937__, new_new_n4938__, new_new_n4939__, new_new_n4940__,
    new_new_n4941__, new_new_n4942__, new_new_n4943__, new_new_n4944__,
    new_new_n4945__, new_new_n4946__, new_new_n4947__, new_new_n4948__,
    new_new_n4949__, new_new_n4950__, new_new_n4951__, new_new_n4952__,
    new_new_n4953__, new_new_n4954__, new_new_n4955__, new_new_n4956__,
    new_new_n4957__, new_new_n4958__, new_new_n4959__, new_new_n4960__,
    new_new_n4961__, new_new_n4962__, new_new_n4963__, new_new_n4964__,
    new_new_n4965__, new_new_n4966__, new_new_n4967__, new_new_n4968__,
    new_new_n4969__, new_new_n4970__, new_new_n4971__, new_new_n4972__,
    new_new_n4973__, new_new_n4974__, new_new_n4975__, new_new_n4976__,
    new_new_n4977__, new_new_n4978__, new_new_n4979__, new_new_n4980__,
    new_new_n4981__, new_new_n4982__, new_new_n4983__, new_new_n4984__,
    new_new_n4985__, new_new_n4986__, new_new_n4987__, new_new_n4988__,
    new_new_n4989__, new_new_n4990__, new_new_n4991__, new_new_n4992__,
    new_new_n4993__, new_new_n4994__, new_new_n4995__, new_new_n4996__,
    new_new_n4997__, new_new_n4998__, new_new_n4999__, new_new_n5000__,
    new_new_n5001__, new_new_n5002__, new_new_n5003__, new_new_n5004__,
    new_new_n5005__, new_new_n5006__, new_new_n5007__, new_new_n5008__,
    new_new_n5009__, new_new_n5010__, new_new_n5011__, new_new_n5012__,
    new_new_n5013__, new_new_n5014__, new_new_n5015__, new_new_n5016__,
    new_new_n5017__, new_new_n5018__, new_new_n5019__, new_new_n5020__,
    new_new_n5021__, new_new_n5022__, new_new_n5023__, new_new_n5024__,
    new_new_n5025__, new_new_n5026__, new_new_n5027__, new_new_n5028__,
    new_new_n5029__, new_new_n5030__, new_new_n5031__, new_new_n5032__,
    new_new_n5033__, new_new_n5034__, new_new_n5035__, new_new_n5036__,
    new_new_n5037__, new_new_n5038__, new_new_n5039__, new_new_n5040__,
    new_new_n5041__, new_new_n5042__, new_new_n5043__, new_new_n5044__,
    new_new_n5045__, new_new_n5046__, new_new_n5047__, new_new_n5048__,
    new_new_n5049__, new_new_n5050__, new_new_n5051__, new_new_n5052__,
    new_new_n5053__, new_new_n5054__, new_new_n5055__, new_new_n5056__,
    new_new_n5057__, new_new_n5058__, new_new_n5059__, new_new_n5060__,
    new_new_n5061__, new_new_n5062__, new_new_n5063__, new_new_n5064__,
    new_new_n5065__, new_new_n5066__, new_new_n5067__, new_new_n5068__,
    new_new_n5069__, new_new_n5070__, new_new_n5071__, new_new_n5072__,
    new_new_n5073__, new_new_n5074__, new_new_n5075__, new_new_n5076__,
    new_new_n5077__, new_new_n5078__, new_new_n5079__, new_new_n5080__,
    new_new_n5081__, new_new_n5082__, new_new_n5083__, new_new_n5084__,
    new_new_n5085__, new_new_n5086__, new_new_n5087__, new_new_n5088__,
    new_new_n5089__, new_new_n5090__, new_new_n5091__, new_new_n5092__,
    new_new_n5093__, new_new_n5094__, new_new_n5095__, new_new_n5096__,
    new_new_n5097__, new_new_n5098__, new_new_n5099__, new_new_n5100__,
    new_new_n5101__, new_new_n5102__, new_new_n5103__, new_new_n5104__,
    new_new_n5105__, new_new_n5106__, new_new_n5107__, new_new_n5108__,
    new_new_n5109__, new_new_n5110__, new_new_n5111__, new_new_n5112__,
    new_new_n5113__, new_new_n5114__, new_new_n5115__, new_new_n5116__,
    new_new_n5117__, new_new_n5118__, new_new_n5119__, new_new_n5120__,
    new_new_n5121__, new_new_n5122__, new_new_n5123__, new_new_n5124__,
    new_new_n5125__, new_new_n5126__, new_new_n5127__, new_new_n5128__,
    new_new_n5129__, new_new_n5130__, new_new_n5131__, new_new_n5132__,
    new_new_n5133__, new_new_n5134__, new_new_n5135__, new_new_n5136__,
    new_new_n5137__, new_new_n5138__, new_new_n5139__, new_new_n5140__,
    new_new_n5141__, new_new_n5142__, new_new_n5143__, new_new_n5144__,
    new_new_n5145__, new_new_n5146__, new_new_n5147__, new_new_n5148__,
    new_new_n5149__, new_new_n5150__, new_new_n5151__, new_new_n5152__,
    new_new_n5153__, new_new_n5154__, new_new_n5155__, new_new_n5156__,
    new_new_n5157__, new_new_n5158__, new_new_n5159__, new_new_n5160__,
    new_new_n5161__, new_new_n5162__, new_new_n5163__, new_new_n5164__,
    new_new_n5165__, new_new_n5166__, new_new_n5167__, new_new_n5168__,
    new_new_n5169__, new_new_n5170__, new_new_n5171__, new_new_n5172__,
    new_new_n5173__, new_new_n5174__, new_new_n5175__, new_new_n5176__,
    new_new_n5177__, new_new_n5178__, new_new_n5179__, new_new_n5180__,
    new_new_n5181__, new_new_n5182__, new_new_n5183__, new_new_n5184__,
    new_new_n5185__, new_new_n5186__, new_new_n5187__, new_new_n5188__,
    new_new_n5189__, new_new_n5190__, new_new_n5191__, new_new_n5192__,
    new_new_n5193__, new_new_n5194__, new_new_n5195__, new_new_n5196__,
    new_new_n5197__, new_new_n5198__, new_new_n5199__, new_new_n5200__,
    new_new_n5201__, new_new_n5202__, new_new_n5203__, new_new_n5204__,
    new_new_n5205__, new_new_n5206__, new_new_n5207__, new_new_n5208__,
    new_new_n5209__, new_new_n5210__, new_new_n5211__, new_new_n5212__,
    new_new_n5213__, new_new_n5214__, new_new_n5215__, new_new_n5216__,
    new_new_n5217__, new_new_n5218__, new_new_n5219__, new_new_n5220__,
    new_new_n5221__, new_new_n5222__, new_new_n5223__, new_new_n5224__,
    new_new_n5225__, new_new_n5226__, new_new_n5227__, new_new_n5228__,
    new_new_n5229__, new_new_n5230__, new_new_n5231__, new_new_n5232__,
    new_new_n5233__, new_new_n5234__, new_new_n5235__, new_new_n5236__,
    new_new_n5237__, new_new_n5238__, new_new_n5239__, new_new_n5240__,
    new_new_n5241__, new_new_n5242__, new_new_n5243__, new_new_n5244__,
    new_new_n5245__, new_new_n5246__, new_new_n5247__, new_new_n5248__,
    new_new_n5249__, new_new_n5250__, new_new_n5251__, new_new_n5252__,
    new_new_n5253__, new_new_n5254__, new_new_n5255__, new_new_n5256__,
    new_new_n5257__, new_new_n5258__, new_new_n5259__, new_new_n5260__,
    new_new_n5261__, new_new_n5262__, new_new_n5263__, new_new_n5264__,
    new_new_n5265__, new_new_n5266__, new_new_n5267__, new_new_n5268__,
    new_new_n5269__, new_new_n5270__, new_new_n5271__, new_new_n5272__,
    new_new_n5273__, new_new_n5274__, new_new_n5275__, new_new_n5276__,
    new_new_n5277__, new_new_n5278__, new_new_n5279__, new_new_n5280__,
    new_new_n5281__, new_new_n5282__, new_new_n5283__, new_new_n5284__,
    new_new_n5285__, new_new_n5286__, new_new_n5287__, new_new_n5288__,
    new_new_n5289__, new_new_n5290__, new_new_n5291__, new_new_n5292__,
    new_new_n5293__, new_new_n5294__, new_new_n5295__, new_new_n5296__,
    new_new_n5297__, new_new_n5298__, new_new_n5299__, new_new_n5300__,
    new_new_n5301__, new_new_n5302__, new_new_n5303__, new_new_n5304__,
    new_new_n5305__, new_new_n5306__, new_new_n5307__, new_new_n5308__,
    new_new_n5309__, new_new_n5310__, new_new_n5311__, new_new_n5312__,
    new_new_n5313__, new_new_n5314__, new_new_n5315__, new_new_n5316__,
    new_new_n5317__, new_new_n5318__, new_new_n5319__, new_new_n5320__,
    new_new_n5321__, new_new_n5322__, new_new_n5323__, new_new_n5324__,
    new_new_n5325__, new_new_n5326__, new_new_n5327__, new_new_n5328__,
    new_new_n5329__, new_new_n5330__, new_new_n5331__, new_new_n5332__,
    new_new_n5333__, new_new_n5334__, new_new_n5335__, new_new_n5336__,
    new_new_n5337__, new_new_n5338__, new_new_n5339__, new_new_n5340__,
    new_new_n5341__, new_new_n5342__, new_new_n5343__, new_new_n5344__,
    new_new_n5345__, new_new_n5346__, new_new_n5347__, new_new_n5348__,
    new_new_n5349__, new_new_n5350__, new_new_n5351__, new_new_n5352__,
    new_new_n5353__, new_new_n5354__, new_new_n5355__, new_new_n5356__,
    new_new_n5357__, new_new_n5358__, new_new_n5359__, new_new_n5360__,
    new_new_n5361__, new_new_n5362__, new_new_n5363__, new_new_n5364__,
    new_new_n5365__, new_new_n5366__, new_new_n5367__, new_new_n5368__,
    new_new_n5369__, new_new_n5370__, new_new_n5371__, new_new_n5372__,
    new_new_n5373__, new_new_n5374__, new_new_n5375__, new_new_n5376__,
    new_new_n5377__, new_new_n5378__, new_new_n5379__, new_new_n5380__,
    new_new_n5381__, new_new_n5382__, new_new_n5383__, new_new_n5384__,
    new_new_n5385__, new_new_n5386__, new_new_n5387__, new_new_n5388__,
    new_new_n5389__, new_new_n5390__, new_new_n5391__, new_new_n5392__,
    new_new_n5393__, new_new_n5394__, new_new_n5395__, new_new_n5396__,
    new_new_n5397__, new_new_n5398__, new_new_n5399__, new_new_n5400__,
    new_new_n5401__, new_new_n5402__, new_new_n5403__, new_new_n5404__,
    new_new_n5405__, new_new_n5406__, new_new_n5407__, new_new_n5408__,
    new_new_n5409__, new_new_n5410__, new_new_n5411__, new_new_n5412__,
    new_new_n5413__, new_new_n5414__, new_new_n5415__, new_new_n5416__,
    new_new_n5417__, new_new_n5418__, new_new_n5419__, new_new_n5420__,
    new_new_n5421__, new_new_n5422__, new_new_n5423__, new_new_n5424__,
    new_new_n5425__, new_new_n5426__, new_new_n5427__, new_new_n5428__,
    new_new_n5429__, new_new_n5430__, new_new_n5431__, new_new_n5432__,
    new_new_n5433__, new_new_n5434__, new_new_n5435__, new_new_n5436__,
    new_new_n5437__, new_new_n5438__, new_new_n5439__, new_new_n5440__,
    new_new_n5441__, new_new_n5442__, new_new_n5443__, new_new_n5444__,
    new_new_n5445__, new_new_n5446__, new_new_n5447__, new_new_n5448__,
    new_new_n5449__, new_new_n5450__, new_new_n5451__, new_new_n5452__,
    new_new_n5453__, new_new_n5454__, new_new_n5455__, new_new_n5456__,
    new_new_n5457__, new_new_n5458__, new_new_n5459__, new_new_n5460__,
    new_new_n5461__, new_new_n5462__, new_new_n5463__, new_new_n5464__,
    new_new_n5465__, new_new_n5466__, new_new_n5467__, new_new_n5468__,
    new_new_n5469__, new_new_n5470__, new_new_n5471__, new_new_n5472__,
    new_new_n5473__, new_new_n5474__, new_new_n5475__, new_new_n5476__,
    new_new_n5477__, new_new_n5478__, new_new_n5479__, new_new_n5480__,
    new_new_n5481__, new_new_n5482__, new_new_n5483__, new_new_n5484__,
    new_new_n5485__, new_new_n5486__, new_new_n5487__, new_new_n5488__,
    new_new_n5489__, new_new_n5490__, new_new_n5491__, new_new_n5492__,
    new_new_n5493__, new_new_n5494__, new_new_n5495__, new_new_n5496__,
    new_new_n5497__, new_new_n5498__, new_new_n5499__, new_new_n5500__,
    new_new_n5501__, new_new_n5502__, new_new_n5503__, new_new_n5504__,
    new_new_n5505__, new_new_n5506__, new_new_n5507__, new_new_n5508__,
    new_new_n5509__, new_new_n5510__, new_new_n5511__, new_new_n5512__,
    new_new_n5513__, new_new_n5514__, new_new_n5515__, new_new_n5516__,
    new_new_n5517__, new_new_n5518__, new_new_n5519__, new_new_n5520__,
    new_new_n5521__, new_new_n5522__, new_new_n5523__, new_new_n5524__,
    new_new_n5525__, new_new_n5526__, new_new_n5527__, new_new_n5528__,
    new_new_n5529__, new_new_n5530__, new_new_n5531__, new_new_n5532__,
    new_new_n5533__, new_new_n5534__, new_new_n5535__, new_new_n5536__,
    new_new_n5537__, new_new_n5538__, new_new_n5539__, new_new_n5540__,
    new_new_n5541__, new_new_n5542__, new_new_n5543__, new_new_n5544__,
    new_new_n5545__, new_new_n5546__, new_new_n5547__, new_new_n5548__,
    new_new_n5549__, new_new_n5550__, new_new_n5551__, new_new_n5552__,
    new_new_n5553__, new_new_n5554__, new_new_n5555__, new_new_n5556__,
    new_new_n5557__, new_new_n5558__, new_new_n5559__, new_new_n5560__,
    new_new_n5561__, new_new_n5562__, new_new_n5563__, new_new_n5564__,
    new_new_n5565__, new_new_n5566__, new_new_n5567__, new_new_n5568__,
    new_new_n5569__, new_new_n5570__, new_new_n5571__, new_new_n5572__,
    new_new_n5573__, new_new_n5574__, new_new_n5575__, new_new_n5576__,
    new_new_n5577__, new_new_n5578__, new_new_n5579__, new_new_n5580__,
    new_new_n5581__, new_new_n5582__, new_new_n5583__, new_new_n5584__,
    new_new_n5585__, new_new_n5586__, new_new_n5587__, new_new_n5588__,
    new_new_n5589__, new_new_n5590__, new_new_n5591__, new_new_n5592__,
    new_new_n5593__, new_new_n5594__, new_new_n5595__, new_new_n5596__,
    new_new_n5597__, new_new_n5598__, new_new_n5599__, new_new_n5600__,
    new_new_n5601__, new_new_n5602__, new_new_n5603__, new_new_n5604__,
    new_new_n5605__, new_new_n5606__, new_new_n5607__, new_new_n5608__,
    new_new_n5609__, new_new_n5610__, new_new_n5611__, new_new_n5612__,
    new_new_n5613__, new_new_n5614__, new_new_n5615__, new_new_n5616__,
    new_new_n5617__, new_new_n5618__, new_new_n5619__, new_new_n5620__,
    new_new_n5621__, new_new_n5622__, new_new_n5623__, new_new_n5624__,
    new_new_n5625__, new_new_n5626__, new_new_n5627__, new_new_n5628__,
    new_new_n5629__, new_new_n5630__, new_new_n5631__, new_new_n5632__,
    new_new_n5633__, new_new_n5634__, new_new_n5635__, new_new_n5636__,
    new_new_n5637__, new_new_n5638__, new_new_n5639__, new_new_n5640__,
    new_new_n5641__, new_new_n5642__, new_new_n5643__, new_new_n5644__,
    new_new_n5645__, new_new_n5646__, new_new_n5647__, new_new_n5648__,
    new_new_n5649__, new_new_n5650__, new_new_n5651__, new_new_n5652__,
    new_new_n5653__, new_new_n5654__, new_new_n5655__, new_new_n5656__,
    new_new_n5657__, new_new_n5658__, new_new_n5659__, new_new_n5660__,
    new_new_n5661__, new_new_n5662__, new_new_n5663__, new_new_n5664__,
    new_new_n5665__, new_new_n5666__, new_new_n5667__, new_new_n5668__,
    new_new_n5669__, new_new_n5670__, new_new_n5671__, new_new_n5672__,
    new_new_n5673__, new_new_n5674__, new_new_n5675__, new_new_n5676__,
    new_new_n5677__, new_new_n5678__, new_new_n5679__, new_new_n5680__,
    new_new_n5681__, new_new_n5682__, new_new_n5683__, new_new_n5684__,
    new_new_n5685__, new_new_n5686__, new_new_n5687__, new_new_n5688__,
    new_new_n5689__, new_new_n5690__, new_new_n5691__, new_new_n5692__,
    new_new_n5693__, new_new_n5694__, new_new_n5695__, new_new_n5696__,
    new_new_n5697__, new_new_n5698__, new_new_n5699__, new_new_n5700__,
    new_new_n5701__, new_new_n5702__, new_new_n5703__, new_new_n5704__,
    new_new_n5705__, new_new_n5706__, new_new_n5707__, new_new_n5708__,
    new_new_n5709__, new_new_n5710__, new_new_n5711__, new_new_n5712__,
    new_new_n5713__, new_new_n5714__, new_new_n5715__, new_new_n5716__,
    new_new_n5717__, new_new_n5718__, new_new_n5719__, new_new_n5720__,
    new_new_n5721__, new_new_n5722__, new_new_n5723__, new_new_n5724__,
    new_new_n5725__, new_new_n5726__, new_new_n5727__, new_new_n5728__,
    new_new_n5729__, new_new_n5730__, new_new_n5731__, new_new_n5732__,
    new_new_n5733__, new_new_n5734__, new_new_n5735__, new_new_n5736__,
    new_new_n5737__, new_new_n5738__, new_new_n5739__, new_new_n5740__,
    new_new_n5741__, new_new_n5742__, new_new_n5743__, new_new_n5744__,
    new_new_n5745__, new_new_n5746__, new_new_n5747__, new_new_n5748__,
    new_new_n5749__, new_new_n5750__, new_new_n5751__, new_new_n5752__,
    new_new_n5753__, new_new_n5754__, new_new_n5755__, new_new_n5756__,
    new_new_n5757__, new_new_n5758__, new_new_n5759__, new_new_n5760__,
    new_new_n5761__, new_new_n5762__, new_new_n5763__, new_new_n5764__,
    new_new_n5765__, new_new_n5766__, new_new_n5767__, new_new_n5768__,
    new_new_n5769__, new_new_n5770__, new_new_n5771__, new_new_n5772__,
    new_new_n5773__, new_new_n5774__, new_new_n5775__, new_new_n5776__,
    new_new_n5777__, new_new_n5778__, new_new_n5779__, new_new_n5780__,
    new_new_n5781__, new_new_n5782__, new_new_n5783__, new_new_n5784__,
    new_new_n5785__, new_new_n5786__, new_new_n5787__, new_new_n5788__,
    new_new_n5789__, new_new_n5790__, new_new_n5791__, new_new_n5792__,
    new_new_n5793__, new_new_n5794__, new_new_n5795__, new_new_n5796__,
    new_new_n5797__, new_new_n5798__, new_new_n5799__, new_new_n5800__,
    new_new_n5801__, new_new_n5802__, new_new_n5803__, new_new_n5804__,
    new_new_n5805__, new_new_n5806__, new_new_n5807__, new_new_n5808__,
    new_new_n5809__, new_new_n5810__, new_new_n5811__, new_new_n5812__,
    new_new_n5813__, new_new_n5814__, new_new_n5815__, new_new_n5816__,
    new_new_n5817__, new_new_n5818__, new_new_n5819__, new_new_n5820__,
    new_new_n5821__, new_new_n5822__, new_new_n5823__, new_new_n5824__,
    new_new_n5825__, new_new_n5826__, new_new_n5827__, new_new_n5828__,
    new_new_n5829__, new_new_n5830__, new_new_n5831__, new_new_n5832__,
    new_new_n5833__, new_new_n5834__, new_new_n5835__, new_new_n5836__,
    new_new_n5837__, new_new_n5838__, new_new_n5839__, new_new_n5840__,
    new_new_n5841__, new_new_n5842__, new_new_n5843__, new_new_n5844__,
    new_new_n5845__, new_new_n5846__, new_new_n5847__, new_new_n5848__,
    new_new_n5849__, new_new_n5850__, new_new_n5851__, new_new_n5852__,
    new_new_n5853__, new_new_n5854__, new_new_n5855__, new_new_n5856__,
    new_new_n5857__, new_new_n5858__, new_new_n5859__, new_new_n5860__,
    new_new_n5861__, new_new_n5862__, new_new_n5863__, new_new_n5864__,
    new_new_n5865__, new_new_n5866__, new_new_n5867__, new_new_n5868__,
    new_new_n5869__, new_new_n5870__, new_new_n5871__, new_new_n5872__,
    new_new_n5873__, new_new_n5874__, new_new_n5875__, new_new_n5876__,
    new_new_n5877__, new_new_n5878__, new_new_n5879__, new_new_n5880__,
    new_new_n5881__, new_new_n5882__, new_new_n5883__, new_new_n5884__,
    new_new_n5885__, new_new_n5886__, new_new_n5887__, new_new_n5888__,
    new_new_n5889__, new_new_n5890__, new_new_n5891__, new_new_n5892__,
    new_new_n5893__, new_new_n5894__, new_new_n5895__, new_new_n5896__,
    new_new_n5897__, new_new_n5898__, new_new_n5899__, new_new_n5900__,
    new_new_n5901__, new_new_n5902__, new_new_n5903__, new_new_n5904__,
    new_new_n5905__, new_new_n5906__, new_new_n5907__, new_new_n5908__,
    new_new_n5909__, new_new_n5910__, new_new_n5911__, new_new_n5912__,
    new_new_n5913__, new_new_n5914__, new_new_n5915__, new_new_n5916__,
    new_new_n5917__, new_new_n5918__, new_new_n5919__, new_new_n5920__,
    new_new_n5921__, new_new_n5922__, new_new_n5923__, new_new_n5924__,
    new_new_n5925__, new_new_n5926__, new_new_n5927__, new_new_n5928__,
    new_new_n5929__, new_new_n5930__, new_new_n5931__, new_new_n5932__,
    new_new_n5933__, new_new_n5934__, new_new_n5935__, new_new_n5936__,
    new_new_n5937__, new_new_n5938__, new_new_n5939__, new_new_n5940__,
    new_new_n5941__, new_new_n5942__, new_new_n5943__, new_new_n5944__,
    new_new_n5945__, new_new_n5946__, new_new_n5947__, new_new_n5948__,
    new_new_n5949__, new_new_n5950__, new_new_n5951__, new_new_n5952__,
    new_new_n5953__, new_new_n5954__, new_new_n5955__, new_new_n5956__,
    new_new_n5957__, new_new_n5958__, new_new_n5959__, new_new_n5960__,
    new_new_n5961__, new_new_n5962__, new_new_n5963__, new_new_n5964__,
    new_new_n5965__, new_new_n5966__, new_new_n5967__, new_new_n5968__,
    new_new_n5969__, new_new_n5970__, new_new_n5971__, new_new_n5972__,
    new_new_n5973__, new_new_n5974__, new_new_n5975__, new_new_n5976__,
    new_new_n5977__, new_new_n5978__, new_new_n5979__, new_new_n5980__,
    new_new_n5981__, new_new_n5982__, new_new_n5983__, new_new_n5984__,
    new_new_n5985__, new_new_n5986__, new_new_n5987__, new_new_n5988__,
    new_new_n5989__, new_new_n5990__, new_new_n5991__, new_new_n5992__,
    new_new_n5993__, new_new_n5994__, new_new_n5995__, new_new_n5996__,
    new_new_n5997__, new_new_n5998__, new_new_n5999__, new_new_n6000__,
    new_new_n6001__, new_new_n6002__, new_new_n6003__, new_new_n6004__,
    new_new_n6005__, new_new_n6006__, new_new_n6007__, new_new_n6008__,
    new_new_n6009__, new_new_n6010__, new_new_n6011__, new_new_n6012__,
    new_new_n6013__, new_new_n6014__, new_new_n6015__, new_new_n6016__,
    new_new_n6017__, new_new_n6018__, new_new_n6019__, new_new_n6020__,
    new_new_n6021__, new_new_n6022__, new_new_n6023__, new_new_n6024__,
    new_new_n6025__, new_new_n6026__, new_new_n6027__, new_new_n6028__,
    new_new_n6029__, new_new_n6030__, new_new_n6031__, new_new_n6032__,
    new_new_n6033__, new_new_n6034__, new_new_n6035__, new_new_n6036__,
    new_new_n6037__, new_new_n6038__, new_new_n6039__, new_new_n6040__,
    new_new_n6041__, new_new_n6042__, new_new_n6043__, new_new_n6044__,
    new_new_n6045__, new_new_n6046__, new_new_n6047__, new_new_n6048__,
    new_new_n6049__, new_new_n6050__, new_new_n6051__, new_new_n6052__,
    new_new_n6053__, new_new_n6054__, new_new_n6055__, new_new_n6056__,
    new_new_n6057__, new_new_n6058__, new_new_n6059__, new_new_n6060__,
    new_new_n6061__, new_new_n6062__, new_new_n6063__, new_new_n6064__,
    new_new_n6065__, new_new_n6066__, new_new_n6067__, new_new_n6068__,
    new_new_n6069__, new_new_n6070__, new_new_n6071__, new_new_n6072__,
    new_new_n6073__, new_new_n6074__, new_new_n6075__, new_new_n6076__,
    new_new_n6077__, new_new_n6078__, new_new_n6079__, new_new_n6080__,
    new_new_n6081__, new_new_n6082__, new_new_n6083__, new_new_n6084__,
    new_new_n6085__, new_new_n6086__, new_new_n6087__, new_new_n6088__,
    new_new_n6089__, new_new_n6090__, new_new_n6091__, new_new_n6092__,
    new_new_n6093__, new_new_n6094__, new_new_n6095__, new_new_n6096__,
    new_new_n6097__, new_new_n6098__, new_new_n6099__, new_new_n6100__,
    new_new_n6101__, new_new_n6102__, new_new_n6103__, new_new_n6104__,
    new_new_n6105__, new_new_n6106__, new_new_n6107__, new_new_n6108__,
    new_new_n6109__, new_new_n6110__, new_new_n6111__, new_new_n6112__,
    new_new_n6113__, new_new_n6114__, new_new_n6115__, new_new_n6116__,
    new_new_n6117__, new_new_n6118__, new_new_n6119__, new_new_n6120__,
    new_new_n6121__, new_new_n6122__, new_new_n6123__, new_new_n6124__,
    new_new_n6125__, new_new_n6126__, new_new_n6127__, new_new_n6128__,
    new_new_n6129__, new_new_n6130__, new_new_n6131__, new_new_n6132__,
    new_new_n6133__, new_new_n6134__, new_new_n6135__, new_new_n6136__,
    new_new_n6137__, new_new_n6138__, new_new_n6139__, new_new_n6140__,
    new_new_n6141__, new_new_n6142__, new_new_n6143__, new_new_n6144__,
    new_new_n6145__, new_new_n6146__, new_new_n6147__, new_new_n6148__,
    new_new_n6149__, new_new_n6150__, new_new_n6151__, new_new_n6152__,
    new_new_n6153__, new_new_n6154__, new_new_n6155__, new_new_n6156__,
    new_new_n6157__, new_new_n6158__, new_new_n6159__, new_new_n6160__,
    new_new_n6161__, new_new_n6162__, new_new_n6163__, new_new_n6164__,
    new_new_n6165__, new_new_n6166__, new_new_n6167__, new_new_n6168__,
    new_new_n6169__, new_new_n6170__, new_new_n6171__, new_new_n6172__,
    new_new_n6173__, new_new_n6174__, new_new_n6175__, new_new_n6176__,
    new_new_n6177__, new_new_n6178__, new_new_n6179__, new_new_n6180__,
    new_new_n6181__, new_new_n6182__, new_new_n6183__, new_new_n6184__,
    new_new_n6185__, new_new_n6186__, new_new_n6187__, new_new_n6188__,
    new_new_n6189__, new_new_n6190__, new_new_n6191__, new_new_n6192__,
    new_new_n6193__, new_new_n6194__, new_new_n6195__, new_new_n6196__,
    new_new_n6197__, new_new_n6198__, new_new_n6199__, new_new_n6200__,
    new_new_n6201__, new_new_n6202__, new_new_n6203__, new_new_n6204__,
    new_new_n6205__, new_new_n6206__, new_new_n6207__, new_new_n6208__,
    new_new_n6209__, new_new_n6210__, new_new_n6211__, new_new_n6212__,
    new_new_n6213__, new_new_n6214__, new_new_n6215__, new_new_n6216__,
    new_new_n6217__, new_new_n6218__, new_new_n6219__, new_new_n6220__,
    new_new_n6221__, new_new_n6222__, new_new_n6223__, new_new_n6224__,
    new_new_n6225__, new_new_n6226__, new_new_n6227__, new_new_n6228__,
    new_new_n6229__, new_new_n6230__, new_new_n6231__, new_new_n6232__,
    new_new_n6233__, new_new_n6234__, new_new_n6235__, new_new_n6236__,
    new_new_n6237__, new_new_n6238__, new_new_n6239__, new_new_n6240__,
    new_new_n6241__, new_new_n6242__, new_new_n6243__, new_new_n6244__,
    new_new_n6245__, new_new_n6246__, new_new_n6247__, new_new_n6248__,
    new_new_n6249__, new_new_n6250__, new_new_n6251__, new_new_n6252__,
    new_new_n6253__, new_new_n6254__, new_new_n6255__, new_new_n6256__,
    new_new_n6257__, new_new_n6258__, new_new_n6259__, new_new_n6260__,
    new_new_n6261__, new_new_n6262__, new_new_n6263__, new_new_n6264__,
    new_new_n6265__, new_new_n6266__, new_new_n6267__, new_new_n6268__,
    new_new_n6269__, new_new_n6270__, new_new_n6271__, new_new_n6272__,
    new_new_n6273__, new_new_n6274__, new_new_n6275__, new_new_n6276__,
    new_new_n6277__, new_new_n6278__, new_new_n6279__, new_new_n6280__,
    new_new_n6281__, new_new_n6282__, new_new_n6283__, new_new_n6284__,
    new_new_n6285__, new_new_n6286__, new_new_n6287__, new_new_n6288__,
    new_new_n6289__, new_new_n6290__, new_new_n6291__, new_new_n6292__,
    new_new_n6293__, new_new_n6294__, new_new_n6295__, new_new_n6296__,
    new_new_n6297__, new_new_n6298__, new_new_n6299__, new_new_n6300__,
    new_new_n6301__, new_new_n6302__, new_new_n6303__, new_new_n6304__,
    new_new_n6305__, new_new_n6306__, new_new_n6307__, new_new_n6308__,
    new_new_n6309__, new_new_n6310__, new_new_n6311__, new_new_n6312__,
    new_new_n6313__, new_new_n6314__, new_new_n6315__, new_new_n6316__,
    new_new_n6317__, new_new_n6318__, new_new_n6319__, new_new_n6320__,
    new_new_n6321__, new_new_n6322__, new_new_n6323__, new_new_n6324__,
    new_new_n6325__, new_new_n6326__, new_new_n6327__, new_new_n6328__,
    new_new_n6329__, new_new_n6330__, new_new_n6331__, new_new_n6332__,
    new_new_n6333__, new_new_n6334__, new_new_n6335__, new_new_n6336__,
    new_new_n6337__, new_new_n6338__, new_new_n6339__, new_new_n6340__,
    new_new_n6341__, new_new_n6342__, new_new_n6343__, new_new_n6344__,
    new_new_n6345__, new_new_n6346__, new_new_n6347__, new_new_n6348__,
    new_new_n6349__, new_new_n6350__, new_new_n6351__, new_new_n6352__,
    new_new_n6353__, new_new_n6354__, new_new_n6355__, new_new_n6356__,
    new_new_n6357__, new_new_n6358__, new_new_n6359__, new_new_n6360__,
    new_new_n6361__, new_new_n6362__, new_new_n6363__, new_new_n6364__,
    new_new_n6365__, new_new_n6366__, new_new_n6367__, new_new_n6368__,
    new_new_n6369__, new_new_n6370__, new_new_n6371__, new_new_n6372__,
    new_new_n6373__, new_new_n6374__, new_new_n6375__, new_new_n6376__,
    new_new_n6377__, new_new_n6378__, new_new_n6379__, new_new_n6380__,
    new_new_n6381__, new_new_n6382__, new_new_n6383__, new_new_n6384__,
    new_new_n6385__, new_new_n6386__, new_new_n6387__, new_new_n6388__,
    new_new_n6389__, new_new_n6390__, new_new_n6391__, new_new_n6392__,
    new_new_n6393__, new_new_n6394__, new_new_n6395__, new_new_n6396__,
    new_new_n6397__, new_new_n6398__, new_new_n6399__, new_new_n6400__,
    new_new_n6401__, new_new_n6402__, new_new_n6403__, new_new_n6404__,
    new_new_n6405__, new_new_n6406__, new_new_n6407__, new_new_n6408__,
    new_new_n6409__, new_new_n6410__, new_new_n6411__, new_new_n6412__,
    new_new_n6413__, new_new_n6414__, new_new_n6415__, new_new_n6416__,
    new_new_n6417__, new_new_n6418__, new_new_n6419__, new_new_n6420__,
    new_new_n6421__, new_new_n6422__, new_new_n6423__, new_new_n6424__,
    new_new_n6425__, new_new_n6426__, new_new_n6427__, new_new_n6428__,
    new_new_n6429__, new_new_n6430__, new_new_n6431__, new_new_n6432__,
    new_new_n6433__, new_new_n6434__, new_new_n6435__, new_new_n6436__,
    new_new_n6437__, new_new_n6438__, new_new_n6439__, new_new_n6440__,
    new_new_n6441__, new_new_n6442__, new_new_n6443__, new_new_n6444__,
    new_new_n6445__, new_new_n6446__, new_new_n6447__, new_new_n6448__,
    new_new_n6449__, new_new_n6450__, new_new_n6451__, new_new_n6452__,
    new_new_n6453__, new_new_n6454__, new_new_n6455__, new_new_n6456__,
    new_new_n6457__, new_new_n6458__, new_new_n6459__, new_new_n6460__,
    new_new_n6461__, new_new_n6462__, new_new_n6463__, new_new_n6464__,
    new_new_n6465__, new_new_n6466__, new_new_n6467__, new_new_n6468__,
    new_new_n6469__, new_new_n6470__, new_new_n6471__, new_new_n6472__,
    new_new_n6473__, new_new_n6474__, new_new_n6475__, new_new_n6476__,
    new_new_n6477__, new_new_n6478__, new_new_n6479__, new_new_n6480__,
    new_new_n6481__, new_new_n6482__, new_new_n6483__, new_new_n6484__,
    new_new_n6485__, new_new_n6486__, new_new_n6487__, new_new_n6488__,
    new_new_n6489__, new_new_n6490__, new_new_n6491__, new_new_n6492__,
    new_new_n6493__, new_new_n6494__, new_new_n6495__, new_new_n6496__,
    new_new_n6497__, new_new_n6498__, new_new_n6499__, new_new_n6500__,
    new_new_n6501__, new_new_n6502__, new_new_n6503__, new_new_n6504__,
    new_new_n6505__, new_new_n6506__, new_new_n6507__, new_new_n6508__,
    new_new_n6509__, new_new_n6510__, new_new_n6511__, new_new_n6512__,
    new_new_n6513__, new_new_n6514__, new_new_n6515__, new_new_n6516__,
    new_new_n6517__, new_new_n6518__, new_new_n6519__, new_new_n6520__,
    new_new_n6521__, new_new_n6522__, new_new_n6523__, new_new_n6524__,
    new_new_n6525__, new_new_n6526__, new_new_n6527__, new_new_n6528__,
    new_new_n6529__, new_new_n6530__, new_new_n6531__, new_new_n6532__,
    new_new_n6533__, new_new_n6534__, new_new_n6535__, new_new_n6536__,
    new_new_n6537__, new_new_n6538__, new_new_n6539__, new_new_n6540__,
    new_new_n6541__, new_new_n6542__, new_new_n6543__, new_new_n6544__,
    new_new_n6545__, new_new_n6546__, new_new_n6547__, new_new_n6548__,
    new_new_n6549__, new_new_n6550__, new_new_n6551__, new_new_n6552__,
    new_new_n6553__, new_new_n6554__, new_new_n6555__, new_new_n6556__,
    new_new_n6557__, new_new_n6558__, new_new_n6559__, new_new_n6560__,
    new_new_n6561__, new_new_n6562__, new_new_n6563__, new_new_n6564__,
    new_new_n6565__, new_new_n6566__, new_new_n6567__, new_new_n6568__,
    new_new_n6569__, new_new_n6570__, new_new_n6571__, new_new_n6572__,
    new_new_n6573__, new_new_n6574__, new_new_n6575__, new_new_n6576__,
    new_new_n6577__, new_new_n6578__, new_new_n6579__, new_new_n6580__,
    new_new_n6581__, new_new_n6582__, new_new_n6583__, new_new_n6584__,
    new_new_n6585__, new_new_n6586__, new_new_n6587__, new_new_n6588__,
    new_new_n6589__, new_new_n6590__, new_new_n6591__, new_new_n6592__,
    new_new_n6593__, new_new_n6594__, new_new_n6595__, new_new_n6596__,
    new_new_n6597__, new_new_n6598__, new_new_n6599__, new_new_n6600__,
    new_new_n6601__, new_new_n6602__, new_new_n6603__, new_new_n6604__,
    new_new_n6605__, new_new_n6606__, new_new_n6607__, new_new_n6608__,
    new_new_n6609__, new_new_n6610__, new_new_n6611__, new_new_n6612__,
    new_new_n6613__, new_new_n6614__, new_new_n6615__, new_new_n6616__,
    new_new_n6617__, new_new_n6618__, new_new_n6619__, new_new_n6620__,
    new_new_n6621__, new_new_n6622__, new_new_n6623__, new_new_n6624__,
    new_new_n6625__, new_new_n6626__, new_new_n6627__, new_new_n6628__,
    new_new_n6629__, new_new_n6630__, new_new_n6631__, new_new_n6632__,
    new_new_n6633__, new_new_n6634__, new_new_n6635__, new_new_n6636__,
    new_new_n6637__, new_new_n6638__, new_new_n6639__, new_new_n6640__,
    new_new_n6641__, new_new_n6642__, new_new_n6643__, new_new_n6644__,
    new_new_n6645__, new_new_n6646__, new_new_n6647__, new_new_n6648__,
    new_new_n6649__, new_new_n6650__, new_new_n6651__, new_new_n6652__,
    new_new_n6653__, new_new_n6654__, new_new_n6655__, new_new_n6656__,
    new_new_n6657__, new_new_n6658__, new_new_n6659__, new_new_n6660__,
    new_new_n6661__, new_new_n6662__, new_new_n6663__, new_new_n6664__,
    new_new_n6665__, new_new_n6666__, new_new_n6667__, new_new_n6668__,
    new_new_n6669__, new_new_n6670__, new_new_n6671__, new_new_n6672__,
    new_new_n6673__, new_new_n6674__, new_new_n6675__, new_new_n6676__,
    new_new_n6677__, new_new_n6678__, new_new_n6679__, new_new_n6680__,
    new_new_n6681__, new_new_n6682__, new_new_n6683__, new_new_n6684__,
    new_new_n6685__, new_new_n6686__, new_new_n6687__, new_new_n6688__,
    new_new_n6689__, new_new_n6690__, new_new_n6691__, new_new_n6692__,
    new_new_n6693__, new_new_n6694__, new_new_n6695__, new_new_n6696__,
    new_new_n6697__, new_new_n6698__, new_new_n6699__, new_new_n6700__,
    new_new_n6701__, new_new_n6702__, new_new_n6703__, new_new_n6704__,
    new_new_n6705__, new_new_n6706__, new_new_n6707__, new_new_n6708__,
    new_new_n6709__, new_new_n6710__, new_new_n6711__, new_new_n6712__,
    new_new_n6713__, new_new_n6714__, new_new_n6715__, new_new_n6716__,
    new_new_n6717__, new_new_n6718__, new_new_n6719__, new_new_n6720__,
    new_new_n6721__, new_new_n6722__, new_new_n6723__, new_new_n6724__,
    new_new_n6725__, new_new_n6726__, new_new_n6727__, new_new_n6728__,
    new_new_n6729__, new_new_n6730__, new_new_n6731__, new_new_n6732__,
    new_new_n6733__, new_new_n6734__, new_new_n6735__, new_new_n6736__,
    new_new_n6737__, new_new_n6738__, new_new_n6739__, new_new_n6740__,
    new_new_n6741__, new_new_n6742__, new_new_n6743__, new_new_n6744__,
    new_new_n6745__, new_new_n6746__, new_new_n6747__, new_new_n6748__,
    new_new_n6749__, new_new_n6750__, new_new_n6751__, new_new_n6752__,
    new_new_n6753__, new_new_n6754__, new_new_n6755__, new_new_n6756__,
    new_new_n6757__, new_new_n6758__, new_new_n6759__, new_new_n6760__,
    new_new_n6761__, new_new_n6762__, new_new_n6763__, new_new_n6764__,
    new_new_n6765__, new_new_n6766__, new_new_n6767__, new_new_n6768__,
    new_new_n6769__, new_new_n6770__, new_new_n6771__, new_new_n6772__,
    new_new_n6773__, new_new_n6774__, new_new_n6775__, new_new_n6776__,
    new_new_n6777__, new_new_n6778__, new_new_n6779__, new_new_n6780__,
    new_new_n6781__, new_new_n6782__, new_new_n6783__, new_new_n6784__,
    new_new_n6785__, new_new_n6786__, new_new_n6787__, new_new_n6788__,
    new_new_n6789__, new_new_n6790__, new_new_n6791__, new_new_n6792__,
    new_new_n6793__, new_new_n6794__, new_new_n6795__, new_new_n6796__,
    new_new_n6797__, new_new_n6798__, new_new_n6799__, new_new_n6800__,
    new_new_n6801__, new_new_n6802__, new_new_n6803__, new_new_n6804__,
    new_new_n6805__, new_new_n6806__, new_new_n6807__, new_new_n6808__,
    new_new_n6809__, new_new_n6810__, new_new_n6811__, new_new_n6812__,
    new_new_n6813__, new_new_n6814__, new_new_n6815__, new_new_n6816__,
    new_new_n6817__, new_new_n6818__, new_new_n6819__, new_new_n6820__,
    new_new_n6821__, new_new_n6822__, new_new_n6823__, new_new_n6824__,
    new_new_n6825__, new_new_n6826__, new_new_n6827__, new_new_n6828__,
    new_new_n6829__, new_new_n6830__, new_new_n6831__, new_new_n6832__,
    new_new_n6833__, new_new_n6834__, new_new_n6835__, new_new_n6836__,
    new_new_n6837__, new_new_n6838__, new_new_n6839__, new_new_n6840__,
    new_new_n6841__, new_new_n6842__, new_new_n6843__, new_new_n6844__,
    new_new_n6845__, new_new_n6846__, new_new_n6847__, new_new_n6848__,
    new_new_n6849__, new_new_n6850__, new_new_n6851__, new_new_n6852__,
    new_new_n6853__, new_new_n6854__, new_new_n6855__, new_new_n6856__,
    new_new_n6857__, new_new_n6858__, new_new_n6859__, new_new_n6860__,
    new_new_n6861__, new_new_n6862__, new_new_n6863__, new_new_n6864__,
    new_new_n6865__, new_new_n6866__, new_new_n6867__, new_new_n6868__,
    new_new_n6869__, new_new_n6870__, new_new_n6871__, new_new_n6872__,
    new_new_n6873__, new_new_n6874__, new_new_n6875__, new_new_n6876__,
    new_new_n6877__, new_new_n6878__, new_new_n6879__, new_new_n6880__,
    new_new_n6881__, new_new_n6882__, new_new_n6883__, new_new_n6884__,
    new_new_n6885__, new_new_n6886__, new_new_n6887__, new_new_n6888__,
    new_new_n6889__, new_new_n6890__, new_new_n6891__, new_new_n6892__,
    new_new_n6893__, new_new_n6894__, new_new_n6895__, new_new_n6896__,
    new_new_n6897__, new_new_n6898__, new_new_n6899__, new_new_n6900__,
    new_new_n6901__, new_new_n6902__, new_new_n6903__, new_new_n6904__,
    new_new_n6905__, new_new_n6906__, new_new_n6907__, new_new_n6908__,
    new_new_n6909__, new_new_n6910__, new_new_n6911__, new_new_n6912__,
    new_new_n6913__, new_new_n6914__, new_new_n6915__, new_new_n6916__,
    new_new_n6917__, new_new_n6918__, new_new_n6919__, new_new_n6920__,
    new_new_n6921__, new_new_n6922__, new_new_n6923__, new_new_n6924__,
    new_new_n6925__, new_new_n6926__, new_new_n6927__, new_new_n6928__,
    new_new_n6929__, new_new_n6930__, new_new_n6931__, new_new_n6932__,
    new_new_n6933__, new_new_n6934__, new_new_n6935__, new_new_n6936__,
    new_new_n6937__, new_new_n6938__, new_new_n6939__, new_new_n6940__,
    new_new_n6941__, new_new_n6942__, new_new_n6943__, new_new_n6944__,
    new_new_n6945__, new_new_n6946__, new_new_n6947__, new_new_n6948__,
    new_new_n6949__, new_new_n6950__, new_new_n6951__, new_new_n6952__,
    new_new_n6953__, new_new_n6954__, new_new_n6955__, new_new_n6956__,
    new_new_n6957__, new_new_n6958__, new_new_n6959__, new_new_n6960__,
    new_new_n6961__, new_new_n6962__, new_new_n6963__, new_new_n6964__,
    new_new_n6965__, new_new_n6966__, new_new_n6967__, new_new_n6968__,
    new_new_n6969__, new_new_n6970__, new_new_n6971__, new_new_n6972__,
    new_new_n6973__, new_new_n6974__, new_new_n6975__, new_new_n6976__,
    new_new_n6977__, new_new_n6978__, new_new_n6979__, new_new_n6980__,
    new_new_n6981__, new_new_n6982__, new_new_n6983__, new_new_n6984__,
    new_new_n6985__, new_new_n6986__, new_new_n6987__, new_new_n6988__,
    new_new_n6989__, new_new_n6990__, new_new_n6991__, new_new_n6992__,
    new_new_n6993__, new_new_n6994__, new_new_n6995__, new_new_n6996__,
    new_new_n6997__, new_new_n6998__, new_new_n6999__, new_new_n7000__,
    new_new_n7001__, new_new_n7002__, new_new_n7003__, new_new_n7004__,
    new_new_n7005__, new_new_n7006__, new_new_n7007__, new_new_n7008__,
    new_new_n7009__, new_new_n7010__, new_new_n7011__, new_new_n7012__,
    new_new_n7013__, new_new_n7014__, new_new_n7015__, new_new_n7016__,
    new_new_n7017__, new_new_n7018__, new_new_n7019__, new_new_n7020__,
    new_new_n7021__, new_new_n7022__, new_new_n7023__, new_new_n7024__,
    new_new_n7025__, new_new_n7026__, new_new_n7027__, new_new_n7028__,
    new_new_n7029__, new_new_n7030__, new_new_n7031__, new_new_n7032__,
    new_new_n7033__, new_new_n7034__, new_new_n7035__, new_new_n7036__,
    new_new_n7037__, new_new_n7038__, new_new_n7039__, new_new_n7040__,
    new_new_n7041__, new_new_n7042__, new_new_n7043__, new_new_n7044__,
    new_new_n7045__, new_new_n7046__, new_new_n7047__, new_new_n7048__,
    new_new_n7049__, new_new_n7050__, new_new_n7051__, new_new_n7052__,
    new_new_n7053__, new_new_n7054__, new_new_n7055__, new_new_n7056__,
    new_new_n7057__, new_new_n7058__, new_new_n7059__, new_new_n7060__,
    new_new_n7061__, new_new_n7062__, new_new_n7063__, new_new_n7064__,
    new_new_n7065__, new_new_n7066__, new_new_n7067__, new_new_n7068__,
    new_new_n7069__, new_new_n7070__, new_new_n7071__, new_new_n7072__,
    new_new_n7073__, new_new_n7074__, new_new_n7075__, new_new_n7076__,
    new_new_n7077__, new_new_n7078__, new_new_n7079__, new_new_n7080__,
    new_new_n7081__, new_new_n7082__, new_new_n7083__, new_new_n7084__,
    new_new_n7085__, new_new_n7086__, new_new_n7087__, new_new_n7088__,
    new_new_n7089__, new_new_n7090__, new_new_n7091__, new_new_n7092__,
    new_new_n7093__, new_new_n7094__, new_new_n7095__, new_new_n7096__,
    new_new_n7097__, new_new_n7098__, new_new_n7099__, new_new_n7100__,
    new_new_n7101__, new_new_n7102__, new_new_n7103__, new_new_n7104__,
    new_new_n7105__, new_new_n7106__, new_new_n7107__, new_new_n7108__,
    new_new_n7109__, new_new_n7110__, new_new_n7111__, new_new_n7112__,
    new_new_n7113__, new_new_n7114__, new_new_n7115__, new_new_n7116__,
    new_new_n7117__, new_new_n7118__, new_new_n7119__, new_new_n7120__,
    new_new_n7121__, new_new_n7122__, new_new_n7123__, new_new_n7124__,
    new_new_n7125__, new_new_n7126__, new_new_n7127__, new_new_n7128__,
    new_new_n7129__, new_new_n7130__, new_new_n7131__, new_new_n7132__,
    new_new_n7133__, new_new_n7134__, new_new_n7135__, new_new_n7136__,
    new_new_n7137__, new_new_n7138__, new_new_n7139__, new_new_n7140__,
    new_new_n7141__, new_new_n7142__, new_new_n7143__, new_new_n7144__,
    new_new_n7145__, new_new_n7146__, new_new_n7147__, new_new_n7148__,
    new_new_n7149__, new_new_n7150__, new_new_n7151__, new_new_n7152__,
    new_new_n7153__, new_new_n7154__, new_new_n7155__, new_new_n7156__,
    new_new_n7157__, new_new_n7158__, new_new_n7159__, new_new_n7160__,
    new_new_n7161__, new_new_n7162__, new_new_n7163__, new_new_n7164__,
    new_new_n7165__, new_new_n7166__, new_new_n7167__, new_new_n7168__,
    new_new_n7169__, new_new_n7170__, new_new_n7171__, new_new_n7172__,
    new_new_n7173__, new_new_n7174__, new_new_n7175__, new_new_n7176__,
    new_new_n7177__, new_new_n7178__, new_new_n7179__, new_new_n7180__,
    new_new_n7181__, new_new_n7182__, new_new_n7183__, new_new_n7184__,
    new_new_n7185__, new_new_n7186__, new_new_n7187__, new_new_n7188__,
    new_new_n7189__, new_new_n7190__, new_new_n7191__, new_new_n7192__,
    new_new_n7193__, new_new_n7194__, new_new_n7195__, new_new_n7196__,
    new_new_n7197__, new_new_n7198__, new_new_n7199__, new_new_n7200__,
    new_new_n7201__, new_new_n7202__, new_new_n7203__, new_new_n7204__,
    new_new_n7205__, new_new_n7206__, new_new_n7207__, new_new_n7208__,
    new_new_n7209__, new_new_n7210__, new_new_n7211__, new_new_n7212__,
    new_new_n7213__, new_new_n7214__, new_new_n7215__, new_new_n7216__,
    new_new_n7217__, new_new_n7218__, new_new_n7219__, new_new_n7220__,
    new_new_n7221__, new_new_n7222__, new_new_n7223__, new_new_n7224__,
    new_new_n7225__, new_new_n7226__, new_new_n7227__, new_new_n7228__,
    new_new_n7229__, new_new_n7230__, new_new_n7231__, new_new_n7232__,
    new_new_n7233__, new_new_n7234__, new_new_n7235__, new_new_n7236__,
    new_new_n7237__, new_new_n7238__, new_new_n7239__, new_new_n7240__,
    new_new_n7241__, new_new_n7242__, new_new_n7243__, new_new_n7244__,
    new_new_n7245__, new_new_n7246__, new_new_n7247__, new_new_n7248__,
    new_new_n7249__, new_new_n7250__, new_new_n7251__, new_new_n7252__,
    new_new_n7253__, new_new_n7254__, new_new_n7255__, new_new_n7256__,
    new_new_n7257__, new_new_n7258__, new_new_n7259__, new_new_n7260__,
    new_new_n7261__, new_new_n7262__, new_new_n7263__, new_new_n7264__,
    new_new_n7265__, new_new_n7266__, new_new_n7267__, new_new_n7268__,
    new_new_n7269__, new_new_n7270__, new_new_n7271__, new_new_n7272__,
    new_new_n7273__, new_new_n7274__, new_new_n7275__, new_new_n7276__,
    new_new_n7277__, new_new_n7278__, new_new_n7279__, new_new_n7280__,
    new_new_n7281__, new_new_n7282__, new_new_n7283__, new_new_n7284__,
    new_new_n7285__, new_new_n7286__, new_new_n7287__, new_new_n7288__,
    new_new_n7289__, new_new_n7290__, new_new_n7291__, new_new_n7292__,
    new_new_n7293__, new_new_n7294__, new_new_n7295__, new_new_n7296__,
    new_new_n7297__, new_new_n7298__, new_new_n7299__, new_new_n7300__,
    new_new_n7301__, new_new_n7302__, new_new_n7303__, new_new_n7304__,
    new_new_n7305__, new_new_n7306__, new_new_n7307__, new_new_n7308__,
    new_new_n7309__, new_new_n7310__, new_new_n7311__, new_new_n7312__,
    new_new_n7313__, new_new_n7314__, new_new_n7315__, new_new_n7316__,
    new_new_n7317__, new_new_n7318__, new_new_n7319__, new_new_n7320__,
    new_new_n7321__, new_new_n7322__, new_new_n7323__, new_new_n7324__,
    new_new_n7325__, new_new_n7326__, new_new_n7327__, new_new_n7328__,
    new_new_n7329__, new_new_n7330__, new_new_n7331__, new_new_n7332__,
    new_new_n7333__, new_new_n7334__, new_new_n7335__, new_new_n7336__,
    new_new_n7337__, new_new_n7338__, new_new_n7339__, new_new_n7340__,
    new_new_n7341__, new_new_n7342__, new_new_n7343__, new_new_n7344__,
    new_new_n7345__, new_new_n7346__, new_new_n7347__, new_new_n7348__,
    new_new_n7349__, new_new_n7350__, new_new_n7351__, new_new_n7352__,
    new_new_n7353__, new_new_n7354__, new_new_n7355__, new_new_n7356__,
    new_new_n7357__, new_new_n7358__, new_new_n7359__, new_new_n7360__,
    new_new_n7361__, new_new_n7362__, new_new_n7363__, new_new_n7364__,
    new_new_n7365__, new_new_n7366__, new_new_n7367__, new_new_n7368__,
    new_new_n7369__, new_new_n7370__, new_new_n7371__, new_new_n7372__,
    new_new_n7373__, new_new_n7374__, new_new_n7375__, new_new_n7376__,
    new_new_n7377__, new_new_n7378__, new_new_n7379__, new_new_n7380__,
    new_new_n7381__, new_new_n7382__, new_new_n7383__, new_new_n7384__,
    new_new_n7385__, new_new_n7386__, new_new_n7387__, new_new_n7388__,
    new_new_n7389__, new_new_n7390__, new_new_n7391__, new_new_n7392__,
    new_new_n7393__, new_new_n7394__, new_new_n7395__, new_new_n7396__,
    new_new_n7397__, new_new_n7398__, new_new_n7399__, new_new_n7400__,
    new_new_n7401__, new_new_n7402__, new_new_n7403__, new_new_n7404__,
    new_new_n7405__, new_new_n7406__, new_new_n7407__, new_new_n7408__,
    new_new_n7409__, new_new_n7410__, new_new_n7411__, new_new_n7412__,
    new_new_n7413__, new_new_n7414__, new_new_n7415__, new_new_n7416__,
    new_new_n7417__, new_new_n7418__, new_new_n7419__, new_new_n7420__,
    new_new_n7421__, new_new_n7422__, new_new_n7423__, new_new_n7424__,
    new_new_n7425__, new_new_n7426__, new_new_n7427__, new_new_n7428__,
    new_new_n7429__, new_new_n7430__, new_new_n7431__, new_new_n7432__,
    new_new_n7433__, new_new_n7434__, new_new_n7435__, new_new_n7436__,
    new_new_n7437__, new_new_n7438__, new_new_n7439__, new_new_n7440__,
    new_new_n7441__, new_new_n7442__, new_new_n7443__, new_new_n7444__,
    new_new_n7445__, new_new_n7446__, new_new_n7447__, new_new_n7448__,
    new_new_n7449__, new_new_n7450__, new_new_n7451__, new_new_n7452__,
    new_new_n7453__, new_new_n7454__, new_new_n7455__, new_new_n7456__,
    new_new_n7457__, new_new_n7458__, new_new_n7459__, new_new_n7460__,
    new_new_n7461__, new_new_n7462__, new_new_n7463__, new_new_n7464__,
    new_new_n7465__, new_new_n7466__, new_new_n7467__, new_new_n7468__,
    new_new_n7469__, new_new_n7470__, new_new_n7471__, new_new_n7472__,
    new_new_n7473__, new_new_n7474__, new_new_n7475__, new_new_n7476__,
    new_new_n7477__, new_new_n7478__, new_new_n7479__, new_new_n7480__,
    new_new_n7481__, new_new_n7482__, new_new_n7483__, new_new_n7484__,
    new_new_n7485__, new_new_n7486__, new_new_n7487__, new_new_n7488__,
    new_new_n7489__, new_new_n7490__, new_new_n7491__, new_new_n7492__,
    new_new_n7493__, new_new_n7494__, new_new_n7495__, new_new_n7496__,
    new_new_n7497__, new_new_n7498__, new_new_n7499__, new_new_n7500__,
    new_new_n7501__, new_new_n7502__, new_new_n7503__, new_new_n7504__,
    new_new_n7505__, new_new_n7506__, new_new_n7507__, new_new_n7508__,
    new_new_n7509__, new_new_n7510__, new_new_n7511__, new_new_n7512__,
    new_new_n7513__, new_new_n7514__, new_new_n7515__, new_new_n7516__,
    new_new_n7517__, new_new_n7518__, new_new_n7519__, new_new_n7520__,
    new_new_n7521__, new_new_n7522__, new_new_n7523__, new_new_n7524__,
    new_new_n7525__, new_new_n7526__, new_new_n7527__, new_new_n7528__,
    new_new_n7529__, new_new_n7530__, new_new_n7531__, new_new_n7532__,
    new_new_n7533__, new_new_n7534__, new_new_n7535__, new_new_n7536__,
    new_new_n7537__, new_new_n7538__, new_new_n7539__, new_new_n7540__,
    new_new_n7541__, new_new_n7542__, new_new_n7543__, new_new_n7544__,
    new_new_n7545__, new_new_n7546__, new_new_n7547__, new_new_n7548__,
    new_new_n7549__, new_new_n7550__, new_new_n7551__, new_new_n7552__,
    new_new_n7553__, new_new_n7554__, new_new_n7555__, new_new_n7556__,
    new_new_n7557__, new_new_n7558__, new_new_n7559__, new_new_n7560__,
    new_new_n7561__, new_new_n7562__, new_new_n7563__, new_new_n7564__,
    new_new_n7565__, new_new_n7566__, new_new_n7567__, new_new_n7568__,
    new_new_n7569__, new_new_n7570__, new_new_n7571__, new_new_n7572__,
    new_new_n7573__, new_new_n7574__, new_new_n7575__, new_new_n7576__,
    new_new_n7577__, new_new_n7578__, new_new_n7579__, new_new_n7580__,
    new_new_n7581__, new_new_n7582__, new_new_n7583__, new_new_n7584__,
    new_new_n7585__, new_new_n7586__, new_new_n7587__, new_new_n7588__,
    new_new_n7589__, new_new_n7590__, new_new_n7591__, new_new_n7592__,
    new_new_n7593__, new_new_n7594__, new_new_n7595__, new_new_n7596__,
    new_new_n7597__, new_new_n7598__, new_new_n7599__, new_new_n7600__,
    new_new_n7601__, new_new_n7602__, new_new_n7603__, new_new_n7604__,
    new_new_n7605__, new_new_n7606__, new_new_n7607__, new_new_n7608__,
    new_new_n7609__, new_new_n7610__, new_new_n7611__, new_new_n7612__,
    new_new_n7613__, new_new_n7614__, new_new_n7615__, new_new_n7616__,
    new_new_n7617__, new_new_n7618__, new_new_n7619__, new_new_n7620__,
    new_new_n7621__, new_new_n7622__, new_new_n7623__, new_new_n7624__,
    new_new_n7625__, new_new_n7626__, new_new_n7627__, new_new_n7628__,
    new_new_n7629__, new_new_n7630__, new_new_n7631__, new_new_n7632__,
    new_new_n7633__, new_new_n7634__, new_new_n7635__, new_new_n7636__,
    new_new_n7637__, new_new_n7638__, new_new_n7639__, new_new_n7640__,
    new_new_n7641__, new_new_n7642__, new_new_n7643__, new_new_n7644__,
    new_new_n7645__, new_new_n7646__, new_new_n7647__, new_new_n7648__,
    new_new_n7649__, new_new_n7650__, new_new_n7651__, new_new_n7652__,
    new_new_n7653__, new_new_n7654__, new_new_n7655__, new_new_n7656__,
    new_new_n7657__, new_new_n7658__, new_new_n7659__, new_new_n7660__,
    new_new_n7661__, new_new_n7662__, new_new_n7663__, new_new_n7664__,
    new_new_n7665__, new_new_n7666__, new_new_n7667__, new_new_n7668__,
    new_new_n7669__, new_new_n7670__, new_new_n7671__, new_new_n7672__,
    new_new_n7673__, new_new_n7674__, new_new_n7675__, new_new_n7676__,
    new_new_n7677__, new_new_n7678__, new_new_n7679__, new_new_n7680__,
    new_new_n7681__, new_new_n7682__, new_new_n7683__, new_new_n7684__,
    new_new_n7685__, new_new_n7686__, new_new_n7687__, new_new_n7688__,
    new_new_n7689__, new_new_n7690__, new_new_n7691__, new_new_n7692__,
    new_new_n7693__, new_new_n7694__, new_new_n7695__, new_new_n7696__,
    new_new_n7697__, new_new_n7698__, new_new_n7699__, new_new_n7700__,
    new_new_n7701__, new_new_n7702__, new_new_n7703__, new_new_n7704__,
    new_new_n7705__, new_new_n7706__, new_new_n7707__, new_new_n7708__,
    new_new_n7709__, new_new_n7710__, new_new_n7711__, new_new_n7712__,
    new_new_n7713__, new_new_n7714__, new_new_n7715__, new_new_n7716__,
    new_new_n7717__, new_new_n7718__, new_new_n7719__, new_new_n7720__,
    new_new_n7721__, new_new_n7722__, new_new_n7723__, new_new_n7724__,
    new_new_n7725__, new_new_n7726__, new_new_n7727__, new_new_n7728__,
    new_new_n7729__, new_new_n7730__, new_new_n7731__, new_new_n7732__,
    new_new_n7733__, new_new_n7734__, new_new_n7735__, new_new_n7736__,
    new_new_n7737__, new_new_n7738__, new_new_n7739__, new_new_n7740__,
    new_new_n7741__, new_new_n7742__, new_new_n7743__, new_new_n7744__,
    new_new_n7745__, new_new_n7746__, new_new_n7747__, new_new_n7748__,
    new_new_n7749__, new_new_n7750__, new_new_n7751__, new_new_n7752__,
    new_new_n7753__, new_new_n7754__, new_new_n7755__, new_new_n7756__,
    new_new_n7757__, new_new_n7758__, new_new_n7759__, new_new_n7760__,
    new_new_n7761__, new_new_n7762__, new_new_n7763__, new_new_n7764__,
    new_new_n7765__, new_new_n7766__, new_new_n7767__, new_new_n7768__,
    new_new_n7769__, new_new_n7770__, new_new_n7771__, new_new_n7772__,
    new_new_n7773__, new_new_n7774__, new_new_n7775__, new_new_n7776__,
    new_new_n7777__, new_new_n7778__, new_new_n7779__, new_new_n7780__,
    new_new_n7781__, new_new_n7782__, new_new_n7783__, new_new_n7784__,
    new_new_n7785__, new_new_n7786__, new_new_n7787__, new_new_n7788__,
    new_new_n7789__, new_new_n7790__, new_new_n7791__, new_new_n7792__,
    new_new_n7793__, new_new_n7794__, new_new_n7795__, new_new_n7796__,
    new_new_n7797__, new_new_n7798__, new_new_n7799__, new_new_n7800__,
    new_new_n7801__, new_new_n7802__, new_new_n7803__, new_new_n7804__,
    new_new_n7805__, new_new_n7806__, new_new_n7807__, new_new_n7808__,
    new_new_n7809__, new_new_n7810__, new_new_n7811__, new_new_n7812__,
    new_new_n7813__, new_new_n7814__, new_new_n7815__, new_new_n7816__,
    new_new_n7817__, new_new_n7818__, new_new_n7819__, new_new_n7820__,
    new_new_n7821__, new_new_n7822__, new_new_n7823__, new_new_n7824__,
    new_new_n7825__, new_new_n7826__, new_new_n7827__, new_new_n7828__,
    new_new_n7829__, new_new_n7830__, new_new_n7831__, new_new_n7832__,
    new_new_n7833__, new_new_n7834__, new_new_n7835__, new_new_n7836__,
    new_new_n7837__, new_new_n7838__, new_new_n7839__, new_new_n7840__,
    new_new_n7841__, new_new_n7842__, new_new_n7843__, new_new_n7844__,
    new_new_n7845__, new_new_n7846__, new_new_n7847__, new_new_n7848__,
    new_new_n7849__, new_new_n7850__, new_new_n7851__, new_new_n7852__,
    new_new_n7853__, new_new_n7854__, new_new_n7855__, new_new_n7856__,
    new_new_n7857__, new_new_n7858__, new_new_n7859__, new_new_n7860__,
    new_new_n7861__, new_new_n7862__, new_new_n7863__, new_new_n7864__,
    new_new_n7865__, new_new_n7866__, new_new_n7867__, new_new_n7868__,
    new_new_n7869__, new_new_n7870__, new_new_n7871__, new_new_n7872__,
    new_new_n7873__, new_new_n7874__, new_new_n7875__, new_new_n7876__,
    new_new_n7877__, new_new_n7878__, new_new_n7879__, new_new_n7880__,
    new_new_n7881__, new_new_n7882__, new_new_n7883__, new_new_n7884__,
    new_new_n7885__, new_new_n7886__, new_new_n7887__, new_new_n7888__,
    new_new_n7889__, new_new_n7890__, new_new_n7891__, new_new_n7892__,
    new_new_n7893__, new_new_n7894__, new_new_n7895__, new_new_n7896__,
    new_new_n7897__, new_new_n7898__, new_new_n7899__, new_new_n7900__,
    new_new_n7901__, new_new_n7902__, new_new_n7903__, new_new_n7904__,
    new_new_n7905__, new_new_n7906__, new_new_n7907__, new_new_n7908__,
    new_new_n7909__, new_new_n7910__, new_new_n7911__, new_new_n7912__,
    new_new_n7913__, new_new_n7914__, new_new_n7915__, new_new_n7916__,
    new_new_n7917__, new_new_n7918__, new_new_n7919__, new_new_n7920__,
    new_new_n7921__, new_new_n7922__, new_new_n7923__, new_new_n7924__,
    new_new_n7925__, new_new_n7926__, new_new_n7927__, new_new_n7928__,
    new_new_n7929__, new_new_n7930__, new_new_n7931__, new_new_n7932__,
    new_new_n7933__, new_new_n7934__, new_new_n7935__, new_new_n7936__,
    new_new_n7937__, new_new_n7938__, new_new_n7939__, new_new_n7940__,
    new_new_n7941__, new_new_n7942__, new_new_n7943__, new_new_n7944__,
    new_new_n7945__, new_new_n7946__, new_new_n7947__, new_new_n7948__,
    new_new_n7949__, new_new_n7950__, new_new_n7951__, new_new_n7952__,
    new_new_n7953__, new_new_n7954__, new_new_n7955__, new_new_n7956__,
    new_new_n7957__, new_new_n7958__, new_new_n7959__, new_new_n7960__,
    new_new_n7961__, new_new_n7962__, new_new_n7963__, new_new_n7964__,
    new_new_n7965__, new_new_n7966__, new_new_n7967__, new_new_n7968__,
    new_new_n7969__, new_new_n7970__, new_new_n7971__, new_new_n7972__,
    new_new_n7973__, new_new_n7974__, new_new_n7975__, new_new_n7976__,
    new_new_n7977__, new_new_n7978__, new_new_n7979__, new_new_n7980__,
    new_new_n7981__, new_new_n7982__, new_new_n7983__, new_new_n7984__,
    new_new_n7985__, new_new_n7986__, new_new_n7987__, new_new_n7988__,
    new_new_n7989__, new_new_n7990__, new_new_n7991__, new_new_n7992__,
    new_new_n7993__, new_new_n7994__, new_new_n7995__, new_new_n7996__,
    new_new_n7997__, new_new_n7998__, new_new_n7999__, new_new_n8000__,
    new_new_n8001__, new_new_n8002__, new_new_n8003__, new_new_n8004__,
    new_new_n8005__, new_new_n8006__, new_new_n8007__, new_new_n8008__,
    new_new_n8009__, new_new_n8010__, new_new_n8011__, new_new_n8012__,
    new_new_n8013__, new_new_n8014__, new_new_n8015__, new_new_n8016__,
    new_new_n8017__, new_new_n8018__, new_new_n8019__, new_new_n8020__,
    new_new_n8021__, new_new_n8022__, new_new_n8023__, new_new_n8024__,
    new_new_n8025__, new_new_n8026__, new_new_n8027__, new_new_n8028__,
    new_new_n8029__, new_new_n8030__, new_new_n8031__, new_new_n8032__,
    new_new_n8033__, new_new_n8034__, new_new_n8035__, new_new_n8036__,
    new_new_n8037__, new_new_n8038__, new_new_n8039__, new_new_n8040__,
    new_new_n8041__, new_new_n8042__, new_new_n8043__, new_new_n8044__,
    new_new_n8045__, new_new_n8046__, new_new_n8047__, new_new_n8048__,
    new_new_n8049__, new_new_n8050__, new_new_n8051__, new_new_n8052__,
    new_new_n8053__, new_new_n8054__, new_new_n8055__, new_new_n8056__,
    new_new_n8057__, new_new_n8058__, new_new_n8059__, new_new_n8060__,
    new_new_n8061__, new_new_n8062__, new_new_n8063__, new_new_n8064__,
    new_new_n8065__, new_new_n8066__, new_new_n8067__, new_new_n8068__,
    new_new_n8069__, new_new_n8070__, new_new_n8071__, new_new_n8072__,
    new_new_n8073__, new_new_n8074__, new_new_n8075__, new_new_n8076__,
    new_new_n8077__, new_new_n8078__, new_new_n8079__, new_new_n8080__,
    new_new_n8081__, new_new_n8082__, new_new_n8083__, new_new_n8084__,
    new_new_n8085__, new_new_n8086__, new_new_n8087__, new_new_n8088__,
    new_new_n8089__, new_new_n8090__, new_new_n8091__, new_new_n8092__,
    new_new_n8093__, new_new_n8094__, new_new_n8095__, new_new_n8096__,
    new_new_n8097__, new_new_n8098__, new_new_n8099__, new_new_n8100__,
    new_new_n8101__, new_new_n8102__, new_new_n8103__, new_new_n8104__,
    new_new_n8105__, new_new_n8106__, new_new_n8107__, new_new_n8108__,
    new_new_n8109__, new_new_n8110__, new_new_n8111__, new_new_n8112__,
    new_new_n8113__, new_new_n8114__, new_new_n8115__, new_new_n8116__,
    new_new_n8117__, new_new_n8118__, new_new_n8119__, new_new_n8120__,
    new_new_n8121__, new_new_n8122__, new_new_n8123__, new_new_n8124__,
    new_new_n8125__, new_new_n8126__, new_new_n8127__, new_new_n8128__,
    new_new_n8129__, new_new_n8130__, new_new_n8131__, new_new_n8132__,
    new_new_n8133__, new_new_n8134__, new_new_n8135__, new_new_n8136__,
    new_new_n8137__, new_new_n8138__, new_new_n8139__, new_new_n8140__,
    new_new_n8141__, new_new_n8142__, new_new_n8143__, new_new_n8144__,
    new_new_n8145__, new_new_n8146__, new_new_n8147__, new_new_n8148__,
    new_new_n8149__, new_new_n8150__, new_new_n8151__, new_new_n8152__,
    new_new_n8153__, new_new_n8154__, new_new_n8155__, new_new_n8156__,
    new_new_n8157__, new_new_n8158__, new_new_n8159__, new_new_n8160__,
    new_new_n8161__, new_new_n8162__, new_new_n8163__, new_new_n8164__,
    new_new_n8165__, new_new_n8166__, new_new_n8167__, new_new_n8168__,
    new_new_n8169__, new_new_n8170__, new_new_n8171__, new_new_n8172__,
    new_new_n8173__, new_new_n8174__, new_new_n8175__, new_new_n8176__,
    new_new_n8177__, new_new_n8178__, new_new_n8179__, new_new_n8180__,
    new_new_n8181__, new_new_n8182__, new_new_n8183__, new_new_n8184__,
    new_new_n8185__, new_new_n8186__, new_new_n8187__, new_new_n8188__,
    new_new_n8189__, new_new_n8190__, new_new_n8191__, new_new_n8192__,
    new_new_n8193__, new_new_n8194__, new_new_n8195__, new_new_n8196__,
    new_new_n8197__, new_new_n8198__, new_new_n8199__, new_new_n8200__,
    new_new_n8201__, new_new_n8202__, new_new_n8203__, new_new_n8204__,
    new_new_n8205__, new_new_n8206__, new_new_n8207__, new_new_n8208__,
    new_new_n8209__, new_new_n8210__, new_new_n8211__, new_new_n8212__,
    new_new_n8213__, new_new_n8214__, new_new_n8215__, new_new_n8216__,
    new_new_n8217__, new_new_n8218__, new_new_n8219__, new_new_n8220__,
    new_new_n8221__, new_new_n8222__, new_new_n8223__, new_new_n8224__,
    new_new_n8225__, new_new_n8226__, new_new_n8227__, new_new_n8228__,
    new_new_n8229__, new_new_n8230__, new_new_n8231__, new_new_n8232__,
    new_new_n8233__, new_new_n8234__, new_new_n8235__, new_new_n8236__,
    new_new_n8237__, new_new_n8238__, new_new_n8239__, new_new_n8240__,
    new_new_n8241__, new_new_n8242__, new_new_n8243__, new_new_n8244__,
    new_new_n8245__, new_new_n8246__, new_new_n8247__, new_new_n8248__,
    new_new_n8249__, new_new_n8250__, new_new_n8251__, new_new_n8252__,
    new_new_n8253__, new_new_n8254__, new_new_n8255__, new_new_n8256__,
    new_new_n8257__, new_new_n8258__, new_new_n8259__, new_new_n8260__,
    new_new_n8261__, new_new_n8262__, new_new_n8263__, new_new_n8264__,
    new_new_n8265__, new_new_n8266__, new_new_n8267__, new_new_n8268__,
    new_new_n8269__, new_new_n8270__, new_new_n8271__, new_new_n8272__,
    new_new_n8273__, new_new_n8274__, new_new_n8275__, new_new_n8276__,
    new_new_n8277__, new_new_n8278__, new_new_n8279__, new_new_n8280__,
    new_new_n8281__, new_new_n8282__, new_new_n8283__, new_new_n8284__,
    new_new_n8285__, new_new_n8286__, new_new_n8287__, new_new_n8288__,
    new_new_n8289__, new_new_n8290__, new_new_n8291__, new_new_n8292__,
    new_new_n8293__, new_new_n8294__, new_new_n8295__, new_new_n8296__,
    new_new_n8297__, new_new_n8298__, new_new_n8299__, new_new_n8300__,
    new_new_n8301__, new_new_n8302__, new_new_n8303__, new_new_n8304__,
    new_new_n8305__, new_new_n8306__, new_new_n8307__, new_new_n8308__,
    new_new_n8309__, new_new_n8310__, new_new_n8311__, new_new_n8312__,
    new_new_n8313__, new_new_n8314__, new_new_n8315__, new_new_n8316__,
    new_new_n8317__, new_new_n8318__, new_new_n8319__, new_new_n8320__,
    new_new_n8321__, new_new_n8322__, new_new_n8323__, new_new_n8324__,
    new_new_n8325__, new_new_n8326__, new_new_n8327__, new_new_n8328__,
    new_new_n8329__, new_new_n8330__, new_new_n8331__, new_new_n8332__,
    new_new_n8333__, new_new_n8334__, new_new_n8335__, new_new_n8336__,
    new_new_n8337__, new_new_n8338__, new_new_n8339__, new_new_n8340__,
    new_new_n8341__, new_new_n8342__, new_new_n8343__, new_new_n8344__,
    new_new_n8345__, new_new_n8346__, new_new_n8347__, new_new_n8348__,
    new_new_n8349__, new_new_n8350__, new_new_n8351__, new_new_n8352__,
    new_new_n8353__, new_new_n8354__, new_new_n8355__, new_new_n8356__,
    new_new_n8357__, new_new_n8358__, new_new_n8359__, new_new_n8360__,
    new_new_n8361__, new_new_n8362__, new_new_n8363__, new_new_n8364__,
    new_new_n8365__, new_new_n8366__, new_new_n8367__, new_new_n8368__,
    new_new_n8369__, new_new_n8370__, new_new_n8371__, new_new_n8372__,
    new_new_n8373__, new_new_n8374__, new_new_n8375__, new_new_n8376__,
    new_new_n8377__, new_new_n8378__, new_new_n8379__, new_new_n8380__,
    new_new_n8381__, new_new_n8382__, new_new_n8383__, new_new_n8384__,
    new_new_n8385__, new_new_n8386__, new_new_n8387__, new_new_n8388__,
    new_new_n8389__, new_new_n8390__, new_new_n8391__, new_new_n8392__,
    new_new_n8393__, new_new_n8394__, new_new_n8395__, new_new_n8396__,
    new_new_n8397__, new_new_n8398__, new_new_n8399__, new_new_n8400__,
    new_new_n8401__, new_new_n8402__, new_new_n8403__, new_new_n8404__,
    new_new_n8405__, new_new_n8406__, new_new_n8407__, new_new_n8408__,
    new_new_n8409__, new_new_n8410__, new_new_n8411__, new_new_n8412__,
    new_new_n8413__, new_new_n8414__, new_new_n8415__, new_new_n8416__,
    new_new_n8417__, new_new_n8418__, new_new_n8419__, new_new_n8420__,
    new_new_n8421__, new_new_n8422__, new_new_n8423__, new_new_n8424__,
    new_new_n8425__, new_new_n8426__, new_new_n8427__, new_new_n8428__,
    new_new_n8429__, new_new_n8430__, new_new_n8431__, new_new_n8432__,
    new_new_n8433__, new_new_n8434__, new_new_n8435__, new_new_n8436__,
    new_new_n8437__, new_new_n8438__, new_new_n8439__, new_new_n8440__,
    new_new_n8441__, new_new_n8442__, new_new_n8443__, new_new_n8444__,
    new_new_n8445__, new_new_n8446__, new_new_n8447__, new_new_n8448__,
    new_new_n8449__, new_new_n8450__, new_new_n8451__, new_new_n8452__,
    new_new_n8453__, new_new_n8454__, new_new_n8455__, new_new_n8456__,
    new_new_n8457__, new_new_n8458__, new_new_n8459__, new_new_n8460__,
    new_new_n8461__, new_new_n8462__, new_new_n8463__, new_new_n8464__,
    new_new_n8465__, new_new_n8466__, new_new_n8467__, new_new_n8468__,
    new_new_n8469__, new_new_n8470__, new_new_n8471__, new_new_n8472__,
    new_new_n8473__, new_new_n8474__, new_new_n8475__, new_new_n8476__,
    new_new_n8477__, new_new_n8478__, new_new_n8479__, new_new_n8480__,
    new_new_n8481__, new_new_n8482__, new_new_n8483__, new_new_n8484__,
    new_new_n8485__, new_new_n8486__, new_new_n8487__, new_new_n8488__,
    new_new_n8489__, new_new_n8490__, new_new_n8491__, new_new_n8492__,
    new_new_n8493__, new_new_n8494__, new_new_n8495__, new_new_n8496__,
    new_new_n8497__, new_new_n8498__, new_new_n8499__, new_new_n8500__,
    new_new_n8501__, new_new_n8502__, new_new_n8503__, new_new_n8504__,
    new_new_n8505__, new_new_n8506__, new_new_n8507__, new_new_n8508__,
    new_new_n8509__, new_new_n8510__, new_new_n8511__, new_new_n8512__,
    new_new_n8513__, new_new_n8514__, new_new_n8515__, new_new_n8516__,
    new_new_n8517__, new_new_n8518__, new_new_n8519__, new_new_n8520__,
    new_new_n8521__, new_new_n8522__, new_new_n8523__, new_new_n8524__,
    new_new_n8525__, new_new_n8526__, new_new_n8527__, new_new_n8528__,
    new_new_n8529__, new_new_n8530__, new_new_n8531__, new_new_n8532__,
    new_new_n8533__, new_new_n8534__, new_new_n8535__, new_new_n8536__,
    new_new_n8537__, new_new_n8538__, new_new_n8539__, new_new_n8540__,
    new_new_n8541__, new_new_n8542__, new_new_n8543__, new_new_n8544__,
    new_new_n8545__, new_new_n8546__, new_new_n8547__, new_new_n8548__,
    new_new_n8549__, new_new_n8550__, new_new_n8551__, new_new_n8552__,
    new_new_n8553__, new_new_n8554__, new_new_n8555__, new_new_n8556__,
    new_new_n8557__, new_new_n8558__, new_new_n8559__, new_new_n8560__,
    new_new_n8561__, new_new_n8562__, new_new_n8563__, new_new_n8564__,
    new_new_n8565__, new_new_n8566__, new_new_n8567__, new_new_n8568__,
    new_new_n8569__, new_new_n8570__, new_new_n8571__, new_new_n8572__,
    new_new_n8573__, new_new_n8574__, new_new_n8575__, new_new_n8576__,
    new_new_n8577__, new_new_n8578__, new_new_n8579__, new_new_n8580__,
    new_new_n8581__, new_new_n8582__, new_new_n8583__, new_new_n8584__,
    new_new_n8585__, new_new_n8586__, new_new_n8587__, new_new_n8588__,
    new_new_n8589__, new_new_n8590__, new_new_n8591__, new_new_n8592__,
    new_new_n8593__, new_new_n8594__, new_new_n8595__, new_new_n8596__,
    new_new_n8597__, new_new_n8598__, new_new_n8599__, new_new_n8600__,
    new_new_n8601__, new_new_n8602__, new_new_n8603__, new_new_n8604__,
    new_new_n8605__, new_new_n8606__, new_new_n8607__, new_new_n8608__,
    new_new_n8609__, new_new_n8610__, new_new_n8611__, new_new_n8612__,
    new_new_n8613__, new_new_n8614__, new_new_n8615__, new_new_n8616__,
    new_new_n8617__, new_new_n8618__, new_new_n8619__, new_new_n8620__,
    new_new_n8621__, new_new_n8622__, new_new_n8623__, new_new_n8624__,
    new_new_n8625__, new_new_n8626__, new_new_n8627__, new_new_n8628__,
    new_new_n8629__, new_new_n8630__, new_new_n8631__, new_new_n8632__,
    new_new_n8633__, new_new_n8634__, new_new_n8635__, new_new_n8636__,
    new_new_n8637__, new_new_n8638__, new_new_n8639__, new_new_n8640__,
    new_new_n8641__, new_new_n8642__, new_new_n8643__, new_new_n8644__,
    new_new_n8645__, new_new_n8646__, new_new_n8647__, new_new_n8648__,
    new_new_n8649__, new_new_n8650__, new_new_n8651__, new_new_n8652__,
    new_new_n8653__, new_new_n8654__, new_new_n8655__, new_new_n8656__,
    new_new_n8657__, new_new_n8658__, new_new_n8659__, new_new_n8660__,
    new_new_n8661__, new_new_n8662__, new_new_n8663__, new_new_n8664__,
    new_new_n8665__, new_new_n8666__, new_new_n8667__, new_new_n8668__,
    new_new_n8669__, new_new_n8670__, new_new_n8671__, new_new_n8672__,
    new_new_n8673__, new_new_n8674__, new_new_n8675__, new_new_n8676__,
    new_new_n8677__, new_new_n8678__, new_new_n8679__, new_new_n8680__,
    new_new_n8681__, new_new_n8682__, new_new_n8683__, new_new_n8684__,
    new_new_n8685__, new_new_n8686__, new_new_n8687__, new_new_n8688__,
    new_new_n8689__, new_new_n8690__, new_new_n8691__, new_new_n8692__,
    new_new_n8693__, new_new_n8694__, new_new_n8695__, new_new_n8696__,
    new_new_n8697__, new_new_n8698__, new_new_n8699__, new_new_n8700__,
    new_new_n8701__, new_new_n8702__, new_new_n8703__, new_new_n8704__,
    new_new_n8705__, new_new_n8706__, new_new_n8707__, new_new_n8708__,
    new_new_n8709__, new_new_n8710__, new_new_n8711__, new_new_n8712__,
    new_new_n8713__, new_new_n8714__, new_new_n8715__, new_new_n8716__,
    new_new_n8717__, new_new_n8718__, new_new_n8719__, new_new_n8720__,
    new_new_n8721__, new_new_n8722__, new_new_n8723__, new_new_n8724__,
    new_new_n8725__, new_new_n8726__, new_new_n8727__, new_new_n8728__,
    new_new_n8729__, new_new_n8730__, new_new_n8731__, new_new_n8732__,
    new_new_n8733__, new_new_n8734__, new_new_n8735__, new_new_n8736__,
    new_new_n8737__, new_new_n8738__, new_new_n8739__, new_new_n8740__,
    new_new_n8741__, new_new_n8742__, new_new_n8743__, new_new_n8744__,
    new_new_n8745__, new_new_n8746__, new_new_n8747__, new_new_n8748__,
    new_new_n8749__, new_new_n8750__, new_new_n8751__, new_new_n8752__,
    new_new_n8753__, new_new_n8754__, new_new_n8755__, new_new_n8756__,
    new_new_n8757__, new_new_n8758__, new_new_n8759__, new_new_n8760__,
    new_new_n8761__, new_new_n8762__, new_new_n8763__, new_new_n8764__,
    new_new_n8765__, new_new_n8766__, new_new_n8767__, new_new_n8768__,
    new_new_n8769__, new_new_n8770__, new_new_n8771__, new_new_n8772__,
    new_new_n8773__, new_new_n8774__, new_new_n8775__, new_new_n8776__,
    new_new_n8777__, new_new_n8778__, new_new_n8779__, new_new_n8780__,
    new_new_n8781__, new_new_n8782__, new_new_n8783__, new_new_n8784__,
    new_new_n8785__, new_new_n8786__, new_new_n8787__, new_new_n8788__,
    new_new_n8789__, new_new_n8790__, new_new_n8791__, new_new_n8792__,
    new_new_n8793__, new_new_n8794__, new_new_n8795__, new_new_n8796__,
    new_new_n8797__, new_new_n8798__, new_new_n8799__, new_new_n8800__,
    new_new_n8801__, new_new_n8802__, new_new_n8803__, new_new_n8804__,
    new_new_n8805__, new_new_n8806__, new_new_n8807__, new_new_n8808__,
    new_new_n8809__, new_new_n8810__, new_new_n8811__, new_new_n8812__,
    new_new_n8813__, new_new_n8814__, new_new_n8815__, new_new_n8816__,
    new_new_n8817__, new_new_n8818__, new_new_n8819__, new_new_n8820__,
    new_new_n8821__, new_new_n8822__, new_new_n8823__, new_new_n8824__,
    new_new_n8825__, new_new_n8826__, new_new_n8827__, new_new_n8828__,
    new_new_n8829__, new_new_n8830__, new_new_n8831__, new_new_n8832__,
    new_new_n8833__, new_new_n8834__, new_new_n8835__, new_new_n8836__,
    new_new_n8837__, new_new_n8838__, new_new_n8839__, new_new_n8840__,
    new_new_n8841__, new_new_n8842__, new_new_n8843__, new_new_n8844__,
    new_new_n8845__, new_new_n8846__, new_new_n8847__, new_new_n8848__,
    new_new_n8849__, new_new_n8850__, new_new_n8851__, new_new_n8852__,
    new_new_n8853__, new_new_n8854__, new_new_n8855__, new_new_n8856__,
    new_new_n8857__, new_new_n8858__, new_new_n8859__, new_new_n8860__,
    new_new_n8861__, new_new_n8862__, new_new_n8863__, new_new_n8864__,
    new_new_n8865__, new_new_n8866__, new_new_n8867__, new_new_n8868__,
    new_new_n8869__, new_new_n8870__, new_new_n8871__, new_new_n8872__,
    new_new_n8873__, new_new_n8874__, new_new_n8875__, new_new_n8876__,
    new_new_n8877__, new_new_n8878__, new_new_n8879__, new_new_n8880__,
    new_new_n8881__, new_new_n8882__, new_new_n8883__, new_new_n8884__,
    new_new_n8885__, new_new_n8886__, new_new_n8887__, new_new_n8888__,
    new_new_n8889__, new_new_n8890__, new_new_n8891__, new_new_n8892__,
    new_new_n8893__, new_new_n8894__, new_new_n8895__, new_new_n8896__,
    new_new_n8897__, new_new_n8898__, new_new_n8899__, new_new_n8900__,
    new_new_n8901__, new_new_n8902__, new_new_n8903__, new_new_n8904__,
    new_new_n8905__, new_new_n8906__, new_new_n8907__, new_new_n8908__,
    new_new_n8909__, new_new_n8910__, new_new_n8911__, new_new_n8912__,
    new_new_n8913__, new_new_n8914__, new_new_n8915__, new_new_n8916__,
    new_new_n8917__, new_new_n8918__, new_new_n8919__, new_new_n8920__,
    new_new_n8921__, new_new_n8922__, new_new_n8923__, new_new_n8924__,
    new_new_n8925__, new_new_n8926__, new_new_n8927__, new_new_n8928__,
    new_new_n8929__, new_new_n8930__, new_new_n8931__, new_new_n8932__,
    new_new_n8933__, new_new_n8934__, new_new_n8935__, new_new_n8936__,
    new_new_n8937__, new_new_n8938__, new_new_n8939__, new_new_n8940__,
    new_new_n8941__, new_new_n8942__, new_new_n8943__, new_new_n8944__,
    new_new_n8945__, new_new_n8946__, new_new_n8947__, new_new_n8948__,
    new_new_n8949__, new_new_n8950__, new_new_n8951__, new_new_n8952__,
    new_new_n8953__, new_new_n8954__, new_new_n8955__, new_new_n8956__,
    new_new_n8957__, new_new_n8958__, new_new_n8959__, new_new_n8960__,
    new_new_n8961__, new_new_n8962__, new_new_n8963__, new_new_n8964__,
    new_new_n8965__, new_new_n8966__, new_new_n8967__, new_new_n8968__,
    new_new_n8969__, new_new_n8970__, new_new_n8971__, new_new_n8972__,
    new_new_n8973__, new_new_n8974__, new_new_n8975__, new_new_n8976__,
    new_new_n8977__, new_new_n8978__, new_new_n8979__, new_new_n8980__,
    new_new_n8981__, new_new_n8982__, new_new_n8983__, new_new_n8984__,
    new_new_n8985__, new_new_n8986__, new_new_n8987__, new_new_n8988__,
    new_new_n8989__, new_new_n8990__, new_new_n8991__, new_new_n8992__,
    new_new_n8993__, new_new_n8994__, new_new_n8995__, new_new_n8996__,
    new_new_n8997__, new_new_n8998__, new_new_n8999__, new_new_n9000__,
    new_new_n9001__, new_new_n9002__, new_new_n9003__, new_new_n9004__,
    new_new_n9005__, new_new_n9006__, new_new_n9007__, new_new_n9008__,
    new_new_n9009__, new_new_n9010__, new_new_n9011__, new_new_n9012__,
    new_new_n9013__, new_new_n9014__, new_new_n9015__, new_new_n9016__,
    new_new_n9017__, new_new_n9018__, new_new_n9019__, new_new_n9020__,
    new_new_n9021__, new_new_n9022__, new_new_n9023__, new_new_n9024__,
    new_new_n9025__, new_new_n9026__, new_new_n9027__, new_new_n9028__,
    new_new_n9029__, new_new_n9030__, new_new_n9031__, new_new_n9032__,
    new_new_n9033__, new_new_n9034__, new_new_n9035__, new_new_n9036__,
    new_new_n9037__, new_new_n9038__, new_new_n9039__, new_new_n9040__,
    new_new_n9041__, new_new_n9042__, new_new_n9043__, new_new_n9044__,
    new_new_n9045__, new_new_n9046__, new_new_n9047__, new_new_n9048__,
    new_new_n9049__, new_new_n9050__, new_new_n9051__, new_new_n9052__,
    new_new_n9053__, new_new_n9054__, new_new_n9055__, new_new_n9056__,
    new_new_n9057__, new_new_n9058__, new_new_n9059__, new_new_n9060__,
    new_new_n9061__, new_new_n9062__, new_new_n9063__, new_new_n9064__,
    new_new_n9065__, new_new_n9066__, new_new_n9067__, new_new_n9068__,
    new_new_n9069__, new_new_n9070__, new_new_n9071__, new_new_n9072__,
    new_new_n9073__, new_new_n9074__, new_new_n9075__, new_new_n9076__,
    new_new_n9077__, new_new_n9078__, new_new_n9079__, new_new_n9080__,
    new_new_n9081__, new_new_n9082__, new_new_n9083__, new_new_n9084__,
    new_new_n9085__, new_new_n9086__, new_new_n9087__, new_new_n9088__,
    new_new_n9089__, new_new_n9090__, new_new_n9091__, new_new_n9092__,
    new_new_n9093__, new_new_n9094__, new_new_n9095__, new_new_n9096__,
    new_new_n9097__, new_new_n9098__, new_new_n9099__, new_new_n9100__,
    new_new_n9101__, new_new_n9102__, new_new_n9103__, new_new_n9104__,
    new_new_n9105__, new_new_n9106__, new_new_n9107__, new_new_n9108__,
    new_new_n9109__, new_new_n9110__, new_new_n9111__, new_new_n9112__,
    new_new_n9113__, new_new_n9114__, new_new_n9115__, new_new_n9116__,
    new_new_n9117__, new_new_n9118__, new_new_n9119__, new_new_n9120__,
    new_new_n9121__, new_new_n9122__, new_new_n9123__, new_new_n9124__,
    new_new_n9125__, new_new_n9126__, new_new_n9127__, new_new_n9128__,
    new_new_n9129__, new_new_n9130__, new_new_n9131__, new_new_n9132__,
    new_new_n9133__, new_new_n9134__, new_new_n9135__, new_new_n9136__,
    new_new_n9137__, new_new_n9138__, new_new_n9139__, new_new_n9140__,
    new_new_n9141__, new_new_n9142__, new_new_n9143__, new_new_n9144__,
    new_new_n9145__, new_new_n9146__, new_new_n9147__, new_new_n9148__,
    new_new_n9149__, new_new_n9150__, new_new_n9151__, new_new_n9152__,
    new_new_n9153__, new_new_n9154__, new_new_n9155__, new_new_n9156__,
    new_new_n9157__, new_new_n9158__, new_new_n9159__, new_new_n9160__,
    new_new_n9161__, new_new_n9162__, new_new_n9163__, new_new_n9164__,
    new_new_n9165__, new_new_n9166__, new_new_n9167__, new_new_n9168__,
    new_new_n9169__, new_new_n9170__, new_new_n9171__, new_new_n9172__,
    new_new_n9173__, new_new_n9174__, new_new_n9175__, new_new_n9176__,
    new_new_n9177__, new_new_n9178__, new_new_n9179__, new_new_n9180__,
    new_new_n9181__, new_new_n9182__, new_new_n9183__, new_new_n9184__,
    new_new_n9185__, new_new_n9186__, new_new_n9187__, new_new_n9188__,
    new_new_n9189__, new_new_n9190__, new_new_n9191__, new_new_n9192__,
    new_new_n9193__, new_new_n9194__, new_new_n9195__, new_new_n9196__,
    new_new_n9197__, new_new_n9198__, new_new_n9199__, new_new_n9200__,
    new_new_n9201__, new_new_n9202__, new_new_n9203__, new_new_n9204__,
    new_new_n9205__, new_new_n9206__, new_new_n9207__, new_new_n9208__,
    new_new_n9209__, new_new_n9210__, new_new_n9211__, new_new_n9212__,
    new_new_n9213__, new_new_n9214__, new_new_n9215__, new_new_n9216__,
    new_new_n9217__, new_new_n9218__, new_new_n9219__, new_new_n9220__,
    new_new_n9221__, new_new_n9222__, new_new_n9223__, new_new_n9224__,
    new_new_n9225__, new_new_n9226__, new_new_n9227__, new_new_n9228__,
    new_new_n9229__, new_new_n9230__, new_new_n9231__, new_new_n9232__,
    new_new_n9233__, new_new_n9234__, new_new_n9235__, new_new_n9236__,
    new_new_n9237__, new_new_n9238__, new_new_n9239__, new_new_n9240__,
    new_new_n9241__, new_new_n9242__, new_new_n9243__, new_new_n9244__,
    new_new_n9245__, new_new_n9246__, new_new_n9247__, new_new_n9248__,
    new_new_n9249__, new_new_n9250__, new_new_n9251__, new_new_n9252__,
    new_new_n9253__, new_new_n9254__, new_new_n9255__, new_new_n9256__,
    new_new_n9257__, new_new_n9258__, new_new_n9259__, new_new_n9260__,
    new_new_n9261__, new_new_n9262__, new_new_n9263__, new_new_n9264__,
    new_new_n9265__, new_new_n9266__, new_new_n9267__, new_new_n9268__,
    new_new_n9269__, new_new_n9270__, new_new_n9271__, new_new_n9272__,
    new_new_n9273__, new_new_n9274__, new_new_n9275__, new_new_n9276__,
    new_new_n9277__, new_new_n9278__, new_new_n9279__, new_new_n9280__,
    new_new_n9281__, new_new_n9282__, new_new_n9283__, new_new_n9284__,
    new_new_n9285__, new_new_n9286__, new_new_n9287__, new_new_n9288__,
    new_new_n9289__, new_new_n9290__, new_new_n9291__, new_new_n9292__,
    new_new_n9293__, new_new_n9294__, new_new_n9295__, new_new_n9296__,
    new_new_n9297__, new_new_n9298__, new_new_n9299__, new_new_n9300__,
    new_new_n9301__, new_new_n9302__, new_new_n9303__, new_new_n9304__,
    new_new_n9305__, new_new_n9306__, new_new_n9307__, new_new_n9308__,
    new_new_n9309__, new_new_n9310__, new_new_n9311__, new_new_n9312__,
    new_new_n9313__, new_new_n9314__, new_new_n9315__, new_new_n9316__,
    new_new_n9317__, new_new_n9318__, new_new_n9319__, new_new_n9320__,
    new_new_n9321__, new_new_n9322__, new_new_n9323__, new_new_n9324__,
    new_new_n9325__, new_new_n9326__, new_new_n9327__, new_new_n9328__,
    new_new_n9329__, new_new_n9330__, new_new_n9331__, new_new_n9332__,
    new_new_n9333__, new_new_n9334__, new_new_n9335__, new_new_n9336__,
    new_new_n9337__, new_new_n9338__, new_new_n9339__, new_new_n9340__,
    new_new_n9341__, new_new_n9342__, new_new_n9343__, new_new_n9344__,
    new_new_n9345__, new_new_n9346__, new_new_n9347__, new_new_n9348__,
    new_new_n9349__, new_new_n9350__, new_new_n9351__, new_new_n9352__,
    new_new_n9353__, new_new_n9354__, new_new_n9355__, new_new_n9356__,
    new_new_n9357__, new_new_n9358__, new_new_n9359__, new_new_n9360__,
    new_new_n9361__, new_new_n9362__, new_new_n9363__, new_new_n9364__,
    new_new_n9365__, new_new_n9366__, new_new_n9367__, new_new_n9368__,
    new_new_n9369__, new_new_n9370__, new_new_n9371__, new_new_n9372__,
    new_new_n9373__, new_new_n9374__, new_new_n9375__, new_new_n9376__,
    new_new_n9377__, new_new_n9378__, new_new_n9379__, new_new_n9380__,
    new_new_n9381__, new_new_n9382__, new_new_n9383__, new_new_n9384__,
    new_new_n9385__, new_new_n9386__, new_new_n9387__, new_new_n9388__,
    new_new_n9389__, new_new_n9390__, new_new_n9391__, new_new_n9392__,
    new_new_n9393__, new_new_n9394__, new_new_n9395__, new_new_n9396__,
    new_new_n9397__, new_new_n9398__, new_new_n9399__, new_new_n9400__,
    new_new_n9401__, new_new_n9402__, new_new_n9403__, new_new_n9404__,
    new_new_n9405__, new_new_n9406__, new_new_n9407__, new_new_n9408__,
    new_new_n9409__, new_new_n9410__, new_new_n9411__, new_new_n9412__,
    new_new_n9413__, new_new_n9414__, new_new_n9415__, new_new_n9416__,
    new_new_n9417__, new_new_n9418__, new_new_n9419__, new_new_n9420__,
    new_new_n9421__, new_new_n9422__, new_new_n9423__, new_new_n9424__,
    new_new_n9425__, new_new_n9426__, new_new_n9427__, new_new_n9428__,
    new_new_n9429__, new_new_n9430__, new_new_n9431__, new_new_n9432__,
    new_new_n9433__, new_new_n9434__, new_new_n9435__, new_new_n9436__,
    new_new_n9437__, new_new_n9438__, new_new_n9439__, new_new_n9440__,
    new_new_n9441__, new_new_n9442__, new_new_n9443__, new_new_n9444__,
    new_new_n9445__, new_new_n9446__, new_new_n9447__, new_new_n9448__,
    new_new_n9449__, new_new_n9450__, new_new_n9451__, new_new_n9452__,
    new_new_n9453__, new_new_n9454__, new_new_n9455__, new_new_n9456__,
    new_new_n9457__, new_new_n9458__, new_new_n9459__, new_new_n9460__,
    new_new_n9461__, new_new_n9462__, new_new_n9463__, new_new_n9464__,
    new_new_n9465__, new_new_n9466__, new_new_n9467__, new_new_n9468__,
    new_new_n9469__, new_new_n9470__, new_new_n9471__, new_new_n9472__,
    new_new_n9473__, new_new_n9474__, new_new_n9475__, new_new_n9476__,
    new_new_n9477__, new_new_n9478__, new_new_n9479__, new_new_n9480__,
    new_new_n9481__, new_new_n9482__, new_new_n9483__, new_new_n9484__,
    new_new_n9485__, new_new_n9486__, new_new_n9487__, new_new_n9488__,
    new_new_n9489__, new_new_n9490__, new_new_n9491__, new_new_n9492__,
    new_new_n9493__, new_new_n9494__, new_new_n9495__, new_new_n9496__,
    new_new_n9497__, new_new_n9498__, new_new_n9499__, new_new_n9500__,
    new_new_n9501__, new_new_n9502__, new_new_n9503__, new_new_n9504__,
    new_new_n9505__, new_new_n9506__, new_new_n9507__, new_new_n9508__,
    new_new_n9509__, new_new_n9510__, new_new_n9511__, new_new_n9512__,
    new_new_n9513__, new_new_n9514__, new_new_n9515__, new_new_n9516__,
    new_new_n9517__, new_new_n9518__, new_new_n9519__, new_new_n9520__,
    new_new_n9521__, new_new_n9522__, new_new_n9523__, new_new_n9524__,
    new_new_n9525__, new_new_n9526__, new_new_n9527__, new_new_n9528__,
    new_new_n9529__, new_new_n9530__, new_new_n9531__, new_new_n9532__,
    new_new_n9533__, new_new_n9534__, new_new_n9535__, new_new_n9536__,
    new_new_n9537__, new_new_n9538__, new_new_n9539__, new_new_n9540__,
    new_new_n9541__, new_new_n9542__, new_new_n9543__, new_new_n9544__,
    new_new_n9545__, new_new_n9546__, new_new_n9547__, new_new_n9548__,
    new_new_n9549__, new_new_n9550__, new_new_n9551__, new_new_n9552__,
    new_new_n9553__, new_new_n9554__, new_new_n9555__, new_new_n9556__,
    new_new_n9557__, new_new_n9558__, new_new_n9559__, new_new_n9560__,
    new_new_n9561__, new_new_n9562__, new_new_n9563__, new_new_n9564__,
    new_new_n9565__, new_new_n9566__, new_new_n9567__, new_new_n9568__,
    new_new_n9569__, new_new_n9570__, new_new_n9571__, new_new_n9572__,
    new_new_n9573__, new_new_n9574__, new_new_n9575__, new_new_n9576__,
    new_new_n9577__, new_new_n9578__, new_new_n9579__, new_new_n9580__,
    new_new_n9581__, new_new_n9582__, new_new_n9583__, new_new_n9584__,
    new_new_n9585__, new_new_n9586__, new_new_n9587__, new_new_n9588__,
    new_new_n9589__, new_new_n9590__, new_new_n9591__, new_new_n9592__,
    new_new_n9593__, new_new_n9594__, new_new_n9595__, new_new_n9596__,
    new_new_n9597__, new_new_n9598__, new_new_n9599__, new_new_n9600__,
    new_new_n9601__, new_new_n9602__, new_new_n9603__, new_new_n9604__,
    new_new_n9605__, new_new_n9606__, new_new_n9607__, new_new_n9608__,
    new_new_n9609__, new_new_n9610__, new_new_n9611__, new_new_n9612__,
    new_new_n9613__, new_new_n9614__, new_new_n9615__, new_new_n9616__,
    new_new_n9617__, new_new_n9618__, new_new_n9619__, new_new_n9620__,
    new_new_n9621__, new_new_n9622__, new_new_n9623__, new_new_n9624__,
    new_new_n9625__, new_new_n9626__, new_new_n9627__, new_new_n9628__,
    new_new_n9629__, new_new_n9630__, new_new_n9631__, new_new_n9632__,
    new_new_n9633__, new_new_n9634__, new_new_n9635__, new_new_n9636__,
    new_new_n9637__, new_new_n9638__, new_new_n9639__, new_new_n9640__,
    new_new_n9641__, new_new_n9642__, new_new_n9643__, new_new_n9644__,
    new_new_n9645__, new_new_n9646__, new_new_n9647__, new_new_n9648__,
    new_new_n9649__, new_new_n9650__, new_new_n9651__, new_new_n9652__,
    new_new_n9653__, new_new_n9654__, new_new_n9655__, new_new_n9656__,
    new_new_n9657__, new_new_n9658__, new_new_n9659__, new_new_n9660__,
    new_new_n9661__, new_new_n9662__, new_new_n9663__, new_new_n9664__,
    new_new_n9665__, new_new_n9666__, new_new_n9667__, new_new_n9668__,
    new_new_n9669__, new_new_n9670__, new_new_n9671__, new_new_n9672__,
    new_new_n9673__, new_new_n9674__, new_new_n9675__, new_new_n9676__,
    new_new_n9677__, new_new_n9678__, new_new_n9679__, new_new_n9680__,
    new_new_n9681__, new_new_n9682__, new_new_n9683__, new_new_n9684__,
    new_new_n9685__, new_new_n9686__, new_new_n9687__, new_new_n9688__,
    new_new_n9689__, new_new_n9690__, new_new_n9691__, new_new_n9692__,
    new_new_n9693__, new_new_n9694__, new_new_n9695__, new_new_n9696__,
    new_new_n9697__, new_new_n9698__, new_new_n9699__, new_new_n9700__,
    new_new_n9701__, new_new_n9702__, new_new_n9703__, new_new_n9704__,
    new_new_n9705__, new_new_n9706__, new_new_n9707__, new_new_n9708__,
    new_new_n9709__, new_new_n9710__, new_new_n9711__, new_new_n9712__,
    new_new_n9713__, new_new_n9714__, new_new_n9715__, new_new_n9716__,
    new_new_n9717__, new_new_n9718__, new_new_n9719__, new_new_n9720__,
    new_new_n9721__, new_new_n9722__, new_new_n9723__, new_new_n9724__,
    new_new_n9725__, new_new_n9726__, new_new_n9727__, new_new_n9728__,
    new_new_n9729__, new_new_n9730__, new_new_n9731__, new_new_n9732__,
    new_new_n9733__, new_new_n9734__, new_new_n9735__, new_new_n9736__,
    new_new_n9737__, new_new_n9738__, new_new_n9739__, new_new_n9740__,
    new_new_n9741__, new_new_n9742__, new_new_n9743__, new_new_n9744__,
    new_new_n9745__, new_new_n9746__, new_new_n9747__, new_new_n9748__,
    new_new_n9749__, new_new_n9750__, new_new_n9751__, new_new_n9752__,
    new_new_n9753__, new_new_n9754__, new_new_n9755__, new_new_n9756__,
    new_new_n9757__, new_new_n9758__, new_new_n9759__, new_new_n9760__,
    new_new_n9761__, new_new_n9762__, new_new_n9763__, new_new_n9764__,
    new_new_n9765__, new_new_n9766__, new_new_n9767__, new_new_n9768__,
    new_new_n9769__, new_new_n9770__, new_new_n9771__, new_new_n9772__,
    new_new_n9773__, new_new_n9774__, new_new_n9775__, new_new_n9776__,
    new_new_n9777__, new_new_n9778__, new_new_n9779__, new_new_n9780__,
    new_new_n9781__, new_new_n9782__, new_new_n9783__, new_new_n9784__,
    new_new_n9785__, new_new_n9786__, new_new_n9787__, new_new_n9788__,
    new_new_n9789__, new_new_n9790__, new_new_n9791__, new_new_n9792__,
    new_new_n9793__, new_new_n9794__, new_new_n9795__, new_new_n9796__,
    new_new_n9797__, new_new_n9798__, new_new_n9799__, new_new_n9800__,
    new_new_n9801__, new_new_n9802__, new_new_n9803__, new_new_n9804__,
    new_new_n9805__, new_new_n9806__, new_new_n9807__, new_new_n9808__,
    new_new_n9809__, new_new_n9810__, new_new_n9811__, new_new_n9812__,
    new_new_n9813__, new_new_n9814__, new_new_n9815__, new_new_n9816__,
    new_new_n9817__, new_new_n9818__, new_new_n9819__, new_new_n9820__,
    new_new_n9821__, new_new_n9822__, new_new_n9823__, new_new_n9824__,
    new_new_n9825__, new_new_n9826__, new_new_n9827__, new_new_n9828__,
    new_new_n9829__, new_new_n9830__, new_new_n9831__, new_new_n9832__,
    new_new_n9833__, new_new_n9834__, new_new_n9835__, new_new_n9836__,
    new_new_n9837__, new_new_n9838__, new_new_n9839__, new_new_n9840__,
    new_new_n9841__, new_new_n9842__, new_new_n9843__, new_new_n9844__,
    new_new_n9845__, new_new_n9846__, new_new_n9847__, new_new_n9848__,
    new_new_n9849__, new_new_n9850__, new_new_n9851__, new_new_n9852__,
    new_new_n9853__, new_new_n9854__, new_new_n9855__, new_new_n9856__,
    new_new_n9857__, new_new_n9858__, new_new_n9859__, new_new_n9860__,
    new_new_n9861__, new_new_n9862__, new_new_n9863__, new_new_n9864__,
    new_new_n9865__, new_new_n9866__, new_new_n9867__, new_new_n9868__,
    new_new_n9869__, new_new_n9870__, new_new_n9871__, new_new_n9872__,
    new_new_n9873__, new_new_n9874__, new_new_n9875__, new_new_n9876__,
    new_new_n9877__, new_new_n9878__, new_new_n9879__, new_new_n9880__,
    new_new_n9881__, new_new_n9882__, new_new_n9883__, new_new_n9884__,
    new_new_n9885__, new_new_n9886__, new_new_n9887__, new_new_n9888__,
    new_new_n9889__, new_new_n9890__, new_new_n9891__, new_new_n9892__,
    new_new_n9893__, new_new_n9894__, new_new_n9895__, new_new_n9896__,
    new_new_n9897__, new_new_n9898__, new_new_n9899__, new_new_n9900__,
    new_new_n9901__, new_new_n9902__, new_new_n9903__, new_new_n9904__,
    new_new_n9905__, new_new_n9906__, new_new_n9907__, new_new_n9908__,
    new_new_n9909__, new_new_n9910__, new_new_n9911__, new_new_n9912__,
    new_new_n9913__, new_new_n9914__, new_new_n9915__, new_new_n9916__,
    new_new_n9917__, new_new_n9918__, new_new_n9919__, new_new_n9920__,
    new_new_n9921__, new_new_n9922__, new_new_n9923__, new_new_n9924__,
    new_new_n9925__, new_new_n9926__, new_new_n9927__, new_new_n9928__,
    new_new_n9929__, new_new_n9930__, new_new_n9931__, new_new_n9932__,
    new_new_n9933__, new_new_n9934__, new_new_n9935__, new_new_n9936__,
    new_new_n9937__, new_new_n9938__, new_new_n9939__, new_new_n9940__,
    new_new_n9941__, new_new_n9942__, new_new_n9943__, new_new_n9944__,
    new_new_n9945__, new_new_n9946__, new_new_n9947__, new_new_n9948__,
    new_new_n9949__, new_new_n9950__, new_new_n9951__, new_new_n9952__,
    new_new_n9953__, new_new_n9954__, new_new_n9955__, new_new_n9956__,
    new_new_n9957__, new_new_n9958__, new_new_n9959__, new_new_n9960__,
    new_new_n9961__, new_new_n9962__, new_new_n9963__, new_new_n9964__,
    new_new_n9965__, new_new_n9966__, new_new_n9967__, new_new_n9968__,
    new_new_n9969__, new_new_n9970__, new_new_n9971__, new_new_n9972__,
    new_new_n9973__, new_new_n9974__, new_new_n9975__, new_new_n9976__,
    new_new_n9977__, new_new_n9978__, new_new_n9979__, new_new_n9980__,
    new_new_n9981__, new_new_n9982__, new_new_n9983__, new_new_n9984__,
    new_new_n9985__, new_new_n9986__, new_new_n9987__, new_new_n9988__,
    new_new_n9989__, new_new_n9990__, new_new_n9991__, new_new_n9992__,
    new_new_n9993__, new_new_n9994__, new_new_n9995__, new_new_n9996__,
    new_new_n9997__, new_new_n9998__, new_new_n9999__, new_new_n10000__,
    new_new_n10001__, new_new_n10002__, new_new_n10003__, new_new_n10004__,
    new_new_n10005__, new_new_n10006__, new_new_n10007__, new_new_n10008__,
    new_new_n10009__, new_new_n10010__, new_new_n10011__, new_new_n10012__,
    new_new_n10013__, new_new_n10014__, new_new_n10015__, new_new_n10016__,
    new_new_n10017__, new_new_n10018__, new_new_n10019__, new_new_n10020__,
    new_new_n10021__, new_new_n10022__, new_new_n10023__, new_new_n10024__,
    new_new_n10025__, new_new_n10026__, new_new_n10027__, new_new_n10028__,
    new_new_n10029__, new_new_n10030__, new_new_n10031__, new_new_n10032__,
    new_new_n10033__, new_new_n10034__, new_new_n10035__, new_new_n10036__,
    new_new_n10037__, new_new_n10038__, new_new_n10039__, new_new_n10040__,
    new_new_n10041__, new_new_n10042__, new_new_n10043__, new_new_n10044__,
    new_new_n10045__, new_new_n10046__, new_new_n10047__, new_new_n10048__,
    new_new_n10049__, new_new_n10050__, new_new_n10051__, new_new_n10052__,
    new_new_n10053__, new_new_n10054__, new_new_n10055__, new_new_n10056__,
    new_new_n10057__, new_new_n10058__, new_new_n10059__, new_new_n10060__,
    new_new_n10061__, new_new_n10062__, new_new_n10063__, new_new_n10064__,
    new_new_n10065__, new_new_n10066__, new_new_n10067__, new_new_n10068__,
    new_new_n10069__, new_new_n10070__, new_new_n10071__, new_new_n10072__,
    new_new_n10073__, new_new_n10074__, new_new_n10075__, new_new_n10076__,
    new_new_n10077__, new_new_n10078__, new_new_n10079__, new_new_n10080__,
    new_new_n10081__, new_new_n10082__, new_new_n10083__, new_new_n10084__,
    new_new_n10085__, new_new_n10086__, new_new_n10087__, new_new_n10088__,
    new_new_n10089__, new_new_n10090__, new_new_n10091__, new_new_n10092__,
    new_new_n10093__, new_new_n10094__, new_new_n10095__, new_new_n10096__,
    new_new_n10097__, new_new_n10098__, new_new_n10099__, new_new_n10100__,
    new_new_n10101__, new_new_n10102__, new_new_n10103__, new_new_n10104__,
    new_new_n10105__, new_new_n10106__, new_new_n10107__, new_new_n10108__,
    new_new_n10109__, new_new_n10110__, new_new_n10111__, new_new_n10112__,
    new_new_n10113__, new_new_n10114__, new_new_n10115__, new_new_n10116__,
    new_new_n10117__, new_new_n10118__, new_new_n10119__, new_new_n10120__,
    new_new_n10121__, new_new_n10122__, new_new_n10123__, new_new_n10124__,
    new_new_n10125__, new_new_n10126__, new_new_n10127__, new_new_n10128__,
    new_new_n10129__, new_new_n10130__, new_new_n10131__, new_new_n10132__,
    new_new_n10133__, new_new_n10134__, new_new_n10135__, new_new_n10136__,
    new_new_n10137__, new_new_n10138__, new_new_n10139__, new_new_n10140__,
    new_new_n10141__, new_new_n10142__, new_new_n10143__, new_new_n10144__,
    new_new_n10145__, new_new_n10146__, new_new_n10147__, new_new_n10148__,
    new_new_n10149__, new_new_n10150__, new_new_n10151__, new_new_n10152__,
    new_new_n10153__, new_new_n10154__, new_new_n10155__, new_new_n10156__,
    new_new_n10157__, new_new_n10158__, new_new_n10159__, new_new_n10160__,
    new_new_n10161__, new_new_n10162__, new_new_n10163__, new_new_n10164__,
    new_new_n10165__, new_new_n10166__, new_new_n10167__, new_new_n10168__,
    new_new_n10169__, new_new_n10170__, new_new_n10171__, new_new_n10172__,
    new_new_n10173__, new_new_n10174__, new_new_n10175__, new_new_n10176__,
    new_new_n10177__, new_new_n10178__, new_new_n10179__, new_new_n10180__,
    new_new_n10181__, new_new_n10182__, new_new_n10183__, new_new_n10184__,
    new_new_n10185__, new_new_n10186__, new_new_n10187__, new_new_n10188__,
    new_new_n10189__, new_new_n10190__, new_new_n10191__, new_new_n10192__,
    new_new_n10193__, new_new_n10194__, new_new_n10195__, new_new_n10196__,
    new_new_n10197__, new_new_n10198__, new_new_n10199__, new_new_n10200__,
    new_new_n10201__, new_new_n10202__, new_new_n10203__, new_new_n10204__,
    new_new_n10205__, new_new_n10206__, new_new_n10207__, new_new_n10208__,
    new_new_n10209__, new_new_n10210__, new_new_n10211__, new_new_n10212__,
    new_new_n10213__, new_new_n10214__, new_new_n10215__, new_new_n10216__,
    new_new_n10217__, new_new_n10218__, new_new_n10219__, new_new_n10220__,
    new_new_n10221__, new_new_n10222__, new_new_n10223__, new_new_n10224__,
    new_new_n10225__, new_new_n10226__, new_new_n10227__, new_new_n10228__,
    new_new_n10229__, new_new_n10230__, new_new_n10231__, new_new_n10232__,
    new_new_n10233__, new_new_n10234__, new_new_n10235__, new_new_n10236__,
    new_new_n10237__, new_new_n10238__, new_new_n10239__, new_new_n10240__,
    new_new_n10241__, new_new_n10242__, new_new_n10243__, new_new_n10244__,
    new_new_n10245__, new_new_n10246__, new_new_n10247__, new_new_n10248__,
    new_new_n10249__, new_new_n10250__, new_new_n10251__, new_new_n10252__,
    new_new_n10253__, new_new_n10254__, new_new_n10255__, new_new_n10256__,
    new_new_n10257__, new_new_n10258__, new_new_n10259__, new_new_n10260__,
    new_new_n10261__, new_new_n10262__, new_new_n10263__, new_new_n10264__,
    new_new_n10265__, new_new_n10266__, new_new_n10267__, new_new_n10268__,
    new_new_n10269__, new_new_n10270__, new_new_n10271__, new_new_n10272__,
    new_new_n10273__, new_new_n10274__, new_new_n10275__, new_new_n10276__,
    new_new_n10277__, new_new_n10278__, new_new_n10279__, new_new_n10280__,
    new_new_n10281__, new_new_n10282__, new_new_n10283__, new_new_n10284__,
    new_new_n10285__, new_new_n10286__, new_new_n10287__, new_new_n10288__,
    new_new_n10289__, new_new_n10290__, new_new_n10291__, new_new_n10292__,
    new_new_n10293__, new_new_n10294__, new_new_n10295__, new_new_n10296__,
    new_new_n10297__, new_new_n10298__, new_new_n10299__, new_new_n10300__,
    new_new_n10301__, new_new_n10302__, new_new_n10303__, new_new_n10304__,
    new_new_n10305__, new_new_n10306__, new_new_n10307__, new_new_n10308__,
    new_new_n10309__, new_new_n10310__, new_new_n10311__, new_new_n10312__,
    new_new_n10313__, new_new_n10314__, new_new_n10315__, new_new_n10316__,
    new_new_n10317__, new_new_n10318__, new_new_n10319__, new_new_n10320__,
    new_new_n10321__, new_new_n10322__, new_new_n10323__, new_new_n10324__,
    new_new_n10325__, new_new_n10326__, new_new_n10327__, new_new_n10328__,
    new_new_n10329__, new_new_n10330__, new_new_n10331__, new_new_n10332__,
    new_new_n10333__, new_new_n10334__, new_new_n10335__, new_new_n10336__,
    new_new_n10337__, new_new_n10338__, new_new_n10339__, new_new_n10340__,
    new_new_n10341__, new_new_n10342__, new_new_n10343__, new_new_n10344__,
    new_new_n10345__, new_new_n10346__, new_new_n10347__, new_new_n10348__,
    new_new_n10349__, new_new_n10350__, new_new_n10351__, new_new_n10352__,
    new_new_n10353__, new_new_n10354__, new_new_n10355__, new_new_n10356__,
    new_new_n10357__, new_new_n10358__, new_new_n10359__, new_new_n10360__,
    new_new_n10361__, new_new_n10362__, new_new_n10363__, new_new_n10364__,
    new_new_n10365__, new_new_n10366__, new_new_n10367__, new_new_n10368__,
    new_new_n10369__, new_new_n10370__, new_new_n10371__, new_new_n10372__,
    new_new_n10373__, new_new_n10374__, new_new_n10375__, new_new_n10376__,
    new_new_n10377__, new_new_n10378__, new_new_n10379__, new_new_n10380__,
    new_new_n10381__, new_new_n10382__, new_new_n10383__, new_new_n10384__,
    new_new_n10385__, new_new_n10386__, new_new_n10387__, new_new_n10388__,
    new_new_n10389__, new_new_n10390__, new_new_n10391__, new_new_n10392__,
    new_new_n10393__, new_new_n10394__, new_new_n10395__, new_new_n10396__,
    new_new_n10397__, new_new_n10398__, new_new_n10399__, new_new_n10400__,
    new_new_n10401__, new_new_n10402__, new_new_n10403__, new_new_n10404__,
    new_new_n10405__, new_new_n10406__, new_new_n10407__, new_new_n10408__,
    new_new_n10409__, new_new_n10410__, new_new_n10411__, new_new_n10412__,
    new_new_n10413__, new_new_n10414__, new_new_n10415__, new_new_n10416__,
    new_new_n10417__, new_new_n10418__, new_new_n10419__, new_new_n10420__,
    new_new_n10421__, new_new_n10422__, new_new_n10423__, new_new_n10424__,
    new_new_n10425__, new_new_n10426__, new_new_n10427__, new_new_n10428__,
    new_new_n10429__, new_new_n10430__, new_new_n10431__, new_new_n10432__,
    new_new_n10433__, new_new_n10434__, new_new_n10435__, new_new_n10436__,
    new_new_n10437__, new_new_n10438__, new_new_n10439__, new_new_n10440__,
    new_new_n10441__, new_new_n10442__, new_new_n10443__, new_new_n10444__,
    new_new_n10445__, new_new_n10446__, new_new_n10447__, new_new_n10448__,
    new_new_n10449__, new_new_n10450__, new_new_n10451__, new_new_n10452__,
    new_new_n10453__, new_new_n10454__, new_new_n10455__, new_new_n10456__,
    new_new_n10457__, new_new_n10458__, new_new_n10459__, new_new_n10460__,
    new_new_n10461__, new_new_n10462__, new_new_n10463__, new_new_n10464__,
    new_new_n10465__, new_new_n10466__, new_new_n10467__, new_new_n10468__,
    new_new_n10469__, new_new_n10470__, new_new_n10471__, new_new_n10472__,
    new_new_n10473__, new_new_n10474__, new_new_n10475__, new_new_n10476__,
    new_new_n10477__, new_new_n10478__, new_new_n10479__, new_new_n10480__,
    new_new_n10481__, new_new_n10482__, new_new_n10483__, new_new_n10484__,
    new_new_n10485__, new_new_n10486__, new_new_n10487__, new_new_n10488__,
    new_new_n10489__, new_new_n10490__, new_new_n10491__, new_new_n10492__,
    new_new_n10493__, new_new_n10494__, new_new_n10495__, new_new_n10496__,
    new_new_n10497__, new_new_n10498__, new_new_n10499__, new_new_n10500__,
    new_new_n10501__, new_new_n10502__, new_new_n10503__, new_new_n10504__,
    new_new_n10505__, new_new_n10506__, new_new_n10507__, new_new_n10508__,
    new_new_n10509__, new_new_n10510__, new_new_n10511__, new_new_n10512__,
    new_new_n10513__, new_new_n10514__, new_new_n10515__, new_new_n10516__,
    new_new_n10517__, new_new_n10518__, new_new_n10519__, new_new_n10520__,
    new_new_n10521__, new_new_n10522__, new_new_n10523__, new_new_n10524__,
    new_new_n10525__, new_new_n10526__, new_new_n10527__, new_new_n10528__,
    new_new_n10529__, new_new_n10530__, new_new_n10531__, new_new_n10532__,
    new_new_n10533__, new_new_n10534__, new_new_n10535__, new_new_n10536__,
    new_new_n10537__, new_new_n10538__, new_new_n10539__, new_new_n10540__,
    new_new_n10541__, new_new_n10542__, new_new_n10543__, new_new_n10544__,
    new_new_n10545__, new_new_n10546__, new_new_n10547__, new_new_n10548__,
    new_new_n10549__, new_new_n10550__, new_new_n10551__, new_new_n10552__,
    new_new_n10553__, new_new_n10554__, new_new_n10555__, new_new_n10556__,
    new_new_n10557__, new_new_n10558__, new_new_n10559__, new_new_n10560__,
    new_new_n10561__, new_new_n10562__, new_new_n10563__, new_new_n10564__,
    new_new_n10565__, new_new_n10566__, new_new_n10567__, new_new_n10568__,
    new_new_n10569__, new_new_n10570__, new_new_n10571__, new_new_n10572__,
    new_new_n10573__, new_new_n10574__, new_new_n10575__, new_new_n10576__,
    new_new_n10577__, new_new_n10578__, new_new_n10579__, new_new_n10580__,
    new_new_n10581__, new_new_n10582__, new_new_n10583__, new_new_n10584__,
    new_new_n10585__, new_new_n10586__, new_new_n10587__, new_new_n10588__,
    new_new_n10589__, new_new_n10590__, new_new_n10591__, new_new_n10592__,
    new_new_n10593__, new_new_n10594__, new_new_n10595__, new_new_n10596__,
    new_new_n10597__, new_new_n10598__, new_new_n10599__, new_new_n10600__,
    new_new_n10601__, new_new_n10602__, new_new_n10603__, new_new_n10604__,
    new_new_n10605__, new_new_n10606__, new_new_n10607__, new_new_n10608__,
    new_new_n10609__, new_new_n10610__, new_new_n10611__, new_new_n10612__,
    new_new_n10613__, new_new_n10614__, new_new_n10615__, new_new_n10616__,
    new_new_n10617__, new_new_n10618__, new_new_n10619__, new_new_n10620__,
    new_new_n10621__, new_new_n10622__, new_new_n10623__, new_new_n10624__,
    new_new_n10625__, new_new_n10626__, new_new_n10627__, new_new_n10628__,
    new_new_n10629__, new_new_n10630__, new_new_n10631__, new_new_n10632__,
    new_new_n10633__, new_new_n10634__, new_new_n10635__, new_new_n10636__,
    new_new_n10637__, new_new_n10638__, new_new_n10639__, new_new_n10640__,
    new_new_n10641__, new_new_n10642__, new_new_n10643__, new_new_n10644__,
    new_new_n10645__, new_new_n10646__, new_new_n10647__, new_new_n10648__,
    new_new_n10649__, new_new_n10650__, new_new_n10651__, new_new_n10652__,
    new_new_n10653__, new_new_n10654__, new_new_n10655__, new_new_n10656__,
    new_new_n10657__, new_new_n10658__, new_new_n10659__, new_new_n10660__,
    new_new_n10661__, new_new_n10662__, new_new_n10663__, new_new_n10664__,
    new_new_n10665__, new_new_n10666__, new_new_n10667__, new_new_n10668__,
    new_new_n10669__, new_new_n10670__, new_new_n10671__, new_new_n10672__,
    new_new_n10673__, new_new_n10674__, new_new_n10675__, new_new_n10676__,
    new_new_n10677__, new_new_n10678__, new_new_n10679__, new_new_n10680__,
    new_new_n10681__, new_new_n10682__, new_new_n10683__, new_new_n10684__,
    new_new_n10685__, new_new_n10686__, new_new_n10687__, new_new_n10688__,
    new_new_n10689__, new_new_n10690__, new_new_n10691__, new_new_n10692__,
    new_new_n10693__, new_new_n10694__, new_new_n10695__, new_new_n10696__,
    new_new_n10697__, new_new_n10698__, new_new_n10699__, new_new_n10700__,
    new_new_n10701__, new_new_n10702__, new_new_n10703__, new_new_n10704__,
    new_new_n10705__, new_new_n10706__, new_new_n10707__, new_new_n10708__,
    new_new_n10709__, new_new_n10710__, new_new_n10711__, new_new_n10712__,
    new_new_n10713__, new_new_n10714__, new_new_n10715__, new_new_n10716__,
    new_new_n10717__, new_new_n10718__, new_new_n10719__, new_new_n10720__,
    new_new_n10721__, new_new_n10722__, new_new_n10723__, new_new_n10724__,
    new_new_n10725__, new_new_n10726__, new_new_n10727__, new_new_n10728__,
    new_new_n10729__, new_new_n10730__, new_new_n10731__, new_new_n10732__,
    new_new_n10733__, new_new_n10734__, new_new_n10735__, new_new_n10736__,
    new_new_n10737__, new_new_n10738__, new_new_n10739__, new_new_n10740__,
    new_new_n10741__, new_new_n10742__, new_new_n10743__, new_new_n10744__,
    new_new_n10745__, new_new_n10746__, new_new_n10747__, new_new_n10748__,
    new_new_n10749__, new_new_n10750__, new_new_n10751__, new_new_n10752__,
    new_new_n10753__, new_new_n10754__, new_new_n10755__, new_new_n10756__,
    new_new_n10757__, new_new_n10758__, new_new_n10759__, new_new_n10760__,
    new_new_n10761__, new_new_n10762__, new_new_n10763__, new_new_n10764__,
    new_new_n10765__, new_new_n10766__, new_new_n10767__, new_new_n10768__,
    new_new_n10769__, new_new_n10770__, new_new_n10771__, new_new_n10772__,
    new_new_n10773__, new_new_n10774__, new_new_n10775__, new_new_n10776__,
    new_new_n10777__, new_new_n10778__, new_new_n10779__, new_new_n10780__,
    new_new_n10781__, new_new_n10782__, new_new_n10783__, new_new_n10784__,
    new_new_n10785__, new_new_n10786__, new_new_n10787__, new_new_n10788__,
    new_new_n10789__, new_new_n10790__, new_new_n10791__, new_new_n10792__,
    new_new_n10793__, new_new_n10794__, new_new_n10795__, new_new_n10796__,
    new_new_n10797__, new_new_n10798__, new_new_n10799__, new_new_n10800__,
    new_new_n10801__, new_new_n10802__, new_new_n10803__, new_new_n10804__,
    new_new_n10805__, new_new_n10806__, new_new_n10807__, new_new_n10808__,
    new_new_n10809__, new_new_n10810__, new_new_n10811__, new_new_n10812__,
    new_new_n10813__, new_new_n10814__, new_new_n10815__, new_new_n10816__,
    new_new_n10817__, new_new_n10818__, new_new_n10819__, new_new_n10820__,
    new_new_n10821__, new_new_n10822__, new_new_n10823__, new_new_n10824__,
    new_new_n10825__, new_new_n10826__, new_new_n10827__, new_new_n10828__,
    new_new_n10829__, new_new_n10830__, new_new_n10831__, new_new_n10832__,
    new_new_n10833__, new_new_n10834__, new_new_n10835__, new_new_n10836__,
    new_new_n10837__, new_new_n10838__, new_new_n10839__, new_new_n10840__,
    new_new_n10841__, new_new_n10842__, new_new_n10843__, new_new_n10844__,
    new_new_n10845__, new_new_n10846__, new_new_n10847__, new_new_n10848__,
    new_new_n10849__, new_new_n10850__, new_new_n10851__, new_new_n10852__,
    new_new_n10853__, new_new_n10854__, new_new_n10855__, new_new_n10856__,
    new_new_n10857__, new_new_n10858__, new_new_n10859__, new_new_n10860__,
    new_new_n10861__, new_new_n10862__, new_new_n10863__, new_new_n10864__,
    new_new_n10865__, new_new_n10866__, new_new_n10867__, new_new_n10868__,
    new_new_n10869__, new_new_n10870__, new_new_n10871__, new_new_n10872__,
    new_new_n10873__, new_new_n10874__, new_new_n10875__, new_new_n10876__,
    new_new_n10877__, new_new_n10878__, new_new_n10879__, new_new_n10880__,
    new_new_n10881__, new_new_n10882__, new_new_n10883__, new_new_n10884__,
    new_new_n10885__, new_new_n10886__, new_new_n10887__, new_new_n10888__,
    new_new_n10889__, new_new_n10890__, new_new_n10891__, new_new_n10892__,
    new_new_n10893__, new_new_n10894__, new_new_n10895__, new_new_n10896__,
    new_new_n10897__, new_new_n10898__, new_new_n10899__, new_new_n10900__,
    new_new_n10901__, new_new_n10902__, new_new_n10903__, new_new_n10904__,
    new_new_n10905__, new_new_n10906__, new_new_n10907__, new_new_n10908__,
    new_new_n10909__, new_new_n10910__, new_new_n10911__, new_new_n10912__,
    new_new_n10913__, new_new_n10914__, new_new_n10915__, new_new_n10916__,
    new_new_n10917__, new_new_n10918__, new_new_n10919__, new_new_n10920__,
    new_new_n10921__, new_new_n10922__, new_new_n10923__, new_new_n10924__,
    new_new_n10925__, new_new_n10926__, new_new_n10927__, new_new_n10928__,
    new_new_n10929__, new_new_n10930__, new_new_n10931__, new_new_n10932__,
    new_new_n10933__, new_new_n10934__, new_new_n10935__, new_new_n10936__,
    new_new_n10937__, new_new_n10938__, new_new_n10939__, new_new_n10940__,
    new_new_n10941__, new_new_n10942__, new_new_n10943__, new_new_n10944__,
    new_new_n10945__, new_new_n10946__, new_new_n10947__, new_new_n10948__,
    new_new_n10949__, new_new_n10950__, new_new_n10951__, new_new_n10952__,
    new_new_n10953__, new_new_n10954__, new_new_n10955__, new_new_n10956__,
    new_new_n10957__, new_new_n10958__, new_new_n10959__, new_new_n10960__,
    new_new_n10961__, new_new_n10962__, new_new_n10963__, new_new_n10964__,
    new_new_n10965__, new_new_n10966__, new_new_n10967__, new_new_n10968__,
    new_new_n10969__, new_new_n10970__, new_new_n10971__, new_new_n10972__,
    new_new_n10973__, new_new_n10974__, new_new_n10975__, new_new_n10976__,
    new_new_n10977__, new_new_n10978__, new_new_n10979__, new_new_n10980__,
    new_new_n10981__, new_new_n10982__, new_new_n10983__, new_new_n10984__,
    new_new_n10985__, new_new_n10986__, new_new_n10987__, new_new_n10988__,
    new_new_n10989__, new_new_n10990__, new_new_n10991__, new_new_n10992__,
    new_new_n10993__, new_new_n10994__, new_new_n10995__, new_new_n10996__,
    new_new_n10997__, new_new_n10998__, new_new_n10999__, new_new_n11000__,
    new_new_n11001__, new_new_n11002__, new_new_n11003__, new_new_n11004__,
    new_new_n11005__, new_new_n11006__, new_new_n11007__, new_new_n11008__,
    new_new_n11009__, new_new_n11010__, new_new_n11011__, new_new_n11012__,
    new_new_n11013__, new_new_n11014__, new_new_n11015__, new_new_n11016__,
    new_new_n11017__, new_new_n11018__, new_new_n11019__, new_new_n11020__,
    new_new_n11021__, new_new_n11022__, new_new_n11023__, new_new_n11024__,
    new_new_n11025__, new_new_n11026__, new_new_n11027__, new_new_n11028__,
    new_new_n11029__, new_new_n11030__, new_new_n11031__, new_new_n11032__,
    new_new_n11033__, new_new_n11034__, new_new_n11035__, new_new_n11036__,
    new_new_n11037__, new_new_n11038__, new_new_n11039__, new_new_n11040__,
    new_new_n11041__, new_new_n11042__, new_new_n11043__, new_new_n11044__,
    new_new_n11045__, new_new_n11046__, new_new_n11047__, new_new_n11048__,
    new_new_n11049__, new_new_n11050__, new_new_n11051__, new_new_n11052__,
    new_new_n11053__, new_new_n11054__, new_new_n11055__, new_new_n11056__,
    new_new_n11057__, new_new_n11058__, new_new_n11059__, new_new_n11060__,
    new_new_n11061__, new_new_n11062__, new_new_n11063__, new_new_n11064__,
    new_new_n11065__, new_new_n11066__, new_new_n11067__, new_new_n11068__,
    new_new_n11069__, new_new_n11070__, new_new_n11071__, new_new_n11072__,
    new_new_n11073__, new_new_n11074__, new_new_n11075__, new_new_n11076__,
    new_new_n11077__, new_new_n11078__, new_new_n11079__, new_new_n11080__,
    new_new_n11081__, new_new_n11082__, new_new_n11083__, new_new_n11084__,
    new_new_n11085__, new_new_n11086__, new_new_n11087__, new_new_n11088__,
    new_new_n11089__, new_new_n11090__, new_new_n11091__, new_new_n11092__,
    new_new_n11093__, new_new_n11094__, new_new_n11095__, new_new_n11096__,
    new_new_n11097__, new_new_n11098__, new_new_n11099__, new_new_n11100__,
    new_new_n11101__, new_new_n11102__, new_new_n11103__, new_new_n11104__,
    new_new_n11105__, new_new_n11106__, new_new_n11107__, new_new_n11108__,
    new_new_n11109__, new_new_n11110__, new_new_n11111__, new_new_n11112__,
    new_new_n11113__, new_new_n11114__, new_new_n11115__, new_new_n11116__,
    new_new_n11117__, new_new_n11118__, new_new_n11119__, new_new_n11120__,
    new_new_n11121__, new_new_n11122__, new_new_n11123__, new_new_n11124__,
    new_new_n11125__, new_new_n11126__, new_new_n11127__, new_new_n11128__,
    new_new_n11129__, new_new_n11130__, new_new_n11131__, new_new_n11132__,
    new_new_n11133__, new_new_n11134__, new_new_n11135__, new_new_n11136__,
    new_new_n11137__, new_new_n11138__, new_new_n11139__, new_new_n11140__,
    new_new_n11141__, new_new_n11142__, new_new_n11143__, new_new_n11144__,
    new_new_n11145__, new_new_n11146__, new_new_n11147__, new_new_n11148__,
    new_new_n11149__, new_new_n11150__, new_new_n11151__, new_new_n11152__,
    new_new_n11153__, new_new_n11154__, new_new_n11155__, new_new_n11156__,
    new_new_n11157__, new_new_n11158__, new_new_n11159__, new_new_n11160__,
    new_new_n11161__, new_new_n11162__, new_new_n11163__, new_new_n11164__,
    new_new_n11165__, new_new_n11166__, new_new_n11167__, new_new_n11168__,
    new_new_n11169__, new_new_n11170__, new_new_n11171__, new_new_n11172__,
    new_new_n11173__, new_new_n11174__, new_new_n11175__, new_new_n11176__,
    new_new_n11177__, new_new_n11178__, new_new_n11179__, new_new_n11180__,
    new_new_n11181__, new_new_n11182__, new_new_n11183__, new_new_n11184__,
    new_new_n11185__, new_new_n11186__, new_new_n11187__, new_new_n11188__,
    new_new_n11189__, new_new_n11190__, new_new_n11191__, new_new_n11192__,
    new_new_n11193__, new_new_n11194__, new_new_n11195__, new_new_n11196__,
    new_new_n11197__, new_new_n11198__, new_new_n11199__, new_new_n11200__,
    new_new_n11201__, new_new_n11202__, new_new_n11203__, new_new_n11204__,
    new_new_n11205__, new_new_n11206__, new_new_n11207__, new_new_n11208__,
    new_new_n11209__, new_new_n11210__, new_new_n11211__, new_new_n11212__,
    new_new_n11213__, new_new_n11214__, new_new_n11215__, new_new_n11216__,
    new_new_n11217__, new_new_n11218__, new_new_n11219__, new_new_n11220__,
    new_new_n11221__, new_new_n11222__, new_new_n11223__, new_new_n11224__,
    new_new_n11225__, new_new_n11226__, new_new_n11227__, new_new_n11228__,
    new_new_n11229__, new_new_n11230__, new_new_n11231__, new_new_n11232__,
    new_new_n11233__, new_new_n11234__, new_new_n11235__, new_new_n11236__,
    new_new_n11237__, new_new_n11238__, new_new_n11239__, new_new_n11240__,
    new_new_n11241__, new_new_n11242__, new_new_n11243__, new_new_n11244__,
    new_new_n11245__, new_new_n11246__, new_new_n11247__, new_new_n11248__,
    new_new_n11249__, new_new_n11250__, new_new_n11251__, new_new_n11252__,
    new_new_n11253__, new_new_n11254__, new_new_n11255__, new_new_n11256__,
    new_new_n11257__, new_new_n11258__, new_new_n11259__, new_new_n11260__,
    new_new_n11261__, new_new_n11262__, new_new_n11263__, new_new_n11264__,
    new_new_n11265__, new_new_n11266__, new_new_n11267__, new_new_n11268__,
    new_new_n11269__, new_new_n11270__, new_new_n11271__, new_new_n11272__,
    new_new_n11273__, new_new_n11274__, new_new_n11275__, new_new_n11276__,
    new_new_n11277__, new_new_n11278__, new_new_n11279__, new_new_n11280__,
    new_new_n11281__, new_new_n11282__, new_new_n11283__, new_new_n11284__,
    new_new_n11285__, new_new_n11286__, new_new_n11287__, new_new_n11288__,
    new_new_n11289__, new_new_n11290__, new_new_n11291__, new_new_n11292__,
    new_new_n11293__, new_new_n11294__, new_new_n11295__, new_new_n11296__,
    new_new_n11297__, new_new_n11298__, new_new_n11299__, new_new_n11300__,
    new_new_n11301__, new_new_n11302__, new_new_n11303__, new_new_n11304__,
    new_new_n11305__, new_new_n11306__, new_new_n11307__, new_new_n11308__,
    new_new_n11309__, new_new_n11310__, new_new_n11311__, new_new_n11312__,
    new_new_n11313__, new_new_n11314__, new_new_n11315__, new_new_n11316__,
    new_new_n11317__, new_new_n11318__, new_new_n11319__, new_new_n11320__,
    new_new_n11321__, new_new_n11322__, new_new_n11323__, new_new_n11324__,
    new_new_n11325__, new_new_n11326__, new_new_n11327__, new_new_n11328__,
    new_new_n11329__, new_new_n11330__, new_new_n11331__, new_new_n11332__,
    new_new_n11333__, new_new_n11334__, new_new_n11335__, new_new_n11336__,
    new_new_n11337__, new_new_n11338__, new_new_n11339__, new_new_n11340__,
    new_new_n11341__, new_new_n11342__, new_new_n11343__, new_new_n11344__,
    new_new_n11345__, new_new_n11346__, new_new_n11347__, new_new_n11348__,
    new_new_n11349__, new_new_n11350__, new_new_n11351__, new_new_n11352__,
    new_new_n11353__, new_new_n11354__, new_new_n11355__, new_new_n11356__,
    new_new_n11357__, new_new_n11358__, new_new_n11359__, new_new_n11360__,
    new_new_n11361__, new_new_n11362__, new_new_n11363__, new_new_n11364__,
    new_new_n11365__, new_new_n11366__, new_new_n11367__, new_new_n11368__,
    new_new_n11369__, new_new_n11370__, new_new_n11371__, new_new_n11372__,
    new_new_n11373__, new_new_n11374__, new_new_n11375__, new_new_n11376__,
    new_new_n11377__, new_new_n11378__, new_new_n11379__, new_new_n11380__,
    new_new_n11381__, new_new_n11382__, new_new_n11383__, new_new_n11384__,
    new_new_n11385__, new_new_n11386__, new_new_n11387__, new_new_n11388__,
    new_new_n11389__, new_new_n11390__, new_new_n11391__, new_new_n11392__,
    new_new_n11393__, new_new_n11394__, new_new_n11395__, new_new_n11396__,
    new_new_n11397__, new_new_n11398__, new_new_n11399__, new_new_n11400__,
    new_new_n11401__, new_new_n11402__, new_new_n11403__, new_new_n11404__,
    new_new_n11405__, new_new_n11406__, new_new_n11407__, new_new_n11408__,
    new_new_n11409__, new_new_n11410__, new_new_n11411__, new_new_n11412__,
    new_new_n11413__, new_new_n11414__, new_new_n11415__, new_new_n11416__,
    new_new_n11417__, new_new_n11418__, new_new_n11419__, new_new_n11420__,
    new_new_n11421__, new_new_n11422__, new_new_n11423__, new_new_n11424__,
    new_new_n11425__, new_new_n11426__, new_new_n11427__, new_new_n11428__,
    new_new_n11429__, new_new_n11430__, new_new_n11431__, new_new_n11432__,
    new_new_n11433__, new_new_n11434__, new_new_n11435__, new_new_n11436__,
    new_new_n11437__, new_new_n11438__, new_new_n11439__, new_new_n11440__,
    new_new_n11441__, new_new_n11442__, new_new_n11443__, new_new_n11444__,
    new_new_n11445__, new_new_n11446__, new_new_n11447__, new_new_n11448__,
    new_new_n11449__, new_new_n11450__, new_new_n11451__, new_new_n11452__,
    new_new_n11453__, new_new_n11454__, new_new_n11455__, new_new_n11456__,
    new_new_n11457__, new_new_n11458__, new_new_n11459__, new_new_n11460__,
    new_new_n11461__, new_new_n11462__, new_new_n11463__, new_new_n11464__,
    new_new_n11465__, new_new_n11466__, new_new_n11467__, new_new_n11468__,
    new_new_n11469__, new_new_n11470__, new_new_n11471__, new_new_n11472__,
    new_new_n11473__, new_new_n11474__, new_new_n11475__, new_new_n11476__,
    new_new_n11477__, new_new_n11478__, new_new_n11479__, new_new_n11480__,
    new_new_n11481__, new_new_n11482__, new_new_n11483__, new_new_n11484__,
    new_new_n11485__, new_new_n11486__, new_new_n11487__, new_new_n11488__,
    new_new_n11489__, new_new_n11490__, new_new_n11491__, new_new_n11492__,
    new_new_n11493__, new_new_n11494__, new_new_n11495__, new_new_n11496__,
    new_new_n11497__, new_new_n11498__, new_new_n11499__, new_new_n11500__,
    new_new_n11501__, new_new_n11502__, new_new_n11503__, new_new_n11504__,
    new_new_n11505__, new_new_n11506__, new_new_n11507__, new_new_n11508__,
    new_new_n11509__, new_new_n11510__, new_new_n11511__, new_new_n11512__,
    new_new_n11513__, new_new_n11514__, new_new_n11515__, new_new_n11516__,
    new_new_n11517__, new_new_n11518__, new_new_n11519__, new_new_n11520__,
    new_new_n11521__, new_new_n11522__, new_new_n11523__, new_new_n11524__,
    new_new_n11525__, new_new_n11526__, new_new_n11527__, new_new_n11528__,
    new_new_n11529__, new_new_n11530__, new_new_n11531__, new_new_n11532__,
    new_new_n11533__, new_new_n11534__, new_new_n11535__, new_new_n11536__,
    new_new_n11537__, new_new_n11538__, new_new_n11539__, new_new_n11540__,
    new_new_n11541__, new_new_n11542__, new_new_n11543__, new_new_n11544__,
    new_new_n11545__, new_new_n11546__, new_new_n11547__, new_new_n11548__,
    new_new_n11549__, new_new_n11550__, new_new_n11551__, new_new_n11552__,
    new_new_n11553__, new_new_n11554__, new_new_n11555__, new_new_n11556__,
    new_new_n11557__, new_new_n11558__, new_new_n11559__, new_new_n11560__,
    new_new_n11561__, new_new_n11562__, new_new_n11563__, new_new_n11564__,
    new_new_n11565__, new_new_n11566__, new_new_n11567__, new_new_n11568__,
    new_new_n11569__, new_new_n11570__, new_new_n11571__, new_new_n11572__,
    new_new_n11573__, new_new_n11574__, new_new_n11575__, new_new_n11576__,
    new_new_n11577__, new_new_n11578__, new_new_n11579__, new_new_n11580__,
    new_new_n11581__, new_new_n11582__, new_new_n11583__, new_new_n11584__,
    new_new_n11585__, new_new_n11586__, new_new_n11587__, new_new_n11588__,
    new_new_n11589__, new_new_n11590__, new_new_n11591__, new_new_n11592__,
    new_new_n11593__, new_new_n11594__, new_new_n11595__, new_new_n11596__,
    new_new_n11597__, new_new_n11598__, new_new_n11599__, new_new_n11600__,
    new_new_n11601__, new_new_n11602__, new_new_n11603__, new_new_n11604__,
    new_new_n11605__, new_new_n11606__, new_new_n11607__, new_new_n11608__,
    new_new_n11609__, new_new_n11610__, new_new_n11611__, new_new_n11612__,
    new_new_n11613__, new_new_n11614__, new_new_n11615__, new_new_n11616__,
    new_new_n11617__, new_new_n11618__, new_new_n11619__, new_new_n11620__,
    new_new_n11621__, new_new_n11622__, new_new_n11623__, new_new_n11624__,
    new_new_n11625__, new_new_n11626__, new_new_n11627__, new_new_n11628__,
    new_new_n11629__, new_new_n11630__, new_new_n11631__, new_new_n11632__,
    new_new_n11633__, new_new_n11634__, new_new_n11635__, new_new_n11636__,
    new_new_n11637__, new_new_n11638__, new_new_n11639__, new_new_n11640__,
    new_new_n11641__, new_new_n11642__, new_new_n11643__, new_new_n11644__,
    new_new_n11645__, new_new_n11646__, new_new_n11647__, new_new_n11648__,
    new_new_n11649__, new_new_n11650__, new_new_n11651__, new_new_n11652__,
    new_new_n11653__, new_new_n11654__, new_new_n11655__, new_new_n11656__,
    new_new_n11657__, new_new_n11658__, new_new_n11659__, new_new_n11660__,
    new_new_n11661__, new_new_n11662__, new_new_n11663__, new_new_n11664__,
    new_new_n11665__, new_new_n11666__, new_new_n11667__, new_new_n11668__,
    new_new_n11669__, new_new_n11670__, new_new_n11671__, new_new_n11672__,
    new_new_n11673__, new_new_n11674__, new_new_n11675__, new_new_n11676__,
    new_new_n11677__, new_new_n11678__, new_new_n11679__, new_new_n11680__,
    new_new_n11681__, new_new_n11682__, new_new_n11683__, new_new_n11684__,
    new_new_n11685__, new_new_n11686__, new_new_n11687__, new_new_n11688__,
    new_new_n11689__, new_new_n11690__, new_new_n11691__, new_new_n11692__,
    new_new_n11693__, new_new_n11694__, new_new_n11695__, new_new_n11696__,
    new_new_n11697__, new_new_n11698__, new_new_n11699__, new_new_n11700__,
    new_new_n11701__, new_new_n11702__, new_new_n11703__, new_new_n11704__,
    new_new_n11705__, new_new_n11706__, new_new_n11707__, new_new_n11708__,
    new_new_n11709__, new_new_n11710__, new_new_n11711__, new_new_n11712__,
    new_new_n11713__, new_new_n11714__, new_new_n11715__, new_new_n11716__,
    new_new_n11717__, new_new_n11718__, new_new_n11719__, new_new_n11720__,
    new_new_n11721__, new_new_n11722__, new_new_n11723__, new_new_n11724__,
    new_new_n11725__, new_new_n11726__, new_new_n11727__, new_new_n11728__,
    new_new_n11729__, new_new_n11730__, new_new_n11731__, new_new_n11732__,
    new_new_n11733__, new_new_n11734__, new_new_n11735__, new_new_n11736__,
    new_new_n11737__, new_new_n11738__, new_new_n11739__, new_new_n11740__,
    new_new_n11741__, new_new_n11742__, new_new_n11743__, new_new_n11744__,
    new_new_n11745__, new_new_n11746__, new_new_n11747__, new_new_n11748__,
    new_new_n11749__, new_new_n11750__, new_new_n11751__, new_new_n11752__,
    new_new_n11753__, new_new_n11754__, new_new_n11755__, new_new_n11756__,
    new_new_n11757__, new_new_n11758__, new_new_n11759__, new_new_n11760__,
    new_new_n11761__, new_new_n11762__, new_new_n11763__, new_new_n11764__,
    new_new_n11765__, new_new_n11766__, new_new_n11767__, new_new_n11768__,
    new_new_n11769__, new_new_n11770__, new_new_n11771__, new_new_n11772__,
    new_new_n11773__, new_new_n11774__, new_new_n11775__, new_new_n11776__,
    new_new_n11777__, new_new_n11778__, new_new_n11779__, new_new_n11780__,
    new_new_n11781__, new_new_n11782__, new_new_n11783__, new_new_n11784__,
    new_new_n11785__, new_new_n11786__, new_new_n11787__, new_new_n11788__,
    new_new_n11789__, new_new_n11790__, new_new_n11791__, new_new_n11792__,
    new_new_n11793__, new_new_n11794__, new_new_n11795__, new_new_n11796__,
    new_new_n11797__, new_new_n11798__, new_new_n11799__, new_new_n11800__,
    new_new_n11801__, new_new_n11802__, new_new_n11803__, new_new_n11804__,
    new_new_n11805__, new_new_n11806__, new_new_n11807__, new_new_n11808__,
    new_new_n11809__, new_new_n11810__, new_new_n11811__, new_new_n11812__,
    new_new_n11813__, new_new_n11814__, new_new_n11815__, new_new_n11816__,
    new_new_n11817__, new_new_n11818__, new_new_n11819__, new_new_n11820__,
    new_new_n11821__, new_new_n11822__, new_new_n11823__, new_new_n11824__,
    new_new_n11825__, new_new_n11826__, new_new_n11827__, new_new_n11828__,
    new_new_n11829__, new_new_n11830__, new_new_n11831__, new_new_n11832__,
    new_new_n11833__, new_new_n11834__, new_new_n11835__, new_new_n11836__,
    new_new_n11837__, new_new_n11838__, new_new_n11839__, new_new_n11840__,
    new_new_n11841__, new_new_n11842__, new_new_n11843__, new_new_n11844__,
    new_new_n11845__, new_new_n11846__, new_new_n11847__, new_new_n11848__,
    new_new_n11849__, new_new_n11850__, new_new_n11851__, new_new_n11852__,
    new_new_n11853__, new_new_n11854__, new_new_n11855__, new_new_n11856__,
    new_new_n11857__, new_new_n11858__, new_new_n11859__, new_new_n11860__,
    new_new_n11861__, new_new_n11862__, new_new_n11863__, new_new_n11864__,
    new_new_n11865__, new_new_n11866__, new_new_n11867__, new_new_n11868__,
    new_new_n11869__, new_new_n11870__, new_new_n11871__, new_new_n11872__,
    new_new_n11873__, new_new_n11874__, new_new_n11875__, new_new_n11876__,
    new_new_n11877__, new_new_n11878__, new_new_n11879__, new_new_n11880__,
    new_new_n11881__, new_new_n11882__, new_new_n11883__, new_new_n11884__,
    new_new_n11885__, new_new_n11886__, new_new_n11887__, new_new_n11888__,
    new_new_n11889__, new_new_n11890__, new_new_n11891__, new_new_n11892__,
    new_new_n11893__, new_new_n11894__, new_new_n11895__, new_new_n11896__,
    new_new_n11897__, new_new_n11898__, new_new_n11899__, new_new_n11900__,
    new_new_n11901__, new_new_n11902__, new_new_n11903__, new_new_n11904__,
    new_new_n11905__, new_new_n11906__, new_new_n11907__, new_new_n11908__,
    new_new_n11909__, new_new_n11910__, new_new_n11911__, new_new_n11912__,
    new_new_n11913__, new_new_n11914__, new_new_n11915__, new_new_n11916__,
    new_new_n11917__, new_new_n11918__, new_new_n11919__, new_new_n11920__,
    new_new_n11921__, new_new_n11922__, new_new_n11923__, new_new_n11924__,
    new_new_n11925__, new_new_n11926__, new_new_n11927__, new_new_n11928__,
    new_new_n11929__, new_new_n11930__, new_new_n11931__, new_new_n11932__,
    new_new_n11933__, new_new_n11934__, new_new_n11935__, new_new_n11936__,
    new_new_n11937__, new_new_n11938__, new_new_n11939__, new_new_n11940__,
    new_new_n11941__, new_new_n11942__, new_new_n11943__, new_new_n11944__,
    new_new_n11945__, new_new_n11946__, new_new_n11947__, new_new_n11948__,
    new_new_n11949__, new_new_n11950__, new_new_n11951__, new_new_n11952__,
    new_new_n11953__, new_new_n11954__, new_new_n11955__, new_new_n11956__,
    new_new_n11957__, new_new_n11958__, new_new_n11959__, new_new_n11960__,
    new_new_n11961__, new_new_n11962__, new_new_n11963__, new_new_n11964__,
    new_new_n11965__, new_new_n11966__, new_new_n11967__, new_new_n11968__,
    new_new_n11969__, new_new_n11970__, new_new_n11971__, new_new_n11972__,
    new_new_n11973__, new_new_n11974__, new_new_n11975__, new_new_n11976__,
    new_new_n11977__, new_new_n11978__, new_new_n11979__, new_new_n11980__,
    new_new_n11981__, new_new_n11982__, new_new_n11983__, new_new_n11984__,
    new_new_n11985__, new_new_n11986__, new_new_n11987__, new_new_n11988__,
    new_new_n11989__, new_new_n11990__, new_new_n11991__, new_new_n11992__,
    new_new_n11993__, new_new_n11994__, new_new_n11995__, new_new_n11996__,
    new_new_n11997__, new_new_n11998__, new_new_n11999__, new_new_n12000__,
    new_new_n12001__, new_new_n12002__, new_new_n12003__, new_new_n12004__,
    new_new_n12005__, new_new_n12006__, new_new_n12007__, new_new_n12008__,
    new_new_n12009__, new_new_n12010__, new_new_n12011__, new_new_n12012__,
    new_new_n12013__, new_new_n12014__, new_new_n12015__, new_new_n12016__,
    new_new_n12017__, new_new_n12018__, new_new_n12019__, new_new_n12020__,
    new_new_n12021__, new_new_n12022__, new_new_n12023__, new_new_n12024__,
    new_new_n12025__, new_new_n12026__, new_new_n12027__, new_new_n12028__,
    new_new_n12029__, new_new_n12030__, new_new_n12031__, new_new_n12032__,
    new_new_n12033__, new_new_n12034__, new_new_n12035__, new_new_n12036__,
    new_new_n12037__, new_new_n12038__, new_new_n12039__, new_new_n12040__,
    new_new_n12041__, new_new_n12042__, new_new_n12043__, new_new_n12044__,
    new_new_n12045__, new_new_n12046__, new_new_n12047__, new_new_n12048__,
    new_new_n12049__, new_new_n12050__, new_new_n12051__, new_new_n12052__,
    new_new_n12053__, new_new_n12054__, new_new_n12055__, new_new_n12056__,
    new_new_n12057__, new_new_n12058__, new_new_n12059__, new_new_n12060__,
    new_new_n12061__, new_new_n12062__, new_new_n12063__, new_new_n12064__,
    new_new_n12065__, new_new_n12066__, new_new_n12067__, new_new_n12068__,
    new_new_n12069__, new_new_n12070__, new_new_n12071__, new_new_n12072__,
    new_new_n12073__, new_new_n12074__, new_new_n12075__, new_new_n12076__,
    new_new_n12077__, new_new_n12078__, new_new_n12079__, new_new_n12080__,
    new_new_n12081__, new_new_n12082__, new_new_n12083__, new_new_n12084__,
    new_new_n12085__, new_new_n12086__, new_new_n12087__, new_new_n12088__,
    new_new_n12089__, new_new_n12090__, new_new_n12091__, new_new_n12092__,
    new_new_n12093__, new_new_n12094__, new_new_n12095__, new_new_n12096__,
    new_new_n12097__, new_new_n12098__, new_new_n12099__, new_new_n12100__,
    new_new_n12101__, new_new_n12102__, new_new_n12103__, new_new_n12104__,
    new_new_n12105__, new_new_n12106__, new_new_n12107__, new_new_n12108__,
    new_new_n12109__, new_new_n12110__, new_new_n12111__, new_new_n12112__,
    new_new_n12113__, new_new_n12114__, new_new_n12115__, new_new_n12116__,
    new_new_n12117__, new_new_n12118__, new_new_n12119__, new_new_n12120__,
    new_new_n12121__, new_new_n12122__, new_new_n12123__, new_new_n12124__,
    new_new_n12125__, new_new_n12126__, new_new_n12127__, new_new_n12128__,
    new_new_n12129__, new_new_n12130__, new_new_n12131__, new_new_n12132__,
    new_new_n12133__, new_new_n12134__, new_new_n12135__, new_new_n12136__,
    new_new_n12137__, new_new_n12138__, new_new_n12139__, new_new_n12140__,
    new_new_n12141__, new_new_n12142__, new_new_n12143__, new_new_n12144__,
    new_new_n12145__, new_new_n12146__, new_new_n12147__, new_new_n12148__,
    new_new_n12149__, new_new_n12150__, new_new_n12151__, new_new_n12152__,
    new_new_n12153__, new_new_n12154__, new_new_n12155__, new_new_n12156__,
    new_new_n12157__, new_new_n12158__, new_new_n12159__, new_new_n12160__,
    new_new_n12161__, new_new_n12162__, new_new_n12163__, new_new_n12164__,
    new_new_n12165__, new_new_n12166__, new_new_n12167__, new_new_n12168__,
    new_new_n12169__, new_new_n12170__, new_new_n12171__, new_new_n12172__,
    new_new_n12173__, new_new_n12174__, new_new_n12175__, new_new_n12176__,
    new_new_n12177__, new_new_n12178__, new_new_n12179__, new_new_n12180__,
    new_new_n12181__, new_new_n12182__, new_new_n12183__, new_new_n12184__,
    new_new_n12185__, new_new_n12186__, new_new_n12187__, new_new_n12188__,
    new_new_n12189__, new_new_n12190__, new_new_n12191__, new_new_n12192__,
    new_new_n12193__, new_new_n12194__, new_new_n12195__, new_new_n12196__,
    new_new_n12197__, new_new_n12198__, new_new_n12199__, new_new_n12200__,
    new_new_n12201__, new_new_n12202__, new_new_n12203__, new_new_n12204__,
    new_new_n12205__, new_new_n12206__, new_new_n12207__, new_new_n12208__,
    new_new_n12209__, new_new_n12210__, new_new_n12211__, new_new_n12212__,
    new_new_n12213__, new_new_n12214__, new_new_n12215__, new_new_n12216__,
    new_new_n12217__, new_new_n12218__, new_new_n12219__, new_new_n12220__,
    new_new_n12221__, new_new_n12222__, new_new_n12223__, new_new_n12224__,
    new_new_n12225__, new_new_n12226__, new_new_n12227__, new_new_n12228__,
    new_new_n12229__, new_new_n12230__, new_new_n12231__, new_new_n12232__,
    new_new_n12233__, new_new_n12234__, new_new_n12235__, new_new_n12236__,
    new_new_n12237__, new_new_n12238__, new_new_n12239__, new_new_n12240__,
    new_new_n12241__, new_new_n12242__, new_new_n12243__, new_new_n12244__,
    new_new_n12245__, new_new_n12246__, new_new_n12247__, new_new_n12248__,
    new_new_n12249__, new_new_n12250__, new_new_n12251__, new_new_n12252__,
    new_new_n12253__, new_new_n12254__, new_new_n12255__, new_new_n12256__,
    new_new_n12257__, new_new_n12258__, new_new_n12259__, new_new_n12260__,
    new_new_n12261__, new_new_n12262__, new_new_n12263__, new_new_n12264__,
    new_new_n12265__, new_new_n12266__, new_new_n12267__, new_new_n12268__,
    new_new_n12269__, new_new_n12270__, new_new_n12271__, new_new_n12272__,
    new_new_n12273__, new_new_n12274__, new_new_n12275__, new_new_n12276__,
    new_new_n12277__, new_new_n12278__, new_new_n12279__, new_new_n12280__,
    new_new_n12281__, new_new_n12282__, new_new_n12283__, new_new_n12284__,
    new_new_n12285__, new_new_n12286__, new_new_n12287__, new_new_n12288__,
    new_new_n12289__, new_new_n12290__, new_new_n12291__, new_new_n12292__,
    new_new_n12293__, new_new_n12294__, new_new_n12295__, new_new_n12296__,
    new_new_n12297__, new_new_n12298__, new_new_n12299__, new_new_n12300__,
    new_new_n12301__, new_new_n12302__, new_new_n12303__, new_new_n12304__,
    new_new_n12305__, new_new_n12306__, new_new_n12307__, new_new_n12308__,
    new_new_n12309__, new_new_n12310__, new_new_n12311__, new_new_n12312__,
    new_new_n12313__, new_new_n12314__, new_new_n12315__, new_new_n12316__,
    new_new_n12317__, new_new_n12318__, new_new_n12319__, new_new_n12320__,
    new_new_n12321__, new_new_n12322__, new_new_n12323__, new_new_n12324__,
    new_new_n12325__, new_new_n12326__, new_new_n12327__, new_new_n12328__,
    new_new_n12329__, new_new_n12330__, new_new_n12331__, new_new_n12332__,
    new_new_n12333__, new_new_n12334__, new_new_n12335__, new_new_n12336__,
    new_new_n12337__, new_new_n12338__, new_new_n12339__, new_new_n12340__,
    new_new_n12341__, new_new_n12342__, new_new_n12343__, new_new_n12344__,
    new_new_n12345__, new_new_n12346__, new_new_n12347__, new_new_n12348__,
    new_new_n12349__, new_new_n12350__, new_new_n12351__, new_new_n12352__,
    new_new_n12353__, new_new_n12354__, new_new_n12355__, new_new_n12356__,
    new_new_n12357__, new_new_n12358__, new_new_n12359__, new_new_n12360__,
    new_new_n12361__, new_new_n12362__, new_new_n12363__, new_new_n12364__,
    new_new_n12365__, new_new_n12366__, new_new_n12367__, new_new_n12368__,
    new_new_n12369__, new_new_n12370__, new_new_n12371__, new_new_n12372__,
    new_new_n12373__, new_new_n12374__, new_new_n12375__, new_new_n12376__,
    new_new_n12377__, new_new_n12378__, new_new_n12379__, new_new_n12380__,
    new_new_n12381__, new_new_n12382__, new_new_n12383__, new_new_n12384__,
    new_new_n12385__, new_new_n12386__, new_new_n12387__, new_new_n12388__,
    new_new_n12389__, new_new_n12390__, new_new_n12391__, new_new_n12392__,
    new_new_n12393__, new_new_n12394__, new_new_n12395__, new_new_n12396__,
    new_new_n12397__, new_new_n12398__, new_new_n12399__, new_new_n12400__,
    new_new_n12401__, new_new_n12402__, new_new_n12403__, new_new_n12404__,
    new_new_n12405__, new_new_n12406__, new_new_n12407__, new_new_n12408__,
    new_new_n12409__, new_new_n12410__, new_new_n12411__, new_new_n12412__,
    new_new_n12413__, new_new_n12414__, new_new_n12415__, new_new_n12416__,
    new_new_n12417__, new_new_n12418__, new_new_n12419__, new_new_n12420__,
    new_new_n12421__, new_new_n12422__, new_new_n12423__, new_new_n12424__,
    new_new_n12425__, new_new_n12426__, new_new_n12427__, new_new_n12428__,
    new_new_n12429__, new_new_n12430__, new_new_n12431__, new_new_n12432__,
    new_new_n12433__, new_new_n12434__, new_new_n12435__, new_new_n12436__,
    new_new_n12437__, new_new_n12438__, new_new_n12439__, new_new_n12440__,
    new_new_n12441__, new_new_n12442__, new_new_n12443__, new_new_n12444__,
    new_new_n12445__, new_new_n12446__, new_new_n12447__, new_new_n12448__,
    new_new_n12449__, new_new_n12450__, new_new_n12451__, new_new_n12452__,
    new_new_n12453__, new_new_n12454__, new_new_n12455__, new_new_n12456__,
    new_new_n12457__, new_new_n12458__, new_new_n12459__, new_new_n12460__,
    new_new_n12461__, new_new_n12462__, new_new_n12463__, new_new_n12464__,
    new_new_n12465__, new_new_n12466__, new_new_n12467__, new_new_n12468__,
    new_new_n12469__, new_new_n12470__, new_new_n12471__, new_new_n12472__,
    new_new_n12473__, new_new_n12474__, new_new_n12475__, new_new_n12476__,
    new_new_n12477__, new_new_n12478__, new_new_n12479__, new_new_n12480__,
    new_new_n12481__, new_new_n12482__, new_new_n12483__, new_new_n12484__,
    new_new_n12485__, new_new_n12486__, new_new_n12487__, new_new_n12488__,
    new_new_n12489__, new_new_n12490__, new_new_n12491__, new_new_n12492__,
    new_new_n12493__, new_new_n12494__, new_new_n12495__, new_new_n12496__,
    new_new_n12497__, new_new_n12498__, new_new_n12499__, new_new_n12500__,
    new_new_n12501__, new_new_n12502__, new_new_n12503__, new_new_n12504__,
    new_new_n12505__, new_new_n12506__, new_new_n12507__, new_new_n12508__,
    new_new_n12509__, new_new_n12510__, new_new_n12511__, new_new_n12512__,
    new_new_n12513__, new_new_n12514__, new_new_n12515__, new_new_n12516__,
    new_new_n12517__, new_new_n12518__, new_new_n12519__, new_new_n12520__,
    new_new_n12521__, new_new_n12522__, new_new_n12523__, new_new_n12524__,
    new_new_n12525__, new_new_n12526__, new_new_n12527__, new_new_n12528__,
    new_new_n12529__, new_new_n12530__, new_new_n12531__, new_new_n12532__,
    new_new_n12533__, new_new_n12534__, new_new_n12535__, new_new_n12536__,
    new_new_n12537__, new_new_n12538__, new_new_n12539__, new_new_n12540__,
    new_new_n12541__, new_new_n12542__, new_new_n12543__, new_new_n12544__,
    new_new_n12545__, new_new_n12546__, new_new_n12547__, new_new_n12548__,
    new_new_n12549__, new_new_n12550__, new_new_n12551__, new_new_n12552__,
    new_new_n12553__, new_new_n12554__, new_new_n12555__, new_new_n12556__,
    new_new_n12557__, new_new_n12558__, new_new_n12559__, new_new_n12560__,
    new_new_n12561__, new_new_n12562__, new_new_n12563__, new_new_n12564__,
    new_new_n12565__, new_new_n12566__, new_new_n12567__, new_new_n12568__,
    new_new_n12569__, new_new_n12570__, new_new_n12571__, new_new_n12572__,
    new_new_n12573__, new_new_n12574__, new_new_n12575__, new_new_n12576__,
    new_new_n12577__, new_new_n12578__, new_new_n12579__, new_new_n12580__,
    new_new_n12581__, new_new_n12582__, new_new_n12583__, new_new_n12584__,
    new_new_n12585__, new_new_n12586__, new_new_n12587__, new_new_n12588__,
    new_new_n12589__, new_new_n12590__, new_new_n12591__, new_new_n12592__,
    new_new_n12593__, new_new_n12594__, new_new_n12595__, new_new_n12596__,
    new_new_n12597__, new_new_n12598__, new_new_n12599__, new_new_n12600__,
    new_new_n12601__, new_new_n12602__, new_new_n12603__, new_new_n12604__,
    new_new_n12605__, new_new_n12606__, new_new_n12607__, new_new_n12608__,
    new_new_n12609__, new_new_n12610__, new_new_n12611__, new_new_n12612__,
    new_new_n12613__, new_new_n12614__, new_new_n12615__, new_new_n12616__,
    new_new_n12617__, new_new_n12618__, new_new_n12619__, new_new_n12620__,
    new_new_n12621__, new_new_n12622__, new_new_n12623__, new_new_n12624__,
    new_new_n12625__, new_new_n12626__, new_new_n12627__, new_new_n12628__,
    new_new_n12629__, new_new_n12630__, new_new_n12631__, new_new_n12632__,
    new_new_n12633__, new_new_n12634__, new_new_n12635__, new_new_n12636__,
    new_new_n12637__, new_new_n12638__, new_new_n12639__, new_new_n12640__,
    new_new_n12641__, new_new_n12642__, new_new_n12643__, new_new_n12644__,
    new_new_n12645__, new_new_n12646__, new_new_n12647__, new_new_n12648__,
    new_new_n12649__, new_new_n12650__, new_new_n12651__, new_new_n12652__,
    new_new_n12653__, new_new_n12654__, new_new_n12655__, new_new_n12656__,
    new_new_n12657__, new_new_n12658__, new_new_n12659__, new_new_n12660__,
    new_new_n12661__, new_new_n12662__, new_new_n12663__, new_new_n12664__,
    new_new_n12665__, new_new_n12666__, new_new_n12667__, new_new_n12668__,
    new_new_n12669__, new_new_n12670__, new_new_n12671__, new_new_n12672__,
    new_new_n12673__, new_new_n12674__, new_new_n12675__, new_new_n12676__,
    new_new_n12677__, new_new_n12678__, new_new_n12679__, new_new_n12680__,
    new_new_n12681__, new_new_n12682__, new_new_n12683__, new_new_n12684__,
    new_new_n12685__, new_new_n12686__, new_new_n12687__, new_new_n12688__,
    new_new_n12689__, new_new_n12690__, new_new_n12691__, new_new_n12692__,
    new_new_n12693__, new_new_n12694__, new_new_n12695__, new_new_n12696__,
    new_new_n12697__, new_new_n12698__, new_new_n12699__, new_new_n12700__,
    new_new_n12701__, new_new_n12702__, new_new_n12703__, new_new_n12704__,
    new_new_n12705__, new_new_n12706__, new_new_n12707__, new_new_n12708__,
    new_new_n12709__, new_new_n12710__, new_new_n12711__, new_new_n12712__,
    new_new_n12713__, new_new_n12714__, new_new_n12715__, new_new_n12716__,
    new_new_n12717__, new_new_n12718__, new_new_n12719__, new_new_n12720__,
    new_new_n12721__, new_new_n12722__, new_new_n12723__, new_new_n12724__,
    new_new_n12725__, new_new_n12726__, new_new_n12727__, new_new_n12728__,
    new_new_n12729__, new_new_n12730__, new_new_n12731__, new_new_n12732__,
    new_new_n12733__, new_new_n12734__, new_new_n12735__, new_new_n12736__,
    new_new_n12737__, new_new_n12738__, new_new_n12739__, new_new_n12740__,
    new_new_n12741__, new_new_n12742__, new_new_n12743__, new_new_n12744__,
    new_new_n12745__, new_new_n12746__, new_new_n12747__, new_new_n12748__,
    new_new_n12749__, new_new_n12750__, new_new_n12751__, new_new_n12752__,
    new_new_n12753__, new_new_n12754__, new_new_n12755__, new_new_n12756__,
    new_new_n12757__, new_new_n12758__, new_new_n12759__, new_new_n12760__,
    new_new_n12761__, new_new_n12762__, new_new_n12763__, new_new_n12764__,
    new_new_n12765__, new_new_n12766__, new_new_n12767__, new_new_n12768__,
    new_new_n12769__, new_new_n12770__, new_new_n12771__, new_new_n12772__,
    new_new_n12773__, new_new_n12774__, new_new_n12775__, new_new_n12776__,
    new_new_n12777__, new_new_n12778__, new_new_n12779__, new_new_n12780__,
    new_new_n12781__, new_new_n12782__, new_new_n12783__, new_new_n12784__,
    new_new_n12785__, new_new_n12786__, new_new_n12787__, new_new_n12788__,
    new_new_n12789__, new_new_n12790__, new_new_n12791__, new_new_n12792__,
    new_new_n12793__, new_new_n12794__, new_new_n12795__, new_new_n12796__,
    new_new_n12797__, new_new_n12798__, new_new_n12799__, new_new_n12800__,
    new_new_n12801__, new_new_n12802__, new_new_n12803__, new_new_n12804__,
    new_new_n12805__, new_new_n12806__, new_new_n12807__, new_new_n12808__,
    new_new_n12809__, new_new_n12810__, new_new_n12811__, new_new_n12812__,
    new_new_n12813__, new_new_n12814__, new_new_n12815__, new_new_n12816__,
    new_new_n12817__, new_new_n12818__, new_new_n12819__, new_new_n12820__,
    new_new_n12821__, new_new_n12822__, new_new_n12823__, new_new_n12824__,
    new_new_n12825__, new_new_n12826__, new_new_n12827__, new_new_n12828__,
    new_new_n12829__, new_new_n12830__, new_new_n12831__, new_new_n12832__,
    new_new_n12833__, new_new_n12834__, new_new_n12835__, new_new_n12836__,
    new_new_n12837__, new_new_n12838__, new_new_n12839__, new_new_n12840__,
    new_new_n12841__, new_new_n12842__, new_new_n12843__, new_new_n12844__,
    new_new_n12845__, new_new_n12846__, new_new_n12847__, new_new_n12848__,
    new_new_n12849__, new_new_n12850__, new_new_n12851__, new_new_n12852__,
    new_new_n12853__, new_new_n12854__, new_new_n12855__, new_new_n12856__,
    new_new_n12857__, new_new_n12858__, new_new_n12859__, new_new_n12860__,
    new_new_n12861__, new_new_n12862__, new_new_n12863__, new_new_n12864__,
    new_new_n12865__, new_new_n12866__, new_new_n12867__, new_new_n12868__,
    new_new_n12869__, new_new_n12870__, new_new_n12871__, new_new_n12872__,
    new_new_n12873__, new_new_n12874__, new_new_n12875__, new_new_n12876__,
    new_new_n12877__, new_new_n12878__, new_new_n12879__, new_new_n12880__,
    new_new_n12881__, new_new_n12882__, new_new_n12883__, new_new_n12884__,
    new_new_n12885__, new_new_n12886__, new_new_n12887__, new_new_n12888__,
    new_new_n12889__, new_new_n12890__, new_new_n12891__, new_new_n12892__,
    new_new_n12893__, new_new_n12894__, new_new_n12895__, new_new_n12896__,
    new_new_n12897__, new_new_n12898__, new_new_n12899__, new_new_n12900__,
    new_new_n12901__, new_new_n12902__, new_new_n12903__, new_new_n12904__,
    new_new_n12905__, new_new_n12906__, new_new_n12907__, new_new_n12908__,
    new_new_n12909__, new_new_n12910__, new_new_n12911__, new_new_n12912__,
    new_new_n12913__, new_new_n12914__, new_new_n12915__, new_new_n12916__,
    new_new_n12917__, new_new_n12918__, new_new_n12919__, new_new_n12920__,
    new_new_n12921__, new_new_n12922__, new_new_n12923__, new_new_n12924__,
    new_new_n12925__, new_new_n12926__, new_new_n12927__, new_new_n12928__,
    new_new_n12929__, new_new_n12930__, new_new_n12931__, new_new_n12932__,
    new_new_n12933__, new_new_n12934__, new_new_n12935__, new_new_n12936__,
    new_new_n12937__, new_new_n12938__, new_new_n12939__, new_new_n12940__,
    new_new_n12941__, new_new_n12942__, new_new_n12943__, new_new_n12944__,
    new_new_n12945__, new_new_n12946__, new_new_n12947__, new_new_n12948__,
    new_new_n12949__, new_new_n12950__, new_new_n12951__, new_new_n12952__,
    new_new_n12953__, new_new_n12954__, new_new_n12955__, new_new_n12956__,
    new_new_n12957__, new_new_n12958__, new_new_n12959__, new_new_n12960__,
    new_new_n12961__, new_new_n12962__, new_new_n12963__, new_new_n12964__,
    new_new_n12965__, new_new_n12966__, new_new_n12967__, new_new_n12968__,
    new_new_n12969__, new_new_n12970__, new_new_n12971__, new_new_n12972__,
    new_new_n12973__, new_new_n12974__, new_new_n12975__, new_new_n12976__,
    new_new_n12977__, new_new_n12978__, new_new_n12979__, new_new_n12980__,
    new_new_n12981__, new_new_n12982__, new_new_n12983__, new_new_n12984__,
    new_new_n12985__, new_new_n12986__, new_new_n12987__, new_new_n12988__,
    new_new_n12989__, new_new_n12990__, new_new_n12991__, new_new_n12992__,
    new_new_n12993__, new_new_n12994__, new_new_n12995__, new_new_n12996__,
    new_new_n12997__, new_new_n12998__, new_new_n12999__, new_new_n13000__,
    new_new_n13001__, new_new_n13002__, new_new_n13003__, new_new_n13004__,
    new_new_n13005__, new_new_n13006__, new_new_n13007__, new_new_n13008__,
    new_new_n13009__, new_new_n13010__, new_new_n13011__, new_new_n13012__,
    new_new_n13013__, new_new_n13014__, new_new_n13015__, new_new_n13016__,
    new_new_n13017__, new_new_n13018__, new_new_n13019__, new_new_n13020__,
    new_new_n13021__, new_new_n13022__, new_new_n13023__, new_new_n13024__,
    new_new_n13025__, new_new_n13026__, new_new_n13027__, new_new_n13028__,
    new_new_n13029__, new_new_n13030__, new_new_n13031__, new_new_n13032__,
    new_new_n13033__, new_new_n13034__, new_new_n13035__, new_new_n13036__,
    new_new_n13037__, new_new_n13038__, new_new_n13039__, new_new_n13040__,
    new_new_n13041__, new_new_n13042__, new_new_n13043__, new_new_n13044__,
    new_new_n13045__, new_new_n13046__, new_new_n13047__, new_new_n13048__,
    new_new_n13049__, new_new_n13050__, new_new_n13051__, new_new_n13052__,
    new_new_n13053__, new_new_n13054__, new_new_n13055__, new_new_n13056__,
    new_new_n13057__, new_new_n13058__, new_new_n13059__, new_new_n13060__,
    new_new_n13061__, new_new_n13062__, new_new_n13063__, new_new_n13064__,
    new_new_n13065__, new_new_n13066__, new_new_n13067__, new_new_n13068__,
    new_new_n13069__, new_new_n13070__, new_new_n13071__, new_new_n13072__,
    new_new_n13073__, new_new_n13074__, new_new_n13075__, new_new_n13076__,
    new_new_n13077__, new_new_n13078__, new_new_n13079__, new_new_n13080__,
    new_new_n13081__, new_new_n13082__, new_new_n13083__, new_new_n13084__,
    new_new_n13085__, new_new_n13086__, new_new_n13087__, new_new_n13088__,
    new_new_n13089__, new_new_n13090__, new_new_n13091__, new_new_n13092__,
    new_new_n13093__, new_new_n13094__, new_new_n13095__, new_new_n13096__,
    new_new_n13097__, new_new_n13098__, new_new_n13099__, new_new_n13100__,
    new_new_n13101__, new_new_n13102__, new_new_n13103__, new_new_n13104__,
    new_new_n13105__, new_new_n13106__, new_new_n13107__, new_new_n13108__,
    new_new_n13109__, new_new_n13110__, new_new_n13111__, new_new_n13112__,
    new_new_n13113__, new_new_n13114__, new_new_n13115__, new_new_n13116__,
    new_new_n13117__, new_new_n13118__, new_new_n13119__, new_new_n13120__,
    new_new_n13121__, new_new_n13122__, new_new_n13123__, new_new_n13124__,
    new_new_n13125__, new_new_n13126__, new_new_n13127__, new_new_n13128__,
    new_new_n13129__, new_new_n13130__, new_new_n13131__, new_new_n13132__,
    new_new_n13133__, new_new_n13134__, new_new_n13135__, new_new_n13136__,
    new_new_n13137__, new_new_n13138__, new_new_n13139__, new_new_n13140__,
    new_new_n13141__, new_new_n13142__, new_new_n13143__, new_new_n13144__,
    new_new_n13145__, new_new_n13146__, new_new_n13147__, new_new_n13148__,
    new_new_n13149__, new_new_n13150__, new_new_n13151__, new_new_n13152__,
    new_new_n13153__, new_new_n13154__, new_new_n13155__, new_new_n13156__,
    new_new_n13157__, new_new_n13158__, new_new_n13159__, new_new_n13160__,
    new_new_n13161__, new_new_n13162__, new_new_n13163__, new_new_n13164__,
    new_new_n13165__, new_new_n13166__, new_new_n13167__, new_new_n13168__,
    new_new_n13169__, new_new_n13170__, new_new_n13171__, new_new_n13172__,
    new_new_n13173__, new_new_n13174__, new_new_n13175__, new_new_n13176__,
    new_new_n13177__, new_new_n13178__, new_new_n13179__, new_new_n13180__,
    new_new_n13181__, new_new_n13182__, new_new_n13183__, new_new_n13184__,
    new_new_n13185__, new_new_n13186__, new_new_n13187__, new_new_n13188__,
    new_new_n13189__, new_new_n13190__, new_new_n13191__, new_new_n13192__,
    new_new_n13193__, new_new_n13194__, new_new_n13195__, new_new_n13196__,
    new_new_n13197__, new_new_n13198__, new_new_n13199__, new_new_n13200__,
    new_new_n13201__, new_new_n13202__, new_new_n13203__, new_new_n13204__,
    new_new_n13205__, new_new_n13206__, new_new_n13207__, new_new_n13208__,
    new_new_n13209__, new_new_n13210__, new_new_n13211__, new_new_n13212__,
    new_new_n13213__, new_new_n13214__, new_new_n13215__, new_new_n13216__,
    new_new_n13217__, new_new_n13218__, new_new_n13219__, new_new_n13220__,
    new_new_n13221__, new_new_n13222__, new_new_n13223__, new_new_n13224__,
    new_new_n13225__, new_new_n13226__, new_new_n13227__, new_new_n13228__,
    new_new_n13229__, new_new_n13230__, new_new_n13231__, new_new_n13232__,
    new_new_n13233__, new_new_n13234__, new_new_n13235__, new_new_n13236__,
    new_new_n13237__, new_new_n13238__, new_new_n13239__, new_new_n13240__,
    new_new_n13241__, new_new_n13242__, new_new_n13243__, new_new_n13244__,
    new_new_n13245__, new_new_n13246__, new_new_n13247__, new_new_n13248__,
    new_new_n13249__, new_new_n13250__, new_new_n13251__, new_new_n13252__,
    new_new_n13253__, new_new_n13254__, new_new_n13255__, new_new_n13256__,
    new_new_n13257__, new_new_n13258__, new_new_n13259__, new_new_n13260__,
    new_new_n13261__, new_new_n13262__, new_new_n13263__, new_new_n13264__,
    new_new_n13265__, new_new_n13266__, new_new_n13267__, new_new_n13268__,
    new_new_n13269__, new_new_n13270__, new_new_n13271__, new_new_n13272__,
    new_new_n13273__, new_new_n13274__, new_new_n13275__, new_new_n13276__,
    new_new_n13277__, new_new_n13278__, new_new_n13279__, new_new_n13280__,
    new_new_n13281__, new_new_n13282__, new_new_n13283__, new_new_n13284__,
    new_new_n13285__, new_new_n13286__, new_new_n13287__, new_new_n13288__,
    new_new_n13289__, new_new_n13290__, new_new_n13291__, new_new_n13292__,
    new_new_n13293__, new_new_n13294__, new_new_n13295__, new_new_n13296__,
    new_new_n13297__, new_new_n13298__, new_new_n13299__, new_new_n13300__,
    new_new_n13301__, new_new_n13302__, new_new_n13303__, new_new_n13304__,
    new_new_n13305__, new_new_n13306__, new_new_n13307__, new_new_n13308__,
    new_new_n13309__, new_new_n13310__, new_new_n13311__, new_new_n13312__,
    new_new_n13313__, new_new_n13314__, new_new_n13315__, new_new_n13316__,
    new_new_n13317__, new_new_n13318__, new_new_n13319__, new_new_n13320__,
    new_new_n13321__, new_new_n13322__, new_new_n13323__, new_new_n13324__,
    new_new_n13325__, new_new_n13326__, new_new_n13327__, new_new_n13328__,
    new_new_n13329__, new_new_n13330__, new_new_n13331__, new_new_n13332__,
    new_new_n13333__, new_new_n13334__, new_new_n13335__, new_new_n13336__,
    new_new_n13337__, new_new_n13338__, new_new_n13339__, new_new_n13340__,
    new_new_n13341__, new_new_n13342__, new_new_n13343__, new_new_n13344__,
    new_new_n13345__, new_new_n13346__, new_new_n13347__, new_new_n13348__,
    new_new_n13349__, new_new_n13350__, new_new_n13351__, new_new_n13352__,
    new_new_n13353__, new_new_n13354__, new_new_n13355__, new_new_n13356__,
    new_new_n13357__, new_new_n13358__, new_new_n13359__, new_new_n13360__,
    new_new_n13361__, new_new_n13362__, new_new_n13363__, new_new_n13364__,
    new_new_n13365__, new_new_n13366__, new_new_n13367__, new_new_n13368__,
    new_new_n13369__, new_new_n13370__, new_new_n13371__, new_new_n13372__,
    new_new_n13373__, new_new_n13374__, new_new_n13375__, new_new_n13376__,
    new_new_n13377__, new_new_n13378__, new_new_n13379__, new_new_n13380__,
    new_new_n13381__, new_new_n13382__, new_new_n13383__, new_new_n13384__,
    new_new_n13385__, new_new_n13386__, new_new_n13387__, new_new_n13388__,
    new_new_n13389__, new_new_n13390__, new_new_n13391__, new_new_n13392__,
    new_new_n13393__, new_new_n13394__, new_new_n13395__, new_new_n13396__,
    new_new_n13397__, new_new_n13398__, new_new_n13399__, new_new_n13400__,
    new_new_n13401__, new_new_n13402__, new_new_n13403__, new_new_n13404__,
    new_new_n13405__, new_new_n13406__, new_new_n13407__, new_new_n13408__,
    new_new_n13409__, new_new_n13410__, new_new_n13411__, new_new_n13412__,
    new_new_n13413__, new_new_n13414__, new_new_n13415__, new_new_n13416__,
    new_new_n13417__, new_new_n13418__, new_new_n13419__, new_new_n13420__,
    new_new_n13421__, new_new_n13422__, new_new_n13423__, new_new_n13424__,
    new_new_n13425__, new_new_n13426__, new_new_n13427__, new_new_n13428__,
    new_new_n13429__, new_new_n13430__, new_new_n13431__, new_new_n13432__,
    new_new_n13433__, new_new_n13434__, new_new_n13435__, new_new_n13436__,
    new_new_n13437__, new_new_n13438__, new_new_n13439__, new_new_n13440__,
    new_new_n13441__, new_new_n13442__, new_new_n13443__, new_new_n13444__,
    new_new_n13445__, new_new_n13446__, new_new_n13447__, new_new_n13448__,
    new_new_n13449__, new_new_n13450__, new_new_n13451__, new_new_n13452__,
    new_new_n13453__, new_new_n13454__, new_new_n13455__, new_new_n13456__,
    new_new_n13457__, new_new_n13458__, new_new_n13459__, new_new_n13460__,
    new_new_n13461__, new_new_n13462__, new_new_n13463__, new_new_n13464__,
    new_new_n13465__, new_new_n13466__, new_new_n13467__, new_new_n13468__,
    new_new_n13469__, new_new_n13470__, new_new_n13471__, new_new_n13472__,
    new_new_n13473__, new_new_n13474__, new_new_n13475__, new_new_n13476__,
    new_new_n13477__, new_new_n13478__, new_new_n13479__, new_new_n13480__,
    new_new_n13481__, new_new_n13482__, new_new_n13483__, new_new_n13484__,
    new_new_n13485__, new_new_n13486__, new_new_n13487__, new_new_n13488__,
    new_new_n13489__, new_new_n13490__, new_new_n13491__, new_new_n13492__,
    new_new_n13493__, new_new_n13494__, new_new_n13495__, new_new_n13496__,
    new_new_n13497__, new_new_n13498__, new_new_n13499__, new_new_n13500__,
    new_new_n13501__, new_new_n13502__, new_new_n13503__, new_new_n13504__,
    new_new_n13505__, new_new_n13506__, new_new_n13507__, new_new_n13508__,
    new_new_n13509__, new_new_n13510__, new_new_n13511__, new_new_n13512__,
    new_new_n13513__, new_new_n13514__, new_new_n13515__, new_new_n13516__,
    new_new_n13517__, new_new_n13518__, new_new_n13519__, new_new_n13520__,
    new_new_n13521__, new_new_n13522__, new_new_n13523__, new_new_n13524__,
    new_new_n13525__, new_new_n13526__, new_new_n13527__, new_new_n13528__,
    new_new_n13529__, new_new_n13530__, new_new_n13531__, new_new_n13532__,
    new_new_n13533__, new_new_n13534__, new_new_n13535__, new_new_n13536__,
    new_new_n13537__, new_new_n13538__, new_new_n13539__, new_new_n13540__,
    new_new_n13541__, new_new_n13542__, new_new_n13543__, new_new_n13544__,
    new_new_n13545__, new_new_n13546__, new_new_n13547__, new_new_n13548__,
    new_new_n13549__, new_new_n13550__, new_new_n13551__, new_new_n13552__,
    new_new_n13553__, new_new_n13554__, new_new_n13555__, new_new_n13556__,
    new_new_n13557__, new_new_n13558__, new_new_n13559__, new_new_n13560__,
    new_new_n13561__, new_new_n13562__, new_new_n13563__, new_new_n13564__,
    new_new_n13565__, new_new_n13566__, new_new_n13567__, new_new_n13568__,
    new_new_n13569__, new_new_n13570__, new_new_n13571__, new_new_n13572__,
    new_new_n13573__, new_new_n13574__, new_new_n13575__, new_new_n13576__,
    new_new_n13577__, new_new_n13578__, new_new_n13579__, new_new_n13580__,
    new_new_n13581__, new_new_n13582__, new_new_n13583__, new_new_n13584__,
    new_new_n13585__, new_new_n13586__, new_new_n13587__, new_new_n13588__,
    new_new_n13589__, new_new_n13590__, new_new_n13591__, new_new_n13592__,
    new_new_n13593__, new_new_n13594__, new_new_n13595__, new_new_n13596__,
    new_new_n13597__, new_new_n13598__, new_new_n13599__, new_new_n13600__,
    new_new_n13601__, new_new_n13602__, new_new_n13603__, new_new_n13604__,
    new_new_n13605__, new_new_n13606__, new_new_n13607__, new_new_n13608__,
    new_new_n13609__, new_new_n13610__, new_new_n13611__, new_new_n13612__,
    new_new_n13613__, new_new_n13614__, new_new_n13615__, new_new_n13616__,
    new_new_n13617__, new_new_n13618__, new_new_n13619__, new_new_n13620__,
    new_new_n13621__, new_new_n13622__, new_new_n13623__, new_new_n13624__,
    new_new_n13625__, new_new_n13626__, new_new_n13627__, new_new_n13628__,
    new_new_n13629__, new_new_n13630__, new_new_n13631__, new_new_n13632__,
    new_new_n13633__, new_new_n13634__, new_new_n13635__, new_new_n13636__,
    new_new_n13637__, new_new_n13638__, new_new_n13639__, new_new_n13640__,
    new_new_n13641__, new_new_n13642__, new_new_n13643__, new_new_n13644__,
    new_new_n13645__, new_new_n13646__, new_new_n13647__, new_new_n13648__,
    new_new_n13649__, new_new_n13650__, new_new_n13651__, new_new_n13652__,
    new_new_n13653__, new_new_n13654__, new_new_n13655__, new_new_n13656__,
    new_new_n13657__, new_new_n13658__, new_new_n13659__, new_new_n13660__,
    new_new_n13661__, new_new_n13662__, new_new_n13663__, new_new_n13664__,
    new_new_n13665__, new_new_n13666__, new_new_n13667__, new_new_n13668__,
    new_new_n13669__, new_new_n13670__, new_new_n13671__, new_new_n13672__,
    new_new_n13673__, new_new_n13674__, new_new_n13675__, new_new_n13676__,
    new_new_n13677__, new_new_n13678__, new_new_n13679__, new_new_n13680__,
    new_new_n13681__, new_new_n13682__, new_new_n13683__, new_new_n13684__,
    new_new_n13685__, new_new_n13686__, new_new_n13687__, new_new_n13688__,
    new_new_n13689__, new_new_n13690__, new_new_n13691__, new_new_n13692__,
    new_new_n13693__, new_new_n13694__, new_new_n13695__, new_new_n13696__,
    new_new_n13697__, new_new_n13698__, new_new_n13699__, new_new_n13700__,
    new_new_n13701__, new_new_n13702__, new_new_n13703__, new_new_n13704__,
    new_new_n13705__, new_new_n13706__, new_new_n13707__, new_new_n13708__,
    new_new_n13709__, new_new_n13710__, new_new_n13711__, new_new_n13712__,
    new_new_n13713__, new_new_n13714__, new_new_n13715__, new_new_n13716__,
    new_new_n13717__, new_new_n13718__, new_new_n13719__, new_new_n13720__,
    new_new_n13721__, new_new_n13722__, new_new_n13723__, new_new_n13724__,
    new_new_n13725__, new_new_n13726__, new_new_n13727__, new_new_n13728__,
    new_new_n13729__, new_new_n13730__, new_new_n13731__, new_new_n13732__,
    new_new_n13733__, new_new_n13734__, new_new_n13735__, new_new_n13736__,
    new_new_n13737__, new_new_n13738__, new_new_n13739__, new_new_n13740__,
    new_new_n13741__, new_new_n13742__, new_new_n13743__, new_new_n13744__,
    new_new_n13745__, new_new_n13746__, new_new_n13747__, new_new_n13748__,
    new_new_n13749__, new_new_n13750__, new_new_n13751__, new_new_n13752__,
    new_new_n13753__, new_new_n13754__, new_new_n13755__, new_new_n13756__,
    new_new_n13757__, new_new_n13758__, new_new_n13759__, new_new_n13760__,
    new_new_n13761__, new_new_n13762__, new_new_n13763__, new_new_n13764__,
    new_new_n13765__, new_new_n13766__, new_new_n13767__, new_new_n13768__,
    new_new_n13769__, new_new_n13770__, new_new_n13771__, new_new_n13772__,
    new_new_n13773__, new_new_n13774__, new_new_n13775__, new_new_n13776__,
    new_new_n13777__, new_new_n13778__, new_new_n13779__, new_new_n13780__,
    new_new_n13781__, new_new_n13782__, new_new_n13783__, new_new_n13784__,
    new_new_n13785__, new_new_n13786__, new_new_n13787__, new_new_n13788__,
    new_new_n13789__, new_new_n13790__, new_new_n13791__, new_new_n13792__,
    new_new_n13793__, new_new_n13794__, new_new_n13795__, new_new_n13796__,
    new_new_n13797__, new_new_n13798__, new_new_n13799__, new_new_n13800__,
    new_new_n13801__, new_new_n13802__, new_new_n13803__, new_new_n13804__,
    new_new_n13805__, new_new_n13806__, new_new_n13807__, new_new_n13808__,
    new_new_n13809__, new_new_n13810__, new_new_n13811__, new_new_n13812__,
    new_new_n13813__, new_new_n13814__, new_new_n13815__, new_new_n13816__,
    new_new_n13817__, new_new_n13818__, new_new_n13819__, new_new_n13820__,
    new_new_n13821__, new_new_n13822__, new_new_n13823__, new_new_n13824__,
    new_new_n13825__, new_new_n13826__, new_new_n13827__, new_new_n13828__,
    new_new_n13829__, new_new_n13830__, new_new_n13831__, new_new_n13832__,
    new_new_n13833__, new_new_n13834__, new_new_n13835__, new_new_n13836__,
    new_new_n13837__, new_new_n13838__, new_new_n13839__, new_new_n13840__,
    new_new_n13841__, new_new_n13842__, new_new_n13843__, new_new_n13844__,
    new_new_n13845__, new_new_n13846__, new_new_n13847__, new_new_n13848__,
    new_new_n13849__, new_new_n13850__, new_new_n13851__, new_new_n13852__,
    new_new_n13853__, new_new_n13854__, new_new_n13855__, new_new_n13856__,
    new_new_n13857__, new_new_n13858__, new_new_n13859__, new_new_n13860__,
    new_new_n13861__, new_new_n13862__, new_new_n13863__, new_new_n13864__,
    new_new_n13865__, new_new_n13866__, new_new_n13867__, new_new_n13868__,
    new_new_n13869__, new_new_n13870__, new_new_n13871__, new_new_n13872__,
    new_new_n13873__, new_new_n13874__, new_new_n13875__, new_new_n13876__,
    new_new_n13877__, new_new_n13878__, new_new_n13879__, new_new_n13880__,
    new_new_n13881__, new_new_n13882__, new_new_n13883__, new_new_n13884__,
    new_new_n13885__, new_new_n13886__, new_new_n13887__, new_new_n13888__,
    new_new_n13889__, new_new_n13890__, new_new_n13891__, new_new_n13892__,
    new_new_n13893__, new_new_n13894__, new_new_n13895__, new_new_n13896__,
    new_new_n13897__, new_new_n13898__, new_new_n13899__, new_new_n13900__,
    new_new_n13901__, new_new_n13902__, new_new_n13903__, new_new_n13904__,
    new_new_n13905__, new_new_n13906__, new_new_n13907__, new_new_n13908__,
    new_new_n13909__, new_new_n13910__, new_new_n13911__, new_new_n13912__,
    new_new_n13913__, new_new_n13914__, new_new_n13915__, new_new_n13916__,
    new_new_n13917__, new_new_n13918__, new_new_n13919__, new_new_n13920__,
    new_new_n13921__, new_new_n13922__, new_new_n13923__, new_new_n13924__,
    new_new_n13925__, new_new_n13926__, new_new_n13927__, new_new_n13928__,
    new_new_n13929__, new_new_n13930__, new_new_n13931__, new_new_n13932__,
    new_new_n13933__, new_new_n13934__, new_new_n13935__, new_new_n13936__,
    new_new_n13937__, new_new_n13938__, new_new_n13939__, new_new_n13940__,
    new_new_n13941__, new_new_n13942__, new_new_n13943__, new_new_n13944__,
    new_new_n13945__, new_new_n13946__, new_new_n13947__, new_new_n13948__,
    new_new_n13949__, new_new_n13950__, new_new_n13951__, new_new_n13952__,
    new_new_n13953__, new_new_n13954__, new_new_n13955__, new_new_n13956__,
    new_new_n13957__, new_new_n13958__, new_new_n13959__, new_new_n13960__,
    new_new_n13961__, new_new_n13962__, new_new_n13963__, new_new_n13964__,
    new_new_n13965__, new_new_n13966__, new_new_n13967__, new_new_n13968__,
    new_new_n13969__, new_new_n13970__, new_new_n13971__, new_new_n13972__,
    new_new_n13973__, new_new_n13974__, new_new_n13975__, new_new_n13976__,
    new_new_n13977__, new_new_n13978__, new_new_n13979__, new_new_n13980__,
    new_new_n13981__, new_new_n13982__, new_new_n13983__, new_new_n13984__,
    new_new_n13985__, new_new_n13986__, new_new_n13987__, new_new_n13988__,
    new_new_n13989__, new_new_n13990__, new_new_n13991__, new_new_n13992__,
    new_new_n13993__, new_new_n13994__, new_new_n13995__, new_new_n13996__,
    new_new_n13997__, new_new_n13998__, new_new_n13999__, new_new_n14000__,
    new_new_n14001__, new_new_n14002__, new_new_n14003__, new_new_n14004__,
    new_new_n14005__, new_new_n14006__, new_new_n14007__, new_new_n14008__,
    new_new_n14009__, new_new_n14010__, new_new_n14011__, new_new_n14012__,
    new_new_n14013__, new_new_n14014__, new_new_n14015__, new_new_n14016__,
    new_new_n14017__, new_new_n14018__, new_new_n14019__, new_new_n14020__,
    new_new_n14021__, new_new_n14022__, new_new_n14023__, new_new_n14024__,
    new_new_n14025__, new_new_n14026__, new_new_n14027__, new_new_n14028__,
    new_new_n14029__, new_new_n14030__, new_new_n14031__, new_new_n14032__,
    new_new_n14033__, new_new_n14034__, new_new_n14035__, new_new_n14036__,
    new_new_n14037__, new_new_n14038__, new_new_n14039__, new_new_n14040__,
    new_new_n14041__, new_new_n14042__, new_new_n14043__, new_new_n14044__,
    new_new_n14045__, new_new_n14046__, new_new_n14047__, new_new_n14048__,
    new_new_n14049__, new_new_n14050__, new_new_n14051__, new_new_n14052__,
    new_new_n14053__, new_new_n14054__, new_new_n14055__, new_new_n14056__,
    new_new_n14057__, new_new_n14058__, new_new_n14059__, new_new_n14060__,
    new_new_n14061__, new_new_n14062__, new_new_n14063__, new_new_n14064__,
    new_new_n14065__, new_new_n14066__, new_new_n14067__, new_new_n14068__,
    new_new_n14069__, new_new_n14070__, new_new_n14071__, new_new_n14072__,
    new_new_n14073__, new_new_n14074__, new_new_n14075__, new_new_n14076__,
    new_new_n14077__, new_new_n14078__, new_new_n14079__, new_new_n14080__,
    new_new_n14081__, new_new_n14082__, new_new_n14083__, new_new_n14084__,
    new_new_n14085__, new_new_n14086__, new_new_n14087__, new_new_n14088__,
    new_new_n14089__, new_new_n14090__, new_new_n14091__, new_new_n14092__,
    new_new_n14093__, new_new_n14094__, new_new_n14095__, new_new_n14096__,
    new_new_n14097__, new_new_n14098__, new_new_n14099__, new_new_n14100__,
    new_new_n14101__, new_new_n14102__, new_new_n14103__, new_new_n14104__,
    new_new_n14105__, new_new_n14106__, new_new_n14107__, new_new_n14108__,
    new_new_n14109__, new_new_n14110__, new_new_n14111__, new_new_n14112__,
    new_new_n14113__, new_new_n14114__, new_new_n14115__, new_new_n14116__,
    new_new_n14117__, new_new_n14118__, new_new_n14119__, new_new_n14120__,
    new_new_n14121__, new_new_n14122__, new_new_n14123__, new_new_n14124__,
    new_new_n14125__, new_new_n14126__, new_new_n14127__, new_new_n14128__,
    new_new_n14129__, new_new_n14130__, new_new_n14131__, new_new_n14132__,
    new_new_n14133__, new_new_n14134__, new_new_n14135__, new_new_n14136__,
    new_new_n14137__, new_new_n14138__, new_new_n14139__, new_new_n14140__,
    new_new_n14141__, new_new_n14142__, new_new_n14143__, new_new_n14144__,
    new_new_n14145__, new_new_n14146__, new_new_n14147__, new_new_n14148__,
    new_new_n14149__, new_new_n14150__, new_new_n14151__, new_new_n14152__,
    new_new_n14153__, new_new_n14154__, new_new_n14155__, new_new_n14156__,
    new_new_n14157__, new_new_n14158__, new_new_n14159__, new_new_n14160__,
    new_new_n14161__, new_new_n14162__, new_new_n14163__, new_new_n14164__,
    new_new_n14165__, new_new_n14166__, new_new_n14167__, new_new_n14168__,
    new_new_n14169__, new_new_n14170__, new_new_n14171__, new_new_n14172__,
    new_new_n14173__, new_new_n14174__, new_new_n14175__, new_new_n14176__,
    new_new_n14177__, new_new_n14178__, new_new_n14179__, new_new_n14180__,
    new_new_n14181__, new_new_n14182__, new_new_n14183__, new_new_n14184__,
    new_new_n14185__, new_new_n14186__, new_new_n14187__, new_new_n14188__,
    new_new_n14189__, new_new_n14190__, new_new_n14191__, new_new_n14192__,
    new_new_n14193__, new_new_n14194__, new_new_n14195__, new_new_n14196__,
    new_new_n14197__, new_new_n14198__, new_new_n14199__, new_new_n14200__,
    new_new_n14201__, new_new_n14202__, new_new_n14203__, new_new_n14204__,
    new_new_n14205__, new_new_n14206__, new_new_n14207__, new_new_n14208__,
    new_new_n14209__, new_new_n14210__, new_new_n14211__, new_new_n14212__,
    new_new_n14213__, new_new_n14214__, new_new_n14215__, new_new_n14216__,
    new_new_n14217__, new_new_n14218__, new_new_n14219__, new_new_n14220__,
    new_new_n14221__, new_new_n14222__, new_new_n14223__, new_new_n14224__,
    new_new_n14225__, new_new_n14226__, new_new_n14227__, new_new_n14228__,
    new_new_n14229__, new_new_n14230__, new_new_n14231__, new_new_n14232__,
    new_new_n14233__, new_new_n14234__, new_new_n14235__, new_new_n14236__,
    new_new_n14237__, new_new_n14238__, new_new_n14239__, new_new_n14240__,
    new_new_n14241__, new_new_n14242__, new_new_n14243__, new_new_n14244__,
    new_new_n14245__, new_new_n14246__, new_new_n14247__, new_new_n14248__,
    new_new_n14249__, new_new_n14250__, new_new_n14251__, new_new_n14252__,
    new_new_n14253__, new_new_n14254__, new_new_n14255__, new_new_n14256__,
    new_new_n14257__, new_new_n14258__, new_new_n14259__, new_new_n14260__,
    new_new_n14261__, new_new_n14262__, new_new_n14263__, new_new_n14264__,
    new_new_n14265__, new_new_n14266__, new_new_n14267__, new_new_n14268__,
    new_new_n14269__, new_new_n14270__, new_new_n14271__, new_new_n14272__,
    new_new_n14273__, new_new_n14274__, new_new_n14275__, new_new_n14276__,
    new_new_n14277__, new_new_n14278__, new_new_n14279__, new_new_n14280__,
    new_new_n14281__, new_new_n14282__, new_new_n14283__, new_new_n14284__,
    new_new_n14285__, new_new_n14286__, new_new_n14287__, new_new_n14288__,
    new_new_n14289__, new_new_n14290__, new_new_n14291__, new_new_n14292__,
    new_new_n14293__, new_new_n14294__, new_new_n14295__, new_new_n14296__,
    new_new_n14297__, new_new_n14298__, new_new_n14299__, new_new_n14300__,
    new_new_n14301__, new_new_n14302__, new_new_n14303__, new_new_n14304__,
    new_new_n14305__, new_new_n14306__, new_new_n14307__, new_new_n14308__,
    new_new_n14309__, new_new_n14310__, new_new_n14311__, new_new_n14312__,
    new_new_n14313__, new_new_n14314__, new_new_n14315__, new_new_n14316__,
    new_new_n14317__, new_new_n14318__, new_new_n14319__, new_new_n14320__,
    new_new_n14321__, new_new_n14322__, new_new_n14323__, new_new_n14324__,
    new_new_n14325__, new_new_n14326__, new_new_n14327__, new_new_n14328__,
    new_new_n14329__, new_new_n14330__, new_new_n14331__, new_new_n14332__,
    new_new_n14333__, new_new_n14334__, new_new_n14335__, new_new_n14336__,
    new_new_n14337__, new_new_n14338__, new_new_n14339__, new_new_n14340__,
    new_new_n14341__, new_new_n14342__, new_new_n14343__, new_new_n14344__,
    new_new_n14345__, new_new_n14346__, new_new_n14347__, new_new_n14348__,
    new_new_n14349__, new_new_n14350__, new_new_n14351__, new_new_n14352__,
    new_new_n14353__, new_new_n14354__, new_new_n14355__, new_new_n14356__,
    new_new_n14357__, new_new_n14358__, new_new_n14359__, new_new_n14360__,
    new_new_n14361__, new_new_n14362__, new_new_n14363__, new_new_n14364__,
    new_new_n14365__, new_new_n14366__, new_new_n14367__, new_new_n14368__,
    new_new_n14369__, new_new_n14370__, new_new_n14371__, new_new_n14372__,
    new_new_n14373__, new_new_n14374__, new_new_n14375__, new_new_n14376__,
    new_new_n14377__, new_new_n14378__, new_new_n14379__, new_new_n14380__,
    new_new_n14381__, new_new_n14382__, new_new_n14383__, new_new_n14384__,
    new_new_n14385__, new_new_n14386__, new_new_n14387__, new_new_n14388__,
    new_new_n14389__, new_new_n14390__, new_new_n14391__, new_new_n14392__,
    new_new_n14393__, new_new_n14394__, new_new_n14395__, new_new_n14396__,
    new_new_n14397__, new_new_n14398__, new_new_n14399__, new_new_n14400__,
    new_new_n14401__, new_new_n14402__, new_new_n14403__, new_new_n14404__,
    new_new_n14405__, new_new_n14406__, new_new_n14407__, new_new_n14408__,
    new_new_n14409__, new_new_n14410__, new_new_n14411__, new_new_n14412__,
    new_new_n14413__, new_new_n14414__, new_new_n14415__, new_new_n14416__,
    new_new_n14417__, new_new_n14418__, new_new_n14419__, new_new_n14420__,
    new_new_n14421__, new_new_n14422__, new_new_n14423__, new_new_n14424__,
    new_new_n14425__, new_new_n14426__, new_new_n14427__, new_new_n14428__,
    new_new_n14429__, new_new_n14430__, new_new_n14431__, new_new_n14432__,
    new_new_n14433__, new_new_n14434__, new_new_n14435__, new_new_n14436__,
    new_new_n14437__, new_new_n14438__, new_new_n14439__, new_new_n14440__,
    new_new_n14441__, new_new_n14442__, new_new_n14443__, new_new_n14444__,
    new_new_n14445__, new_new_n14446__, new_new_n14447__, new_new_n14448__,
    new_new_n14449__, new_new_n14450__, new_new_n14451__, new_new_n14452__,
    new_new_n14453__, new_new_n14454__, new_new_n14455__, new_new_n14456__,
    new_new_n14457__, new_new_n14458__, new_new_n14459__, new_new_n14460__,
    new_new_n14461__, new_new_n14462__, new_new_n14463__, new_new_n14464__,
    new_new_n14465__, new_new_n14466__, new_new_n14467__, new_new_n14468__,
    new_new_n14469__, new_new_n14470__, new_new_n14471__, new_new_n14472__,
    new_new_n14473__, new_new_n14474__, new_new_n14475__, new_new_n14476__,
    new_new_n14477__, new_new_n14478__, new_new_n14479__, new_new_n14480__,
    new_new_n14481__, new_new_n14482__, new_new_n14483__, new_new_n14484__,
    new_new_n14485__, new_new_n14486__, new_new_n14487__, new_new_n14488__,
    new_new_n14489__, new_new_n14490__, new_new_n14491__, new_new_n14492__,
    new_new_n14493__, new_new_n14494__, new_new_n14495__, new_new_n14496__,
    new_new_n14497__, new_new_n14498__, new_new_n14499__, new_new_n14500__,
    new_new_n14501__, new_new_n14502__, new_new_n14503__, new_new_n14504__,
    new_new_n14505__, new_new_n14506__, new_new_n14507__, new_new_n14508__,
    new_new_n14509__, new_new_n14510__, new_new_n14511__, new_new_n14512__,
    new_new_n14513__, new_new_n14514__, new_new_n14515__, new_new_n14516__,
    new_new_n14517__, new_new_n14518__, new_new_n14519__, new_new_n14520__,
    new_new_n14521__, new_new_n14522__, new_new_n14523__, new_new_n14524__,
    new_new_n14525__, new_new_n14526__, new_new_n14527__, new_new_n14528__,
    new_new_n14529__, new_new_n14530__, new_new_n14531__, new_new_n14532__,
    new_new_n14533__, new_new_n14534__, new_new_n14535__, new_new_n14536__,
    new_new_n14537__, new_new_n14538__, new_new_n14539__, new_new_n14540__,
    new_new_n14541__, new_new_n14542__, new_new_n14543__, new_new_n14544__,
    new_new_n14545__, new_new_n14546__, new_new_n14547__, new_new_n14548__,
    new_new_n14549__, new_new_n14550__, new_new_n14551__, new_new_n14552__,
    new_new_n14553__, new_new_n14554__, new_new_n14555__, new_new_n14556__,
    new_new_n14557__, new_new_n14558__, new_new_n14559__, new_new_n14560__,
    new_new_n14561__, new_new_n14562__, new_new_n14563__, new_new_n14564__,
    new_new_n14565__, new_new_n14566__, new_new_n14567__, new_new_n14568__,
    new_new_n14569__, new_new_n14570__, new_new_n14571__, new_new_n14572__,
    new_new_n14573__, new_new_n14574__, new_new_n14575__, new_new_n14576__,
    new_new_n14577__, new_new_n14578__, new_new_n14579__, new_new_n14580__,
    new_new_n14581__, new_new_n14582__, new_new_n14583__, new_new_n14584__,
    new_new_n14585__, new_new_n14586__, new_new_n14587__, new_new_n14588__,
    new_new_n14589__, new_new_n14590__, new_new_n14591__, new_new_n14592__,
    new_new_n14593__, new_new_n14594__, new_new_n14595__, new_new_n14596__,
    new_new_n14597__, new_new_n14598__, new_new_n14599__, new_new_n14600__,
    new_new_n14601__, new_new_n14602__, new_new_n14603__, new_new_n14604__,
    new_new_n14605__, new_new_n14606__, new_new_n14607__, new_new_n14608__,
    new_new_n14609__, new_new_n14610__, new_new_n14611__, new_new_n14612__,
    new_new_n14613__, new_new_n14614__, new_new_n14615__, new_new_n14616__,
    new_new_n14617__, new_new_n14618__, new_new_n14619__, new_new_n14620__,
    new_new_n14621__, new_new_n14622__, new_new_n14623__, new_new_n14624__,
    new_new_n14625__, new_new_n14626__, new_new_n14627__, new_new_n14628__,
    new_new_n14629__, new_new_n14630__, new_new_n14631__, new_new_n14632__,
    new_new_n14633__, new_new_n14634__, new_new_n14635__, new_new_n14636__,
    new_new_n14637__, new_new_n14638__, new_new_n14639__, new_new_n14640__,
    new_new_n14641__, new_new_n14642__, new_new_n14643__, new_new_n14644__,
    new_new_n14645__, new_new_n14646__, new_new_n14647__, new_new_n14648__,
    new_new_n14649__, new_new_n14650__, new_new_n14651__, new_new_n14652__,
    new_new_n14653__, new_new_n14654__, new_new_n14655__, new_new_n14656__,
    new_new_n14657__, new_new_n14658__, new_new_n14659__, new_new_n14660__,
    new_new_n14661__, new_new_n14662__, new_new_n14663__, new_new_n14664__,
    new_new_n14665__, new_new_n14666__, new_new_n14667__, new_new_n14668__,
    new_new_n14669__, new_new_n14670__, new_new_n14671__, new_new_n14672__,
    new_new_n14673__, new_new_n14674__, new_new_n14675__, new_new_n14676__,
    new_new_n14677__, new_new_n14678__, new_new_n14679__, new_new_n14680__,
    new_new_n14681__, new_new_n14682__, new_new_n14683__, new_new_n14684__,
    new_new_n14685__, new_new_n14686__, new_new_n14687__, new_new_n14688__,
    new_new_n14689__, new_new_n14690__, new_new_n14691__, new_new_n14692__,
    new_new_n14693__, new_new_n14694__, new_new_n14695__, new_new_n14696__,
    new_new_n14697__, new_new_n14698__, new_new_n14699__, new_new_n14700__,
    new_new_n14701__, new_new_n14702__, new_new_n14703__, new_new_n14704__,
    new_new_n14705__, new_new_n14706__, new_new_n14707__, new_new_n14708__,
    new_new_n14709__, new_new_n14710__, new_new_n14711__, new_new_n14712__,
    new_new_n14713__, new_new_n14714__, new_new_n14715__, new_new_n14716__,
    new_new_n14717__, new_new_n14718__, new_new_n14719__, new_new_n14720__,
    new_new_n14721__, new_new_n14722__, new_new_n14723__, new_new_n14724__,
    new_new_n14725__, new_new_n14726__, new_new_n14727__, new_new_n14728__,
    new_new_n14729__, new_new_n14730__, new_new_n14731__, new_new_n14732__,
    new_new_n14733__, new_new_n14734__, new_new_n14735__, new_new_n14736__,
    new_new_n14737__, new_new_n14738__, new_new_n14739__, new_new_n14740__,
    new_new_n14741__, new_new_n14742__, new_new_n14743__, new_new_n14744__,
    new_new_n14745__, new_new_n14746__, new_new_n14747__, new_new_n14748__,
    new_new_n14749__, new_new_n14750__, new_new_n14751__, new_new_n14752__,
    new_new_n14753__, new_new_n14754__, new_new_n14755__, new_new_n14756__,
    new_new_n14757__, new_new_n14758__, new_new_n14759__, new_new_n14760__,
    new_new_n14761__, new_new_n14762__, new_new_n14763__, new_new_n14764__,
    new_new_n14765__, new_new_n14766__, new_new_n14767__, new_new_n14768__,
    new_new_n14769__, new_new_n14770__, new_new_n14771__, new_new_n14772__,
    new_new_n14773__, new_new_n14774__, new_new_n14775__, new_new_n14776__,
    new_new_n14777__, new_new_n14778__, new_new_n14779__, new_new_n14780__,
    new_new_n14781__, new_new_n14782__, new_new_n14783__, new_new_n14784__,
    new_new_n14785__, new_new_n14786__, new_new_n14787__, new_new_n14788__,
    new_new_n14789__, new_new_n14790__, new_new_n14791__, new_new_n14792__,
    new_new_n14793__, new_new_n14794__, new_new_n14795__, new_new_n14796__,
    new_new_n14797__, new_new_n14798__, new_new_n14799__, new_new_n14800__,
    new_new_n14801__, new_new_n14802__, new_new_n14803__, new_new_n14804__,
    new_new_n14805__, new_new_n14806__, new_new_n14807__, new_new_n14808__,
    new_new_n14809__, new_new_n14810__, new_new_n14811__, new_new_n14812__,
    new_new_n14813__, new_new_n14814__, new_new_n14815__, new_new_n14816__,
    new_new_n14817__, new_new_n14818__, new_new_n14819__, new_new_n14820__,
    new_new_n14821__, new_new_n14822__, new_new_n14823__, new_new_n14824__,
    new_new_n14825__, new_new_n14826__, new_new_n14827__, new_new_n14828__,
    new_new_n14829__, new_new_n14830__, new_new_n14831__, new_new_n14832__,
    new_new_n14833__, new_new_n14834__, new_new_n14835__, new_new_n14836__,
    new_new_n14837__, new_new_n14838__, new_new_n14839__, new_new_n14840__,
    new_new_n14841__, new_new_n14842__, new_new_n14843__, new_new_n14844__,
    new_new_n14845__, new_new_n14846__, new_new_n14847__, new_new_n14848__,
    new_new_n14849__, new_new_n14850__, new_new_n14851__, new_new_n14852__,
    new_new_n14853__, new_new_n14854__, new_new_n14855__, new_new_n14856__,
    new_new_n14857__, new_new_n14858__, new_new_n14859__, new_new_n14860__,
    new_new_n14861__, new_new_n14862__, new_new_n14863__, new_new_n14864__,
    new_new_n14865__, new_new_n14866__, new_new_n14867__, new_new_n14868__,
    new_new_n14869__, new_new_n14870__, new_new_n14871__, new_new_n14872__,
    new_new_n14873__, new_new_n14874__, new_new_n14875__, new_new_n14876__,
    new_new_n14877__, new_new_n14878__, new_new_n14879__, new_new_n14880__,
    new_new_n14881__, new_new_n14882__, new_new_n14883__, new_new_n14884__,
    new_new_n14885__, new_new_n14886__, new_new_n14887__, new_new_n14888__,
    new_new_n14889__, new_new_n14890__, new_new_n14891__, new_new_n14892__,
    new_new_n14893__, new_new_n14894__, new_new_n14895__, new_new_n14896__,
    new_new_n14897__, new_new_n14898__, new_new_n14899__, new_new_n14900__,
    new_new_n14901__, new_new_n14902__, new_new_n14903__, new_new_n14904__,
    new_new_n14905__, new_new_n14906__, new_new_n14907__, new_new_n14908__,
    new_new_n14909__, new_new_n14910__, new_new_n14911__, new_new_n14912__,
    new_new_n14913__, new_new_n14914__, new_new_n14915__, new_new_n14916__,
    new_new_n14917__, new_new_n14918__, new_new_n14919__, new_new_n14920__,
    new_new_n14921__, new_new_n14922__, new_new_n14923__, new_new_n14924__,
    new_new_n14925__, new_new_n14926__, new_new_n14927__, new_new_n14928__,
    new_new_n14929__, new_new_n14930__, new_new_n14931__, new_new_n14932__,
    new_new_n14933__, new_new_n14934__, new_new_n14935__, new_new_n14936__,
    new_new_n14937__, new_new_n14938__, new_new_n14939__, new_new_n14940__,
    new_new_n14941__, new_new_n14942__, new_new_n14943__, new_new_n14944__,
    new_new_n14945__, new_new_n14946__, new_new_n14947__, new_new_n14948__,
    new_new_n14949__, new_new_n14950__, new_new_n14951__, new_new_n14952__,
    new_new_n14953__, new_new_n14954__, new_new_n14955__, new_new_n14956__,
    new_new_n14957__, new_new_n14958__, new_new_n14959__, new_new_n14960__,
    new_new_n14961__, new_new_n14962__, new_new_n14963__, new_new_n14964__,
    new_new_n14965__, new_new_n14966__, new_new_n14967__, new_new_n14968__,
    new_new_n14969__, new_new_n14970__, new_new_n14971__, new_new_n14972__,
    new_new_n14973__, new_new_n14974__, new_new_n14975__, new_new_n14976__,
    new_new_n14977__, new_new_n14978__, new_new_n14979__, new_new_n14980__,
    new_new_n14981__, new_new_n14982__, new_new_n14983__, new_new_n14984__,
    new_new_n14985__, new_new_n14986__, new_new_n14987__, new_new_n14988__,
    new_new_n14989__, new_new_n14990__, new_new_n14991__, new_new_n14992__,
    new_new_n14993__, new_new_n14994__, new_new_n14995__, new_new_n14996__,
    new_new_n14997__, new_new_n14998__, new_new_n14999__, new_new_n15000__,
    new_new_n15001__, new_new_n15002__, new_new_n15003__, new_new_n15004__,
    new_new_n15005__, new_new_n15006__, new_new_n15007__, new_new_n15008__,
    new_new_n15009__, new_new_n15010__, new_new_n15011__, new_new_n15012__,
    new_new_n15013__, new_new_n15014__, new_new_n15015__, new_new_n15016__,
    new_new_n15017__, new_new_n15018__, new_new_n15019__, new_new_n15020__,
    new_new_n15021__, new_new_n15022__, new_new_n15023__, new_new_n15024__,
    new_new_n15025__, new_new_n15026__, new_new_n15027__, new_new_n15028__,
    new_new_n15029__, new_new_n15030__, new_new_n15031__, new_new_n15032__,
    new_new_n15033__, new_new_n15034__, new_new_n15035__, new_new_n15036__,
    new_new_n15037__, new_new_n15038__, new_new_n15039__, new_new_n15040__,
    new_new_n15041__, new_new_n15042__, new_new_n15043__, new_new_n15044__,
    new_new_n15045__, new_new_n15046__, new_new_n15047__, new_new_n15048__,
    new_new_n15049__, new_new_n15050__, new_new_n15051__, new_new_n15052__,
    new_new_n15053__, new_new_n15054__, new_new_n15055__, new_new_n15056__,
    new_new_n15057__, new_new_n15058__, new_new_n15059__, new_new_n15060__,
    new_new_n15061__, new_new_n15062__, new_new_n15063__, new_new_n15064__,
    new_new_n15065__, new_new_n15066__, new_new_n15067__, new_new_n15068__,
    new_new_n15069__, new_new_n15070__, new_new_n15071__, new_new_n15072__,
    new_new_n15073__, new_new_n15074__, new_new_n15075__, new_new_n15076__,
    new_new_n15077__, new_new_n15078__, new_new_n15079__, new_new_n15080__,
    new_new_n15081__, new_new_n15082__, new_new_n15083__, new_new_n15084__,
    new_new_n15085__, new_new_n15086__, new_new_n15087__, new_new_n15088__,
    new_new_n15089__, new_new_n15090__, new_new_n15091__, new_new_n15092__,
    new_new_n15093__, new_new_n15094__, new_new_n15095__, new_new_n15096__,
    new_new_n15097__, new_new_n15098__, new_new_n15099__, new_new_n15100__,
    new_new_n15101__, new_new_n15102__, new_new_n15103__, new_new_n15104__,
    new_new_n15105__, new_new_n15106__, new_new_n15107__, new_new_n15108__,
    new_new_n15109__, new_new_n15110__, new_new_n15111__, new_new_n15112__,
    new_new_n15113__, new_new_n15114__, new_new_n15115__, new_new_n15116__,
    new_new_n15117__, new_new_n15118__, new_new_n15119__, new_new_n15120__,
    new_new_n15121__, new_new_n15122__, new_new_n15123__, new_new_n15124__,
    new_new_n15125__, new_new_n15126__, new_new_n15127__, new_new_n15128__,
    new_new_n15129__, new_new_n15130__, new_new_n15131__, new_new_n15132__,
    new_new_n15133__, new_new_n15134__, new_new_n15135__, new_new_n15136__,
    new_new_n15137__, new_new_n15138__, new_new_n15139__, new_new_n15140__,
    new_new_n15141__, new_new_n15142__, new_new_n15143__, new_new_n15144__,
    new_new_n15145__, new_new_n15146__, new_new_n15147__, new_new_n15148__,
    new_new_n15149__, new_new_n15150__, new_new_n15151__, new_new_n15152__,
    new_new_n15153__, new_new_n15154__, new_new_n15155__, new_new_n15156__,
    new_new_n15157__, new_new_n15158__, new_new_n15159__, new_new_n15160__,
    new_new_n15161__, new_new_n15162__, new_new_n15163__, new_new_n15164__,
    new_new_n15165__, new_new_n15166__, new_new_n15167__, new_new_n15168__,
    new_new_n15169__, new_new_n15170__, new_new_n15171__, new_new_n15172__,
    new_new_n15173__, new_new_n15174__, new_new_n15175__, new_new_n15176__,
    new_new_n15177__, new_new_n15178__, new_new_n15179__, new_new_n15180__,
    new_new_n15181__, new_new_n15182__, new_new_n15183__, new_new_n15184__,
    new_new_n15185__, new_new_n15186__, new_new_n15187__, new_new_n15188__,
    new_new_n15189__, new_new_n15190__, new_new_n15191__, new_new_n15192__,
    new_new_n15193__, new_new_n15194__, new_new_n15195__, new_new_n15196__,
    new_new_n15197__, new_new_n15198__, new_new_n15199__, new_new_n15200__,
    new_new_n15201__, new_new_n15202__, new_new_n15203__, new_new_n15204__,
    new_new_n15205__, new_new_n15206__, new_new_n15207__, new_new_n15208__,
    new_new_n15209__, new_new_n15210__, new_new_n15211__, new_new_n15212__,
    new_new_n15213__, new_new_n15214__, new_new_n15215__, new_new_n15216__,
    new_new_n15217__, new_new_n15218__, new_new_n15219__, new_new_n15220__,
    new_new_n15221__, new_new_n15222__, new_new_n15223__, new_new_n15224__,
    new_new_n15225__, new_new_n15226__, new_new_n15227__, new_new_n15228__,
    new_new_n15229__, new_new_n15230__, new_new_n15231__, new_new_n15232__,
    new_new_n15233__, new_new_n15234__, new_new_n15235__, new_new_n15236__,
    new_new_n15237__, new_new_n15238__, new_new_n15239__, new_new_n15240__,
    new_new_n15241__, new_new_n15242__, new_new_n15243__, new_new_n15244__,
    new_new_n15245__, new_new_n15246__, new_new_n15247__, new_new_n15248__,
    new_new_n15249__, new_new_n15250__, new_new_n15251__, new_new_n15252__,
    new_new_n15253__, new_new_n15254__, new_new_n15255__, new_new_n15256__,
    new_new_n15257__, new_new_n15258__, new_new_n15259__, new_new_n15260__,
    new_new_n15261__, new_new_n15262__, new_new_n15263__, new_new_n15264__,
    new_new_n15265__, new_new_n15266__, new_new_n15267__, new_new_n15268__,
    new_new_n15269__, new_new_n15270__, new_new_n15271__, new_new_n15272__,
    new_new_n15273__, new_new_n15274__, new_new_n15275__, new_new_n15276__,
    new_new_n15277__, new_new_n15278__, new_new_n15279__, new_new_n15280__,
    new_new_n15281__, new_new_n15282__, new_new_n15283__, new_new_n15284__,
    new_new_n15285__, new_new_n15286__, new_new_n15287__, new_new_n15288__,
    new_new_n15289__, new_new_n15290__, new_new_n15291__, new_new_n15292__,
    new_new_n15293__, new_new_n15294__, new_new_n15295__, new_new_n15296__,
    new_new_n15297__, new_new_n15298__, new_new_n15299__, new_new_n15300__,
    new_new_n15301__, new_new_n15302__, new_new_n15303__, new_new_n15304__,
    new_new_n15305__, new_new_n15306__, new_new_n15307__, new_new_n15308__,
    new_new_n15309__, new_new_n15310__, new_new_n15311__, new_new_n15312__,
    new_new_n15313__, new_new_n15314__, new_new_n15315__, new_new_n15316__,
    new_new_n15317__, new_new_n15318__, new_new_n15319__, new_new_n15320__,
    new_new_n15321__, new_new_n15322__, new_new_n15323__, new_new_n15324__,
    new_new_n15325__, new_new_n15326__, new_new_n15327__, new_new_n15328__,
    new_new_n15329__, new_new_n15330__, new_new_n15331__, new_new_n15332__,
    new_new_n15333__, new_new_n15334__, new_new_n15335__, new_new_n15336__,
    new_new_n15337__, new_new_n15338__, new_new_n15339__, new_new_n15340__,
    new_new_n15341__, new_new_n15342__, new_new_n15343__, new_new_n15344__,
    new_new_n15345__, new_new_n15346__, new_new_n15347__, new_new_n15348__,
    new_new_n15349__, new_new_n15350__, new_new_n15351__, new_new_n15352__,
    new_new_n15353__, new_new_n15354__, new_new_n15355__, new_new_n15356__,
    new_new_n15357__, new_new_n15358__, new_new_n15359__, new_new_n15360__,
    new_new_n15361__, new_new_n15362__, new_new_n15363__, new_new_n15364__,
    new_new_n15365__, new_new_n15366__, new_new_n15367__, new_new_n15368__,
    new_new_n15369__, new_new_n15370__, new_new_n15371__, new_new_n15372__,
    new_new_n15373__, new_new_n15374__, new_new_n15375__, new_new_n15376__,
    new_new_n15377__, new_new_n15378__, new_new_n15379__, new_new_n15380__,
    new_new_n15381__, new_new_n15382__, new_new_n15383__, new_new_n15384__,
    new_new_n15385__, new_new_n15386__, new_new_n15387__, new_new_n15388__,
    new_new_n15389__, new_new_n15390__, new_new_n15391__, new_new_n15392__,
    new_new_n15393__, new_new_n15394__, new_new_n15395__, new_new_n15396__,
    new_new_n15397__, new_new_n15398__, new_new_n15399__, new_new_n15400__,
    new_new_n15401__, new_new_n15402__, new_new_n15403__, new_new_n15404__,
    new_new_n15405__, new_new_n15406__, new_new_n15407__, new_new_n15408__,
    new_new_n15409__, new_new_n15410__, new_new_n15411__, new_new_n15412__,
    new_new_n15413__, new_new_n15414__, new_new_n15415__, new_new_n15416__,
    new_new_n15417__, new_new_n15418__, new_new_n15419__, new_new_n15420__,
    new_new_n15421__, new_new_n15422__, new_new_n15423__, new_new_n15424__,
    new_new_n15425__, new_new_n15426__, new_new_n15427__, new_new_n15428__,
    new_new_n15429__, new_new_n15430__, new_new_n15431__, new_new_n15432__,
    new_new_n15433__, new_new_n15434__, new_new_n15435__, new_new_n15436__,
    new_new_n15437__, new_new_n15438__, new_new_n15439__, new_new_n15440__,
    new_new_n15441__, new_new_n15442__, new_new_n15443__, new_new_n15444__,
    new_new_n15445__, new_new_n15446__, new_new_n15447__, new_new_n15448__,
    new_new_n15449__, new_new_n15450__, new_new_n15451__, new_new_n15452__,
    new_new_n15453__, new_new_n15454__, new_new_n15455__, new_new_n15456__,
    new_new_n15457__, new_new_n15458__, new_new_n15459__, new_new_n15460__,
    new_new_n15461__, new_new_n15462__, new_new_n15463__, new_new_n15464__,
    new_new_n15465__, new_new_n15466__, new_new_n15467__, new_new_n15468__,
    new_new_n15469__, new_new_n15470__, new_new_n15471__, new_new_n15472__,
    new_new_n15473__, new_new_n15474__, new_new_n15475__, new_new_n15476__,
    new_new_n15477__, new_new_n15478__, new_new_n15479__, new_new_n15480__,
    new_new_n15481__, new_new_n15482__, new_new_n15483__, new_new_n15484__,
    new_new_n15485__, new_new_n15486__, new_new_n15487__, new_new_n15488__,
    new_new_n15489__, new_new_n15490__, new_new_n15491__, new_new_n15492__,
    new_new_n15493__, new_new_n15494__, new_new_n15495__, new_new_n15496__,
    new_new_n15497__, new_new_n15498__, new_new_n15499__, new_new_n15500__,
    new_new_n15501__, new_new_n15502__, new_new_n15503__, new_new_n15504__,
    new_new_n15505__, new_new_n15506__, new_new_n15507__, new_new_n15508__,
    new_new_n15509__, new_new_n15510__, new_new_n15511__, new_new_n15512__,
    new_new_n15513__, new_new_n15514__, new_new_n15515__, new_new_n15516__,
    new_new_n15517__, new_new_n15518__, new_new_n15519__, new_new_n15520__,
    new_new_n15521__, new_new_n15522__, new_new_n15523__, new_new_n15524__,
    new_new_n15525__, new_new_n15526__, new_new_n15527__, new_new_n15528__,
    new_new_n15529__, new_new_n15530__, new_new_n15531__, new_new_n15532__,
    new_new_n15533__, new_new_n15534__, new_new_n15535__, new_new_n15536__,
    new_new_n15537__, new_new_n15538__, new_new_n15539__, new_new_n15540__,
    new_new_n15541__, new_new_n15542__, new_new_n15543__, new_new_n15544__,
    new_new_n15545__, new_new_n15546__, new_new_n15547__, new_new_n15548__,
    new_new_n15549__, new_new_n15550__, new_new_n15551__, new_new_n15552__,
    new_new_n15553__, new_new_n15554__, new_new_n15555__, new_new_n15556__,
    new_new_n15557__, new_new_n15558__, new_new_n15559__, new_new_n15560__,
    new_new_n15561__, new_new_n15562__, new_new_n15563__, new_new_n15564__,
    new_new_n15565__, new_new_n15566__, new_new_n15567__, new_new_n15568__,
    new_new_n15569__, new_new_n15570__, new_new_n15571__, new_new_n15572__,
    new_new_n15573__, new_new_n15574__, new_new_n15575__, new_new_n15576__,
    new_new_n15577__, new_new_n15578__, new_new_n15579__, new_new_n15580__,
    new_new_n15581__, new_new_n15582__, new_new_n15583__, new_new_n15584__,
    new_new_n15585__, new_new_n15586__, new_new_n15587__, new_new_n15588__,
    new_new_n15589__, new_new_n15590__, new_new_n15591__, new_new_n15592__,
    new_new_n15593__, new_new_n15594__, new_new_n15595__, new_new_n15596__,
    new_new_n15597__, new_new_n15598__, new_new_n15599__, new_new_n15600__,
    new_new_n15601__, new_new_n15602__, new_new_n15603__, new_new_n15604__,
    new_new_n15605__, new_new_n15606__, new_new_n15607__, new_new_n15608__,
    new_new_n15609__, new_new_n15610__, new_new_n15611__, new_new_n15612__,
    new_new_n15613__, new_new_n15614__, new_new_n15615__, new_new_n15616__,
    new_new_n15617__, new_new_n15618__, new_new_n15619__, new_new_n15620__,
    new_new_n15621__, new_new_n15622__, new_new_n15623__, new_new_n15624__,
    new_new_n15625__, new_new_n15626__, new_new_n15627__, new_new_n15628__,
    new_new_n15629__, new_new_n15630__, new_new_n15631__, new_new_n15632__,
    new_new_n15633__, new_new_n15634__, new_new_n15635__, new_new_n15636__,
    new_new_n15637__, new_new_n15638__, new_new_n15639__, new_new_n15640__,
    new_new_n15641__, new_new_n15642__, new_new_n15643__, new_new_n15644__,
    new_new_n15645__, new_new_n15646__, new_new_n15647__, new_new_n15648__,
    new_new_n15649__, new_new_n15650__, new_new_n15651__, new_new_n15652__,
    new_new_n15653__, new_new_n15654__, new_new_n15655__, new_new_n15656__,
    new_new_n15657__, new_new_n15658__, new_new_n15659__, new_new_n15660__,
    new_new_n15661__, new_new_n15662__, new_new_n15663__, new_new_n15664__,
    new_new_n15665__, new_new_n15666__, new_new_n15667__, new_new_n15668__,
    new_new_n15669__, new_new_n15670__, new_new_n15671__, new_new_n15672__,
    new_new_n15673__, new_new_n15674__, new_new_n15675__, new_new_n15676__,
    new_new_n15677__, new_new_n15678__, new_new_n15679__, new_new_n15680__,
    new_new_n15681__, new_new_n15682__, new_new_n15683__, new_new_n15684__,
    new_new_n15685__, new_new_n15686__, new_new_n15687__, new_new_n15688__,
    new_new_n15689__, new_new_n15690__, new_new_n15691__, new_new_n15692__,
    new_new_n15693__, new_new_n15694__, new_new_n15695__, new_new_n15696__,
    new_new_n15697__, new_new_n15698__, new_new_n15699__, new_new_n15700__,
    new_new_n15701__, new_new_n15702__, new_new_n15703__, new_new_n15704__,
    new_new_n15705__, new_new_n15706__, new_new_n15707__, new_new_n15708__,
    new_new_n15709__, new_new_n15710__, new_new_n15711__, new_new_n15712__,
    new_new_n15713__, new_new_n15714__, new_new_n15715__, new_new_n15716__,
    new_new_n15717__, new_new_n15718__, new_new_n15719__, new_new_n15720__,
    new_new_n15721__, new_new_n15722__, new_new_n15723__, new_new_n15724__,
    new_new_n15725__, new_new_n15726__, new_new_n15727__, new_new_n15728__,
    new_new_n15729__, new_new_n15730__, new_new_n15731__, new_new_n15732__,
    new_new_n15733__, new_new_n15734__, new_new_n15735__, new_new_n15736__,
    new_new_n15737__, new_new_n15738__, new_new_n15739__, new_new_n15740__,
    new_new_n15741__, new_new_n15742__, new_new_n15743__, new_new_n15744__,
    new_new_n15745__, new_new_n15746__, new_new_n15747__, new_new_n15748__,
    new_new_n15749__, new_new_n15750__, new_new_n15751__, new_new_n15752__,
    new_new_n15753__, new_new_n15754__, new_new_n15755__, new_new_n15756__,
    new_new_n15757__, new_new_n15758__, new_new_n15759__, new_new_n15760__,
    new_new_n15761__, new_new_n15762__, new_new_n15763__, new_new_n15764__,
    new_new_n15765__, new_new_n15766__, new_new_n15767__, new_new_n15768__,
    new_new_n15769__, new_new_n15770__, new_new_n15771__, new_new_n15772__,
    new_new_n15773__, new_new_n15774__, new_new_n15775__, new_new_n15776__,
    new_new_n15777__, new_new_n15778__, new_new_n15779__, new_new_n15780__,
    new_new_n15781__, new_new_n15782__, new_new_n15783__, new_new_n15784__,
    new_new_n15785__, new_new_n15786__, new_new_n15787__, new_new_n15788__,
    new_new_n15789__, new_new_n15790__, new_new_n15791__, new_new_n15792__,
    new_new_n15793__, new_new_n15794__, new_new_n15795__, new_new_n15796__,
    new_new_n15797__, new_new_n15798__, new_new_n15799__, new_new_n15800__,
    new_new_n15801__, new_new_n15802__, new_new_n15803__, new_new_n15804__,
    new_new_n15805__, new_new_n15806__, new_new_n15807__, new_new_n15808__,
    new_new_n15809__, new_new_n15810__, new_new_n15811__, new_new_n15812__,
    new_new_n15813__, new_new_n15814__, new_new_n15815__, new_new_n15816__,
    new_new_n15817__, new_new_n15818__, new_new_n15819__, new_new_n15820__,
    new_new_n15821__, new_new_n15822__, new_new_n15823__, new_new_n15824__,
    new_new_n15825__, new_new_n15826__, new_new_n15827__, new_new_n15828__,
    new_new_n15829__, new_new_n15830__, new_new_n15831__, new_new_n15832__,
    new_new_n15833__, new_new_n15834__, new_new_n15835__, new_new_n15836__,
    new_new_n15837__, new_new_n15838__, new_new_n15839__, new_new_n15840__,
    new_new_n15841__, new_new_n15842__, new_new_n15843__, new_new_n15844__,
    new_new_n15845__, new_new_n15846__, new_new_n15847__, new_new_n15848__,
    new_new_n15849__, new_new_n15850__, new_new_n15851__, new_new_n15852__,
    new_new_n15853__, new_new_n15854__, new_new_n15855__, new_new_n15856__,
    new_new_n15857__, new_new_n15858__, new_new_n15859__, new_new_n15860__,
    new_new_n15861__, new_new_n15862__, new_new_n15863__, new_new_n15864__,
    new_new_n15865__, new_new_n15866__, new_new_n15867__, new_new_n15868__,
    new_new_n15869__, new_new_n15870__, new_new_n15871__, new_new_n15872__,
    new_new_n15873__, new_new_n15874__, new_new_n15875__, new_new_n15876__,
    new_new_n15877__, new_new_n15878__, new_new_n15879__, new_new_n15880__,
    new_new_n15881__, new_new_n15882__, new_new_n15883__, new_new_n15884__,
    new_new_n15885__, new_new_n15886__, new_new_n15887__, new_new_n15888__,
    new_new_n15889__, new_new_n15890__, new_new_n15891__, new_new_n15892__,
    new_new_n15893__, new_new_n15894__, new_new_n15895__, new_new_n15896__,
    new_new_n15897__, new_new_n15898__, new_new_n15899__, new_new_n15900__,
    new_new_n15901__, new_new_n15902__, new_new_n15903__, new_new_n15904__,
    new_new_n15905__, new_new_n15906__, new_new_n15907__, new_new_n15908__,
    new_new_n15909__, new_new_n15910__, new_new_n15911__, new_new_n15912__,
    new_new_n15913__, new_new_n15914__, new_new_n15915__, new_new_n15916__,
    new_new_n15917__, new_new_n15918__, new_new_n15919__, new_new_n15920__,
    new_new_n15921__, new_new_n15922__, new_new_n15923__, new_new_n15924__,
    new_new_n15925__, new_new_n15926__, new_new_n15927__, new_new_n15928__,
    new_new_n15929__, new_new_n15930__, new_new_n15931__, new_new_n15932__,
    new_new_n15933__, new_new_n15934__, new_new_n15935__, new_new_n15936__,
    new_new_n15937__, new_new_n15938__, new_new_n15939__, new_new_n15940__,
    new_new_n15941__, new_new_n15942__, new_new_n15943__, new_new_n15944__,
    new_new_n15945__, new_new_n15946__, new_new_n15947__, new_new_n15948__,
    new_new_n15949__, new_new_n15950__, new_new_n15951__, new_new_n15952__,
    new_new_n15953__, new_new_n15954__, new_new_n15955__, new_new_n15956__,
    new_new_n15957__, new_new_n15958__, new_new_n15959__, new_new_n15960__,
    new_new_n15961__, new_new_n15962__, new_new_n15963__, new_new_n15964__,
    new_new_n15965__, new_new_n15966__, new_new_n15967__, new_new_n15968__,
    new_new_n15969__, new_new_n15970__, new_new_n15971__, new_new_n15972__,
    new_new_n15973__, new_new_n15974__, new_new_n15975__, new_new_n15976__,
    new_new_n15977__, new_new_n15978__, new_new_n15979__, new_new_n15980__,
    new_new_n15981__, new_new_n15982__, new_new_n15983__, new_new_n15984__,
    new_new_n15985__, new_new_n15986__, new_new_n15987__, new_new_n15988__,
    new_new_n15989__, new_new_n15990__, new_new_n15991__, new_new_n15992__,
    new_new_n15993__, new_new_n15994__, new_new_n15995__, new_new_n15996__,
    new_new_n15997__, new_new_n15998__, new_new_n15999__, new_new_n16000__,
    new_new_n16001__, new_new_n16002__, new_new_n16003__, new_new_n16004__,
    new_new_n16005__, new_new_n16006__, new_new_n16007__, new_new_n16008__,
    new_new_n16009__, new_new_n16010__, new_new_n16011__, new_new_n16012__,
    new_new_n16013__, new_new_n16014__, new_new_n16015__, new_new_n16016__,
    new_new_n16017__, new_new_n16018__, new_new_n16019__, new_new_n16020__,
    new_new_n16021__, new_new_n16022__, new_new_n16023__, new_new_n16024__,
    new_new_n16025__, new_new_n16026__, new_new_n16027__, new_new_n16028__,
    new_new_n16029__, new_new_n16030__, new_new_n16031__, new_new_n16032__,
    new_new_n16033__, new_new_n16034__, new_new_n16035__, new_new_n16036__,
    new_new_n16037__, new_new_n16038__, new_new_n16039__, new_new_n16040__,
    new_new_n16041__, new_new_n16042__, new_new_n16043__, new_new_n16044__,
    new_new_n16045__, new_new_n16046__, new_new_n16047__, new_new_n16048__,
    new_new_n16049__, new_new_n16050__, new_new_n16051__, new_new_n16052__,
    new_new_n16053__, new_new_n16054__, new_new_n16055__, new_new_n16056__,
    new_new_n16057__, new_new_n16058__, new_new_n16059__, new_new_n16060__,
    new_new_n16061__, new_new_n16062__, new_new_n16063__, new_new_n16064__,
    new_new_n16065__, new_new_n16066__, new_new_n16067__, new_new_n16068__,
    new_new_n16069__, new_new_n16070__, new_new_n16071__, new_new_n16072__,
    new_new_n16073__, new_new_n16074__, new_new_n16075__, new_new_n16076__,
    new_new_n16077__, new_new_n16078__, new_new_n16079__, new_new_n16080__,
    new_new_n16081__, new_new_n16082__, new_new_n16083__, new_new_n16084__,
    new_new_n16085__, new_new_n16086__, new_new_n16087__, new_new_n16088__,
    new_new_n16089__, new_new_n16090__, new_new_n16091__, new_new_n16092__,
    new_new_n16093__, new_new_n16094__, new_new_n16095__, new_new_n16096__,
    new_new_n16097__, new_new_n16098__, new_new_n16099__, new_new_n16100__,
    new_new_n16101__, new_new_n16102__, new_new_n16103__, new_new_n16104__,
    new_new_n16105__, new_new_n16106__, new_new_n16107__, new_new_n16108__,
    new_new_n16109__, new_new_n16110__, new_new_n16111__, new_new_n16112__,
    new_new_n16113__, new_new_n16114__, new_new_n16115__, new_new_n16116__,
    new_new_n16117__, new_new_n16118__, new_new_n16119__, new_new_n16120__,
    new_new_n16121__, new_new_n16122__, new_new_n16123__, new_new_n16124__,
    new_new_n16125__, new_new_n16126__, new_new_n16127__, new_new_n16128__,
    new_new_n16129__, new_new_n16130__, new_new_n16131__, new_new_n16132__,
    new_new_n16133__, new_new_n16134__, new_new_n16135__, new_new_n16136__,
    new_new_n16137__, new_new_n16138__, new_new_n16139__, new_new_n16140__,
    new_new_n16141__, new_new_n16142__, new_new_n16143__, new_new_n16144__,
    new_new_n16145__, new_new_n16146__, new_new_n16147__, new_new_n16148__,
    new_new_n16149__, new_new_n16150__, new_new_n16151__, new_new_n16152__,
    new_new_n16153__, new_new_n16154__, new_new_n16155__, new_new_n16156__,
    new_new_n16157__, new_new_n16158__, new_new_n16159__, new_new_n16160__,
    new_new_n16161__, new_new_n16162__, new_new_n16163__, new_new_n16164__,
    new_new_n16165__, new_new_n16166__, new_new_n16167__, new_new_n16168__,
    new_new_n16169__, new_new_n16170__, new_new_n16171__, new_new_n16172__,
    new_new_n16173__, new_new_n16174__, new_new_n16175__, new_new_n16176__,
    new_new_n16177__, new_new_n16178__, new_new_n16179__, new_new_n16180__,
    new_new_n16181__, new_new_n16182__, new_new_n16183__, new_new_n16184__,
    new_new_n16185__, new_new_n16186__, new_new_n16187__, new_new_n16188__,
    new_new_n16189__, new_new_n16190__, new_new_n16191__, new_new_n16192__,
    new_new_n16193__, new_new_n16194__, new_new_n16195__, new_new_n16196__,
    new_new_n16197__, new_new_n16198__, new_new_n16199__, new_new_n16200__,
    new_new_n16201__, new_new_n16202__, new_new_n16203__, new_new_n16204__,
    new_new_n16205__, new_new_n16206__, new_new_n16207__, new_new_n16208__,
    new_new_n16209__, new_new_n16210__, new_new_n16211__, new_new_n16212__,
    new_new_n16213__, new_new_n16214__, new_new_n16215__, new_new_n16216__,
    new_new_n16217__, new_new_n16218__, new_new_n16219__, new_new_n16220__,
    new_new_n16221__, new_new_n16222__, new_new_n16223__, new_new_n16224__,
    new_new_n16225__, new_new_n16226__, new_new_n16227__, new_new_n16228__,
    new_new_n16229__, new_new_n16230__, new_new_n16231__, new_new_n16232__,
    new_new_n16233__, new_new_n16234__, new_new_n16235__, new_new_n16236__,
    new_new_n16237__, new_new_n16238__, new_new_n16239__, new_new_n16240__,
    new_new_n16241__, new_new_n16242__, new_new_n16243__, new_new_n16244__,
    new_new_n16245__, new_new_n16246__, new_new_n16247__, new_new_n16248__,
    new_new_n16249__, new_new_n16250__, new_new_n16251__, new_new_n16252__,
    new_new_n16253__, new_new_n16254__, new_new_n16255__, new_new_n16256__,
    new_new_n16257__, new_new_n16258__, new_new_n16259__, new_new_n16260__,
    new_new_n16261__, new_new_n16262__, new_new_n16263__, new_new_n16264__,
    new_new_n16265__, new_new_n16266__, new_new_n16267__, new_new_n16268__,
    new_new_n16269__, new_new_n16270__, new_new_n16271__, new_new_n16272__,
    new_new_n16273__, new_new_n16274__, new_new_n16275__, new_new_n16276__,
    new_new_n16277__, new_new_n16278__, new_new_n16279__, new_new_n16280__,
    new_new_n16281__, new_new_n16282__, new_new_n16283__, new_new_n16284__,
    new_new_n16285__, new_new_n16286__, new_new_n16287__, new_new_n16288__,
    new_new_n16289__, new_new_n16290__, new_new_n16291__, new_new_n16292__,
    new_new_n16293__, new_new_n16294__, new_new_n16295__, new_new_n16296__,
    new_new_n16297__, new_new_n16298__, new_new_n16299__, new_new_n16300__,
    new_new_n16301__, new_new_n16302__, new_new_n16303__, new_new_n16304__,
    new_new_n16305__, new_new_n16306__, new_new_n16307__, new_new_n16308__,
    new_new_n16309__, new_new_n16310__, new_new_n16311__, new_new_n16312__,
    new_new_n16313__, new_new_n16314__, new_new_n16315__, new_new_n16316__,
    new_new_n16317__, new_new_n16318__, new_new_n16319__, new_new_n16320__,
    new_new_n16321__, new_new_n16322__, new_new_n16323__, new_new_n16324__,
    new_new_n16325__, new_new_n16326__, new_new_n16327__, new_new_n16328__,
    new_new_n16329__, new_new_n16330__, new_new_n16331__, new_new_n16332__,
    new_new_n16333__, new_new_n16334__, new_new_n16335__, new_new_n16336__,
    new_new_n16337__, new_new_n16338__, new_new_n16339__, new_new_n16340__,
    new_new_n16341__, new_new_n16342__, new_new_n16343__, new_new_n16344__,
    new_new_n16345__, new_new_n16346__, new_new_n16347__, new_new_n16348__,
    new_new_n16349__, new_new_n16350__, new_new_n16351__, new_new_n16352__,
    new_new_n16353__, new_new_n16354__, new_new_n16355__, new_new_n16356__,
    new_new_n16357__, new_new_n16358__, new_new_n16359__, new_new_n16360__,
    new_new_n16361__, new_new_n16362__, new_new_n16363__, new_new_n16364__,
    new_new_n16365__, new_new_n16366__, new_new_n16367__, new_new_n16368__,
    new_new_n16369__, new_new_n16370__, new_new_n16371__, new_new_n16372__,
    new_new_n16373__, new_new_n16374__, new_new_n16375__, new_new_n16376__,
    new_new_n16377__, new_new_n16378__, new_new_n16379__, new_new_n16380__,
    new_new_n16381__, new_new_n16382__, new_new_n16383__, new_new_n16384__,
    new_new_n16385__, new_new_n16386__, new_new_n16387__, new_new_n16388__,
    new_new_n16389__, new_new_n16390__, new_new_n16391__, new_new_n16392__,
    new_new_n16393__, new_new_n16394__, new_new_n16395__, new_new_n16396__,
    new_new_n16397__, new_new_n16398__, new_new_n16399__, new_new_n16400__,
    new_new_n16401__, new_new_n16402__, new_new_n16403__, new_new_n16404__,
    new_new_n16405__, new_new_n16406__, new_new_n16407__, new_new_n16408__,
    new_new_n16409__, new_new_n16410__, new_new_n16411__, new_new_n16412__,
    new_new_n16413__, new_new_n16414__, new_new_n16415__, new_new_n16416__,
    new_new_n16417__, new_new_n16418__, new_new_n16419__, new_new_n16420__,
    new_new_n16421__, new_new_n16422__, new_new_n16423__, new_new_n16424__,
    new_new_n16425__, new_new_n16426__, new_new_n16427__, new_new_n16428__,
    new_new_n16429__, new_new_n16430__, new_new_n16431__, new_new_n16432__,
    new_new_n16433__, new_new_n16434__, new_new_n16435__, new_new_n16436__,
    new_new_n16437__, new_new_n16438__, new_new_n16439__, new_new_n16440__,
    new_new_n16441__, new_new_n16442__, new_new_n16443__, new_new_n16444__,
    new_new_n16445__, new_new_n16446__, new_new_n16447__, new_new_n16448__,
    new_new_n16449__, new_new_n16450__, new_new_n16451__, new_new_n16452__,
    new_new_n16453__, new_new_n16454__, new_new_n16455__, new_new_n16456__,
    new_new_n16457__, new_new_n16458__, new_new_n16459__, new_new_n16460__,
    new_new_n16461__, new_new_n16462__, new_new_n16463__, new_new_n16464__,
    new_new_n16465__, new_new_n16466__, new_new_n16467__, new_new_n16468__,
    new_new_n16469__, new_new_n16470__, new_new_n16471__, new_new_n16472__,
    new_new_n16473__, new_new_n16474__, new_new_n16475__, new_new_n16476__,
    new_new_n16477__, new_new_n16478__, new_new_n16479__, new_new_n16480__,
    new_new_n16481__, new_new_n16482__, new_new_n16483__, new_new_n16484__,
    new_new_n16485__, new_new_n16486__, new_new_n16487__, new_new_n16488__,
    new_new_n16489__, new_new_n16490__, new_new_n16491__, new_new_n16492__,
    new_new_n16493__, new_new_n16494__, new_new_n16495__, new_new_n16496__,
    new_new_n16497__, new_new_n16498__, new_new_n16499__, new_new_n16500__,
    new_new_n16501__, new_new_n16502__, new_new_n16503__, new_new_n16504__,
    new_new_n16505__, new_new_n16506__, new_new_n16507__, new_new_n16508__,
    new_new_n16509__, new_new_n16510__, new_new_n16511__, new_new_n16512__,
    new_new_n16513__, new_new_n16514__, new_new_n16515__, new_new_n16516__,
    new_new_n16517__, new_new_n16518__, new_new_n16519__, new_new_n16520__,
    new_new_n16521__, new_new_n16522__, new_new_n16523__, new_new_n16524__,
    new_new_n16525__, new_new_n16526__, new_new_n16527__, new_new_n16528__,
    new_new_n16529__, new_new_n16530__, new_new_n16531__, new_new_n16532__,
    new_new_n16533__, new_new_n16534__, new_new_n16535__, new_new_n16536__,
    new_new_n16537__, new_new_n16538__, new_new_n16539__, new_new_n16540__,
    new_new_n16541__, new_new_n16542__, new_new_n16543__, new_new_n16544__,
    new_new_n16545__, new_new_n16546__, new_new_n16547__, new_new_n16548__,
    new_new_n16549__, new_new_n16550__, new_new_n16551__, new_new_n16552__,
    new_new_n16553__, new_new_n16554__, new_new_n16555__, new_new_n16556__,
    new_new_n16557__, new_new_n16558__, new_new_n16559__, new_new_n16560__,
    new_new_n16561__, new_new_n16562__, new_new_n16563__, new_new_n16564__,
    new_new_n16565__, new_new_n16566__, new_new_n16567__, new_new_n16568__,
    new_new_n16569__, new_new_n16570__, new_new_n16571__, new_new_n16572__,
    new_new_n16573__, new_new_n16574__, new_new_n16575__, new_new_n16576__,
    new_new_n16577__, new_new_n16578__, new_new_n16579__, new_new_n16580__,
    new_new_n16581__, new_new_n16582__, new_new_n16583__, new_new_n16584__,
    new_new_n16585__, new_new_n16586__, new_new_n16587__, new_new_n16588__,
    new_new_n16589__, new_new_n16590__, new_new_n16591__, new_new_n16592__,
    new_new_n16593__, new_new_n16594__, new_new_n16595__, new_new_n16596__,
    new_new_n16597__, new_new_n16598__, new_new_n16599__, new_new_n16600__,
    new_new_n16601__, new_new_n16602__, new_new_n16603__, new_new_n16604__,
    new_new_n16605__, new_new_n16606__, new_new_n16607__, new_new_n16608__,
    new_new_n16609__, new_new_n16610__, new_new_n16611__, new_new_n16612__,
    new_new_n16613__, new_new_n16614__, new_new_n16615__, new_new_n16616__,
    new_new_n16617__, new_new_n16618__, new_new_n16619__, new_new_n16620__,
    new_new_n16621__, new_new_n16622__, new_new_n16623__, new_new_n16624__,
    new_new_n16625__, new_new_n16626__, new_new_n16627__, new_new_n16628__,
    new_new_n16629__, new_new_n16630__, new_new_n16631__, new_new_n16632__,
    new_new_n16633__, new_new_n16634__, new_new_n16635__, new_new_n16636__,
    new_new_n16637__, new_new_n16638__, new_new_n16639__, new_new_n16640__,
    new_new_n16641__, new_new_n16642__, new_new_n16643__, new_new_n16644__,
    new_new_n16645__, new_new_n16646__, new_new_n16647__, new_new_n16648__,
    new_new_n16649__, new_new_n16650__, new_new_n16651__, new_new_n16652__,
    new_new_n16653__, new_new_n16654__, new_new_n16655__, new_new_n16656__,
    new_new_n16657__, new_new_n16658__, new_new_n16659__, new_new_n16660__,
    new_new_n16661__, new_new_n16662__, new_new_n16663__, new_new_n16664__,
    new_new_n16665__, new_new_n16666__, new_new_n16667__, new_new_n16668__,
    new_new_n16669__, new_new_n16670__, new_new_n16671__, new_new_n16672__,
    new_new_n16673__, new_new_n16674__, new_new_n16675__, new_new_n16676__,
    new_new_n16677__, new_new_n16678__, new_new_n16679__, new_new_n16680__,
    new_new_n16681__, new_new_n16682__, new_new_n16683__, new_new_n16684__,
    new_new_n16685__, new_new_n16686__, new_new_n16687__, new_new_n16688__,
    new_new_n16689__, new_new_n16690__, new_new_n16691__, new_new_n16692__,
    new_new_n16693__, new_new_n16694__, new_new_n16695__, new_new_n16696__,
    new_new_n16697__, new_new_n16698__, new_new_n16699__, new_new_n16700__,
    new_new_n16701__, new_new_n16702__, new_new_n16703__, new_new_n16704__,
    new_new_n16705__, new_new_n16706__, new_new_n16707__, new_new_n16708__,
    new_new_n16709__, new_new_n16710__, new_new_n16711__, new_new_n16712__,
    new_new_n16713__, new_new_n16714__, new_new_n16715__, new_new_n16716__,
    new_new_n16717__, new_new_n16718__, new_new_n16719__, new_new_n16720__,
    new_new_n16721__, new_new_n16722__, new_new_n16723__, new_new_n16724__,
    new_new_n16725__, new_new_n16726__, new_new_n16727__, new_new_n16728__,
    new_new_n16729__, new_new_n16730__, new_new_n16731__, new_new_n16732__,
    new_new_n16733__, new_new_n16734__, new_new_n16735__, new_new_n16736__,
    new_new_n16737__, new_new_n16738__, new_new_n16739__, new_new_n16740__,
    new_new_n16741__, new_new_n16742__, new_new_n16743__, new_new_n16744__,
    new_new_n16745__, new_new_n16746__, new_new_n16747__, new_new_n16748__,
    new_new_n16749__, new_new_n16750__, new_new_n16751__, new_new_n16752__,
    new_new_n16753__, new_new_n16754__, new_new_n16755__, new_new_n16756__,
    new_new_n16757__, new_new_n16758__, new_new_n16759__, new_new_n16760__,
    new_new_n16761__, new_new_n16762__, new_new_n16763__, new_new_n16764__,
    new_new_n16765__, new_new_n16766__, new_new_n16767__, new_new_n16768__,
    new_new_n16769__, new_new_n16770__, new_new_n16771__, new_new_n16772__,
    new_new_n16773__, new_new_n16774__, new_new_n16775__, new_new_n16776__,
    new_new_n16777__, new_new_n16778__, new_new_n16779__, new_new_n16780__,
    new_new_n16781__, new_new_n16782__, new_new_n16783__, new_new_n16784__,
    new_new_n16785__, new_new_n16786__, new_new_n16787__, new_new_n16788__,
    new_new_n16789__, new_new_n16790__, new_new_n16791__, new_new_n16792__,
    new_new_n16793__, new_new_n16794__, new_new_n16795__, new_new_n16796__,
    new_new_n16797__, new_new_n16798__, new_new_n16799__, new_new_n16800__,
    new_new_n16801__, new_new_n16802__, new_new_n16803__, new_new_n16804__,
    new_new_n16805__, new_new_n16806__, new_new_n16807__, new_new_n16808__,
    new_new_n16809__, new_new_n16810__, new_new_n16811__, new_new_n16812__,
    new_new_n16813__, new_new_n16814__, new_new_n16815__, new_new_n16816__,
    new_new_n16817__, new_new_n16818__, new_new_n16819__, new_new_n16820__,
    new_new_n16821__, new_new_n16822__, new_new_n16823__, new_new_n16824__,
    new_new_n16825__, new_new_n16826__, new_new_n16827__, new_new_n16828__,
    new_new_n16829__, new_new_n16830__, new_new_n16831__, new_new_n16832__,
    new_new_n16833__, new_new_n16834__, new_new_n16835__, new_new_n16836__,
    new_new_n16837__, new_new_n16838__, new_new_n16839__, new_new_n16840__,
    new_new_n16841__, new_new_n16842__, new_new_n16843__, new_new_n16844__,
    new_new_n16845__, new_new_n16846__, new_new_n16847__, new_new_n16848__,
    new_new_n16849__, new_new_n16850__, new_new_n16851__, new_new_n16852__,
    new_new_n16853__, new_new_n16854__, new_new_n16855__, new_new_n16856__,
    new_new_n16857__, new_new_n16858__, new_new_n16859__, new_new_n16860__,
    new_new_n16861__, new_new_n16862__, new_new_n16863__, new_new_n16864__,
    new_new_n16865__, new_new_n16866__, new_new_n16867__, new_new_n16868__,
    new_new_n16869__, new_new_n16870__, new_new_n16871__, new_new_n16872__,
    new_new_n16873__, new_new_n16874__, new_new_n16875__, new_new_n16876__,
    new_new_n16877__, new_new_n16878__, new_new_n16879__, new_new_n16880__,
    new_new_n16881__, new_new_n16882__, new_new_n16883__, new_new_n16884__,
    new_new_n16885__, new_new_n16886__, new_new_n16887__, new_new_n16888__,
    new_new_n16889__, new_new_n16890__, new_new_n16891__, new_new_n16892__,
    new_new_n16893__, new_new_n16894__, new_new_n16895__, new_new_n16896__,
    new_new_n16897__, new_new_n16898__, new_new_n16899__, new_new_n16900__,
    new_new_n16901__, new_new_n16902__, new_new_n16903__, new_new_n16904__,
    new_new_n16905__, new_new_n16906__, new_new_n16907__, new_new_n16908__,
    new_new_n16909__, new_new_n16910__, new_new_n16911__, new_new_n16912__,
    new_new_n16913__, new_new_n16914__, new_new_n16915__, new_new_n16916__,
    new_new_n16917__, new_new_n16918__, new_new_n16919__, new_new_n16920__,
    new_new_n16921__, new_new_n16922__, new_new_n16923__, new_new_n16924__,
    new_new_n16925__, new_new_n16926__, new_new_n16927__, new_new_n16928__,
    new_new_n16929__, new_new_n16930__, new_new_n16931__, new_new_n16932__,
    new_new_n16933__, new_new_n16934__, new_new_n16935__, new_new_n16936__,
    new_new_n16937__, new_new_n16938__, new_new_n16939__, new_new_n16940__,
    new_new_n16941__, new_new_n16942__, new_new_n16943__, new_new_n16944__,
    new_new_n16945__, new_new_n16946__, new_new_n16947__, new_new_n16948__,
    new_new_n16949__, new_new_n16950__, new_new_n16951__, new_new_n16952__,
    new_new_n16953__, new_new_n16954__, new_new_n16955__, new_new_n16956__,
    new_new_n16957__, new_new_n16958__, new_new_n16959__, new_new_n16960__,
    new_new_n16961__, new_new_n16962__, new_new_n16963__, new_new_n16964__,
    new_new_n16965__, new_new_n16966__, new_new_n16967__, new_new_n16968__,
    new_new_n16969__, new_new_n16970__, new_new_n16971__, new_new_n16972__,
    new_new_n16973__, new_new_n16974__, new_new_n16975__, new_new_n16976__,
    new_new_n16977__, new_new_n16978__, new_new_n16979__, new_new_n16980__,
    new_new_n16981__, new_new_n16982__, new_new_n16983__, new_new_n16984__,
    new_new_n16985__, new_new_n16986__, new_new_n16987__, new_new_n16988__,
    new_new_n16989__, new_new_n16990__, new_new_n16991__, new_new_n16992__,
    new_new_n16993__, new_new_n16994__, new_new_n16995__, new_new_n16996__,
    new_new_n16997__, new_new_n16998__, new_new_n16999__, new_new_n17000__,
    new_new_n17001__, new_new_n17002__, new_new_n17003__, new_new_n17004__,
    new_new_n17005__, new_new_n17006__, new_new_n17007__, new_new_n17008__,
    new_new_n17009__, new_new_n17010__, new_new_n17011__, new_new_n17012__,
    new_new_n17013__, new_new_n17014__, new_new_n17015__, new_new_n17016__,
    new_new_n17017__, new_new_n17018__, new_new_n17019__, new_new_n17020__,
    new_new_n17021__, new_new_n17022__, new_new_n17023__, new_new_n17024__,
    new_new_n17025__, new_new_n17026__, new_new_n17027__, new_new_n17028__,
    new_new_n17029__, new_new_n17030__, new_new_n17031__, new_new_n17032__,
    new_new_n17033__, new_new_n17034__, new_new_n17035__, new_new_n17036__,
    new_new_n17037__, new_new_n17038__, new_new_n17039__, new_new_n17040__,
    new_new_n17041__, new_new_n17042__, new_new_n17043__, new_new_n17044__,
    new_new_n17045__, new_new_n17046__, new_new_n17047__, new_new_n17048__,
    new_new_n17049__, new_new_n17050__, new_new_n17051__, new_new_n17052__,
    new_new_n17053__, new_new_n17054__, new_new_n17055__, new_new_n17056__,
    new_new_n17057__, new_new_n17058__, new_new_n17059__, new_new_n17060__,
    new_new_n17061__, new_new_n17062__, new_new_n17063__, new_new_n17064__,
    new_new_n17065__, new_new_n17066__, new_new_n17067__, new_new_n17068__,
    new_new_n17069__, new_new_n17070__, new_new_n17071__, new_new_n17072__,
    new_new_n17073__, new_new_n17074__, new_new_n17075__, new_new_n17076__,
    new_new_n17077__, new_new_n17078__, new_new_n17079__, new_new_n17080__,
    new_new_n17081__, new_new_n17082__, new_new_n17083__, new_new_n17084__,
    new_new_n17085__, new_new_n17086__, new_new_n17087__, new_new_n17088__,
    new_new_n17089__, new_new_n17090__, new_new_n17091__, new_new_n17092__,
    new_new_n17093__, new_new_n17094__, new_new_n17095__, new_new_n17096__,
    new_new_n17097__, new_new_n17098__, new_new_n17099__, new_new_n17100__,
    new_new_n17101__, new_new_n17102__, new_new_n17103__, new_new_n17104__,
    new_new_n17105__, new_new_n17106__, new_new_n17107__, new_new_n17108__,
    new_new_n17109__, new_new_n17110__, new_new_n17111__, new_new_n17112__,
    new_new_n17113__, new_new_n17114__, new_new_n17115__, new_new_n17116__,
    new_new_n17117__, new_new_n17118__, new_new_n17119__, new_new_n17120__,
    new_new_n17121__, new_new_n17122__, new_new_n17123__, new_new_n17124__,
    new_new_n17125__, new_new_n17126__, new_new_n17127__, new_new_n17128__,
    new_new_n17129__, new_new_n17130__, new_new_n17131__, new_new_n17132__,
    new_new_n17133__, new_new_n17134__, new_new_n17135__, new_new_n17136__,
    new_new_n17137__, new_new_n17138__, new_new_n17139__, new_new_n17140__,
    new_new_n17141__, new_new_n17142__, new_new_n17143__, new_new_n17144__,
    new_new_n17145__, new_new_n17146__, new_new_n17147__, new_new_n17148__,
    new_new_n17149__, new_new_n17150__, new_new_n17151__, new_new_n17152__,
    new_new_n17153__, new_new_n17154__, new_new_n17155__, new_new_n17156__,
    new_new_n17157__, new_new_n17158__, new_new_n17159__, new_new_n17160__,
    new_new_n17161__, new_new_n17162__, new_new_n17163__, new_new_n17164__,
    new_new_n17165__, new_new_n17166__, new_new_n17167__, new_new_n17168__,
    new_new_n17169__, new_new_n17170__, new_new_n17171__, new_new_n17172__,
    new_new_n17173__, new_new_n17174__, new_new_n17175__, new_new_n17176__,
    new_new_n17177__, new_new_n17178__, new_new_n17179__, new_new_n17180__,
    new_new_n17181__, new_new_n17182__, new_new_n17183__, new_new_n17184__,
    new_new_n17185__, new_new_n17186__, new_new_n17187__, new_new_n17188__,
    new_new_n17189__, new_new_n17190__, new_new_n17191__, new_new_n17192__,
    new_new_n17193__, new_new_n17194__, new_new_n17195__, new_new_n17196__,
    new_new_n17197__, new_new_n17198__, new_new_n17199__, new_new_n17200__,
    new_new_n17201__, new_new_n17202__, new_new_n17203__, new_new_n17204__,
    new_new_n17205__, new_new_n17206__, new_new_n17207__, new_new_n17208__,
    new_new_n17209__, new_new_n17210__, new_new_n17211__, new_new_n17212__,
    new_new_n17213__, new_new_n17214__, new_new_n17215__, new_new_n17216__,
    new_new_n17217__, new_new_n17218__, new_new_n17219__, new_new_n17220__,
    new_new_n17221__, new_new_n17222__, new_new_n17223__, new_new_n17224__,
    new_new_n17225__, new_new_n17226__, new_new_n17227__, new_new_n17228__,
    new_new_n17229__, new_new_n17230__, new_new_n17231__, new_new_n17232__,
    new_new_n17233__, new_new_n17234__, new_new_n17235__, new_new_n17236__,
    new_new_n17237__, new_new_n17238__, new_new_n17239__, new_new_n17240__,
    new_new_n17241__, new_new_n17242__, new_new_n17243__, new_new_n17244__,
    new_new_n17245__, new_new_n17246__, new_new_n17247__, new_new_n17248__,
    new_new_n17249__, new_new_n17250__, new_new_n17251__, new_new_n17252__,
    new_new_n17253__, new_new_n17254__, new_new_n17255__, new_new_n17256__,
    new_new_n17257__, new_new_n17258__, new_new_n17259__, new_new_n17260__,
    new_new_n17261__, new_new_n17262__, new_new_n17263__, new_new_n17264__,
    new_new_n17265__, new_new_n17266__, new_new_n17267__, new_new_n17268__,
    new_new_n17269__, new_new_n17270__, new_new_n17271__, new_new_n17272__,
    new_new_n17273__, new_new_n17274__, new_new_n17275__, new_new_n17276__,
    new_new_n17277__, new_new_n17278__, new_new_n17279__, new_new_n17280__,
    new_new_n17281__, new_new_n17282__, new_new_n17283__, new_new_n17284__,
    new_new_n17285__, new_new_n17286__, new_new_n17287__, new_new_n17288__,
    new_new_n17289__, new_new_n17290__, new_new_n17291__, new_new_n17292__,
    new_new_n17293__, new_new_n17294__, new_new_n17295__, new_new_n17296__,
    new_new_n17297__, new_new_n17298__, new_new_n17299__, new_new_n17300__,
    new_new_n17301__, new_new_n17302__, new_new_n17303__, new_new_n17304__,
    new_new_n17305__, new_new_n17306__, new_new_n17307__, new_new_n17308__,
    new_new_n17309__, new_new_n17310__, new_new_n17311__, new_new_n17312__,
    new_new_n17313__, new_new_n17314__, new_new_n17315__, new_new_n17316__,
    new_new_n17317__, new_new_n17318__, new_new_n17319__, new_new_n17320__,
    new_new_n17321__, new_new_n17322__, new_new_n17323__, new_new_n17324__,
    new_new_n17325__, new_new_n17326__, new_new_n17327__, new_new_n17328__,
    new_new_n17329__, new_new_n17330__, new_new_n17331__, new_new_n17332__,
    new_new_n17333__, new_new_n17334__, new_new_n17335__, new_new_n17336__,
    new_new_n17337__, new_new_n17338__, new_new_n17339__, new_new_n17340__,
    new_new_n17341__, new_new_n17342__, new_new_n17343__, new_new_n17344__,
    new_new_n17345__, new_new_n17346__, new_new_n17347__, new_new_n17348__,
    new_new_n17349__, new_new_n17350__, new_new_n17351__, new_new_n17352__,
    new_new_n17353__, new_new_n17354__, new_new_n17355__, new_new_n17356__,
    new_new_n17357__, new_new_n17358__, new_new_n17359__, new_new_n17360__,
    new_new_n17361__, new_new_n17362__, new_new_n17363__, new_new_n17364__,
    new_new_n17365__, new_new_n17366__, new_new_n17367__, new_new_n17368__,
    new_new_n17369__, new_new_n17370__, new_new_n17371__, new_new_n17372__,
    new_new_n17373__, new_new_n17374__, new_new_n17375__, new_new_n17376__,
    new_new_n17377__, new_new_n17378__, new_new_n17379__, new_new_n17380__,
    new_new_n17381__, new_new_n17382__, new_new_n17383__, new_new_n17384__,
    new_new_n17385__, new_new_n17386__, new_new_n17387__, new_new_n17388__,
    new_new_n17389__, new_new_n17390__, new_new_n17391__, new_new_n17392__,
    new_new_n17393__, new_new_n17394__, new_new_n17395__, new_new_n17396__,
    new_new_n17397__, new_new_n17398__, new_new_n17399__, new_new_n17400__,
    new_new_n17401__, new_new_n17402__, new_new_n17403__, new_new_n17404__,
    new_new_n17405__, new_new_n17406__, new_new_n17407__, new_new_n17408__,
    new_new_n17409__, new_new_n17410__, new_new_n17411__, new_new_n17412__,
    new_new_n17413__, new_new_n17414__, new_new_n17415__, new_new_n17416__,
    new_new_n17417__, new_new_n17418__, new_new_n17419__, new_new_n17420__,
    new_new_n17421__, new_new_n17422__, new_new_n17423__, new_new_n17424__,
    new_new_n17425__, new_new_n17426__, new_new_n17427__, new_new_n17428__,
    new_new_n17429__, new_new_n17430__, new_new_n17431__, new_new_n17432__,
    new_new_n17433__, new_new_n17434__, new_new_n17435__, new_new_n17436__,
    new_new_n17437__, new_new_n17438__, new_new_n17439__, new_new_n17440__,
    new_new_n17441__, new_new_n17442__, new_new_n17443__, new_new_n17444__,
    new_new_n17445__, new_new_n17446__, new_new_n17447__, new_new_n17448__,
    new_new_n17449__, new_new_n17450__, new_new_n17451__, new_new_n17452__,
    new_new_n17453__, new_new_n17454__, new_new_n17455__, new_new_n17456__,
    new_new_n17457__, new_new_n17458__, new_new_n17459__, new_new_n17460__,
    new_new_n17461__, new_new_n17462__, new_new_n17463__, new_new_n17464__,
    new_new_n17465__, new_new_n17466__, new_new_n17467__, new_new_n17468__,
    new_new_n17469__, new_new_n17470__, new_new_n17471__, new_new_n17472__,
    new_new_n17473__, new_new_n17474__, new_new_n17475__, new_new_n17476__,
    new_new_n17477__, new_new_n17478__, new_new_n17479__, new_new_n17480__,
    new_new_n17481__, new_new_n17482__, new_new_n17483__, new_new_n17484__,
    new_new_n17485__, new_new_n17486__, new_new_n17487__, new_new_n17488__,
    new_new_n17489__, new_new_n17490__, new_new_n17491__, new_new_n17492__,
    new_new_n17493__, new_new_n17494__, new_new_n17495__, new_new_n17496__,
    new_new_n17497__, new_new_n17498__, new_new_n17499__, new_new_n17500__,
    new_new_n17501__, new_new_n17502__, new_new_n17503__, new_new_n17504__,
    new_new_n17505__, new_new_n17506__, new_new_n17507__, new_new_n17508__,
    new_new_n17509__, new_new_n17510__, new_new_n17511__, new_new_n17512__,
    new_new_n17513__, new_new_n17514__, new_new_n17515__, new_new_n17516__,
    new_new_n17517__, new_new_n17518__, new_new_n17519__, new_new_n17520__,
    new_new_n17521__, new_new_n17522__, new_new_n17523__, new_new_n17524__,
    new_new_n17525__, new_new_n17526__, new_new_n17527__, new_new_n17528__,
    new_new_n17529__, new_new_n17530__, new_new_n17531__, new_new_n17532__,
    new_new_n17533__, new_new_n17534__, new_new_n17535__, new_new_n17536__,
    new_new_n17537__, new_new_n17538__, new_new_n17539__, new_new_n17540__,
    new_new_n17541__, new_new_n17542__, new_new_n17543__, new_new_n17544__,
    new_new_n17545__, new_new_n17546__, new_new_n17547__, new_new_n17548__,
    new_new_n17549__, new_new_n17550__, new_new_n17551__, new_new_n17552__,
    new_new_n17553__, new_new_n17554__, new_new_n17555__, new_new_n17556__,
    new_new_n17557__, new_new_n17558__, new_new_n17559__, new_new_n17560__,
    new_new_n17561__, new_new_n17562__, new_new_n17563__, new_new_n17564__,
    new_new_n17565__, new_new_n17566__, new_new_n17567__, new_new_n17568__,
    new_new_n17569__, new_new_n17570__, new_new_n17571__, new_new_n17572__,
    new_new_n17573__, new_new_n17574__, new_new_n17575__, new_new_n17576__,
    new_new_n17577__, new_new_n17578__, new_new_n17579__, new_new_n17580__,
    new_new_n17581__, new_new_n17582__, new_new_n17583__, new_new_n17584__,
    new_new_n17585__, new_new_n17586__, new_new_n17587__, new_new_n17588__,
    new_new_n17589__, new_new_n17590__, new_new_n17591__, new_new_n17592__,
    new_new_n17593__, new_new_n17594__, new_new_n17595__, new_new_n17596__,
    new_new_n17597__, new_new_n17598__, new_new_n17599__, new_new_n17600__,
    new_new_n17601__, new_new_n17602__, new_new_n17603__, new_new_n17604__,
    new_new_n17605__, new_new_n17606__, new_new_n17607__, new_new_n17608__,
    new_new_n17609__, new_new_n17610__, new_new_n17611__, new_new_n17612__,
    new_new_n17613__, new_new_n17614__, new_new_n17615__, new_new_n17616__,
    new_new_n17617__, new_new_n17618__, new_new_n17619__, new_new_n17620__,
    new_new_n17621__, new_new_n17622__, new_new_n17623__, new_new_n17624__,
    new_new_n17625__, new_new_n17626__, new_new_n17627__, new_new_n17628__,
    new_new_n17629__, new_new_n17630__, new_new_n17631__, new_new_n17632__,
    new_new_n17633__, new_new_n17634__, new_new_n17635__, new_new_n17636__,
    new_new_n17637__, new_new_n17638__, new_new_n17639__, new_new_n17640__,
    new_new_n17641__, new_new_n17642__, new_new_n17643__, new_new_n17644__,
    new_new_n17645__, new_new_n17646__, new_new_n17647__, new_new_n17648__,
    new_new_n17649__, new_new_n17650__, new_new_n17651__, new_new_n17652__,
    new_new_n17653__, new_new_n17654__, new_new_n17655__, new_new_n17656__,
    new_new_n17657__, new_new_n17658__, new_new_n17659__, new_new_n17660__,
    new_new_n17661__, new_new_n17662__, new_new_n17663__, new_new_n17664__,
    new_new_n17665__, new_new_n17666__, new_new_n17667__, new_new_n17668__,
    new_new_n17669__, new_new_n17670__, new_new_n17671__, new_new_n17672__,
    new_new_n17673__, new_new_n17674__, new_new_n17675__, new_new_n17676__,
    new_new_n17677__, new_new_n17678__, new_new_n17679__, new_new_n17680__,
    new_new_n17681__, new_new_n17682__, new_new_n17683__, new_new_n17684__,
    new_new_n17685__, new_new_n17686__, new_new_n17687__, new_new_n17688__,
    new_new_n17689__, new_new_n17690__, new_new_n17691__, new_new_n17692__,
    new_new_n17693__, new_new_n17694__, new_new_n17695__, new_new_n17696__,
    new_new_n17697__, new_new_n17698__, new_new_n17699__, new_new_n17700__,
    new_new_n17701__, new_new_n17702__, new_new_n17703__, new_new_n17704__,
    new_new_n17705__, new_new_n17706__, new_new_n17707__, new_new_n17708__,
    new_new_n17709__, new_new_n17710__, new_new_n17711__, new_new_n17712__,
    new_new_n17713__, new_new_n17714__, new_new_n17715__, new_new_n17716__,
    new_new_n17717__, new_new_n17718__, new_new_n17719__, new_new_n17720__,
    new_new_n17721__, new_new_n17722__, new_new_n17723__, new_new_n17724__,
    new_new_n17725__, new_new_n17726__, new_new_n17727__, new_new_n17728__,
    new_new_n17729__, new_new_n17730__, new_new_n17731__, new_new_n17732__,
    new_new_n17733__, new_new_n17734__, new_new_n17735__, new_new_n17736__,
    new_new_n17737__, new_new_n17738__, new_new_n17739__, new_new_n17740__,
    new_new_n17741__, new_new_n17742__, new_new_n17743__, new_new_n17744__,
    new_new_n17745__, new_new_n17746__, new_new_n17747__, new_new_n17748__,
    new_new_n17749__, new_new_n17750__, new_new_n17751__, new_new_n17752__,
    new_new_n17753__, new_new_n17754__, new_new_n17755__, new_new_n17756__,
    new_new_n17757__, new_new_n17758__, new_new_n17759__, new_new_n17760__,
    new_new_n17761__, new_new_n17762__, new_new_n17763__, new_new_n17764__,
    new_new_n17765__, new_new_n17766__, new_new_n17767__, new_new_n17768__,
    new_new_n17769__, new_new_n17770__, new_new_n17771__, new_new_n17772__,
    new_new_n17773__, new_new_n17774__, new_new_n17775__, new_new_n17776__,
    new_new_n17777__, new_new_n17778__, new_new_n17779__, new_new_n17780__,
    new_new_n17781__, new_new_n17782__, new_new_n17783__, new_new_n17784__,
    new_new_n17785__, new_new_n17786__, new_new_n17787__, new_new_n17788__,
    new_new_n17789__, new_new_n17790__, new_new_n17791__, new_new_n17792__,
    new_new_n17793__, new_new_n17794__, new_new_n17795__, new_new_n17796__,
    new_new_n17797__, new_new_n17798__, new_new_n17799__, new_new_n17800__,
    new_new_n17801__, new_new_n17802__, new_new_n17803__, new_new_n17804__,
    new_new_n17805__, new_new_n17806__, new_new_n17807__, new_new_n17808__,
    new_new_n17809__, new_new_n17810__, new_new_n17811__, new_new_n17812__,
    new_new_n17813__, new_new_n17814__, new_new_n17815__, new_new_n17816__,
    new_new_n17817__, new_new_n17818__, new_new_n17819__, new_new_n17820__,
    new_new_n17821__, new_new_n17822__, new_new_n17823__, new_new_n17824__,
    new_new_n17825__, new_new_n17826__, new_new_n17827__, new_new_n17828__,
    new_new_n17829__, new_new_n17830__, new_new_n17831__, new_new_n17832__,
    new_new_n17833__, new_new_n17834__, new_new_n17835__, new_new_n17836__,
    new_new_n17837__, new_new_n17838__, new_new_n17839__, new_new_n17840__,
    new_new_n17841__, new_new_n17842__, new_new_n17843__, new_new_n17844__,
    new_new_n17845__, new_new_n17846__, new_new_n17847__, new_new_n17848__,
    new_new_n17849__, new_new_n17850__, new_new_n17851__, new_new_n17852__,
    new_new_n17853__, new_new_n17854__, new_new_n17855__, new_new_n17856__,
    new_new_n17857__, new_new_n17858__, new_new_n17859__, new_new_n17860__,
    new_new_n17861__, new_new_n17862__, new_new_n17863__, new_new_n17864__,
    new_new_n17865__, new_new_n17866__, new_new_n17867__, new_new_n17868__,
    new_new_n17869__, new_new_n17870__, new_new_n17871__, new_new_n17872__,
    new_new_n17873__, new_new_n17874__, new_new_n17875__, new_new_n17876__,
    new_new_n17877__, new_new_n17878__, new_new_n17879__, new_new_n17880__,
    new_new_n17881__, new_new_n17882__, new_new_n17883__, new_new_n17884__,
    new_new_n17885__, new_new_n17886__, new_new_n17887__, new_new_n17888__,
    new_new_n17889__, new_new_n17890__, new_new_n17891__, new_new_n17892__,
    new_new_n17893__, new_new_n17894__, new_new_n17895__, new_new_n17896__,
    new_new_n17897__, new_new_n17898__, new_new_n17899__, new_new_n17900__,
    new_new_n17901__, new_new_n17902__, new_new_n17903__, new_new_n17904__,
    new_new_n17905__, new_new_n17906__, new_new_n17907__, new_new_n17908__,
    new_new_n17909__, new_new_n17910__, new_new_n17911__, new_new_n17912__,
    new_new_n17913__, new_new_n17914__, new_new_n17915__, new_new_n17916__,
    new_new_n17917__, new_new_n17918__, new_new_n17919__, new_new_n17920__,
    new_new_n17921__, new_new_n17922__, new_new_n17923__, new_new_n17924__,
    new_new_n17925__, new_new_n17926__, new_new_n17927__, new_new_n17928__,
    new_new_n17929__, new_new_n17930__, new_new_n17931__, new_new_n17932__,
    new_new_n17933__, new_new_n17934__, new_new_n17935__, new_new_n17936__,
    new_new_n17937__, new_new_n17938__, new_new_n17939__, new_new_n17940__,
    new_new_n17941__, new_new_n17942__, new_new_n17943__, new_new_n17944__,
    new_new_n17945__, new_new_n17946__, new_new_n17947__, new_new_n17948__,
    new_new_n17949__, new_new_n17950__, new_new_n17951__, new_new_n17952__,
    new_new_n17953__, new_new_n17954__, new_new_n17955__, new_new_n17956__,
    new_new_n17957__, new_new_n17958__, new_new_n17959__, new_new_n17960__,
    new_new_n17961__, new_new_n17962__, new_new_n17963__, new_new_n17964__,
    new_new_n17965__, new_new_n17966__, new_new_n17967__, new_new_n17968__,
    new_new_n17969__, new_new_n17970__, new_new_n17971__, new_new_n17972__,
    new_new_n17973__, new_new_n17974__, new_new_n17975__, new_new_n17976__,
    new_new_n17977__, new_new_n17978__, new_new_n17979__, new_new_n17980__,
    new_new_n17981__, new_new_n17982__, new_new_n17983__, new_new_n17984__,
    new_new_n17985__, new_new_n17986__, new_new_n17987__, new_new_n17988__,
    new_new_n17989__, new_new_n17990__, new_new_n17991__, new_new_n17992__,
    new_new_n17993__, new_new_n17994__, new_new_n17995__, new_new_n17996__,
    new_new_n17997__, new_new_n17998__, new_new_n17999__, new_new_n18000__,
    new_new_n18001__, new_new_n18002__, new_new_n18003__, new_new_n18004__,
    new_new_n18005__, new_new_n18006__, new_new_n18007__, new_new_n18008__,
    new_new_n18009__, new_new_n18010__, new_new_n18011__, new_new_n18012__,
    new_new_n18013__, new_new_n18014__, new_new_n18015__, new_new_n18016__,
    new_new_n18017__, new_new_n18018__, new_new_n18019__, new_new_n18020__,
    new_new_n18021__, new_new_n18022__, new_new_n18023__, new_new_n18024__,
    new_new_n18025__, new_new_n18026__, new_new_n18027__, new_new_n18028__,
    new_new_n18029__, new_new_n18030__, new_new_n18031__, new_new_n18032__,
    new_new_n18033__, new_new_n18034__, new_new_n18035__, new_new_n18036__,
    new_new_n18037__, new_new_n18038__, new_new_n18039__, new_new_n18040__,
    new_new_n18041__, new_new_n18042__, new_new_n18043__, new_new_n18044__,
    new_new_n18045__, new_new_n18046__, new_new_n18047__, new_new_n18048__,
    new_new_n18049__, new_new_n18050__, new_new_n18051__, new_new_n18052__,
    new_new_n18053__, new_new_n18054__, new_new_n18055__, new_new_n18056__,
    new_new_n18057__, new_new_n18058__, new_new_n18059__, new_new_n18060__,
    new_new_n18061__, new_new_n18062__, new_new_n18063__, new_new_n18064__,
    new_new_n18065__, new_new_n18066__, new_new_n18067__, new_new_n18068__,
    new_new_n18069__, new_new_n18070__, new_new_n18071__, new_new_n18072__,
    new_new_n18073__, new_new_n18074__, new_new_n18075__, new_new_n18076__,
    new_new_n18077__, new_new_n18078__, new_new_n18079__, new_new_n18080__,
    new_new_n18081__, new_new_n18082__, new_new_n18083__, new_new_n18084__,
    new_new_n18085__, new_new_n18086__, new_new_n18087__, new_new_n18088__,
    new_new_n18089__, new_new_n18090__, new_new_n18091__, new_new_n18092__,
    new_new_n18093__, new_new_n18094__, new_new_n18095__, new_new_n18096__,
    new_new_n18097__, new_new_n18098__, new_new_n18099__, new_new_n18100__,
    new_new_n18101__, new_new_n18102__, new_new_n18103__, new_new_n18104__,
    new_new_n18105__, new_new_n18106__, new_new_n18107__, new_new_n18108__,
    new_new_n18109__, new_new_n18110__, new_new_n18111__, new_new_n18112__,
    new_new_n18113__, new_new_n18114__, new_new_n18115__, new_new_n18116__,
    new_new_n18117__, new_new_n18118__, new_new_n18119__, new_new_n18120__,
    new_new_n18121__, new_new_n18122__, new_new_n18123__, new_new_n18124__,
    new_new_n18125__, new_new_n18126__, new_new_n18127__, new_new_n18128__,
    new_new_n18129__, new_new_n18130__, new_new_n18131__, new_new_n18132__,
    new_new_n18133__, new_new_n18134__, new_new_n18135__, new_new_n18136__,
    new_new_n18137__, new_new_n18138__, new_new_n18139__, new_new_n18140__,
    new_new_n18141__, new_new_n18142__, new_new_n18143__, new_new_n18144__,
    new_new_n18145__, new_new_n18146__, new_new_n18147__, new_new_n18148__,
    new_new_n18149__, new_new_n18150__, new_new_n18151__, new_new_n18152__,
    new_new_n18153__, new_new_n18154__, new_new_n18155__, new_new_n18156__,
    new_new_n18157__, new_new_n18158__, new_new_n18159__, new_new_n18160__,
    new_new_n18161__, new_new_n18162__, new_new_n18163__, new_new_n18164__,
    new_new_n18165__, new_new_n18166__, new_new_n18167__, new_new_n18168__,
    new_new_n18169__, new_new_n18170__, new_new_n18171__, new_new_n18172__,
    new_new_n18173__, new_new_n18174__, new_new_n18175__, new_new_n18176__,
    new_new_n18177__, new_new_n18178__, new_new_n18179__, new_new_n18180__,
    new_new_n18181__, new_new_n18182__, new_new_n18183__, new_new_n18184__,
    new_new_n18185__, new_new_n18186__, new_new_n18187__, new_new_n18188__,
    new_new_n18189__, new_new_n18190__, new_new_n18191__, new_new_n18192__,
    new_new_n18193__, new_new_n18194__, new_new_n18195__, new_new_n18196__,
    new_new_n18197__, new_new_n18198__, new_new_n18199__, new_new_n18200__,
    new_new_n18201__, new_new_n18202__, new_new_n18203__, new_new_n18204__,
    new_new_n18205__, new_new_n18206__, new_new_n18207__, new_new_n18208__,
    new_new_n18209__, new_new_n18210__, new_new_n18211__, new_new_n18212__,
    new_new_n18213__, new_new_n18214__, new_new_n18215__, new_new_n18216__,
    new_new_n18217__, new_new_n18218__, new_new_n18219__, new_new_n18220__,
    new_new_n18221__, new_new_n18222__, new_new_n18223__, new_new_n18224__,
    new_new_n18225__, new_new_n18226__, new_new_n18227__, new_new_n18228__,
    new_new_n18229__, new_new_n18230__, new_new_n18231__, new_new_n18232__,
    new_new_n18233__, new_new_n18234__, new_new_n18235__, new_new_n18236__,
    new_new_n18237__, new_new_n18238__, new_new_n18239__, new_new_n18240__,
    new_new_n18241__, new_new_n18242__, new_new_n18243__, new_new_n18244__,
    new_new_n18245__, new_new_n18246__, new_new_n18247__, new_new_n18248__,
    new_new_n18249__, new_new_n18250__, new_new_n18251__, new_new_n18252__,
    new_new_n18253__, new_new_n18254__, new_new_n18255__, new_new_n18256__,
    new_new_n18257__, new_new_n18258__, new_new_n18259__, new_new_n18260__,
    new_new_n18261__, new_new_n18262__, new_new_n18263__, new_new_n18264__,
    new_new_n18265__, new_new_n18266__, new_new_n18267__, new_new_n18268__,
    new_new_n18269__, new_new_n18270__, new_new_n18271__, new_new_n18272__,
    new_new_n18273__, new_new_n18274__, new_new_n18275__, new_new_n18276__,
    new_new_n18277__, new_new_n18278__, new_new_n18279__, new_new_n18280__,
    new_new_n18281__, new_new_n18282__, new_new_n18283__, new_new_n18284__,
    new_new_n18285__, new_new_n18286__, new_new_n18287__, new_new_n18288__,
    new_new_n18289__, new_new_n18290__, new_new_n18291__, new_new_n18292__,
    new_new_n18293__, new_new_n18294__, new_new_n18295__, new_new_n18296__,
    new_new_n18297__, new_new_n18298__, new_new_n18299__, new_new_n18300__,
    new_new_n18301__, new_new_n18302__, new_new_n18303__, new_new_n18304__,
    new_new_n18305__, new_new_n18306__, new_new_n18307__, new_new_n18308__,
    new_new_n18309__, new_new_n18310__, new_new_n18311__, new_new_n18312__,
    new_new_n18313__, new_new_n18314__, new_new_n18315__, new_new_n18316__,
    new_new_n18317__, new_new_n18318__, new_new_n18319__, new_new_n18320__,
    new_new_n18321__, new_new_n18322__, new_new_n18323__, new_new_n18324__,
    new_new_n18325__, new_new_n18326__, new_new_n18327__, new_new_n18328__,
    new_new_n18329__, new_new_n18330__, new_new_n18331__, new_new_n18332__,
    new_new_n18333__, new_new_n18334__, new_new_n18335__, new_new_n18336__,
    new_new_n18337__, new_new_n18338__, new_new_n18339__, new_new_n18340__,
    new_new_n18341__, new_new_n18342__, new_new_n18343__, new_new_n18344__,
    new_new_n18345__, new_new_n18346__, new_new_n18347__, new_new_n18348__,
    new_new_n18349__, new_new_n18350__, new_new_n18351__, new_new_n18352__,
    new_new_n18353__, new_new_n18354__, new_new_n18355__, new_new_n18356__,
    new_new_n18357__, new_new_n18358__, new_new_n18359__, new_new_n18360__,
    new_new_n18361__, new_new_n18362__, new_new_n18363__, new_new_n18364__,
    new_new_n18365__, new_new_n18366__, new_new_n18367__, new_new_n18368__,
    new_new_n18369__, new_new_n18370__, new_new_n18371__, new_new_n18372__,
    new_new_n18373__, new_new_n18374__, new_new_n18375__, new_new_n18376__,
    new_new_n18377__, new_new_n18378__, new_new_n18379__, new_new_n18380__,
    new_new_n18381__, new_new_n18382__, new_new_n18383__, new_new_n18384__,
    new_new_n18385__, new_new_n18386__, new_new_n18387__, new_new_n18388__,
    new_new_n18389__, new_new_n18390__, new_new_n18391__, new_new_n18392__,
    new_new_n18393__, new_new_n18394__, new_new_n18395__, new_new_n18396__,
    new_new_n18397__, new_new_n18398__, new_new_n18399__, new_new_n18400__,
    new_new_n18401__, new_new_n18402__, new_new_n18403__, new_new_n18404__,
    new_new_n18405__, new_new_n18406__, new_new_n18407__, new_new_n18408__,
    new_new_n18409__, new_new_n18410__, new_new_n18411__, new_new_n18412__,
    new_new_n18413__, new_new_n18414__, new_new_n18415__, new_new_n18416__,
    new_new_n18417__, new_new_n18418__, new_new_n18419__, new_new_n18420__,
    new_new_n18421__, new_new_n18422__, new_new_n18423__, new_new_n18424__,
    new_new_n18425__, new_new_n18426__, new_new_n18427__, new_new_n18428__,
    new_new_n18429__, new_new_n18430__, new_new_n18431__, new_new_n18432__,
    new_new_n18433__, new_new_n18434__, new_new_n18435__, new_new_n18436__,
    new_new_n18437__, new_new_n18438__, new_new_n18439__, new_new_n18440__,
    new_new_n18441__, new_new_n18442__, new_new_n18443__, new_new_n18444__,
    new_new_n18445__, new_new_n18446__, new_new_n18447__, new_new_n18448__,
    new_new_n18449__, new_new_n18450__, new_new_n18451__, new_new_n18452__,
    new_new_n18453__, new_new_n18454__, new_new_n18455__, new_new_n18456__,
    new_new_n18457__, new_new_n18458__, new_new_n18459__, new_new_n18460__,
    new_new_n18461__, new_new_n18462__, new_new_n18463__, new_new_n18464__,
    new_new_n18465__, new_new_n18466__, new_new_n18467__, new_new_n18468__,
    new_new_n18469__, new_new_n18470__, new_new_n18471__, new_new_n18472__,
    new_new_n18473__, new_new_n18474__, new_new_n18475__, new_new_n18476__,
    new_new_n18477__, new_new_n18478__, new_new_n18479__, new_new_n18480__,
    new_new_n18481__, new_new_n18482__, new_new_n18483__, new_new_n18484__,
    new_new_n18485__, new_new_n18486__, new_new_n18487__, new_new_n18488__,
    new_new_n18489__, new_new_n18490__, new_new_n18491__, new_new_n18492__,
    new_new_n18493__, new_new_n18494__, new_new_n18495__, new_new_n18496__,
    new_new_n18497__, new_new_n18498__, new_new_n18499__, new_new_n18500__,
    new_new_n18501__, new_new_n18502__, new_new_n18503__, new_new_n18504__,
    new_new_n18505__, new_new_n18506__, new_new_n18507__, new_new_n18508__,
    new_new_n18509__, new_new_n18510__, new_new_n18511__, new_new_n18512__,
    new_new_n18513__, new_new_n18514__, new_new_n18515__, new_new_n18516__,
    new_new_n18517__, new_new_n18518__, new_new_n18519__, new_new_n18520__,
    new_new_n18521__, new_new_n18522__, new_new_n18523__, new_new_n18524__,
    new_new_n18525__, new_new_n18526__, new_new_n18527__, new_new_n18528__,
    new_new_n18529__, new_new_n18530__, new_new_n18531__, new_new_n18532__,
    new_new_n18533__, new_new_n18534__, new_new_n18535__, new_new_n18536__,
    new_new_n18537__, new_new_n18538__, new_new_n18539__, new_new_n18540__,
    new_new_n18541__, new_new_n18542__, new_new_n18543__, new_new_n18544__,
    new_new_n18545__, new_new_n18546__, new_new_n18547__, new_new_n18548__,
    new_new_n18549__, new_new_n18550__, new_new_n18551__, new_new_n18552__,
    new_new_n18553__, new_new_n18554__, new_new_n18555__, new_new_n18556__,
    new_new_n18557__, new_new_n18558__, new_new_n18559__, new_new_n18560__,
    new_new_n18561__, new_new_n18562__, new_new_n18563__, new_new_n18564__,
    new_new_n18565__, new_new_n18566__, new_new_n18567__, new_new_n18568__,
    new_new_n18569__, new_new_n18570__, new_new_n18571__, new_new_n18572__,
    new_new_n18573__, new_new_n18574__, new_new_n18575__, new_new_n18576__,
    new_new_n18577__, new_new_n18578__, new_new_n18579__, new_new_n18580__,
    new_new_n18581__, new_new_n18582__, new_new_n18583__, new_new_n18584__,
    new_new_n18585__, new_new_n18586__, new_new_n18587__, new_new_n18588__,
    new_new_n18589__, new_new_n18590__, new_new_n18591__, new_new_n18592__,
    new_new_n18593__, new_new_n18594__, new_new_n18595__, new_new_n18596__,
    new_new_n18597__, new_new_n18598__, new_new_n18599__, new_new_n18600__,
    new_new_n18601__, new_new_n18602__, new_new_n18603__, new_new_n18604__,
    new_new_n18605__, new_new_n18606__, new_new_n18607__, new_new_n18608__,
    new_new_n18609__, new_new_n18610__, new_new_n18611__, new_new_n18612__,
    new_new_n18613__, new_new_n18614__, new_new_n18615__, new_new_n18616__,
    new_new_n18617__, new_new_n18618__, new_new_n18619__, new_new_n18620__,
    new_new_n18621__, new_new_n18622__, new_new_n18623__, new_new_n18624__,
    new_new_n18625__, new_new_n18626__, new_new_n18627__, new_new_n18628__,
    new_new_n18629__, new_new_n18630__, new_new_n18631__, new_new_n18632__,
    new_new_n18633__, new_new_n18634__, new_new_n18635__, new_new_n18636__,
    new_new_n18637__, new_new_n18638__, new_new_n18639__, new_new_n18640__,
    new_new_n18641__, new_new_n18642__, new_new_n18643__, new_new_n18644__,
    new_new_n18645__, new_new_n18646__, new_new_n18647__, new_new_n18648__,
    new_new_n18649__, new_new_n18650__, new_new_n18651__, new_new_n18652__,
    new_new_n18653__, new_new_n18654__, new_new_n18655__, new_new_n18656__,
    new_new_n18657__, new_new_n18658__, new_new_n18659__, new_new_n18660__,
    new_new_n18661__, new_new_n18662__, new_new_n18663__, new_new_n18664__,
    new_new_n18665__, new_new_n18666__, new_new_n18667__, new_new_n18668__,
    new_new_n18669__, new_new_n18670__, new_new_n18671__, new_new_n18672__,
    new_new_n18673__, new_new_n18674__, new_new_n18675__, new_new_n18676__,
    new_new_n18677__, new_new_n18678__, new_new_n18679__, new_new_n18680__,
    new_new_n18681__, new_new_n18682__, new_new_n18683__, new_new_n18684__,
    new_new_n18685__, new_new_n18686__, new_new_n18687__, new_new_n18688__,
    new_new_n18689__, new_new_n18690__, new_new_n18691__, new_new_n18692__,
    new_new_n18693__, new_new_n18694__, new_new_n18695__, new_new_n18696__,
    new_new_n18697__, new_new_n18698__, new_new_n18699__, new_new_n18700__,
    new_new_n18701__, new_new_n18702__, new_new_n18703__, new_new_n18704__,
    new_new_n18705__, new_new_n18706__, new_new_n18707__, new_new_n18708__,
    new_new_n18709__, new_new_n18710__, new_new_n18711__, new_new_n18712__,
    new_new_n18713__, new_new_n18714__, new_new_n18715__, new_new_n18716__,
    new_new_n18717__, new_new_n18718__, new_new_n18719__, new_new_n18720__,
    new_new_n18721__, new_new_n18722__, new_new_n18723__, new_new_n18724__,
    new_new_n18725__, new_new_n18726__, new_new_n18727__, new_new_n18728__,
    new_new_n18729__, new_new_n18730__, new_new_n18731__, new_new_n18732__,
    new_new_n18733__, new_new_n18734__, new_new_n18735__, new_new_n18736__,
    new_new_n18737__, new_new_n18738__, new_new_n18739__, new_new_n18740__,
    new_new_n18741__, new_new_n18742__, new_new_n18743__, new_new_n18744__,
    new_new_n18745__, new_new_n18746__, new_new_n18747__, new_new_n18748__,
    new_new_n18749__, new_new_n18750__, new_new_n18751__, new_new_n18752__,
    new_new_n18753__, new_new_n18754__, new_new_n18755__, new_new_n18756__,
    new_new_n18757__, new_new_n18758__, new_new_n18759__, new_new_n18760__,
    new_new_n18761__, new_new_n18762__, new_new_n18763__, new_new_n18764__,
    new_new_n18765__, new_new_n18766__, new_new_n18767__, new_new_n18768__,
    new_new_n18769__, new_new_n18770__, new_new_n18771__, new_new_n18772__,
    new_new_n18773__, new_new_n18774__, new_new_n18775__, new_new_n18776__,
    new_new_n18777__, new_new_n18778__, new_new_n18779__, new_new_n18780__,
    new_new_n18781__, new_new_n18782__, new_new_n18783__, new_new_n18784__,
    new_new_n18785__, new_new_n18786__, new_new_n18787__, new_new_n18788__,
    new_new_n18789__, new_new_n18790__, new_new_n18791__, new_new_n18792__,
    new_new_n18793__, new_new_n18794__, new_new_n18795__, new_new_n18796__,
    new_new_n18797__, new_new_n18798__, new_new_n18799__, new_new_n18800__,
    new_new_n18801__, new_new_n18802__, new_new_n18803__, new_new_n18804__,
    new_new_n18805__, new_new_n18806__, new_new_n18807__, new_new_n18808__,
    new_new_n18809__, new_new_n18810__, new_new_n18811__, new_new_n18812__,
    new_new_n18813__, new_new_n18814__, new_new_n18815__, new_new_n18816__,
    new_new_n18817__, new_new_n18818__, new_new_n18819__, new_new_n18820__,
    new_new_n18821__, new_new_n18822__, new_new_n18823__, new_new_n18824__,
    new_new_n18825__, new_new_n18826__, new_new_n18827__, new_new_n18828__,
    new_new_n18829__, new_new_n18830__, new_new_n18831__, new_new_n18832__,
    new_new_n18833__, new_new_n18834__, new_new_n18835__, new_new_n18836__,
    new_new_n18837__, new_new_n18838__, new_new_n18839__, new_new_n18840__,
    new_new_n18841__, new_new_n18842__, new_new_n18843__, new_new_n18844__,
    new_new_n18845__, new_new_n18846__, new_new_n18847__, new_new_n18848__,
    new_new_n18849__, new_new_n18850__, new_new_n18851__, new_new_n18852__,
    new_new_n18853__, new_new_n18854__, new_new_n18855__, new_new_n18856__,
    new_new_n18857__, new_new_n18858__, new_new_n18859__, new_new_n18860__,
    new_new_n18861__, new_new_n18862__, new_new_n18863__, new_new_n18864__,
    new_new_n18865__, new_new_n18866__, new_new_n18867__, new_new_n18868__,
    new_new_n18869__, new_new_n18870__, new_new_n18871__, new_new_n18872__,
    new_new_n18873__, new_new_n18874__, new_new_n18875__, new_new_n18876__,
    new_new_n18877__, new_new_n18878__, new_new_n18879__, new_new_n18880__,
    new_new_n18881__, new_new_n18882__, new_new_n18883__, new_new_n18884__,
    new_new_n18885__, new_new_n18886__, new_new_n18887__, new_new_n18888__,
    new_new_n18889__, new_new_n18890__, new_new_n18891__, new_new_n18892__,
    new_new_n18893__, new_new_n18894__, new_new_n18895__, new_new_n18896__,
    new_new_n18897__, new_new_n18898__, new_new_n18899__, new_new_n18900__,
    new_new_n18901__, new_new_n18902__, new_new_n18903__, new_new_n18904__,
    new_new_n18905__, new_new_n18906__, new_new_n18907__, new_new_n18908__,
    new_new_n18909__, new_new_n18910__, new_new_n18911__, new_new_n18912__,
    new_new_n18913__, new_new_n18914__, new_new_n18915__, new_new_n18916__,
    new_new_n18917__, new_new_n18918__, new_new_n18919__, new_new_n18920__,
    new_new_n18921__, new_new_n18922__, new_new_n18923__, new_new_n18924__,
    new_new_n18925__, new_new_n18926__, new_new_n18927__, new_new_n18928__,
    new_new_n18929__, new_new_n18930__, new_new_n18931__, new_new_n18932__,
    new_new_n18933__, new_new_n18934__, new_new_n18935__, new_new_n18936__,
    new_new_n18937__, new_new_n18938__, new_new_n18939__, new_new_n18940__,
    new_new_n18941__, new_new_n18942__, new_new_n18943__, new_new_n18944__,
    new_new_n18945__, new_new_n18946__, new_new_n18947__, new_new_n18948__,
    new_new_n18949__, new_new_n18950__, new_new_n18951__, new_new_n18952__,
    new_new_n18953__, new_new_n18954__, new_new_n18955__, new_new_n18956__,
    new_new_n18957__, new_new_n18958__, new_new_n18959__, new_new_n18960__,
    new_new_n18961__, new_new_n18962__, new_new_n18963__, new_new_n18964__,
    new_new_n18965__, new_new_n18966__, new_new_n18967__, new_new_n18968__,
    new_new_n18969__, new_new_n18970__, new_new_n18971__, new_new_n18972__,
    new_new_n18973__, new_new_n18974__, new_new_n18975__, new_new_n18976__,
    new_new_n18977__, new_new_n18978__, new_new_n18979__, new_new_n18980__,
    new_new_n18981__, new_new_n18982__, new_new_n18983__, new_new_n18984__,
    new_new_n18985__, new_new_n18986__, new_new_n18987__, new_new_n18988__,
    new_new_n18989__, new_new_n18990__, new_new_n18991__, new_new_n18992__,
    new_new_n18993__, new_new_n18994__, new_new_n18995__, new_new_n18996__,
    new_new_n18997__, new_new_n18998__, new_new_n18999__, new_new_n19000__,
    new_new_n19001__, new_new_n19002__, new_new_n19003__, new_new_n19004__,
    new_new_n19005__, new_new_n19006__, new_new_n19007__, new_new_n19008__,
    new_new_n19009__, new_new_n19010__, new_new_n19011__, new_new_n19012__,
    new_new_n19013__, new_new_n19014__, new_new_n19015__, new_new_n19016__,
    new_new_n19017__, new_new_n19018__, new_new_n19019__, new_new_n19020__,
    new_new_n19021__, new_new_n19022__, new_new_n19023__, new_new_n19024__,
    new_new_n19025__, new_new_n19026__, new_new_n19027__, new_new_n19028__,
    new_new_n19029__, new_new_n19030__, new_new_n19031__, new_new_n19032__,
    new_new_n19033__, new_new_n19034__, new_new_n19035__, new_new_n19036__,
    new_new_n19037__, new_new_n19038__, new_new_n19039__, new_new_n19040__,
    new_new_n19041__, new_new_n19042__, new_new_n19043__, new_new_n19044__,
    new_new_n19045__, new_new_n19046__, new_new_n19047__, new_new_n19048__,
    new_new_n19049__, new_new_n19050__, new_new_n19051__, new_new_n19052__,
    new_new_n19053__, new_new_n19054__, new_new_n19055__, new_new_n19056__,
    new_new_n19057__, new_new_n19058__, new_new_n19059__, new_new_n19060__,
    new_new_n19061__, new_new_n19062__, new_new_n19063__, new_new_n19064__,
    new_new_n19065__, new_new_n19066__, new_new_n19067__, new_new_n19068__,
    new_new_n19069__, new_new_n19070__, new_new_n19071__, new_new_n19072__,
    new_new_n19073__, new_new_n19074__, new_new_n19075__, new_new_n19076__,
    new_new_n19077__, new_new_n19078__, new_new_n19079__, new_new_n19080__,
    new_new_n19081__, new_new_n19082__, new_new_n19083__, new_new_n19084__,
    new_new_n19085__, new_new_n19086__, new_new_n19087__, new_new_n19088__,
    new_new_n19089__, new_new_n19090__, new_new_n19091__, new_new_n19092__,
    new_new_n19093__, new_new_n19094__, new_new_n19095__, new_new_n19096__,
    new_new_n19097__, new_new_n19098__, new_new_n19099__, new_new_n19100__,
    new_new_n19101__, new_new_n19102__, new_new_n19103__, new_new_n19104__,
    new_new_n19105__, new_new_n19106__, new_new_n19107__, new_new_n19108__,
    new_new_n19109__, new_new_n19110__, new_new_n19111__, new_new_n19112__,
    new_new_n19113__, new_new_n19114__, new_new_n19115__, new_new_n19116__,
    new_new_n19117__, new_new_n19118__, new_new_n19119__, new_new_n19120__,
    new_new_n19121__, new_new_n19122__, new_new_n19123__, new_new_n19124__,
    new_new_n19125__, new_new_n19126__, new_new_n19127__, new_new_n19128__,
    new_new_n19129__, new_new_n19130__, new_new_n19131__, new_new_n19132__,
    new_new_n19133__, new_new_n19134__, new_new_n19135__, new_new_n19136__,
    new_new_n19137__, new_new_n19138__, new_new_n19139__, new_new_n19140__,
    new_new_n19141__, new_new_n19142__, new_new_n19143__, new_new_n19144__,
    new_new_n19145__, new_new_n19146__, new_new_n19147__, new_new_n19148__,
    new_new_n19149__, new_new_n19150__, new_new_n19151__, new_new_n19152__,
    new_new_n19153__, new_new_n19154__, new_new_n19155__, new_new_n19156__,
    new_new_n19157__, new_new_n19158__, new_new_n19159__, new_new_n19160__,
    new_new_n19161__, new_new_n19162__, new_new_n19163__, new_new_n19164__,
    new_new_n19165__, new_new_n19166__, new_new_n19167__, new_new_n19168__,
    new_new_n19169__, new_new_n19170__, new_new_n19171__, new_new_n19172__,
    new_new_n19173__, new_new_n19174__, new_new_n19175__, new_new_n19176__,
    new_new_n19177__, new_new_n19178__, new_new_n19179__, new_new_n19180__,
    new_new_n19181__, new_new_n19182__, new_new_n19183__, new_new_n19184__,
    new_new_n19185__, new_new_n19186__, new_new_n19187__, new_new_n19188__,
    new_new_n19189__, new_new_n19190__, new_new_n19191__, new_new_n19192__,
    new_new_n19193__, new_new_n19194__, new_new_n19195__, new_new_n19196__,
    new_new_n19197__, new_new_n19198__, new_new_n19199__, new_new_n19200__,
    new_new_n19201__, new_new_n19202__, new_new_n19203__, new_new_n19204__,
    new_new_n19205__, new_new_n19206__, new_new_n19207__, new_new_n19208__,
    new_new_n19209__, new_new_n19210__, new_new_n19211__, new_new_n19212__,
    new_new_n19213__, new_new_n19214__, new_new_n19215__, new_new_n19216__,
    new_new_n19217__, new_new_n19218__, new_new_n19219__, new_new_n19220__,
    new_new_n19221__, new_new_n19222__, new_new_n19223__, new_new_n19224__,
    new_new_n19225__, new_new_n19226__, new_new_n19227__, new_new_n19228__,
    new_new_n19229__, new_new_n19230__, new_new_n19231__, new_new_n19232__,
    new_new_n19233__, new_new_n19234__, new_new_n19235__, new_new_n19236__,
    new_new_n19237__, new_new_n19238__, new_new_n19239__, new_new_n19240__,
    new_new_n19241__, new_new_n19242__, new_new_n19243__, new_new_n19244__,
    new_new_n19245__, new_new_n19246__, new_new_n19247__, new_new_n19248__,
    new_new_n19249__, new_new_n19250__, new_new_n19251__, new_new_n19252__,
    new_new_n19253__, new_new_n19254__, new_new_n19255__, new_new_n19256__,
    new_new_n19257__, new_new_n19258__, new_new_n19259__, new_new_n19260__,
    new_new_n19261__, new_new_n19262__, new_new_n19263__, new_new_n19264__,
    new_new_n19265__, new_new_n19266__, new_new_n19267__, new_new_n19268__,
    new_new_n19269__, new_new_n19270__, new_new_n19271__, new_new_n19272__,
    new_new_n19273__, new_new_n19274__, new_new_n19275__, new_new_n19276__,
    new_new_n19277__, new_new_n19278__, new_new_n19279__, new_new_n19280__,
    new_new_n19281__, new_new_n19282__, new_new_n19283__, new_new_n19284__,
    new_new_n19285__, new_new_n19286__, new_new_n19287__, new_new_n19288__,
    new_new_n19289__, new_new_n19290__, new_new_n19291__, new_new_n19292__,
    new_new_n19293__, new_new_n19294__, new_new_n19295__, new_new_n19296__,
    new_new_n19297__, new_new_n19298__, new_new_n19299__, new_new_n19300__,
    new_new_n19301__, new_new_n19302__, new_new_n19303__, new_new_n19304__,
    new_new_n19305__, new_new_n19306__, new_new_n19307__, new_new_n19308__,
    new_new_n19309__, new_new_n19310__, new_new_n19311__, new_new_n19312__,
    new_new_n19313__, new_new_n19314__, new_new_n19315__, new_new_n19316__,
    new_new_n19317__, new_new_n19318__, new_new_n19319__, new_new_n19320__,
    new_new_n19321__, new_new_n19322__, new_new_n19323__, new_new_n19324__,
    new_new_n19325__, new_new_n19326__, new_new_n19327__, new_new_n19328__,
    new_new_n19329__, new_new_n19330__, new_new_n19331__, new_new_n19332__,
    new_new_n19333__, new_new_n19334__, new_new_n19335__, new_new_n19336__,
    new_new_n19337__, new_new_n19338__, new_new_n19339__, new_new_n19340__,
    new_new_n19341__, new_new_n19342__, new_new_n19343__, new_new_n19344__,
    new_new_n19345__, new_new_n19346__, new_new_n19347__, new_new_n19348__,
    new_new_n19349__, new_new_n19350__, new_new_n19351__, new_new_n19352__,
    new_new_n19353__, new_new_n19354__, new_new_n19355__, new_new_n19356__,
    new_new_n19357__, new_new_n19358__, new_new_n19359__, new_new_n19360__,
    new_new_n19361__, new_new_n19362__, new_new_n19363__, new_new_n19364__,
    new_new_n19365__, new_new_n19366__, new_new_n19367__, new_new_n19368__,
    new_new_n19369__, new_new_n19370__, new_new_n19371__, new_new_n19372__,
    new_new_n19373__, new_new_n19374__, new_new_n19375__, new_new_n19376__,
    new_new_n19377__, new_new_n19378__, new_new_n19379__, new_new_n19380__,
    new_new_n19381__, new_new_n19382__, new_new_n19383__, new_new_n19384__,
    new_new_n19385__, new_new_n19386__, new_new_n19387__, new_new_n19388__,
    new_new_n19389__, new_new_n19390__, new_new_n19391__, new_new_n19392__,
    new_new_n19393__, new_new_n19394__, new_new_n19395__, new_new_n19396__,
    new_new_n19397__, new_new_n19398__, new_new_n19399__, new_new_n19400__,
    new_new_n19401__, new_new_n19402__, new_new_n19403__, new_new_n19404__,
    new_new_n19405__, new_new_n19406__, new_new_n19407__, new_new_n19408__,
    new_new_n19409__, new_new_n19410__, new_new_n19411__, new_new_n19412__,
    new_new_n19413__, new_new_n19414__, new_new_n19415__, new_new_n19416__,
    new_new_n19417__, new_new_n19418__, new_new_n19419__, new_new_n19420__,
    new_new_n19421__, new_new_n19422__, new_new_n19423__, new_new_n19424__,
    new_new_n19425__, new_new_n19426__, new_new_n19427__, new_new_n19428__,
    new_new_n19429__, new_new_n19430__, new_new_n19431__, new_new_n19432__,
    new_new_n19433__, new_new_n19434__, new_new_n19435__, new_new_n19436__,
    new_new_n19437__, new_new_n19438__, new_new_n19439__, new_new_n19440__,
    new_new_n19441__, new_new_n19442__, new_new_n19443__, new_new_n19444__,
    new_new_n19445__, new_new_n19446__, new_new_n19447__, new_new_n19448__,
    new_new_n19449__, new_new_n19450__, new_new_n19451__, new_new_n19452__,
    new_new_n19453__, new_new_n19454__, new_new_n19455__, new_new_n19456__,
    new_new_n19457__, new_new_n19458__, new_new_n19459__, new_new_n19460__,
    new_new_n19461__, new_new_n19462__, new_new_n19463__, new_new_n19464__,
    new_new_n19465__, new_new_n19466__, new_new_n19467__, new_new_n19468__,
    new_new_n19469__, new_new_n19470__, new_new_n19471__, new_new_n19472__,
    new_new_n19473__, new_new_n19474__, new_new_n19475__, new_new_n19476__,
    new_new_n19477__, new_new_n19478__, new_new_n19479__, new_new_n19480__,
    new_new_n19481__, new_new_n19482__, new_new_n19483__, new_new_n19484__,
    new_new_n19485__, new_new_n19486__, new_new_n19487__, new_new_n19488__,
    new_new_n19489__, new_new_n19490__, new_new_n19491__, new_new_n19492__,
    new_new_n19493__, new_new_n19494__, new_new_n19495__, new_new_n19496__,
    new_new_n19497__, new_new_n19498__, new_new_n19499__, new_new_n19500__,
    new_new_n19501__, new_new_n19502__, new_new_n19503__, new_new_n19504__,
    new_new_n19505__, new_new_n19506__, new_new_n19507__, new_new_n19508__,
    new_new_n19509__, new_new_n19510__, new_new_n19511__, new_new_n19512__,
    new_new_n19513__, new_new_n19514__, new_new_n19515__, new_new_n19516__,
    new_new_n19517__, new_new_n19518__, new_new_n19519__, new_new_n19520__,
    new_new_n19521__, new_new_n19522__, new_new_n19523__, new_new_n19524__,
    new_new_n19525__, new_new_n19526__, new_new_n19527__, new_new_n19528__,
    new_new_n19529__, new_new_n19530__, new_new_n19531__, new_new_n19532__,
    new_new_n19533__, new_new_n19534__, new_new_n19535__, new_new_n19536__,
    new_new_n19537__, new_new_n19538__, new_new_n19539__, new_new_n19540__,
    new_new_n19541__, new_new_n19542__, new_new_n19543__, new_new_n19544__,
    new_new_n19545__, new_new_n19546__, new_new_n19547__, new_new_n19548__,
    new_new_n19549__, new_new_n19550__, new_new_n19551__, new_new_n19552__,
    new_new_n19553__, new_new_n19554__, new_new_n19555__, new_new_n19556__,
    new_new_n19557__, new_new_n19558__, new_new_n19559__, new_new_n19560__,
    new_new_n19561__, new_new_n19562__, new_new_n19563__, new_new_n19564__,
    new_new_n19565__, new_new_n19566__, new_new_n19567__, new_new_n19568__,
    new_new_n19569__, new_new_n19570__, new_new_n19571__, new_new_n19572__,
    new_new_n19573__, new_new_n19574__, new_new_n19575__, new_new_n19576__,
    new_new_n19577__, new_new_n19578__, new_new_n19579__, new_new_n19580__,
    new_new_n19581__, new_new_n19582__, new_new_n19583__, new_new_n19584__,
    new_new_n19585__, new_new_n19586__, new_new_n19587__, new_new_n19588__,
    new_new_n19589__, new_new_n19590__, new_new_n19591__, new_new_n19592__,
    new_new_n19593__, new_new_n19594__, new_new_n19595__, new_new_n19596__,
    new_new_n19597__, new_new_n19598__, new_new_n19599__, new_new_n19600__,
    new_new_n19601__, new_new_n19602__, new_new_n19603__, new_new_n19604__,
    new_new_n19605__, new_new_n19606__, new_new_n19607__, new_new_n19608__,
    new_new_n19609__, new_new_n19610__, new_new_n19611__, new_new_n19612__,
    new_new_n19613__, new_new_n19614__, new_new_n19615__, new_new_n19616__,
    new_new_n19617__, new_new_n19618__, new_new_n19619__, new_new_n19620__,
    new_new_n19621__, new_new_n19622__, new_new_n19623__, new_new_n19624__,
    new_new_n19625__, new_new_n19626__, new_new_n19627__, new_new_n19628__,
    new_new_n19629__, new_new_n19630__, new_new_n19631__, new_new_n19632__,
    new_new_n19633__, new_new_n19634__, new_new_n19635__, new_new_n19636__,
    new_new_n19637__, new_new_n19638__, new_new_n19639__, new_new_n19640__,
    new_new_n19641__, new_new_n19642__, new_new_n19643__, new_new_n19644__,
    new_new_n19645__, new_new_n19646__, new_new_n19647__, new_new_n19648__,
    new_new_n19649__, new_new_n19650__, new_new_n19651__, new_new_n19652__,
    new_new_n19653__, new_new_n19654__, new_new_n19655__, new_new_n19656__,
    new_new_n19657__, new_new_n19658__, new_new_n19659__, new_new_n19660__,
    new_new_n19661__, new_new_n19662__, new_new_n19663__, new_new_n19664__,
    new_new_n19665__, new_new_n19666__, new_new_n19667__, new_new_n19668__,
    new_new_n19669__, new_new_n19670__, new_new_n19671__, new_new_n19672__,
    new_new_n19673__, new_new_n19674__, new_new_n19675__, new_new_n19676__,
    new_new_n19677__, new_new_n19678__, new_new_n19679__, new_new_n19680__,
    new_new_n19681__, new_new_n19682__, new_new_n19683__, new_new_n19684__,
    new_new_n19685__, new_new_n19686__, new_new_n19687__, new_new_n19688__,
    new_new_n19689__, new_new_n19690__, new_new_n19691__, new_new_n19692__,
    new_new_n19693__, new_new_n19694__, new_new_n19695__, new_new_n19696__,
    new_new_n19697__, new_new_n19698__, new_new_n19699__, new_new_n19700__,
    new_new_n19701__, new_new_n19702__, new_new_n19703__, new_new_n19704__,
    new_new_n19705__, new_new_n19706__, new_new_n19707__, new_new_n19708__,
    new_new_n19709__, new_new_n19710__, new_new_n19711__, new_new_n19712__,
    new_new_n19713__, new_new_n19714__, new_new_n19715__, new_new_n19716__,
    new_new_n19717__, new_new_n19718__, new_new_n19719__, new_new_n19720__,
    new_new_n19721__, new_new_n19722__, new_new_n19723__, new_new_n19724__,
    new_new_n19725__, new_new_n19726__, new_new_n19727__, new_new_n19728__,
    new_new_n19729__, new_new_n19730__, new_new_n19731__, new_new_n19732__,
    new_new_n19733__, new_new_n19734__, new_new_n19735__, new_new_n19736__,
    new_new_n19737__, new_new_n19738__, new_new_n19739__, new_new_n19740__,
    new_new_n19741__, new_new_n19742__, new_new_n19743__, new_new_n19744__,
    new_new_n19745__, new_new_n19746__, new_new_n19747__, new_new_n19748__,
    new_new_n19749__, new_new_n19750__, new_new_n19751__, new_new_n19752__,
    new_new_n19753__, new_new_n19754__, new_new_n19755__, new_new_n19756__,
    new_new_n19757__, new_new_n19758__, new_new_n19759__, new_new_n19760__,
    new_new_n19761__, new_new_n19762__, new_new_n19763__, new_new_n19764__,
    new_new_n19765__, new_new_n19766__, new_new_n19767__, new_new_n19768__,
    new_new_n19769__, new_new_n19770__, new_new_n19771__, new_new_n19772__,
    new_new_n19773__, new_new_n19774__, new_new_n19775__, new_new_n19776__,
    new_new_n19777__, new_new_n19778__, new_new_n19779__, new_new_n19780__,
    new_new_n19781__, new_new_n19782__, new_new_n19783__, new_new_n19784__,
    new_new_n19785__, new_new_n19786__, new_new_n19787__, new_new_n19788__,
    new_new_n19789__, new_new_n19790__, new_new_n19791__, new_new_n19792__,
    new_new_n19793__, new_new_n19794__, new_new_n19795__, new_new_n19796__,
    new_new_n19797__, new_new_n19798__, new_new_n19799__, new_new_n19800__,
    new_new_n19801__, new_new_n19802__, new_new_n19803__, new_new_n19804__,
    new_new_n19805__, new_new_n19806__, new_new_n19807__, new_new_n19808__,
    new_new_n19809__, new_new_n19810__, new_new_n19811__, new_new_n19812__,
    new_new_n19813__, new_new_n19814__, new_new_n19815__, new_new_n19816__,
    new_new_n19817__, new_new_n19818__, new_new_n19819__, new_new_n19820__,
    new_new_n19821__, new_new_n19822__, new_new_n19823__, new_new_n19824__,
    new_new_n19825__, new_new_n19826__, new_new_n19827__, new_new_n19828__,
    new_new_n19829__, new_new_n19830__, new_new_n19831__, new_new_n19832__,
    new_new_n19833__, new_new_n19834__, new_new_n19835__, new_new_n19836__,
    new_new_n19837__, new_new_n19838__, new_new_n19839__, new_new_n19840__,
    new_new_n19841__, new_new_n19842__, new_new_n19843__, new_new_n19844__,
    new_new_n19845__, new_new_n19846__, new_new_n19847__, new_new_n19848__,
    new_new_n19849__, new_new_n19850__, new_new_n19851__, new_new_n19852__,
    new_new_n19853__, new_new_n19854__, new_new_n19855__, new_new_n19856__,
    new_new_n19857__, new_new_n19858__, new_new_n19859__, new_new_n19860__,
    new_new_n19861__, new_new_n19862__, new_new_n19863__, new_new_n19864__,
    new_new_n19865__, new_new_n19866__, new_new_n19867__, new_new_n19868__,
    new_new_n19869__, new_new_n19870__, new_new_n19871__, new_new_n19872__,
    new_new_n19873__, new_new_n19874__, new_new_n19875__, new_new_n19876__,
    new_new_n19877__, new_new_n19878__, new_new_n19879__, new_new_n19880__,
    new_new_n19881__, new_new_n19882__, new_new_n19883__, new_new_n19884__,
    new_new_n19885__, new_new_n19886__, new_new_n19887__, new_new_n19888__,
    new_new_n19889__, new_new_n19890__, new_new_n19891__, new_new_n19892__,
    new_new_n19893__, new_new_n19894__, new_new_n19895__, new_new_n19896__,
    new_new_n19897__, new_new_n19898__, new_new_n19899__, new_new_n19900__,
    new_new_n19901__, new_new_n19902__, new_new_n19903__, new_new_n19904__,
    new_new_n19905__, new_new_n19906__, new_new_n19907__, new_new_n19908__,
    new_new_n19909__, new_new_n19910__, new_new_n19911__, new_new_n19912__,
    new_new_n19913__, new_new_n19914__, new_new_n19915__, new_new_n19916__,
    new_new_n19917__, new_new_n19918__, new_new_n19919__, new_new_n19920__,
    new_new_n19921__, new_new_n19922__, new_new_n19923__, new_new_n19924__,
    new_new_n19925__, new_new_n19926__, new_new_n19927__, new_new_n19928__,
    new_new_n19929__, new_new_n19930__, new_new_n19931__, new_new_n19932__,
    new_new_n19933__, new_new_n19934__, new_new_n19935__, new_new_n19936__,
    new_new_n19937__, new_new_n19938__, new_new_n19939__, new_new_n19940__,
    new_new_n19941__, new_new_n19942__, new_new_n19943__, new_new_n19944__,
    new_new_n19945__, new_new_n19946__, new_new_n19947__, new_new_n19948__,
    new_new_n19949__, new_new_n19950__, new_new_n19951__, new_new_n19952__,
    new_new_n19953__, new_new_n19954__, new_new_n19955__, new_new_n19956__,
    new_new_n19957__, new_new_n19958__, new_new_n19959__, new_new_n19960__,
    new_new_n19961__, new_new_n19962__, new_new_n19963__, new_new_n19964__,
    new_new_n19965__, new_new_n19966__, new_new_n19967__, new_new_n19968__,
    new_new_n19969__, new_new_n19970__, new_new_n19971__, new_new_n19972__,
    new_new_n19973__, new_new_n19974__, new_new_n19975__, new_new_n19976__,
    new_new_n19977__, new_new_n19978__, new_new_n19979__, new_new_n19980__,
    new_new_n19981__, new_new_n19982__, new_new_n19983__, new_new_n19984__,
    new_new_n19985__, new_new_n19986__, new_new_n19987__, new_new_n19988__,
    new_new_n19989__, new_new_n19990__, new_new_n19991__, new_new_n19992__,
    new_new_n19993__, new_new_n19994__, new_new_n19995__, new_new_n19996__,
    new_new_n19997__, new_new_n19998__, new_new_n19999__, new_new_n20000__,
    new_new_n20001__, new_new_n20002__, new_new_n20003__, new_new_n20004__,
    new_new_n20005__, new_new_n20006__, new_new_n20007__, new_new_n20008__,
    new_new_n20009__, new_new_n20010__, new_new_n20011__, new_new_n20012__,
    new_new_n20013__, new_new_n20014__, new_new_n20015__, new_new_n20016__,
    new_new_n20017__, new_new_n20018__, new_new_n20019__, new_new_n20020__,
    new_new_n20021__, new_new_n20022__, new_new_n20023__, new_new_n20024__,
    new_new_n20025__, new_new_n20026__, new_new_n20027__, new_new_n20028__,
    new_new_n20029__, new_new_n20030__, new_new_n20031__, new_new_n20032__,
    new_new_n20033__, new_new_n20034__, new_new_n20035__, new_new_n20036__,
    new_new_n20037__, new_new_n20038__, new_new_n20039__, new_new_n20040__,
    new_new_n20041__, new_new_n20042__, new_new_n20043__, new_new_n20044__,
    new_new_n20045__, new_new_n20046__, new_new_n20047__, new_new_n20048__,
    new_new_n20049__, new_new_n20050__, new_new_n20051__, new_new_n20052__,
    new_new_n20053__, new_new_n20054__, new_new_n20055__, new_new_n20056__,
    new_new_n20057__, new_new_n20058__, new_new_n20059__, new_new_n20060__,
    new_new_n20061__, new_new_n20062__, new_new_n20063__, new_new_n20064__,
    new_new_n20065__, new_new_n20066__, new_new_n20067__, new_new_n20068__,
    new_new_n20069__, new_new_n20070__, new_new_n20071__, new_new_n20072__,
    new_new_n20073__, new_new_n20074__, new_new_n20075__, new_new_n20076__,
    new_new_n20077__, new_new_n20078__, new_new_n20079__, new_new_n20080__,
    new_new_n20081__, new_new_n20082__, new_new_n20083__, new_new_n20084__,
    new_new_n20085__, new_new_n20086__, new_new_n20087__, new_new_n20088__,
    new_new_n20089__, new_new_n20090__, new_new_n20091__, new_new_n20092__,
    new_new_n20093__, new_new_n20094__, new_new_n20095__, new_new_n20096__,
    new_new_n20097__, new_new_n20098__, new_new_n20099__, new_new_n20100__,
    new_new_n20101__, new_new_n20102__, new_new_n20103__, new_new_n20104__,
    new_new_n20105__, new_new_n20106__, new_new_n20107__, new_new_n20108__,
    new_new_n20109__, new_new_n20110__, new_new_n20111__, new_new_n20112__,
    new_new_n20113__, new_new_n20114__, new_new_n20115__, new_new_n20116__,
    new_new_n20117__, new_new_n20118__, new_new_n20119__, new_new_n20120__,
    new_new_n20121__, new_new_n20122__, new_new_n20123__, new_new_n20124__,
    new_new_n20125__, new_new_n20126__, new_new_n20127__, new_new_n20128__,
    new_new_n20129__, new_new_n20130__, new_new_n20131__, new_new_n20132__,
    new_new_n20133__, new_new_n20134__, new_new_n20135__, new_new_n20136__,
    new_new_n20137__, new_new_n20138__, new_new_n20139__, new_new_n20140__,
    new_new_n20141__, new_new_n20142__, new_new_n20143__, new_new_n20144__,
    new_new_n20145__, new_new_n20146__, new_new_n20147__, new_new_n20148__,
    new_new_n20149__, new_new_n20150__, new_new_n20151__, new_new_n20152__,
    new_new_n20153__, new_new_n20154__, new_new_n20155__, new_new_n20156__,
    new_new_n20157__, new_new_n20158__, new_new_n20159__, new_new_n20160__,
    new_new_n20161__, new_new_n20162__, new_new_n20163__, new_new_n20164__,
    new_new_n20165__, new_new_n20166__, new_new_n20167__, new_new_n20168__,
    new_new_n20169__, new_new_n20170__, new_new_n20171__, new_new_n20172__,
    new_new_n20173__, new_new_n20174__, new_new_n20175__, new_new_n20176__,
    new_new_n20177__, new_new_n20178__, new_new_n20179__, new_new_n20180__,
    new_new_n20181__, new_new_n20182__, new_new_n20183__, new_new_n20184__,
    new_new_n20185__, new_new_n20186__, new_new_n20187__, new_new_n20188__,
    new_new_n20189__, new_new_n20190__, new_new_n20191__, new_new_n20192__,
    new_new_n20193__, new_new_n20194__, new_new_n20195__, new_new_n20196__,
    new_new_n20197__, new_new_n20198__, new_new_n20199__, new_new_n20200__,
    new_new_n20201__, new_new_n20202__, new_new_n20203__, new_new_n20204__,
    new_new_n20205__, new_new_n20206__, new_new_n20207__, new_new_n20208__,
    new_new_n20209__, new_new_n20210__, new_new_n20211__, new_new_n20212__,
    new_new_n20213__, new_new_n20214__, new_new_n20215__, new_new_n20216__,
    new_new_n20217__, new_new_n20218__, new_new_n20219__, new_new_n20220__,
    new_new_n20221__, new_new_n20222__, new_new_n20223__, new_new_n20224__,
    new_new_n20225__, new_new_n20226__, new_new_n20227__, new_new_n20228__,
    new_new_n20229__, new_new_n20230__, new_new_n20231__, new_new_n20232__,
    new_new_n20233__, new_new_n20234__, new_new_n20235__, new_new_n20236__,
    new_new_n20237__, new_new_n20238__, new_new_n20239__, new_new_n20240__,
    new_new_n20241__, new_new_n20242__, new_new_n20243__, new_new_n20244__,
    new_new_n20245__, new_new_n20246__, new_new_n20247__, new_new_n20248__,
    new_new_n20249__, new_new_n20250__, new_new_n20251__, new_new_n20252__,
    new_new_n20253__, new_new_n20254__, new_new_n20255__, new_new_n20256__,
    new_new_n20257__, new_new_n20258__, new_new_n20259__, new_new_n20260__,
    new_new_n20261__, new_new_n20262__, new_new_n20263__, new_new_n20264__,
    new_new_n20265__, new_new_n20266__, new_new_n20267__, new_new_n20268__,
    new_new_n20269__, new_new_n20270__, new_new_n20271__, new_new_n20272__,
    new_new_n20273__, new_new_n20274__, new_new_n20275__, new_new_n20276__,
    new_new_n20277__, new_new_n20278__, new_new_n20279__, new_new_n20280__,
    new_new_n20281__, new_new_n20282__, new_new_n20283__, new_new_n20284__,
    new_new_n20285__, new_new_n20286__, new_new_n20287__, new_new_n20288__,
    new_new_n20289__, new_new_n20290__, new_new_n20291__, new_new_n20292__,
    new_new_n20293__, new_new_n20294__, new_new_n20295__, new_new_n20296__,
    new_new_n20297__, new_new_n20298__, new_new_n20299__, new_new_n20300__,
    new_new_n20301__, new_new_n20302__, new_new_n20303__, new_new_n20304__,
    new_new_n20305__, new_new_n20306__, new_new_n20307__, new_new_n20308__,
    new_new_n20309__, new_new_n20310__, new_new_n20311__, new_new_n20312__,
    new_new_n20313__, new_new_n20314__, new_new_n20315__, new_new_n20316__,
    new_new_n20317__, new_new_n20318__, new_new_n20319__, new_new_n20320__,
    new_new_n20321__, new_new_n20322__, new_new_n20323__, new_new_n20324__,
    new_new_n20325__, new_new_n20326__, new_new_n20327__, new_new_n20328__,
    new_new_n20329__, new_new_n20330__, new_new_n20331__, new_new_n20332__,
    new_new_n20333__, new_new_n20334__, new_new_n20335__, new_new_n20336__,
    new_new_n20337__, new_new_n20338__, new_new_n20339__, new_new_n20340__,
    new_new_n20341__, new_new_n20342__, new_new_n20343__, new_new_n20344__,
    new_new_n20345__, new_new_n20346__, new_new_n20347__, new_new_n20348__,
    new_new_n20349__, new_new_n20350__, new_new_n20351__, new_new_n20352__,
    new_new_n20353__, new_new_n20354__, new_new_n20355__, new_new_n20356__,
    new_new_n20357__, new_new_n20358__, new_new_n20359__, new_new_n20360__,
    new_new_n20361__, new_new_n20362__, new_new_n20363__, new_new_n20364__,
    new_new_n20365__, new_new_n20366__, new_new_n20367__, new_new_n20368__,
    new_new_n20369__, new_new_n20370__, new_new_n20371__, new_new_n20372__,
    new_new_n20373__, new_new_n20374__, new_new_n20375__, new_new_n20376__,
    new_new_n20377__, new_new_n20378__, new_new_n20379__, new_new_n20380__,
    new_new_n20381__, new_new_n20382__, new_new_n20383__, new_new_n20384__,
    new_new_n20385__, new_new_n20386__, new_new_n20387__, new_new_n20388__,
    new_new_n20389__, new_new_n20390__, new_new_n20391__, new_new_n20392__,
    new_new_n20393__, new_new_n20394__, new_new_n20395__, new_new_n20396__,
    new_new_n20397__, new_new_n20398__, new_new_n20399__, new_new_n20400__,
    new_new_n20401__, new_new_n20402__, new_new_n20403__, new_new_n20404__,
    new_new_n20405__, new_new_n20406__, new_new_n20407__, new_new_n20408__,
    new_new_n20409__, new_new_n20410__, new_new_n20411__, new_new_n20412__,
    new_new_n20413__, new_new_n20414__, new_new_n20415__, new_new_n20416__,
    new_new_n20417__, new_new_n20418__, new_new_n20419__, new_new_n20420__,
    new_new_n20421__, new_new_n20422__, new_new_n20423__, new_new_n20424__,
    new_new_n20425__, new_new_n20426__, new_new_n20427__, new_new_n20428__,
    new_new_n20429__, new_new_n20430__, new_new_n20431__, new_new_n20432__,
    new_new_n20433__, new_new_n20434__, new_new_n20435__, new_new_n20436__,
    new_new_n20437__, new_new_n20438__, new_new_n20439__, new_new_n20440__,
    new_new_n20441__, new_new_n20442__, new_new_n20443__, new_new_n20444__,
    new_new_n20445__, new_new_n20446__, new_new_n20447__, new_new_n20448__,
    new_new_n20449__, new_new_n20450__, new_new_n20451__, new_new_n20452__,
    new_new_n20453__, new_new_n20454__, new_new_n20455__, new_new_n20456__,
    new_new_n20457__, new_new_n20458__, new_new_n20459__, new_new_n20460__,
    new_new_n20461__, new_new_n20462__, new_new_n20463__, new_new_n20464__,
    new_new_n20465__, new_new_n20466__, new_new_n20467__, new_new_n20468__,
    new_new_n20469__, new_new_n20470__, new_new_n20471__, new_new_n20472__,
    new_new_n20473__, new_new_n20474__, new_new_n20475__, new_new_n20476__,
    new_new_n20477__, new_new_n20478__, new_new_n20479__, new_new_n20480__,
    new_new_n20481__, new_new_n20482__, new_new_n20483__, new_new_n20484__,
    new_new_n20485__, new_new_n20486__, new_new_n20487__, new_new_n20488__,
    new_new_n20489__, new_new_n20490__, new_new_n20491__, new_new_n20492__,
    new_new_n20493__, new_new_n20494__, new_new_n20495__, new_new_n20496__,
    new_new_n20497__, new_new_n20498__, new_new_n20499__, new_new_n20500__,
    new_new_n20501__, new_new_n20502__, new_new_n20503__, new_new_n20504__,
    new_new_n20505__, new_new_n20506__, new_new_n20507__, new_new_n20508__,
    new_new_n20509__, new_new_n20510__, new_new_n20511__, new_new_n20512__,
    new_new_n20513__, new_new_n20514__, new_new_n20515__, new_new_n20516__,
    new_new_n20517__, new_new_n20518__, new_new_n20519__, new_new_n20520__,
    new_new_n20521__, new_new_n20522__, new_new_n20523__, new_new_n20524__,
    new_new_n20525__, new_new_n20526__, new_new_n20527__, new_new_n20528__,
    new_new_n20529__, new_new_n20530__, new_new_n20531__, new_new_n20532__,
    new_new_n20533__, new_new_n20534__, new_new_n20535__, new_new_n20536__,
    new_new_n20537__, new_new_n20538__, new_new_n20539__, new_new_n20540__,
    new_new_n20541__, new_new_n20542__, new_new_n20543__, new_new_n20544__,
    new_new_n20545__, new_new_n20546__, new_new_n20547__, new_new_n20548__,
    new_new_n20549__, new_new_n20550__, new_new_n20551__, new_new_n20552__,
    new_new_n20553__, new_new_n20554__, new_new_n20555__, new_new_n20556__,
    new_new_n20557__, new_new_n20558__, new_new_n20559__, new_new_n20560__,
    new_new_n20561__, new_new_n20562__, new_new_n20563__, new_new_n20564__,
    new_new_n20565__, new_new_n20566__, new_new_n20567__, new_new_n20568__,
    new_new_n20569__, new_new_n20570__, new_new_n20571__, new_new_n20572__,
    new_new_n20573__, new_new_n20574__, new_new_n20575__, new_new_n20576__,
    new_new_n20577__, new_new_n20578__, new_new_n20579__, new_new_n20580__,
    new_new_n20581__, new_new_n20582__, new_new_n20583__, new_new_n20584__,
    new_new_n20585__, new_new_n20586__, new_new_n20587__, new_new_n20588__,
    new_new_n20589__, new_new_n20590__, new_new_n20591__, new_new_n20592__,
    new_new_n20593__, new_new_n20594__, new_new_n20595__, new_new_n20596__,
    new_new_n20597__, new_new_n20598__, new_new_n20599__, new_new_n20600__,
    new_new_n20601__, new_new_n20602__, new_new_n20603__, new_new_n20604__,
    new_new_n20605__, new_new_n20606__, new_new_n20607__, new_new_n20608__,
    new_new_n20609__, new_new_n20610__, new_new_n20611__, new_new_n20612__,
    new_new_n20613__, new_new_n20614__, new_new_n20615__, new_new_n20616__,
    new_new_n20617__, new_new_n20618__, new_new_n20619__, new_new_n20620__,
    new_new_n20621__, new_new_n20622__, new_new_n20623__, new_new_n20624__,
    new_new_n20625__, new_new_n20626__, new_new_n20627__, new_new_n20628__,
    new_new_n20629__, new_new_n20630__, new_new_n20631__, new_new_n20632__,
    new_new_n20633__, new_new_n20634__, new_new_n20635__, new_new_n20636__,
    new_new_n20637__, new_new_n20638__, new_new_n20639__, new_new_n20640__,
    new_new_n20641__, new_new_n20642__, new_new_n20643__, new_new_n20644__,
    new_new_n20645__, new_new_n20646__, new_new_n20647__, new_new_n20648__,
    new_new_n20649__, new_new_n20650__, new_new_n20651__, new_new_n20652__,
    new_new_n20653__, new_new_n20654__, new_new_n20655__, new_new_n20656__,
    new_new_n20657__, new_new_n20658__, new_new_n20659__, new_new_n20660__,
    new_new_n20661__, new_new_n20662__, new_new_n20663__, new_new_n20664__,
    new_new_n20665__, new_new_n20666__, new_new_n20667__, new_new_n20668__,
    new_new_n20669__, new_new_n20670__, new_new_n20671__, new_new_n20672__,
    new_new_n20673__, new_new_n20674__, new_new_n20675__, new_new_n20676__,
    new_new_n20677__, new_new_n20678__, new_new_n20679__, new_new_n20680__,
    new_new_n20681__, new_new_n20682__, new_new_n20683__, new_new_n20684__,
    new_new_n20685__, new_new_n20686__, new_new_n20687__, new_new_n20688__,
    new_new_n20689__, new_new_n20690__, new_new_n20691__, new_new_n20692__,
    new_new_n20693__, new_new_n20694__, new_new_n20695__, new_new_n20696__,
    new_new_n20697__, new_new_n20698__, new_new_n20699__, new_new_n20700__,
    new_new_n20701__, new_new_n20702__, new_new_n20703__, new_new_n20704__,
    new_new_n20705__, new_new_n20706__, new_new_n20707__, new_new_n20708__,
    new_new_n20709__, new_new_n20710__, new_new_n20711__, new_new_n20712__,
    new_new_n20713__, new_new_n20714__, new_new_n20715__, new_new_n20716__,
    new_new_n20717__, new_new_n20718__, new_new_n20719__, new_new_n20720__,
    new_new_n20721__, new_new_n20722__, new_new_n20723__, new_new_n20724__,
    new_new_n20725__, new_new_n20726__, new_new_n20727__, new_new_n20728__,
    new_new_n20729__, new_new_n20730__, new_new_n20731__, new_new_n20732__,
    new_new_n20733__, new_new_n20734__, new_new_n20735__, new_new_n20736__,
    new_new_n20737__, new_new_n20738__, new_new_n20739__, new_new_n20740__,
    new_new_n20741__, new_new_n20742__, new_new_n20743__, new_new_n20744__,
    new_new_n20745__, new_new_n20746__, new_new_n20747__, new_new_n20748__,
    new_new_n20749__, new_new_n20750__, new_new_n20751__, new_new_n20752__,
    new_new_n20753__, new_new_n20754__, new_new_n20755__, new_new_n20756__,
    new_new_n20757__, new_new_n20758__, new_new_n20759__, new_new_n20760__,
    new_new_n20761__, new_new_n20762__, new_new_n20763__, new_new_n20764__,
    new_new_n20765__, new_new_n20766__, new_new_n20767__, new_new_n20768__,
    new_new_n20769__, new_new_n20770__, new_new_n20771__, new_new_n20772__,
    new_new_n20773__, new_new_n20774__, new_new_n20775__, new_new_n20776__,
    new_new_n20777__, new_new_n20778__, new_new_n20779__, new_new_n20780__,
    new_new_n20781__, new_new_n20782__, new_new_n20783__, new_new_n20784__,
    new_new_n20785__, new_new_n20786__, new_new_n20787__, new_new_n20788__,
    new_new_n20789__, new_new_n20790__, new_new_n20791__, new_new_n20792__,
    new_new_n20793__, new_new_n20794__, new_new_n20795__, new_new_n20796__,
    new_new_n20797__, new_new_n20798__, new_new_n20799__, new_new_n20800__,
    new_new_n20801__, new_new_n20802__, new_new_n20803__, new_new_n20804__,
    new_new_n20805__, new_new_n20806__, new_new_n20807__, new_new_n20808__,
    new_new_n20809__, new_new_n20810__, new_new_n20811__, new_new_n20812__,
    new_new_n20813__, new_new_n20814__, new_new_n20815__, new_new_n20816__,
    new_new_n20817__, new_new_n20818__, new_new_n20819__, new_new_n20820__,
    new_new_n20821__, new_new_n20822__, new_new_n20823__, new_new_n20824__,
    new_new_n20825__, new_new_n20826__, new_new_n20827__, new_new_n20828__,
    new_new_n20829__, new_new_n20830__, new_new_n20831__, new_new_n20832__,
    new_new_n20833__, new_new_n20834__, new_new_n20835__, new_new_n20836__,
    new_new_n20837__, new_new_n20838__, new_new_n20839__, new_new_n20840__,
    new_new_n20841__, new_new_n20842__, new_new_n20843__, new_new_n20844__,
    new_new_n20845__, new_new_n20846__, new_new_n20847__, new_new_n20848__,
    new_new_n20849__, new_new_n20850__, new_new_n20851__, new_new_n20852__,
    new_new_n20853__, new_new_n20854__, new_new_n20855__, new_new_n20856__,
    new_new_n20857__, new_new_n20858__, new_new_n20859__, new_new_n20860__,
    new_new_n20861__, new_new_n20862__, new_new_n20863__, new_new_n20864__,
    new_new_n20865__, new_new_n20866__, new_new_n20867__, new_new_n20868__,
    new_new_n20869__, new_new_n20870__, new_new_n20871__, new_new_n20872__,
    new_new_n20873__, new_new_n20874__, new_new_n20875__, new_new_n20876__,
    new_new_n20877__, new_new_n20878__, new_new_n20879__, new_new_n20880__,
    new_new_n20881__, new_new_n20882__, new_new_n20883__, new_new_n20884__,
    new_new_n20885__, new_new_n20886__, new_new_n20887__, new_new_n20888__,
    new_new_n20889__, new_new_n20890__, new_new_n20891__, new_new_n20892__,
    new_new_n20893__, new_new_n20894__, new_new_n20895__, new_new_n20896__,
    new_new_n20897__, new_new_n20898__, new_new_n20899__, new_new_n20900__,
    new_new_n20901__, new_new_n20902__, new_new_n20903__, new_new_n20904__,
    new_new_n20905__, new_new_n20906__, new_new_n20907__, new_new_n20908__,
    new_new_n20909__, new_new_n20910__, new_new_n20911__, new_new_n20912__,
    new_new_n20913__, new_new_n20914__, new_new_n20915__, new_new_n20916__,
    new_new_n20917__, new_new_n20918__, new_new_n20919__, new_new_n20920__,
    new_new_n20921__, new_new_n20922__, new_new_n20923__, new_new_n20924__,
    new_new_n20925__, new_new_n20926__, new_new_n20927__, new_new_n20928__,
    new_new_n20929__, new_new_n20930__, new_new_n20931__, new_new_n20932__,
    new_new_n20933__, new_new_n20934__, new_new_n20935__, new_new_n20936__,
    new_new_n20937__, new_new_n20938__, new_new_n20939__, new_new_n20940__,
    new_new_n20941__, new_new_n20942__, new_new_n20943__, new_new_n20944__,
    new_new_n20945__, new_new_n20946__, new_new_n20947__, new_new_n20948__,
    new_new_n20949__, new_new_n20950__, new_new_n20951__, new_new_n20952__,
    new_new_n20953__, new_new_n20954__, new_new_n20955__, new_new_n20956__,
    new_new_n20957__, new_new_n20958__, new_new_n20959__, new_new_n20960__,
    new_new_n20961__, new_new_n20962__, new_new_n20963__, new_new_n20964__,
    new_new_n20965__, new_new_n20966__, new_new_n20967__, new_new_n20968__,
    new_new_n20969__, new_new_n20970__, new_new_n20971__, new_new_n20972__,
    new_new_n20973__, new_new_n20974__, new_new_n20975__, new_new_n20976__,
    new_new_n20977__, new_new_n20978__, new_new_n20979__, new_new_n20980__,
    new_new_n20981__, new_new_n20982__, new_new_n20983__, new_new_n20984__,
    new_new_n20985__, new_new_n20986__, new_new_n20987__, new_new_n20988__,
    new_new_n20989__, new_new_n20990__, new_new_n20991__, new_new_n20992__,
    new_new_n20993__, new_new_n20994__, new_new_n20995__, new_new_n20996__,
    new_new_n20997__, new_new_n20998__, new_new_n20999__, new_new_n21000__,
    new_new_n21001__, new_new_n21002__, new_new_n21003__, new_new_n21004__,
    new_new_n21005__, new_new_n21006__, new_new_n21007__, new_new_n21008__,
    new_new_n21009__, new_new_n21010__, new_new_n21011__, new_new_n21012__,
    new_new_n21013__, new_new_n21014__, new_new_n21015__, new_new_n21016__,
    new_new_n21017__, new_new_n21018__, new_new_n21019__, new_new_n21020__,
    new_new_n21021__, new_new_n21022__, new_new_n21023__, new_new_n21024__,
    new_new_n21025__, new_new_n21026__, new_new_n21027__, new_new_n21028__,
    new_new_n21029__, new_new_n21030__, new_new_n21031__, new_new_n21032__,
    new_new_n21033__, new_new_n21034__, new_new_n21035__, new_new_n21036__,
    new_new_n21037__, new_new_n21038__, new_new_n21039__, new_new_n21040__,
    new_new_n21041__, new_new_n21042__, new_new_n21043__, new_new_n21044__,
    new_new_n21045__, new_new_n21046__, new_new_n21047__, new_new_n21048__,
    new_new_n21049__, new_new_n21050__, new_new_n21051__, new_new_n21052__,
    new_new_n21053__, new_new_n21054__, new_new_n21055__, new_new_n21056__,
    new_new_n21057__, new_new_n21058__, new_new_n21059__, new_new_n21060__,
    new_new_n21061__, new_new_n21062__, new_new_n21063__, new_new_n21064__,
    new_new_n21065__, new_new_n21066__, new_new_n21067__, new_new_n21068__,
    new_new_n21069__, new_new_n21070__, new_new_n21071__, new_new_n21072__,
    new_new_n21073__, new_new_n21074__, new_new_n21075__, new_new_n21076__,
    new_new_n21077__, new_new_n21078__, new_new_n21079__, new_new_n21080__,
    new_new_n21081__, new_new_n21082__, new_new_n21083__, new_new_n21084__,
    new_new_n21085__, new_new_n21086__, new_new_n21087__, new_new_n21088__,
    new_new_n21089__, new_new_n21090__, new_new_n21091__, new_new_n21092__,
    new_new_n21093__, new_new_n21094__, new_new_n21095__, new_new_n21096__,
    new_new_n21097__, new_new_n21098__, new_new_n21099__, new_new_n21100__,
    new_new_n21101__, new_new_n21102__, new_new_n21103__, new_new_n21104__,
    new_new_n21105__, new_new_n21106__, new_new_n21107__, new_new_n21108__,
    new_new_n21109__, new_new_n21110__, new_new_n21111__, new_new_n21112__,
    new_new_n21113__, new_new_n21114__, new_new_n21115__, new_new_n21116__,
    new_new_n21117__, new_new_n21118__, new_new_n21119__, new_new_n21120__,
    new_new_n21121__, new_new_n21122__, new_new_n21123__, new_new_n21124__,
    new_new_n21125__, new_new_n21126__, new_new_n21127__, new_new_n21128__,
    new_new_n21129__, new_new_n21130__, new_new_n21131__, new_new_n21132__,
    new_new_n21133__, new_new_n21134__, new_new_n21135__, new_new_n21136__,
    new_new_n21137__, new_new_n21138__, new_new_n21139__, new_new_n21140__,
    new_new_n21141__, new_new_n21142__, new_new_n21143__, new_new_n21144__,
    new_new_n21145__, new_new_n21146__, new_new_n21147__, new_new_n21148__,
    new_new_n21149__, new_new_n21150__, new_new_n21151__, new_new_n21152__,
    new_new_n21153__, new_new_n21154__, new_new_n21155__, new_new_n21156__,
    new_new_n21157__, new_new_n21158__, new_new_n21159__, new_new_n21160__,
    new_new_n21161__, new_new_n21162__, new_new_n21163__, new_new_n21164__,
    new_new_n21165__, new_new_n21166__, new_new_n21167__, new_new_n21168__,
    new_new_n21169__, new_new_n21170__, new_new_n21171__, new_new_n21172__,
    new_new_n21173__, new_new_n21174__, new_new_n21175__, new_new_n21176__,
    new_new_n21177__, new_new_n21178__, new_new_n21179__, new_new_n21180__,
    new_new_n21181__, new_new_n21182__, new_new_n21183__, new_new_n21184__,
    new_new_n21185__, new_new_n21186__, new_new_n21187__, new_new_n21188__,
    new_new_n21189__, new_new_n21190__, new_new_n21191__, new_new_n21192__,
    new_new_n21193__, new_new_n21194__, new_new_n21195__, new_new_n21196__,
    new_new_n21197__, new_new_n21198__, new_new_n21199__, new_new_n21200__,
    new_new_n21201__, new_new_n21202__, new_new_n21203__, new_new_n21204__,
    new_new_n21205__, new_new_n21206__, new_new_n21207__, new_new_n21208__,
    new_new_n21209__, new_new_n21210__, new_new_n21211__, new_new_n21212__,
    new_new_n21213__, new_new_n21214__, new_new_n21215__, new_new_n21216__,
    new_new_n21217__, new_new_n21218__, new_new_n21219__, new_new_n21220__,
    new_new_n21221__, new_new_n21222__, new_new_n21223__, new_new_n21224__,
    new_new_n21225__, new_new_n21226__, new_new_n21227__, new_new_n21228__,
    new_new_n21229__, new_new_n21230__, new_new_n21231__, new_new_n21232__,
    new_new_n21233__, new_new_n21234__, new_new_n21235__, new_new_n21236__,
    new_new_n21237__, new_new_n21238__, new_new_n21239__, new_new_n21240__,
    new_new_n21241__, new_new_n21242__, new_new_n21243__, new_new_n21244__,
    new_new_n21245__, new_new_n21246__, new_new_n21247__, new_new_n21248__,
    new_new_n21249__, new_new_n21250__, new_new_n21251__, new_new_n21252__,
    new_new_n21253__, new_new_n21254__, new_new_n21255__, new_new_n21256__,
    new_new_n21257__, new_new_n21258__, new_new_n21259__, new_new_n21260__,
    new_new_n21261__, new_new_n21262__, new_new_n21263__, new_new_n21264__,
    new_new_n21265__, new_new_n21266__, new_new_n21267__, new_new_n21268__,
    new_new_n21269__, new_new_n21270__, new_new_n21271__, new_new_n21272__,
    new_new_n21273__, new_new_n21274__, new_new_n21275__, new_new_n21276__,
    new_new_n21277__, new_new_n21278__, new_new_n21279__, new_new_n21280__,
    new_new_n21281__, new_new_n21282__, new_new_n21283__, new_new_n21284__,
    new_new_n21285__, new_new_n21286__, new_new_n21287__, new_new_n21288__,
    new_new_n21289__, new_new_n21290__, new_new_n21291__, new_new_n21292__,
    new_new_n21293__, new_new_n21294__, new_new_n21295__, new_new_n21296__,
    new_new_n21297__, new_new_n21298__, new_new_n21299__, new_new_n21300__,
    new_new_n21301__, new_new_n21302__, new_new_n21303__, new_new_n21304__,
    new_new_n21305__, new_new_n21306__, new_new_n21307__, new_new_n21308__,
    new_new_n21309__, new_new_n21310__, new_new_n21311__, new_new_n21312__,
    new_new_n21313__, new_new_n21314__, new_new_n21315__, new_new_n21316__,
    new_new_n21317__, new_new_n21318__, new_new_n21319__, new_new_n21320__,
    new_new_n21321__, new_new_n21322__, new_new_n21323__, new_new_n21324__,
    new_new_n21325__, new_new_n21326__, new_new_n21327__, new_new_n21328__,
    new_new_n21329__, new_new_n21330__, new_new_n21331__, new_new_n21332__,
    new_new_n21333__, new_new_n21334__, new_new_n21335__, new_new_n21336__,
    new_new_n21337__, new_new_n21338__, new_new_n21339__, new_new_n21340__,
    new_new_n21341__, new_new_n21342__, new_new_n21343__, new_new_n21344__,
    new_new_n21345__, new_new_n21346__, new_new_n21347__, new_new_n21348__,
    new_new_n21349__, new_new_n21350__, new_new_n21351__, new_new_n21352__,
    new_new_n21353__, new_new_n21354__, new_new_n21355__, new_new_n21356__,
    new_new_n21357__, new_new_n21358__, new_new_n21359__, new_new_n21360__,
    new_new_n21361__, new_new_n21362__, new_new_n21363__, new_new_n21364__,
    new_new_n21365__, new_new_n21366__, new_new_n21367__, new_new_n21368__,
    new_new_n21369__, new_new_n21370__, new_new_n21371__, new_new_n21372__,
    new_new_n21373__, new_new_n21374__, new_new_n21375__, new_new_n21376__,
    new_new_n21377__, new_new_n21378__, new_new_n21379__, new_new_n21380__,
    new_new_n21381__, new_new_n21382__, new_new_n21383__, new_new_n21384__,
    new_new_n21385__, new_new_n21386__, new_new_n21387__, new_new_n21388__,
    new_new_n21389__, new_new_n21390__, new_new_n21391__, new_new_n21392__,
    new_new_n21393__, new_new_n21394__, new_new_n21395__, new_new_n21396__,
    new_new_n21397__, new_new_n21398__, new_new_n21399__, new_new_n21400__,
    new_new_n21401__, new_new_n21402__, new_new_n21403__, new_new_n21404__,
    new_new_n21405__, new_new_n21406__, new_new_n21407__, new_new_n21408__,
    new_new_n21409__, new_new_n21410__, new_new_n21411__, new_new_n21412__,
    new_new_n21413__, new_new_n21414__, new_new_n21415__, new_new_n21416__,
    new_new_n21417__, new_new_n21418__, new_new_n21419__, new_new_n21420__,
    new_new_n21421__, new_new_n21422__, new_new_n21423__, new_new_n21424__,
    new_new_n21425__, new_new_n21426__, new_new_n21427__, new_new_n21428__,
    new_new_n21429__, new_new_n21430__, new_new_n21431__, new_new_n21432__,
    new_new_n21433__, new_new_n21434__, new_new_n21435__, new_new_n21436__,
    new_new_n21437__, new_new_n21438__, new_new_n21439__, new_new_n21440__,
    new_new_n21441__, new_new_n21442__, new_new_n21443__, new_new_n21444__,
    new_new_n21445__, new_new_n21446__, new_new_n21447__, new_new_n21448__,
    new_new_n21449__, new_new_n21450__, new_new_n21451__, new_new_n21452__,
    new_new_n21453__, new_new_n21454__, new_new_n21455__, new_new_n21456__,
    new_new_n21457__, new_new_n21458__, new_new_n21459__, new_new_n21460__,
    new_new_n21461__, new_new_n21462__, new_new_n21463__, new_new_n21464__,
    new_new_n21465__, new_new_n21466__, new_new_n21467__, new_new_n21468__,
    new_new_n21469__, new_new_n21470__, new_new_n21471__, new_new_n21472__,
    new_new_n21473__, new_new_n21474__, new_new_n21475__, new_new_n21476__,
    new_new_n21477__, new_new_n21478__, new_new_n21479__, new_new_n21480__,
    new_new_n21481__, new_new_n21482__, new_new_n21483__, new_new_n21484__,
    new_new_n21485__, new_new_n21486__, new_new_n21487__, new_new_n21488__,
    new_new_n21489__, new_new_n21490__, new_new_n21491__, new_new_n21492__,
    new_new_n21493__, new_new_n21494__, new_new_n21495__, new_new_n21496__,
    new_new_n21497__, new_new_n21498__, new_new_n21499__, new_new_n21500__,
    new_new_n21501__, new_new_n21502__, new_new_n21503__, new_new_n21504__,
    new_new_n21505__, new_new_n21506__, new_new_n21507__, new_new_n21508__,
    new_new_n21509__, new_new_n21510__, new_new_n21511__, new_new_n21512__,
    new_new_n21513__, new_new_n21514__, new_new_n21515__, new_new_n21516__,
    new_new_n21517__, new_new_n21518__, new_new_n21519__, new_new_n21520__,
    new_new_n21521__, new_new_n21522__, new_new_n21523__, new_new_n21524__,
    new_new_n21525__, new_new_n21526__, new_new_n21527__, new_new_n21528__,
    new_new_n21529__, new_new_n21530__, new_new_n21531__, new_new_n21532__,
    new_new_n21533__, new_new_n21534__, new_new_n21535__, new_new_n21536__,
    new_new_n21537__, new_new_n21538__, new_new_n21539__, new_new_n21540__,
    new_new_n21541__, new_new_n21542__, new_new_n21543__, new_new_n21544__,
    new_new_n21545__, new_new_n21546__, new_new_n21547__, new_new_n21548__,
    new_new_n21549__, new_new_n21550__, new_new_n21551__, new_new_n21552__,
    new_new_n21553__, new_new_n21554__, new_new_n21555__, new_new_n21556__,
    new_new_n21557__, new_new_n21558__, new_new_n21559__, new_new_n21560__,
    new_new_n21561__, new_new_n21562__, new_new_n21563__, new_new_n21564__,
    new_new_n21565__, new_new_n21566__, new_new_n21567__, new_new_n21568__,
    new_new_n21569__, new_new_n21570__, new_new_n21571__, new_new_n21572__,
    new_new_n21573__, new_new_n21574__, new_new_n21575__, new_new_n21576__,
    new_new_n21577__, new_new_n21578__, new_new_n21579__, new_new_n21580__,
    new_new_n21581__, new_new_n21582__, new_new_n21583__, new_new_n21584__,
    new_new_n21585__, new_new_n21586__, new_new_n21587__, new_new_n21588__,
    new_new_n21589__, new_new_n21590__, new_new_n21591__, new_new_n21592__,
    new_new_n21593__, new_new_n21594__, new_new_n21595__, new_new_n21596__,
    new_new_n21597__, new_new_n21598__, new_new_n21599__, new_new_n21600__,
    new_new_n21601__, new_new_n21602__, new_new_n21603__, new_new_n21604__,
    new_new_n21605__, new_new_n21606__, new_new_n21607__, new_new_n21608__,
    new_new_n21609__, new_new_n21610__, new_new_n21611__, new_new_n21612__,
    new_new_n21613__, new_new_n21614__, new_new_n21615__, new_new_n21616__,
    new_new_n21617__, new_new_n21618__, new_new_n21619__, new_new_n21620__,
    new_new_n21621__, new_new_n21622__, new_new_n21623__, new_new_n21624__,
    new_new_n21625__, new_new_n21626__, new_new_n21627__, new_new_n21628__,
    new_new_n21629__, new_new_n21630__, new_new_n21631__, new_new_n21632__,
    new_new_n21633__, new_new_n21634__, new_new_n21635__, new_new_n21636__,
    new_new_n21637__, new_new_n21638__, new_new_n21639__, new_new_n21640__,
    new_new_n21641__, new_new_n21642__, new_new_n21643__, new_new_n21644__,
    new_new_n21645__, new_new_n21646__, new_new_n21647__, new_new_n21648__,
    new_new_n21649__, new_new_n21650__, new_new_n21651__, new_new_n21652__,
    new_new_n21653__, new_new_n21654__, new_new_n21655__, new_new_n21656__,
    new_new_n21657__, new_new_n21658__, new_new_n21659__, new_new_n21660__,
    new_new_n21661__, new_new_n21662__, new_new_n21663__, new_new_n21664__,
    new_new_n21665__, new_new_n21666__, new_new_n21667__, new_new_n21668__,
    new_new_n21669__, new_new_n21670__, new_new_n21671__, new_new_n21672__,
    new_new_n21673__, new_new_n21674__, new_new_n21675__, new_new_n21676__,
    new_new_n21677__, new_new_n21678__, new_new_n21679__, new_new_n21680__,
    new_new_n21681__, new_new_n21682__, new_new_n21683__, new_new_n21684__,
    new_new_n21685__, new_new_n21686__, new_new_n21687__, new_new_n21688__,
    new_new_n21689__, new_new_n21690__, new_new_n21691__, new_new_n21692__,
    new_new_n21693__, new_new_n21694__, new_new_n21695__, new_new_n21696__,
    new_new_n21697__, new_new_n21698__, new_new_n21699__, new_new_n21700__,
    new_new_n21701__, new_new_n21702__, new_new_n21703__, new_new_n21704__,
    new_new_n21705__, new_new_n21706__, new_new_n21707__, new_new_n21708__,
    new_new_n21709__, new_new_n21710__, new_new_n21711__, new_new_n21712__,
    new_new_n21713__, new_new_n21714__, new_new_n21715__, new_new_n21716__,
    new_new_n21717__, new_new_n21718__, new_new_n21719__, new_new_n21720__,
    new_new_n21721__, new_new_n21722__, new_new_n21723__, new_new_n21724__,
    new_new_n21725__, new_new_n21726__, new_new_n21727__, new_new_n21728__,
    new_new_n21729__, new_new_n21730__, new_new_n21731__, new_new_n21732__,
    new_new_n21733__, new_new_n21734__, new_new_n21735__, new_new_n21736__,
    new_new_n21737__, new_new_n21738__, new_new_n21739__, new_new_n21740__,
    new_new_n21741__, new_new_n21742__, new_new_n21743__, new_new_n21744__,
    new_new_n21745__, new_new_n21746__, new_new_n21747__, new_new_n21748__,
    new_new_n21749__, new_new_n21750__, new_new_n21751__, new_new_n21752__,
    new_new_n21753__, new_new_n21754__, new_new_n21755__, new_new_n21756__,
    new_new_n21757__, new_new_n21758__, new_new_n21759__, new_new_n21760__,
    new_new_n21761__, new_new_n21762__, new_new_n21763__, new_new_n21764__,
    new_new_n21765__, new_new_n21766__, new_new_n21767__, new_new_n21768__,
    new_new_n21769__, new_new_n21770__, new_new_n21771__, new_new_n21772__,
    new_new_n21773__, new_new_n21774__, new_new_n21775__, new_new_n21776__,
    new_new_n21777__, new_new_n21778__, new_new_n21779__, new_new_n21780__,
    new_new_n21781__, new_new_n21782__, new_new_n21783__, new_new_n21784__,
    new_new_n21785__, new_new_n21786__, new_new_n21787__, new_new_n21788__,
    new_new_n21789__, new_new_n21790__, new_new_n21791__, new_new_n21792__,
    new_new_n21793__, new_new_n21794__, new_new_n21795__, new_new_n21796__,
    new_new_n21797__, new_new_n21798__, new_new_n21799__, new_new_n21800__,
    new_new_n21801__, new_new_n21802__, new_new_n21803__, new_new_n21804__,
    new_new_n21805__, new_new_n21806__, new_new_n21807__, new_new_n21808__,
    new_new_n21809__, new_new_n21810__, new_new_n21811__, new_new_n21812__,
    new_new_n21813__, new_new_n21814__, new_new_n21815__, new_new_n21816__,
    new_new_n21817__, new_new_n21818__, new_new_n21819__, new_new_n21820__,
    new_new_n21821__, new_new_n21822__, new_new_n21823__, new_new_n21824__,
    new_new_n21825__, new_new_n21826__, new_new_n21827__, new_new_n21828__,
    new_new_n21829__, new_new_n21830__, new_new_n21831__, new_new_n21832__,
    new_new_n21833__, new_new_n21834__, new_new_n21835__, new_new_n21836__,
    new_new_n21837__, new_new_n21838__, new_new_n21839__, new_new_n21840__,
    new_new_n21841__, new_new_n21842__, new_new_n21843__, new_new_n21844__,
    new_new_n21845__, new_new_n21846__, new_new_n21847__, new_new_n21848__,
    new_new_n21849__, new_new_n21850__, new_new_n21851__, new_new_n21852__,
    new_new_n21853__, new_new_n21854__, new_new_n21855__, new_new_n21856__,
    new_new_n21857__, new_new_n21858__, new_new_n21859__, new_new_n21860__,
    new_new_n21861__, new_new_n21862__, new_new_n21863__, new_new_n21864__,
    new_new_n21865__, new_new_n21866__, new_new_n21867__, new_new_n21868__,
    new_new_n21869__, new_new_n21870__, new_new_n21871__, new_new_n21872__,
    new_new_n21873__, new_new_n21874__, new_new_n21875__, new_new_n21876__,
    new_new_n21877__, new_new_n21878__, new_new_n21879__, new_new_n21880__,
    new_new_n21881__, new_new_n21882__, new_new_n21883__, new_new_n21884__,
    new_new_n21885__, new_new_n21886__, new_new_n21887__, new_new_n21888__,
    new_new_n21889__, new_new_n21890__, new_new_n21891__, new_new_n21892__,
    new_new_n21893__, new_new_n21894__, new_new_n21895__, new_new_n21896__,
    new_new_n21897__, new_new_n21898__, new_new_n21899__, new_new_n21900__,
    new_new_n21901__, new_new_n21902__, new_new_n21903__, new_new_n21904__,
    new_new_n21905__, new_new_n21906__, new_new_n21907__, new_new_n21908__,
    new_new_n21909__, new_new_n21910__, new_new_n21911__, new_new_n21912__,
    new_new_n21913__, new_new_n21914__, new_new_n21915__, new_new_n21916__,
    new_new_n21917__, new_new_n21918__, new_new_n21919__, new_new_n21920__,
    new_new_n21921__, new_new_n21922__, new_new_n21923__, new_new_n21924__,
    new_new_n21925__, new_new_n21926__, new_new_n21927__, new_new_n21928__,
    new_new_n21929__, new_new_n21930__, new_new_n21931__, new_new_n21932__,
    new_new_n21933__, new_new_n21934__, new_new_n21935__, new_new_n21936__,
    new_new_n21937__, new_new_n21938__, new_new_n21939__, new_new_n21940__,
    new_new_n21941__, new_new_n21942__, new_new_n21943__, new_new_n21944__,
    new_new_n21945__, new_new_n21946__, new_new_n21947__, new_new_n21948__,
    new_new_n21949__, new_new_n21950__, new_new_n21951__, new_new_n21952__,
    new_new_n21953__, new_new_n21954__, new_new_n21955__, new_new_n21956__,
    new_new_n21957__, new_new_n21958__, new_new_n21959__, new_new_n21960__,
    new_new_n21961__, new_new_n21962__, new_new_n21963__, new_new_n21964__,
    new_new_n21965__, new_new_n21966__, new_new_n21967__, new_new_n21968__,
    new_new_n21969__, new_new_n21970__, new_new_n21971__, new_new_n21972__,
    new_new_n21973__, new_new_n21974__, new_new_n21975__, new_new_n21976__,
    new_new_n21977__, new_new_n21978__, new_new_n21979__, new_new_n21980__,
    new_new_n21981__, new_new_n21982__, new_new_n21983__, new_new_n21984__,
    new_new_n21985__, new_new_n21986__, new_new_n21987__, new_new_n21988__,
    new_new_n21989__, new_new_n21990__, new_new_n21991__, new_new_n21992__,
    new_new_n21993__, new_new_n21994__, new_new_n21995__, new_new_n21996__,
    new_new_n21997__, new_new_n21998__, new_new_n21999__, new_new_n22000__,
    new_new_n22001__, new_new_n22002__, new_new_n22003__, new_new_n22004__,
    new_new_n22005__, new_new_n22006__, new_new_n22007__, new_new_n22008__,
    new_new_n22009__, new_new_n22010__, new_new_n22011__, new_new_n22012__,
    new_new_n22013__, new_new_n22014__, new_new_n22015__, new_new_n22016__,
    new_new_n22017__, new_new_n22018__, new_new_n22019__, new_new_n22020__,
    new_new_n22021__, new_new_n22022__, new_new_n22023__, new_new_n22024__,
    new_new_n22025__, new_new_n22026__, new_new_n22027__, new_new_n22028__,
    new_new_n22029__, new_new_n22030__, new_new_n22031__, new_new_n22032__,
    new_new_n22033__, new_new_n22034__, new_new_n22035__, new_new_n22036__,
    new_new_n22037__, new_new_n22038__, new_new_n22039__, new_new_n22040__,
    new_new_n22041__, new_new_n22042__, new_new_n22043__, new_new_n22044__,
    new_new_n22045__, new_new_n22046__, new_new_n22047__, new_new_n22048__,
    new_new_n22049__, new_new_n22050__, new_new_n22051__, new_new_n22052__,
    new_new_n22053__, new_new_n22054__, new_new_n22055__, new_new_n22056__,
    new_new_n22057__, new_new_n22058__, new_new_n22059__, new_new_n22060__,
    new_new_n22061__, new_new_n22062__, new_new_n22063__, new_new_n22064__,
    new_new_n22065__, new_new_n22066__, new_new_n22067__, new_new_n22068__,
    new_new_n22069__, new_new_n22070__, new_new_n22071__, new_new_n22072__,
    new_new_n22073__, new_new_n22074__, new_new_n22075__, new_new_n22076__,
    new_new_n22077__, new_new_n22078__, new_new_n22079__, new_new_n22080__,
    new_new_n22081__, new_new_n22082__, new_new_n22083__, new_new_n22084__,
    new_new_n22085__, new_new_n22086__, new_new_n22087__, new_new_n22088__,
    new_new_n22089__, new_new_n22090__, new_new_n22091__, new_new_n22092__,
    new_new_n22093__, new_new_n22094__, new_new_n22095__, new_new_n22096__,
    new_new_n22097__, new_new_n22098__, new_new_n22099__, new_new_n22100__,
    new_new_n22101__, new_new_n22102__, new_new_n22103__, new_new_n22104__,
    new_new_n22105__, new_new_n22106__, new_new_n22107__, new_new_n22108__,
    new_new_n22109__, new_new_n22110__, new_new_n22111__, new_new_n22112__,
    new_new_n22113__, new_new_n22114__, new_new_n22115__, new_new_n22116__,
    new_new_n22117__, new_new_n22118__, new_new_n22119__, new_new_n22120__,
    new_new_n22121__, new_new_n22122__, new_new_n22123__, new_new_n22124__,
    new_new_n22125__, new_new_n22126__, new_new_n22127__, new_new_n22128__,
    new_new_n22129__, new_new_n22130__, new_new_n22131__, new_new_n22132__,
    new_new_n22133__, new_new_n22134__, new_new_n22135__, new_new_n22136__,
    new_new_n22137__, new_new_n22138__, new_new_n22139__, new_new_n22140__,
    new_new_n22141__, new_new_n22142__, new_new_n22143__, new_new_n22144__,
    new_new_n22145__, new_new_n22146__, new_new_n22147__, new_new_n22148__,
    new_new_n22149__, new_new_n22150__, new_new_n22151__, new_new_n22152__,
    new_new_n22153__, new_new_n22154__, new_new_n22155__, new_new_n22156__,
    new_new_n22157__, new_new_n22158__, new_new_n22159__, new_new_n22160__,
    new_new_n22161__, new_new_n22162__, new_new_n22163__, new_new_n22164__,
    new_new_n22165__, new_new_n22166__, new_new_n22167__, new_new_n22168__,
    new_new_n22169__, new_new_n22170__, new_new_n22171__, new_new_n22172__,
    new_new_n22173__, new_new_n22174__, new_new_n22175__, new_new_n22176__,
    new_new_n22177__, new_new_n22178__, new_new_n22179__, new_new_n22180__,
    new_new_n22181__, new_new_n22182__, new_new_n22183__, new_new_n22184__,
    new_new_n22185__, new_new_n22186__, new_new_n22187__, new_new_n22188__,
    new_new_n22189__, new_new_n22190__, new_new_n22191__, new_new_n22192__,
    new_new_n22193__, new_new_n22194__, new_new_n22195__, new_new_n22196__,
    new_new_n22197__, new_new_n22198__, new_new_n22199__, new_new_n22200__,
    new_new_n22201__, new_new_n22202__, new_new_n22203__, new_new_n22204__,
    new_new_n22205__, new_new_n22206__, new_new_n22207__, new_new_n22208__,
    new_new_n22209__, new_new_n22210__, new_new_n22211__, new_new_n22212__,
    new_new_n22213__, new_new_n22214__, new_new_n22215__, new_new_n22216__,
    new_new_n22217__, new_new_n22218__, new_new_n22219__, new_new_n22220__,
    new_new_n22221__, new_new_n22222__, new_new_n22223__, new_new_n22224__,
    new_new_n22225__, new_new_n22226__, new_new_n22227__, new_new_n22228__,
    new_new_n22229__, new_new_n22230__, new_new_n22231__, new_new_n22232__,
    new_new_n22233__, new_new_n22234__, new_new_n22235__, new_new_n22236__,
    new_new_n22237__, new_new_n22238__, new_new_n22239__, new_new_n22240__,
    new_new_n22241__, new_new_n22242__, new_new_n22243__, new_new_n22244__,
    new_new_n22245__, new_new_n22246__, new_new_n22247__, new_new_n22248__,
    new_new_n22249__, new_new_n22250__, new_new_n22251__, new_new_n22252__,
    new_new_n22253__, new_new_n22254__, new_new_n22255__, new_new_n22256__,
    new_new_n22257__, new_new_n22258__, new_new_n22259__, new_new_n22260__,
    new_new_n22261__, new_new_n22262__, new_new_n22263__, new_new_n22264__,
    new_new_n22265__, new_new_n22266__, new_new_n22267__, new_new_n22268__,
    new_new_n22269__, new_new_n22270__, new_new_n22271__, new_new_n22272__,
    new_new_n22273__, new_new_n22274__, new_new_n22275__, new_new_n22276__,
    new_new_n22277__, new_new_n22278__, new_new_n22279__, new_new_n22280__,
    new_new_n22281__, new_new_n22282__, new_new_n22283__, new_new_n22284__,
    new_new_n22285__, new_new_n22286__, new_new_n22287__, new_new_n22288__,
    new_new_n22289__, new_new_n22290__, new_new_n22291__, new_new_n22292__,
    new_new_n22293__, new_new_n22294__, new_new_n22295__, new_new_n22296__,
    new_new_n22297__, new_new_n22298__, new_new_n22299__, new_new_n22300__,
    new_new_n22301__, new_new_n22302__, new_new_n22303__, new_new_n22304__,
    new_new_n22305__, new_new_n22306__, new_new_n22307__, new_new_n22308__,
    new_new_n22309__, new_new_n22310__, new_new_n22311__, new_new_n22312__,
    new_new_n22313__, new_new_n22314__, new_new_n22315__, new_new_n22316__,
    new_new_n22317__, new_new_n22318__, new_new_n22319__, new_new_n22320__,
    new_new_n22321__, new_new_n22322__, new_new_n22323__, new_new_n22324__,
    new_new_n22325__, new_new_n22326__, new_new_n22327__, new_new_n22328__,
    new_new_n22329__, new_new_n22330__, new_new_n22331__, new_new_n22332__,
    new_new_n22333__, new_new_n22334__, new_new_n22335__, new_new_n22336__,
    new_new_n22337__, new_new_n22338__, new_new_n22339__, new_new_n22340__,
    new_new_n22341__, new_new_n22342__, new_new_n22343__, new_new_n22344__,
    new_new_n22345__, new_new_n22346__, new_new_n22347__, new_new_n22348__,
    new_new_n22349__, new_new_n22350__, new_new_n22351__, new_new_n22352__,
    new_new_n22353__, new_new_n22354__, new_new_n22355__, new_new_n22356__,
    new_new_n22357__, new_new_n22358__, new_new_n22359__, new_new_n22360__,
    new_new_n22361__, new_new_n22362__, new_new_n22363__, new_new_n22364__,
    new_new_n22365__, new_new_n22366__, new_new_n22367__, new_new_n22368__,
    new_new_n22369__, new_new_n22370__, new_new_n22371__, new_new_n22372__,
    new_new_n22373__, new_new_n22374__, new_new_n22375__, new_new_n22376__,
    new_new_n22377__, new_new_n22378__, new_new_n22379__, new_new_n22380__,
    new_new_n22381__, new_new_n22382__, new_new_n22383__, new_new_n22384__,
    new_new_n22385__, new_new_n22386__, new_new_n22387__, new_new_n22388__,
    new_new_n22389__, new_new_n22390__, new_new_n22391__, new_new_n22392__,
    new_new_n22393__, new_new_n22394__, new_new_n22395__, new_new_n22396__,
    new_new_n22397__, new_new_n22398__, new_new_n22399__, new_new_n22400__,
    new_new_n22401__, new_new_n22402__, new_new_n22403__, new_new_n22404__,
    new_new_n22405__, new_new_n22406__, new_new_n22407__, new_new_n22408__,
    new_new_n22409__, new_new_n22410__, new_new_n22411__, new_new_n22412__,
    new_new_n22413__, new_new_n22414__, new_new_n22415__, new_new_n22416__,
    new_new_n22417__, new_new_n22418__, new_new_n22419__, new_new_n22420__,
    new_new_n22421__, new_new_n22422__, new_new_n22423__, new_new_n22424__,
    new_new_n22425__, new_new_n22426__, new_new_n22427__, new_new_n22428__,
    new_new_n22429__, new_new_n22430__, new_new_n22431__, new_new_n22432__,
    new_new_n22433__, new_new_n22434__, new_new_n22435__, new_new_n22436__,
    new_new_n22437__, new_new_n22438__, new_new_n22439__, new_new_n22440__,
    new_new_n22441__, new_new_n22442__, new_new_n22443__, new_new_n22444__,
    new_new_n22445__, new_new_n22446__, new_new_n22447__, new_new_n22448__,
    new_new_n22449__, new_new_n22450__, new_new_n22451__, new_new_n22452__,
    new_new_n22453__, new_new_n22454__, new_new_n22455__, new_new_n22456__,
    new_new_n22457__, new_new_n22458__, new_new_n22459__, new_new_n22460__,
    new_new_n22461__, new_new_n22462__, new_new_n22463__, new_new_n22464__,
    new_new_n22465__, new_new_n22466__, new_new_n22467__, new_new_n22468__,
    new_new_n22469__, new_new_n22470__, new_new_n22471__, new_new_n22472__,
    new_new_n22473__, new_new_n22474__, new_new_n22475__, new_new_n22476__,
    new_new_n22477__, new_new_n22478__, new_new_n22479__, new_new_n22480__,
    new_new_n22481__, new_new_n22482__, new_new_n22483__, new_new_n22484__,
    new_new_n22485__, new_new_n22486__, new_new_n22487__, new_new_n22488__,
    new_new_n22489__, new_new_n22490__, new_new_n22491__, new_new_n22492__,
    new_new_n22493__, new_new_n22494__, new_new_n22495__, new_new_n22496__,
    new_new_n22497__, new_new_n22498__, new_new_n22499__, new_new_n22500__,
    new_new_n22501__, new_new_n22502__, new_new_n22503__, new_new_n22504__,
    new_new_n22505__, new_new_n22506__, new_new_n22507__, new_new_n22508__,
    new_new_n22509__, new_new_n22510__, new_new_n22511__, new_new_n22512__,
    new_new_n22513__, new_new_n22514__, new_new_n22515__, new_new_n22516__,
    new_new_n22517__, new_new_n22518__, new_new_n22519__, new_new_n22520__,
    new_new_n22521__, new_new_n22522__, new_new_n22523__, new_new_n22524__,
    new_new_n22525__, new_new_n22526__, new_new_n22527__, new_new_n22528__,
    new_new_n22529__, new_new_n22530__, new_new_n22531__, new_new_n22532__,
    new_new_n22533__, new_new_n22534__, new_new_n22535__, new_new_n22536__,
    new_new_n22537__, new_new_n22538__, new_new_n22539__, new_new_n22540__,
    new_new_n22541__, new_new_n22542__, new_new_n22543__, new_new_n22544__,
    new_new_n22545__, new_new_n22546__, new_new_n22547__, new_new_n22548__,
    new_new_n22549__, new_new_n22550__, new_new_n22551__, new_new_n22552__,
    new_new_n22553__, new_new_n22554__, new_new_n22555__, new_new_n22556__,
    new_new_n22557__, new_new_n22558__, new_new_n22559__, new_new_n22560__,
    new_new_n22561__, new_new_n22562__, new_new_n22563__, new_new_n22564__,
    new_new_n22565__, new_new_n22566__, new_new_n22567__, new_new_n22568__,
    new_new_n22569__, new_new_n22570__, new_new_n22571__, new_new_n22572__,
    new_new_n22573__, new_new_n22574__, new_new_n22575__, new_new_n22576__,
    new_new_n22577__, new_new_n22578__, new_new_n22579__, new_new_n22580__,
    new_new_n22581__, new_new_n22582__, new_new_n22583__, new_new_n22584__,
    new_new_n22585__, new_new_n22586__, new_new_n22587__, new_new_n22588__,
    new_new_n22589__, new_new_n22590__, new_new_n22591__, new_new_n22592__,
    new_new_n22593__, new_new_n22594__, new_new_n22595__, new_new_n22596__,
    new_new_n22597__, new_new_n22598__, new_new_n22599__, new_new_n22600__,
    new_new_n22601__, new_new_n22602__, new_new_n22603__, new_new_n22604__,
    new_new_n22605__, new_new_n22606__, new_new_n22607__, new_new_n22608__,
    new_new_n22609__, new_new_n22610__, new_new_n22611__, new_new_n22612__,
    new_new_n22613__, new_new_n22614__, new_new_n22615__, new_new_n22616__,
    new_new_n22617__, new_new_n22618__, new_new_n22619__, new_new_n22620__,
    new_new_n22621__, new_new_n22622__, new_new_n22623__, new_new_n22624__,
    new_new_n22625__, new_new_n22626__, new_new_n22627__, new_new_n22628__,
    new_new_n22629__, new_new_n22630__, new_new_n22631__, new_new_n22632__,
    new_new_n22633__, new_new_n22634__, new_new_n22635__, new_new_n22636__,
    new_new_n22637__, new_new_n22638__, new_new_n22639__, new_new_n22640__,
    new_new_n22641__, new_new_n22642__, new_new_n22643__, new_new_n22644__,
    new_new_n22645__, new_new_n22646__, new_new_n22647__, new_new_n22648__,
    new_new_n22649__, new_new_n22650__, new_new_n22651__, new_new_n22652__,
    new_new_n22653__, new_new_n22654__, new_new_n22655__, new_new_n22656__,
    new_new_n22657__, new_new_n22658__, new_new_n22659__, new_new_n22660__,
    new_new_n22661__, new_new_n22662__, new_new_n22663__, new_new_n22664__,
    new_new_n22665__, new_new_n22666__, new_new_n22667__, new_new_n22668__,
    new_new_n22669__, new_new_n22670__, new_new_n22671__, new_new_n22672__,
    new_new_n22673__, new_new_n22674__, new_new_n22675__, new_new_n22676__,
    new_new_n22677__, new_new_n22678__, new_new_n22679__, new_new_n22680__,
    new_new_n22681__, new_new_n22682__, new_new_n22683__, new_new_n22684__,
    new_new_n22685__, new_new_n22686__, new_new_n22687__, new_new_n22688__,
    new_new_n22689__, new_new_n22690__, new_new_n22691__, new_new_n22692__,
    new_new_n22693__, new_new_n22694__, new_new_n22695__, new_new_n22696__,
    new_new_n22697__, new_new_n22698__, new_new_n22699__, new_new_n22700__,
    new_new_n22701__, new_new_n22702__, new_new_n22703__, new_new_n22704__,
    new_new_n22705__, new_new_n22706__, new_new_n22707__, new_new_n22708__,
    new_new_n22709__, new_new_n22710__, new_new_n22711__, new_new_n22712__,
    new_new_n22713__, new_new_n22714__, new_new_n22715__, new_new_n22716__,
    new_new_n22717__, new_new_n22718__, new_new_n22719__, new_new_n22720__,
    new_new_n22721__, new_new_n22722__, new_new_n22723__, new_new_n22724__,
    new_new_n22725__, new_new_n22726__, new_new_n22727__, new_new_n22728__,
    new_new_n22729__, new_new_n22730__, new_new_n22731__, new_new_n22732__,
    new_new_n22733__, new_new_n22734__, new_new_n22735__, new_new_n22736__,
    new_new_n22737__, new_new_n22738__, new_new_n22739__, new_new_n22740__,
    new_new_n22741__, new_new_n22742__, new_new_n22743__, new_new_n22744__,
    new_new_n22745__, new_new_n22746__, new_new_n22747__, new_new_n22748__,
    new_new_n22749__, new_new_n22750__, new_new_n22751__, new_new_n22752__,
    new_new_n22753__, new_new_n22754__, new_new_n22755__, new_new_n22756__,
    new_new_n22757__, new_new_n22758__, new_new_n22759__, new_new_n22760__,
    new_new_n22761__, new_new_n22762__, new_new_n22763__, new_new_n22764__,
    new_new_n22765__, new_new_n22766__, new_new_n22767__, new_new_n22768__,
    new_new_n22769__, new_new_n22770__, new_new_n22771__, new_new_n22772__,
    new_new_n22773__, new_new_n22774__, new_new_n22775__, new_new_n22776__,
    new_new_n22777__, new_new_n22778__, new_new_n22779__, new_new_n22780__,
    new_new_n22781__, new_new_n22782__, new_new_n22783__, new_new_n22784__,
    new_new_n22785__, new_new_n22786__, new_new_n22787__, new_new_n22788__,
    new_new_n22789__, new_new_n22790__, new_new_n22791__, new_new_n22792__,
    new_new_n22793__, new_new_n22794__, new_new_n22795__, new_new_n22796__,
    new_new_n22797__, new_new_n22798__, new_new_n22799__, new_new_n22800__,
    new_new_n22801__, new_new_n22802__, new_new_n22803__, new_new_n22804__,
    new_new_n22805__, new_new_n22806__, new_new_n22807__, new_new_n22808__,
    new_new_n22809__, new_new_n22810__, new_new_n22811__, new_new_n22812__,
    new_new_n22813__, new_new_n22814__, new_new_n22815__, new_new_n22816__,
    new_new_n22817__, new_new_n22818__, new_new_n22819__, new_new_n22820__,
    new_new_n22821__, new_new_n22822__, new_new_n22823__, new_new_n22824__,
    new_new_n22825__, new_new_n22826__, new_new_n22827__, new_new_n22828__,
    new_new_n22829__, new_new_n22830__, new_new_n22831__, new_new_n22832__,
    new_new_n22833__, new_new_n22834__, new_new_n22835__, new_new_n22836__,
    new_new_n22837__, new_new_n22838__, new_new_n22839__, new_new_n22840__,
    new_new_n22841__, new_new_n22842__, new_new_n22843__, new_new_n22844__,
    new_new_n22845__, new_new_n22846__, new_new_n22847__, new_new_n22848__,
    new_new_n22849__, new_new_n22850__, new_new_n22851__, new_new_n22852__,
    new_new_n22853__, new_new_n22854__, new_new_n22855__, new_new_n22856__,
    new_new_n22857__, new_new_n22858__, new_new_n22859__, new_new_n22860__,
    new_new_n22861__, new_new_n22862__, new_new_n22863__, new_new_n22864__,
    new_new_n22865__, new_new_n22866__, new_new_n22867__, new_new_n22868__,
    new_new_n22869__, new_new_n22870__, new_new_n22871__, new_new_n22872__,
    new_new_n22873__, new_new_n22874__, new_new_n22875__, new_new_n22876__,
    new_new_n22877__, new_new_n22878__, new_new_n22879__, new_new_n22880__,
    new_new_n22881__, new_new_n22882__, new_new_n22883__, new_new_n22884__,
    new_new_n22885__, new_new_n22886__, new_new_n22887__, new_new_n22888__,
    new_new_n22889__, new_new_n22890__, new_new_n22891__, new_new_n22892__,
    new_new_n22893__, new_new_n22894__, new_new_n22895__, new_new_n22896__,
    new_new_n22897__, new_new_n22898__, new_new_n22899__, new_new_n22900__,
    new_new_n22901__, new_new_n22902__, new_new_n22903__, new_new_n22904__,
    new_new_n22905__, new_new_n22906__, new_new_n22907__, new_new_n22908__,
    new_new_n22909__, new_new_n22910__, new_new_n22911__, new_new_n22912__,
    new_new_n22913__, new_new_n22914__, new_new_n22915__, new_new_n22916__,
    new_new_n22917__, new_new_n22918__, new_new_n22919__, new_new_n22920__,
    new_new_n22921__, new_new_n22922__, new_new_n22923__, new_new_n22924__,
    new_new_n22925__, new_new_n22926__, new_new_n22927__, new_new_n22928__,
    new_new_n22929__, new_new_n22930__, new_new_n22931__, new_new_n22932__,
    new_new_n22933__, new_new_n22934__, new_new_n22935__, new_new_n22936__,
    new_new_n22937__, new_new_n22938__, new_new_n22939__, new_new_n22940__,
    new_new_n22941__, new_new_n22942__, new_new_n22943__, new_new_n22944__,
    new_new_n22945__, new_new_n22946__, new_new_n22947__, new_new_n22948__,
    new_new_n22949__, new_new_n22950__, new_new_n22951__, new_new_n22952__,
    new_new_n22953__, new_new_n22954__, new_new_n22955__, new_new_n22956__,
    new_new_n22957__, new_new_n22958__, new_new_n22959__, new_new_n22960__,
    new_new_n22961__, new_new_n22962__, new_new_n22963__, new_new_n22964__,
    new_new_n22965__, new_new_n22966__, new_new_n22967__, new_new_n22968__,
    new_new_n22969__, new_new_n22970__, new_new_n22971__, new_new_n22972__,
    new_new_n22973__, new_new_n22974__, new_new_n22975__, new_new_n22976__,
    new_new_n22977__, new_new_n22978__, new_new_n22979__, new_new_n22980__,
    new_new_n22981__, new_new_n22982__, new_new_n22983__, new_new_n22984__,
    new_new_n22985__, new_new_n22986__, new_new_n22987__, new_new_n22988__,
    new_new_n22989__, new_new_n22990__, new_new_n22991__, new_new_n22992__,
    new_new_n22993__, new_new_n22994__, new_new_n22995__, new_new_n22996__,
    new_new_n22997__, new_new_n22998__, new_new_n22999__, new_new_n23000__,
    new_new_n23001__, new_new_n23002__, new_new_n23003__, new_new_n23004__,
    new_new_n23005__, new_new_n23006__, new_new_n23007__, new_new_n23008__,
    new_new_n23009__, new_new_n23010__, new_new_n23011__, new_new_n23012__,
    new_new_n23013__, new_new_n23014__, new_new_n23015__, new_new_n23016__,
    new_new_n23017__, new_new_n23018__, new_new_n23019__, new_new_n23020__,
    new_new_n23021__, new_new_n23022__, new_new_n23023__, new_new_n23024__,
    new_new_n23025__, new_new_n23026__, new_new_n23027__, new_new_n23028__,
    new_new_n23029__, new_new_n23030__, new_new_n23031__, new_new_n23032__,
    new_new_n23033__, new_new_n23034__, new_new_n23035__, new_new_n23036__,
    new_new_n23037__, new_new_n23038__, new_new_n23039__, new_new_n23040__,
    new_new_n23041__, new_new_n23042__, new_new_n23043__, new_new_n23044__,
    new_new_n23045__, new_new_n23046__, new_new_n23047__, new_new_n23048__,
    new_new_n23049__, new_new_n23050__, new_new_n23051__, new_new_n23052__,
    new_new_n23053__, new_new_n23054__, new_new_n23055__, new_new_n23056__,
    new_new_n23057__, new_new_n23058__, new_new_n23059__, new_new_n23060__,
    new_new_n23061__, new_new_n23062__, new_new_n23063__, new_new_n23064__,
    new_new_n23065__, new_new_n23066__, new_new_n23067__, new_new_n23068__,
    new_new_n23069__, new_new_n23070__, new_new_n23071__, new_new_n23072__,
    new_new_n23073__, new_new_n23074__, new_new_n23075__, new_new_n23076__,
    new_new_n23077__, new_new_n23078__, new_new_n23079__, new_new_n23080__,
    new_new_n23081__, new_new_n23082__, new_new_n23083__, new_new_n23084__,
    new_new_n23085__, new_new_n23086__, new_new_n23087__, new_new_n23088__,
    new_new_n23089__, new_new_n23090__, new_new_n23091__, new_new_n23092__,
    new_new_n23093__, new_new_n23094__, new_new_n23095__, new_new_n23096__,
    new_new_n23097__, new_new_n23098__, new_new_n23099__, new_new_n23100__,
    new_new_n23101__, new_new_n23102__, new_new_n23103__, new_new_n23104__,
    new_new_n23105__, new_new_n23106__, new_new_n23107__, new_new_n23108__,
    new_new_n23109__, new_new_n23110__, new_new_n23111__, new_new_n23112__,
    new_new_n23113__, new_new_n23114__, new_new_n23115__, new_new_n23116__,
    new_new_n23117__, new_new_n23118__, new_new_n23119__, new_new_n23120__,
    new_new_n23121__, new_new_n23122__, new_new_n23123__, new_new_n23124__,
    new_new_n23125__, new_new_n23126__, new_new_n23127__, new_new_n23128__,
    new_new_n23129__, new_new_n23130__, new_new_n23131__, new_new_n23132__,
    new_new_n23133__, new_new_n23134__, new_new_n23135__, new_new_n23136__,
    new_new_n23137__, new_new_n23138__, new_new_n23139__, new_new_n23140__,
    new_new_n23141__, new_new_n23142__, new_new_n23143__, new_new_n23144__,
    new_new_n23145__, new_new_n23146__, new_new_n23147__, new_new_n23148__,
    new_new_n23149__, new_new_n23150__, new_new_n23151__, new_new_n23152__,
    new_new_n23153__, new_new_n23154__, new_new_n23155__, new_new_n23156__,
    new_new_n23157__, new_new_n23158__, new_new_n23159__, new_new_n23160__,
    new_new_n23161__, new_new_n23162__, new_new_n23163__, new_new_n23164__,
    new_new_n23165__, new_new_n23166__, new_new_n23167__, new_new_n23168__,
    new_new_n23169__, new_new_n23170__, new_new_n23171__, new_new_n23172__,
    new_new_n23173__, new_new_n23174__, new_new_n23175__, new_new_n23176__,
    new_new_n23177__, new_new_n23178__, new_new_n23179__, new_new_n23180__,
    new_new_n23181__, new_new_n23182__, new_new_n23183__, new_new_n23184__,
    new_new_n23185__, new_new_n23186__, new_new_n23187__, new_new_n23188__,
    new_new_n23189__, new_new_n23190__, new_new_n23191__, new_new_n23192__,
    new_new_n23193__, new_new_n23194__, new_new_n23195__, new_new_n23196__,
    new_new_n23197__, new_new_n23198__, new_new_n23199__, new_new_n23200__,
    new_new_n23201__, new_new_n23202__, new_new_n23203__, new_new_n23204__,
    new_new_n23205__, new_new_n23206__, new_new_n23207__, new_new_n23208__,
    new_new_n23209__, new_new_n23210__, new_new_n23211__, new_new_n23212__,
    new_new_n23213__, new_new_n23214__, new_new_n23215__, new_new_n23216__,
    new_new_n23217__, new_new_n23218__, new_new_n23219__, new_new_n23220__,
    new_new_n23221__, new_new_n23222__, new_new_n23223__, new_new_n23224__,
    new_new_n23225__, new_new_n23226__, new_new_n23227__, new_new_n23228__,
    new_new_n23229__, new_new_n23230__, new_new_n23231__, new_new_n23232__,
    new_new_n23233__, new_new_n23234__, new_new_n23235__, new_new_n23236__,
    new_new_n23237__, new_new_n23238__, new_new_n23239__, new_new_n23240__,
    new_new_n23241__, new_new_n23242__, new_new_n23243__, new_new_n23244__,
    new_new_n23245__, new_new_n23246__, new_new_n23247__, new_new_n23248__,
    new_new_n23249__, new_new_n23250__, new_new_n23251__, new_new_n23252__,
    new_new_n23253__, new_new_n23254__, new_new_n23255__, new_new_n23256__,
    new_new_n23257__, new_new_n23258__, new_new_n23259__, new_new_n23260__,
    new_new_n23261__, new_new_n23262__, new_new_n23263__, new_new_n23264__,
    new_new_n23265__, new_new_n23266__, new_new_n23267__, new_new_n23268__,
    new_new_n23269__, new_new_n23270__, new_new_n23271__, new_new_n23272__,
    new_new_n23273__, new_new_n23274__, new_new_n23275__, new_new_n23276__,
    new_new_n23277__, new_new_n23278__, new_new_n23279__, new_new_n23280__,
    new_new_n23281__, new_new_n23282__, new_new_n23283__, new_new_n23284__,
    new_new_n23285__, new_new_n23286__, new_new_n23287__, new_new_n23288__,
    new_new_n23289__, new_new_n23290__, new_new_n23291__, new_new_n23292__,
    new_new_n23293__, new_new_n23294__, new_new_n23295__, new_new_n23296__,
    new_new_n23297__, new_new_n23298__, new_new_n23299__, new_new_n23300__,
    new_new_n23301__, new_new_n23302__, new_new_n23303__, new_new_n23304__,
    new_new_n23305__, new_new_n23306__, new_new_n23307__, new_new_n23308__,
    new_new_n23309__, new_new_n23310__, new_new_n23311__, new_new_n23312__,
    new_new_n23313__, new_new_n23314__, new_new_n23315__, new_new_n23316__,
    new_new_n23317__, new_new_n23318__, new_new_n23319__, new_new_n23320__,
    new_new_n23321__, new_new_n23322__, new_new_n23323__, new_new_n23324__,
    new_new_n23325__, new_new_n23326__, new_new_n23327__, new_new_n23328__,
    new_new_n23329__, new_new_n23330__, new_new_n23331__, new_new_n23332__,
    new_new_n23333__, new_new_n23334__, new_new_n23335__, new_new_n23336__,
    new_new_n23337__, new_new_n23338__, new_new_n23339__, new_new_n23340__,
    new_new_n23341__, new_new_n23342__, new_new_n23343__, new_new_n23344__,
    new_new_n23345__, new_new_n23346__, new_new_n23347__, new_new_n23348__,
    new_new_n23349__, new_new_n23350__, new_new_n23351__, new_new_n23352__,
    new_new_n23353__, new_new_n23354__, new_new_n23355__, new_new_n23356__,
    new_new_n23357__, new_new_n23358__, new_new_n23359__, new_new_n23360__,
    new_new_n23361__, new_new_n23362__, new_new_n23363__, new_new_n23364__,
    new_new_n23365__, new_new_n23366__, new_new_n23367__, new_new_n23368__,
    new_new_n23369__, new_new_n23370__, new_new_n23371__, new_new_n23372__,
    new_new_n23373__, new_new_n23374__, new_new_n23375__, new_new_n23376__,
    new_new_n23377__, new_new_n23378__, new_new_n23379__, new_new_n23380__,
    new_new_n23381__, new_new_n23382__, new_new_n23383__, new_new_n23384__,
    new_new_n23385__, new_new_n23386__, new_new_n23387__, new_new_n23388__,
    new_new_n23389__, new_new_n23390__, new_new_n23391__, new_new_n23392__,
    new_new_n23393__, new_new_n23394__, new_new_n23395__, new_new_n23396__,
    new_new_n23397__, new_new_n23398__, new_new_n23399__, new_new_n23400__,
    new_new_n23401__, new_new_n23402__, new_new_n23403__, new_new_n23404__,
    new_new_n23405__, new_new_n23406__, new_new_n23407__, new_new_n23408__,
    new_new_n23409__, new_new_n23410__, new_new_n23411__, new_new_n23412__,
    new_new_n23413__, new_new_n23414__, new_new_n23415__, new_new_n23416__,
    new_new_n23417__, new_new_n23418__, new_new_n23419__, new_new_n23420__,
    new_new_n23421__, new_new_n23422__, new_new_n23423__, new_new_n23424__,
    new_new_n23425__, new_new_n23426__, new_new_n23427__, new_new_n23428__,
    new_new_n23429__, new_new_n23430__, new_new_n23431__, new_new_n23432__,
    new_new_n23433__, new_new_n23434__, new_new_n23435__, new_new_n23436__,
    new_new_n23437__, new_new_n23438__, new_new_n23439__, new_new_n23440__,
    new_new_n23441__, new_new_n23442__, new_new_n23443__, new_new_n23444__,
    new_new_n23445__, new_new_n23446__, new_new_n23447__, new_new_n23448__,
    new_new_n23449__, new_new_n23450__, new_new_n23451__, new_new_n23452__,
    new_new_n23453__, new_new_n23454__, new_new_n23455__, new_new_n23456__,
    new_new_n23457__, new_new_n23458__, new_new_n23459__, new_new_n23460__,
    new_new_n23461__, new_new_n23462__, new_new_n23463__, new_new_n23464__,
    new_new_n23465__, new_new_n23466__, new_new_n23467__, new_new_n23468__,
    new_new_n23469__, new_new_n23470__, new_new_n23471__, new_new_n23472__,
    new_new_n23473__, new_new_n23474__, new_new_n23475__, new_new_n23476__,
    new_new_n23477__, new_new_n23478__, new_new_n23479__, new_new_n23480__,
    new_new_n23481__, new_new_n23482__, new_new_n23483__, new_new_n23484__,
    new_new_n23485__, new_new_n23486__, new_new_n23487__, new_new_n23488__,
    new_new_n23489__, new_new_n23490__, new_new_n23491__, new_new_n23492__,
    new_new_n23493__, new_new_n23494__, new_new_n23495__, new_new_n23496__,
    new_new_n23497__, new_new_n23498__, new_new_n23499__, new_new_n23500__,
    new_new_n23501__, new_new_n23502__, new_new_n23503__, new_new_n23504__,
    new_new_n23505__, new_new_n23506__, new_new_n23507__, new_new_n23508__,
    new_new_n23509__, new_new_n23510__, new_new_n23511__, new_new_n23512__,
    new_new_n23513__, new_new_n23514__, new_new_n23515__, new_new_n23516__,
    new_new_n23517__, new_new_n23518__, new_new_n23519__, new_new_n23520__,
    new_new_n23521__, new_new_n23522__, new_new_n23523__, new_new_n23524__,
    new_new_n23525__, new_new_n23526__, new_new_n23527__, new_new_n23528__,
    new_new_n23529__, new_new_n23530__, new_new_n23531__, new_new_n23532__,
    new_new_n23533__, new_new_n23534__, new_new_n23535__, new_new_n23536__,
    new_new_n23537__, new_new_n23538__, new_new_n23539__, new_new_n23540__,
    new_new_n23541__, new_new_n23542__, new_new_n23543__, new_new_n23544__,
    new_new_n23545__, new_new_n23546__, new_new_n23547__, new_new_n23548__,
    new_new_n23549__, new_new_n23550__, new_new_n23551__, new_new_n23552__,
    new_new_n23553__, new_new_n23554__, new_new_n23555__, new_new_n23556__,
    new_new_n23557__, new_new_n23558__, new_new_n23559__, new_new_n23560__,
    new_new_n23561__, new_new_n23562__, new_new_n23563__, new_new_n23564__,
    new_new_n23565__, new_new_n23566__, new_new_n23567__, new_new_n23568__,
    new_new_n23569__, new_new_n23570__, new_new_n23571__, new_new_n23572__,
    new_new_n23573__, new_new_n23574__, new_new_n23575__, new_new_n23576__,
    new_new_n23577__, new_new_n23578__, new_new_n23579__, new_new_n23580__,
    new_new_n23581__, new_new_n23582__, new_new_n23583__, new_new_n23584__,
    new_new_n23585__, new_new_n23586__, new_new_n23587__, new_new_n23588__,
    new_new_n23589__, new_new_n23590__, new_new_n23591__, new_new_n23592__,
    new_new_n23593__, new_new_n23594__, new_new_n23595__, new_new_n23596__,
    new_new_n23597__, new_new_n23598__, new_new_n23599__, new_new_n23600__,
    new_new_n23601__, new_new_n23602__, new_new_n23603__, new_new_n23604__,
    new_new_n23605__, new_new_n23606__, new_new_n23607__, new_new_n23608__,
    new_new_n23609__, new_new_n23610__, new_new_n23611__, new_new_n23612__,
    new_new_n23613__, new_new_n23614__, new_new_n23615__, new_new_n23616__,
    new_new_n23617__, new_new_n23618__, new_new_n23619__, new_new_n23620__,
    new_new_n23621__, new_new_n23622__, new_new_n23623__, new_new_n23624__,
    new_new_n23625__, new_new_n23626__, new_new_n23627__, new_new_n23628__,
    new_new_n23629__, new_new_n23630__, new_new_n23631__, new_new_n23632__,
    new_new_n23633__, new_new_n23634__, new_new_n23635__, new_new_n23636__,
    new_new_n23637__, new_new_n23638__, new_new_n23639__, new_new_n23640__,
    new_new_n23641__, new_new_n23642__, new_new_n23643__, new_new_n23644__,
    new_new_n23645__, new_new_n23646__, new_new_n23647__, new_new_n23648__,
    new_new_n23649__, new_new_n23650__, new_new_n23651__, new_new_n23652__,
    new_new_n23653__, new_new_n23654__, new_new_n23655__, new_new_n23656__,
    new_new_n23657__, new_new_n23658__, new_new_n23659__, new_new_n23660__,
    new_new_n23661__, new_new_n23662__, new_new_n23663__, new_new_n23664__,
    new_new_n23665__, new_new_n23666__, new_new_n23667__, new_new_n23668__,
    new_new_n23669__, new_new_n23670__, new_new_n23671__, new_new_n23672__,
    new_new_n23673__, new_new_n23674__, new_new_n23675__, new_new_n23676__,
    new_new_n23677__, new_new_n23678__, new_new_n23679__, new_new_n23680__,
    new_new_n23681__, new_new_n23682__, new_new_n23683__, new_new_n23684__,
    new_new_n23685__, new_new_n23686__, new_new_n23687__, new_new_n23688__,
    new_new_n23689__, new_new_n23690__, new_new_n23691__, new_new_n23692__,
    new_new_n23693__, new_new_n23694__, new_new_n23695__, new_new_n23696__,
    new_new_n23697__, new_new_n23698__, new_new_n23699__, new_new_n23700__,
    new_new_n23701__, new_new_n23702__, new_new_n23703__, new_new_n23704__,
    new_new_n23705__, new_new_n23706__, new_new_n23707__, new_new_n23708__,
    new_new_n23709__, new_new_n23710__, new_new_n23711__, new_new_n23712__,
    new_new_n23713__, new_new_n23714__, new_new_n23715__, new_new_n23716__,
    new_new_n23717__, new_new_n23718__, new_new_n23719__, new_new_n23720__,
    new_new_n23721__, new_new_n23722__, new_new_n23723__, new_new_n23724__,
    new_new_n23725__, new_new_n23726__, new_new_n23727__, new_new_n23728__,
    new_new_n23729__, new_new_n23730__, new_new_n23731__, new_new_n23732__,
    new_new_n23733__, new_new_n23734__, new_new_n23735__, new_new_n23736__,
    new_new_n23737__, new_new_n23738__, new_new_n23739__, new_new_n23740__,
    new_new_n23741__, new_new_n23742__, new_new_n23743__, new_new_n23744__,
    new_new_n23745__, new_new_n23746__, new_new_n23747__, new_new_n23748__,
    new_new_n23749__, new_new_n23750__, new_new_n23751__, new_new_n23752__,
    new_new_n23753__, new_new_n23754__, new_new_n23755__, new_new_n23756__,
    new_new_n23757__, new_new_n23758__, new_new_n23759__, new_new_n23760__,
    new_new_n23761__, new_new_n23762__, new_new_n23763__, new_new_n23764__,
    new_new_n23765__, new_new_n23766__, new_new_n23767__, new_new_n23768__,
    new_new_n23769__, new_new_n23770__, new_new_n23771__, new_new_n23772__,
    new_new_n23773__, new_new_n23774__, new_new_n23775__, new_new_n23776__,
    new_new_n23777__, new_new_n23778__, new_new_n23779__, new_new_n23780__,
    new_new_n23781__, new_new_n23782__, new_new_n23783__, new_new_n23784__,
    new_new_n23785__, new_new_n23786__, new_new_n23787__, new_new_n23788__,
    new_new_n23789__, new_new_n23790__, new_new_n23791__, new_new_n23792__,
    new_new_n23793__, new_new_n23794__, new_new_n23795__, new_new_n23796__,
    new_new_n23797__, new_new_n23798__, new_new_n23799__, new_new_n23800__,
    new_new_n23801__, new_new_n23802__, new_new_n23803__, new_new_n23804__,
    new_new_n23805__, new_new_n23806__, new_new_n23807__, new_new_n23808__,
    new_new_n23809__, new_new_n23810__, new_new_n23811__, new_new_n23812__,
    new_new_n23813__, new_new_n23814__, new_new_n23815__, new_new_n23816__,
    new_new_n23817__, new_new_n23818__, new_new_n23819__, new_new_n23820__,
    new_new_n23821__, new_new_n23822__, new_new_n23823__, new_new_n23824__,
    new_new_n23825__, new_new_n23826__, new_new_n23827__, new_new_n23828__,
    new_new_n23829__, new_new_n23830__, new_new_n23831__, new_new_n23832__,
    new_new_n23833__, new_new_n23834__, new_new_n23835__, new_new_n23836__,
    new_new_n23837__, new_new_n23838__, new_new_n23839__, new_new_n23840__,
    new_new_n23841__, new_new_n23842__, new_new_n23843__, new_new_n23844__,
    new_new_n23845__, new_new_n23846__, new_new_n23847__, new_new_n23848__,
    new_new_n23849__, new_new_n23850__, new_new_n23851__, new_new_n23852__,
    new_new_n23853__, new_new_n23854__, new_new_n23855__, new_new_n23856__,
    new_new_n23857__, new_new_n23858__, new_new_n23859__, new_new_n23860__,
    new_new_n23861__, new_new_n23862__, new_new_n23863__, new_new_n23864__,
    new_new_n23865__, new_new_n23866__, new_new_n23867__, new_new_n23868__,
    new_new_n23869__, new_new_n23870__, new_new_n23871__, new_new_n23872__,
    new_new_n23873__, new_new_n23874__, new_new_n23875__, new_new_n23876__,
    new_new_n23877__, new_new_n23878__, new_new_n23879__, new_new_n23880__,
    new_new_n23881__, new_new_n23882__, new_new_n23883__, new_new_n23884__,
    new_new_n23885__, new_new_n23886__, new_new_n23887__, new_new_n23888__,
    new_new_n23889__, new_new_n23890__, new_new_n23891__, new_new_n23892__,
    new_new_n23893__, new_new_n23894__, new_new_n23895__, new_new_n23896__,
    new_new_n23897__, new_new_n23898__, new_new_n23899__, new_new_n23900__,
    new_new_n23901__, new_new_n23902__, new_new_n23903__, new_new_n23904__,
    new_new_n23905__, new_new_n23906__, new_new_n23907__, new_new_n23908__,
    new_new_n23909__, new_new_n23910__, new_new_n23911__, new_new_n23912__,
    new_new_n23913__, new_new_n23914__, new_new_n23915__, new_new_n23916__,
    new_new_n23917__, new_new_n23918__, new_new_n23919__, new_new_n23920__,
    new_new_n23921__, new_new_n23922__, new_new_n23923__, new_new_n23924__,
    new_new_n23925__, new_new_n23926__, new_new_n23927__, new_new_n23928__,
    new_new_n23929__, new_new_n23930__, new_new_n23931__, new_new_n23932__,
    new_new_n23933__, new_new_n23934__, new_new_n23935__, new_new_n23936__,
    new_new_n23937__, new_new_n23938__, new_new_n23939__, new_new_n23940__,
    new_new_n23941__, new_new_n23942__, new_new_n23943__, new_new_n23944__,
    new_new_n23945__, new_new_n23946__, new_new_n23947__, new_new_n23948__,
    new_new_n23949__, new_new_n23950__, new_new_n23951__, new_new_n23952__,
    new_new_n23953__, new_new_n23954__, new_new_n23955__, new_new_n23956__,
    new_new_n23957__, new_new_n23958__, new_new_n23959__, new_new_n23960__,
    new_new_n23961__, new_new_n23962__, new_new_n23963__, new_new_n23964__,
    new_new_n23965__, new_new_n23966__, new_new_n23967__, new_new_n23968__,
    new_new_n23969__, new_new_n23970__, new_new_n23971__, new_new_n23972__,
    new_new_n23973__, new_new_n23974__, new_new_n23975__, new_new_n23976__,
    new_new_n23977__, new_new_n23978__, new_new_n23979__, new_new_n23980__,
    new_new_n23981__, new_new_n23982__, new_new_n23983__, new_new_n23984__,
    new_new_n23985__, new_new_n23986__, new_new_n23987__, new_new_n23988__,
    new_new_n23989__, new_new_n23990__, new_new_n23991__, new_new_n23992__,
    new_new_n23993__, new_new_n23994__, new_new_n23995__, new_new_n23996__,
    new_new_n23997__, new_new_n23998__, new_new_n23999__, new_new_n24000__,
    new_new_n24001__, new_new_n24002__, new_new_n24003__, new_new_n24004__,
    new_new_n24005__, new_new_n24006__, new_new_n24007__, new_new_n24008__,
    new_new_n24009__, new_new_n24010__, new_new_n24011__, new_new_n24012__,
    new_new_n24013__, new_new_n24014__, new_new_n24015__, new_new_n24016__,
    new_new_n24017__, new_new_n24018__, new_new_n24019__, new_new_n24020__,
    new_new_n24021__, new_new_n24022__, new_new_n24023__, new_new_n24024__,
    new_new_n24025__, new_new_n24026__, new_new_n24027__, new_new_n24028__,
    new_new_n24029__, new_new_n24030__, new_new_n24031__, new_new_n24032__,
    new_new_n24033__, new_new_n24034__, new_new_n24035__, new_new_n24036__,
    new_new_n24037__, new_new_n24038__, new_new_n24039__, new_new_n24040__,
    new_new_n24041__, new_new_n24042__, new_new_n24043__, new_new_n24044__,
    new_new_n24045__, new_new_n24046__, new_new_n24047__, new_new_n24048__,
    new_new_n24049__, new_new_n24050__, new_new_n24051__, new_new_n24052__,
    new_new_n24053__, new_new_n24054__, new_new_n24055__, new_new_n24056__,
    new_new_n24057__, new_new_n24058__, new_new_n24059__, new_new_n24060__,
    new_new_n24061__, new_new_n24062__, new_new_n24063__, new_new_n24064__,
    new_new_n24065__, new_new_n24066__, new_new_n24067__, new_new_n24068__,
    new_new_n24069__, new_new_n24070__, new_new_n24071__, new_new_n24072__,
    new_new_n24073__, new_new_n24074__, new_new_n24075__, new_new_n24076__,
    new_new_n24077__, new_new_n24078__, new_new_n24079__, new_new_n24080__,
    new_new_n24081__, new_new_n24082__, new_new_n24083__, new_new_n24084__,
    new_new_n24085__, new_new_n24086__, new_new_n24087__, new_new_n24088__,
    new_new_n24089__, new_new_n24090__, new_new_n24091__, new_new_n24092__,
    new_new_n24093__, new_new_n24094__, new_new_n24095__, new_new_n24096__,
    new_new_n24097__, new_new_n24098__, new_new_n24099__, new_new_n24100__,
    new_new_n24101__, new_new_n24102__, new_new_n24103__, new_new_n24104__,
    new_new_n24105__, new_new_n24106__, new_new_n24107__, new_new_n24108__,
    new_new_n24109__, new_new_n24110__, new_new_n24111__, new_new_n24112__,
    new_new_n24113__, new_new_n24114__, new_new_n24115__, new_new_n24116__,
    new_new_n24117__, new_new_n24118__, new_new_n24119__, new_new_n24120__,
    new_new_n24121__, new_new_n24122__, new_new_n24123__, new_new_n24124__,
    new_new_n24125__, new_new_n24126__, new_new_n24127__, new_new_n24128__,
    new_new_n24129__, new_new_n24130__, new_new_n24131__, new_new_n24132__,
    new_new_n24133__, new_new_n24134__, new_new_n24135__, new_new_n24136__,
    new_new_n24137__, new_new_n24138__, new_new_n24139__, new_new_n24140__,
    new_new_n24141__, new_new_n24142__, new_new_n24143__, new_new_n24144__,
    new_new_n24145__, new_new_n24146__, new_new_n24147__, new_new_n24148__,
    new_new_n24149__, new_new_n24150__, new_new_n24151__, new_new_n24152__,
    new_new_n24153__, new_new_n24154__, new_new_n24155__, new_new_n24156__,
    new_new_n24157__, new_new_n24158__, new_new_n24159__, new_new_n24160__,
    new_new_n24161__, new_new_n24162__, new_new_n24163__, new_new_n24164__,
    new_new_n24165__, new_new_n24166__, new_new_n24167__, new_new_n24168__,
    new_new_n24169__, new_new_n24170__, new_new_n24171__, new_new_n24172__,
    new_new_n24173__, new_new_n24174__, new_new_n24175__, new_new_n24176__,
    new_new_n24177__, new_new_n24178__, new_new_n24179__, new_new_n24180__,
    new_new_n24181__, new_new_n24182__, new_new_n24183__, new_new_n24184__,
    new_new_n24185__, new_new_n24186__, new_new_n24187__, new_new_n24188__,
    new_new_n24189__, new_new_n24190__, new_new_n24191__, new_new_n24192__,
    new_new_n24193__, new_new_n24194__, new_new_n24195__, new_new_n24196__,
    new_new_n24197__, new_new_n24198__, new_new_n24199__, new_new_n24200__,
    new_new_n24201__, new_new_n24202__, new_new_n24203__, new_new_n24204__,
    new_new_n24205__, new_new_n24206__, new_new_n24207__, new_new_n24208__,
    new_new_n24209__, new_new_n24210__, new_new_n24211__, new_new_n24212__,
    new_new_n24213__, new_new_n24214__, new_new_n24215__, new_new_n24216__,
    new_new_n24217__, new_new_n24218__, new_new_n24219__, new_new_n24220__,
    new_new_n24221__, new_new_n24222__, new_new_n24223__, new_new_n24224__,
    new_new_n24225__, new_new_n24226__, new_new_n24227__, new_new_n24228__,
    new_new_n24229__, new_new_n24230__, new_new_n24231__, new_new_n24232__,
    new_new_n24233__, new_new_n24234__, new_new_n24235__, new_new_n24236__,
    new_new_n24237__, new_new_n24238__, new_new_n24239__, new_new_n24240__,
    new_new_n24241__, new_new_n24242__, new_new_n24243__, new_new_n24244__,
    new_new_n24245__, new_new_n24246__, new_new_n24247__, new_new_n24248__,
    new_new_n24249__, new_new_n24250__, new_new_n24251__, new_new_n24252__,
    new_new_n24253__, new_new_n24254__, new_new_n24255__, new_new_n24256__,
    new_new_n24257__, new_new_n24258__, new_new_n24259__, new_new_n24260__,
    new_new_n24261__, new_new_n24262__, new_new_n24263__, new_new_n24264__,
    new_new_n24265__, new_new_n24266__, new_new_n24267__, new_new_n24268__,
    new_new_n24269__, new_new_n24270__, new_new_n24271__, new_new_n24272__,
    new_new_n24273__, new_new_n24274__, new_new_n24275__, new_new_n24276__,
    new_new_n24277__, new_new_n24278__, new_new_n24279__, new_new_n24280__,
    new_new_n24281__, new_new_n24282__, new_new_n24283__, new_new_n24284__,
    new_new_n24285__, new_new_n24286__, new_new_n24287__, new_new_n24288__,
    new_new_n24289__, new_new_n24290__, new_new_n24291__, new_new_n24292__,
    new_new_n24293__, new_new_n24294__, new_new_n24295__, new_new_n24296__,
    new_new_n24297__, new_new_n24298__, new_new_n24299__, new_new_n24300__,
    new_new_n24301__, new_new_n24302__, new_new_n24303__, new_new_n24304__,
    new_new_n24305__, new_new_n24306__, new_new_n24307__, new_new_n24308__,
    new_new_n24309__, new_new_n24310__, new_new_n24311__, new_new_n24312__,
    new_new_n24313__, new_new_n24314__, new_new_n24315__, new_new_n24316__,
    new_new_n24317__, new_new_n24318__, new_new_n24319__, new_new_n24320__,
    new_new_n24321__, new_new_n24322__, new_new_n24323__, new_new_n24324__,
    new_new_n24325__, new_new_n24326__, new_new_n24327__, new_new_n24328__,
    new_new_n24329__, new_new_n24330__, new_new_n24331__, new_new_n24332__,
    new_new_n24333__, new_new_n24334__, new_new_n24335__, new_new_n24336__,
    new_new_n24337__, new_new_n24338__, new_new_n24339__, new_new_n24340__,
    new_new_n24341__, new_new_n24342__, new_new_n24343__, new_new_n24344__,
    new_new_n24345__, new_new_n24346__, new_new_n24347__, new_new_n24348__,
    new_new_n24349__, new_new_n24350__, new_new_n24351__, new_new_n24352__,
    new_new_n24353__, new_new_n24354__, new_new_n24355__, new_new_n24356__,
    new_new_n24357__, new_new_n24358__, new_new_n24359__, new_new_n24360__,
    new_new_n24361__, new_new_n24362__, new_new_n24363__, new_new_n24364__,
    new_new_n24365__, new_new_n24366__, new_new_n24367__, new_new_n24368__,
    new_new_n24369__, new_new_n24370__, new_new_n24371__, new_new_n24372__,
    new_new_n24373__, new_new_n24374__, new_new_n24375__, new_new_n24376__,
    new_new_n24377__, new_new_n24378__, new_new_n24379__, new_new_n24380__,
    new_new_n24381__, new_new_n24382__, new_new_n24383__, new_new_n24384__,
    new_new_n24385__, new_new_n24386__, new_new_n24387__, new_new_n24388__,
    new_new_n24389__, new_new_n24390__, new_new_n24391__, new_new_n24392__,
    new_new_n24393__, new_new_n24394__, new_new_n24395__, new_new_n24396__,
    new_new_n24397__, new_new_n24398__, new_new_n24399__, new_new_n24400__,
    new_new_n24401__, new_new_n24402__, new_new_n24403__, new_new_n24404__,
    new_new_n24405__, new_new_n24406__, new_new_n24407__, new_new_n24408__,
    new_new_n24409__, new_new_n24410__, new_new_n24411__, new_new_n24412__,
    new_new_n24413__, new_new_n24414__, new_new_n24415__, new_new_n24416__,
    new_new_n24417__, new_new_n24418__, new_new_n24419__, new_new_n24420__,
    new_new_n24421__, new_new_n24422__, new_new_n24423__, new_new_n24424__,
    new_new_n24425__, new_new_n24426__, new_new_n24427__, new_new_n24428__,
    new_new_n24429__, new_new_n24430__, new_new_n24431__, new_new_n24432__,
    new_new_n24433__, new_new_n24434__, new_new_n24435__, new_new_n24436__,
    new_new_n24437__, new_new_n24438__, new_new_n24439__, new_new_n24440__,
    new_new_n24441__, new_new_n24442__, new_new_n24443__, new_new_n24444__,
    new_new_n24445__, new_new_n24446__, new_new_n24447__, new_new_n24448__,
    new_new_n24449__, new_new_n24450__, new_new_n24451__, new_new_n24452__,
    new_new_n24453__, new_new_n24454__, new_new_n24455__, new_new_n24456__,
    new_new_n24457__, new_new_n24458__, new_new_n24459__, new_new_n24460__,
    new_new_n24461__, new_new_n24462__, new_new_n24463__, new_new_n24464__,
    new_new_n24465__, new_new_n24466__, new_new_n24467__, new_new_n24468__,
    new_new_n24469__, new_new_n24470__, new_new_n24471__, new_new_n24472__,
    new_new_n24473__, new_new_n24474__, new_new_n24475__, new_new_n24476__,
    new_new_n24477__, new_new_n24478__, new_new_n24479__, new_new_n24480__,
    new_new_n24481__, new_new_n24482__, new_new_n24483__, new_new_n24484__,
    new_new_n24485__, new_new_n24486__, new_new_n24487__, new_new_n24488__,
    new_new_n24489__, new_new_n24490__, new_new_n24491__, new_new_n24492__,
    new_new_n24493__, new_new_n24494__, new_new_n24495__, new_new_n24496__,
    new_new_n24497__, new_new_n24498__, new_new_n24499__, new_new_n24500__,
    new_new_n24501__, new_new_n24502__, new_new_n24503__, new_new_n24504__,
    new_new_n24505__, new_new_n24506__, new_new_n24507__, new_new_n24508__,
    new_new_n24509__, new_new_n24510__, new_new_n24511__, new_new_n24512__,
    new_new_n24513__, new_new_n24514__, new_new_n24515__, new_new_n24516__,
    new_new_n24517__, new_new_n24518__, new_new_n24519__, new_new_n24520__,
    new_new_n24521__, new_new_n24522__, new_new_n24523__, new_new_n24524__,
    new_new_n24525__, new_new_n24526__, new_new_n24527__, new_new_n24528__,
    new_new_n24529__, new_new_n24530__, new_new_n24531__, new_new_n24532__,
    new_new_n24533__, new_new_n24534__, new_new_n24535__, new_new_n24536__,
    new_new_n24537__, new_new_n24538__, new_new_n24539__, new_new_n24540__,
    new_new_n24541__, new_new_n24542__, new_new_n24543__, new_new_n24544__,
    new_new_n24545__, new_new_n24546__, new_new_n24547__, new_new_n24548__,
    new_new_n24549__, new_new_n24550__, new_new_n24551__, new_new_n24552__,
    new_new_n24553__, new_new_n24554__, new_new_n24555__, new_new_n24556__,
    new_new_n24557__, new_new_n24558__, new_new_n24559__, new_new_n24560__,
    new_new_n24561__, new_new_n24562__, new_new_n24563__, new_new_n24564__,
    new_new_n24565__, new_new_n24566__, new_new_n24567__, new_new_n24568__,
    new_new_n24569__, new_new_n24570__, new_new_n24571__, new_new_n24572__,
    new_new_n24573__, new_new_n24574__, new_new_n24575__, new_new_n24576__,
    new_new_n24577__, new_new_n24578__, new_new_n24579__, new_new_n24580__,
    new_new_n24581__, new_new_n24582__, new_new_n24583__, new_new_n24584__,
    new_new_n24585__, new_new_n24586__, new_new_n24587__, new_new_n24588__,
    new_new_n24589__, new_new_n24590__, new_new_n24591__, new_new_n24592__,
    new_new_n24593__, new_new_n24594__, new_new_n24595__, new_new_n24596__,
    new_new_n24597__, new_new_n24598__, new_new_n24599__, new_new_n24600__,
    new_new_n24601__, new_new_n24602__, new_new_n24603__, new_new_n24604__,
    new_new_n24605__, new_new_n24606__, new_new_n24607__, new_new_n24608__,
    new_new_n24609__, new_new_n24610__, new_new_n24611__, new_new_n24612__,
    new_new_n24613__, new_new_n24614__, new_new_n24615__, new_new_n24616__,
    new_new_n24617__, new_new_n24618__, new_new_n24619__, new_new_n24620__,
    new_new_n24621__, new_new_n24622__, new_new_n24623__, new_new_n24624__,
    new_new_n24625__, new_new_n24626__, new_new_n24627__, new_new_n24628__,
    new_new_n24629__, new_new_n24630__, new_new_n24631__, new_new_n24632__,
    new_new_n24633__, new_new_n24634__, new_new_n24635__, new_new_n24636__,
    new_new_n24637__, new_new_n24638__, new_new_n24639__, new_new_n24640__,
    new_new_n24641__, new_new_n24642__, new_new_n24643__, new_new_n24644__,
    new_new_n24645__, new_new_n24646__, new_new_n24647__, new_new_n24648__,
    new_new_n24649__, new_new_n24650__, new_new_n24651__, new_new_n24652__,
    new_new_n24653__, new_new_n24654__, new_new_n24655__, new_new_n24656__,
    new_new_n24657__, new_new_n24658__, new_new_n24659__, new_new_n24660__,
    new_new_n24661__, new_new_n24662__, new_new_n24663__, new_new_n24664__,
    new_new_n24665__, new_new_n24666__, new_new_n24667__, new_new_n24668__,
    new_new_n24669__, new_new_n24670__, new_new_n24671__, new_new_n24672__,
    new_new_n24673__, new_new_n24674__, new_new_n24675__, new_new_n24676__,
    new_new_n24677__, new_new_n24678__, new_new_n24679__, new_new_n24680__,
    new_new_n24681__, new_new_n24682__, new_new_n24683__, new_new_n24684__,
    new_new_n24685__, new_new_n24686__, new_new_n24687__, new_new_n24688__,
    new_new_n24689__, new_new_n24690__, new_new_n24691__, new_new_n24692__,
    new_new_n24693__, new_new_n24694__, new_new_n24695__, new_new_n24696__,
    new_new_n24697__, new_new_n24698__, new_new_n24699__, new_new_n24700__,
    new_new_n24701__, new_new_n24702__, new_new_n24703__, new_new_n24704__,
    new_new_n24705__, new_new_n24706__, new_new_n24707__, new_new_n24708__,
    new_new_n24709__, new_new_n24710__, new_new_n24711__, new_new_n24712__,
    new_new_n24713__, new_new_n24714__, new_new_n24715__, new_new_n24716__,
    new_new_n24717__, new_new_n24718__, new_new_n24719__, new_new_n24720__,
    new_new_n24721__, new_new_n24722__, new_new_n24723__, new_new_n24724__,
    new_new_n24725__, new_new_n24726__, new_new_n24727__, new_new_n24728__,
    new_new_n24729__, new_new_n24730__, new_new_n24731__, new_new_n24732__,
    new_new_n24733__, new_new_n24734__, new_new_n24735__, new_new_n24736__,
    new_new_n24737__, new_new_n24738__, new_new_n24739__, new_new_n24740__,
    new_new_n24741__, new_new_n24742__, new_new_n24743__, new_new_n24744__,
    new_new_n24745__, new_new_n24746__, new_new_n24747__, new_new_n24748__,
    new_new_n24749__, new_new_n24750__, new_new_n24751__, new_new_n24752__,
    new_new_n24753__, new_new_n24754__, new_new_n24755__, new_new_n24756__,
    new_new_n24757__, new_new_n24758__, new_new_n24759__, new_new_n24760__,
    new_new_n24761__, new_new_n24762__, new_new_n24763__, new_new_n24764__,
    new_new_n24765__, new_new_n24766__, new_new_n24767__, new_new_n24768__,
    new_new_n24769__, new_new_n24770__, new_new_n24771__, new_new_n24772__,
    new_new_n24773__, new_new_n24774__, new_new_n24775__, new_new_n24776__,
    new_new_n24777__, new_new_n24778__, new_new_n24779__, new_new_n24780__,
    new_new_n24781__, new_new_n24782__, new_new_n24783__, new_new_n24784__,
    new_new_n24785__, new_new_n24786__, new_new_n24787__, new_new_n24788__,
    new_new_n24789__, new_new_n24790__, new_new_n24791__, new_new_n24792__,
    new_new_n24793__, new_new_n24794__, new_new_n24795__, new_new_n24796__,
    new_new_n24797__, new_new_n24798__, new_new_n24799__, new_new_n24800__,
    new_new_n24801__, new_new_n24802__, new_new_n24803__, new_new_n24804__,
    new_new_n24805__, new_new_n24806__, new_new_n24807__, new_new_n24808__,
    new_new_n24809__, new_new_n24810__, new_new_n24811__, new_new_n24812__,
    new_new_n24813__, new_new_n24814__, new_new_n24815__, new_new_n24816__,
    new_new_n24817__, new_new_n24818__, new_new_n24819__, new_new_n24820__,
    new_new_n24821__, new_new_n24822__, new_new_n24823__, new_new_n24824__,
    new_new_n24825__, new_new_n24826__, new_new_n24827__, new_new_n24828__,
    new_new_n24829__, new_new_n24830__, new_new_n24831__, new_new_n24832__,
    new_new_n24833__, new_new_n24834__, new_new_n24835__, new_new_n24836__,
    new_new_n24837__, new_new_n24838__, new_new_n24839__, new_new_n24840__,
    new_new_n24841__, new_new_n24842__, new_new_n24843__, new_new_n24844__,
    new_new_n24845__, new_new_n24846__, new_new_n24847__, new_new_n24848__,
    new_new_n24849__, new_new_n24850__, new_new_n24851__, new_new_n24852__,
    new_new_n24853__, new_new_n24854__, new_new_n24855__, new_new_n24856__,
    new_new_n24857__, new_new_n24858__, new_new_n24859__, new_new_n24860__,
    new_new_n24861__, new_new_n24862__, new_new_n24863__, new_new_n24864__,
    new_new_n24865__, new_new_n24866__, new_new_n24867__, new_new_n24868__,
    new_new_n24869__, new_new_n24870__, new_new_n24871__, new_new_n24872__,
    new_new_n24873__, new_new_n24874__, new_new_n24875__, new_new_n24876__,
    new_new_n24877__, new_new_n24878__, new_new_n24879__, new_new_n24880__,
    new_new_n24881__, new_new_n24882__, new_new_n24883__, new_new_n24884__,
    new_new_n24885__, new_new_n24886__, new_new_n24887__, new_new_n24888__,
    new_new_n24889__, new_new_n24890__, new_new_n24891__, new_new_n24892__,
    new_new_n24893__, new_new_n24894__, new_new_n24895__, new_new_n24896__,
    new_new_n24897__, new_new_n24898__, new_new_n24899__, new_new_n24900__,
    new_new_n24901__, new_new_n24902__, new_new_n24903__, new_new_n24904__,
    new_new_n24905__, new_new_n24906__, new_new_n24907__, new_new_n24908__,
    new_new_n24909__, new_new_n24910__, new_new_n24911__, new_new_n24912__,
    new_new_n24913__, new_new_n24914__, new_new_n24915__, new_new_n24916__,
    new_new_n24917__, new_new_n24918__, new_new_n24919__, new_new_n24920__,
    new_new_n24921__, new_new_n24922__, new_new_n24923__, new_new_n24924__,
    new_new_n24925__, new_new_n24926__, new_new_n24927__, new_new_n24928__,
    new_new_n24929__, new_new_n24930__, new_new_n24931__, new_new_n24932__,
    new_new_n24933__, new_new_n24934__, new_new_n24935__, new_new_n24936__,
    new_new_n24937__, new_new_n24938__, new_new_n24939__, new_new_n24940__,
    new_new_n24941__, new_new_n24942__, new_new_n24943__, new_new_n24944__,
    new_new_n24945__, new_new_n24946__, new_new_n24947__, new_new_n24948__,
    new_new_n24949__, new_new_n24950__, new_new_n24951__, new_new_n24952__,
    new_new_n24953__, new_new_n24954__, new_new_n24955__, new_new_n24956__,
    new_new_n24957__, new_new_n24958__, new_new_n24959__, new_new_n24960__,
    new_new_n24961__, new_new_n24962__, new_new_n24963__, new_new_n24964__,
    new_new_n24965__, new_new_n24966__, new_new_n24967__, new_new_n24968__,
    new_new_n24969__, new_new_n24970__, new_new_n24971__, new_new_n24972__,
    new_new_n24973__, new_new_n24974__, new_new_n24975__, new_new_n24976__,
    new_new_n24977__, new_new_n24978__, new_new_n24979__, new_new_n24980__,
    new_new_n24981__, new_new_n24982__, new_new_n24983__, new_new_n24984__,
    new_new_n24985__, new_new_n24986__, new_new_n24987__, new_new_n24988__,
    new_new_n24989__, new_new_n24990__, new_new_n24991__, new_new_n24992__,
    new_new_n24993__, new_new_n24994__, new_new_n24995__, new_new_n24996__,
    new_new_n24997__, new_new_n24998__, new_new_n24999__, new_new_n25000__,
    new_new_n25001__, new_new_n25002__, new_new_n25003__, new_new_n25004__,
    new_new_n25005__, new_new_n25006__, new_new_n25007__, new_new_n25008__,
    new_new_n25009__, new_new_n25010__, new_new_n25011__, new_new_n25012__,
    new_new_n25013__, new_new_n25014__, new_new_n25015__, new_new_n25016__,
    new_new_n25017__, new_new_n25018__, new_new_n25019__, new_new_n25020__,
    new_new_n25021__, new_new_n25022__, new_new_n25023__, new_new_n25024__,
    new_new_n25025__, new_new_n25026__, new_new_n25027__, new_new_n25028__,
    new_new_n25029__, new_new_n25030__, new_new_n25031__, new_new_n25032__,
    new_new_n25033__, new_new_n25034__, new_new_n25035__, new_new_n25036__,
    new_new_n25037__, new_new_n25038__, new_new_n25039__, new_new_n25040__,
    new_new_n25041__, new_new_n25042__, new_new_n25043__, new_new_n25044__,
    new_new_n25045__, new_new_n25046__, new_new_n25047__, new_new_n25048__,
    new_new_n25049__, new_new_n25050__, new_new_n25051__, new_new_n25052__,
    new_new_n25053__, new_new_n25054__, new_new_n25055__, new_new_n25056__,
    new_new_n25057__, new_new_n25058__, new_new_n25059__, new_new_n25060__,
    new_new_n25061__, new_new_n25062__, new_new_n25063__, new_new_n25064__,
    new_new_n25065__, new_new_n25066__, new_new_n25067__, new_new_n25068__,
    new_new_n25069__, new_new_n25070__, new_new_n25071__, new_new_n25072__,
    new_new_n25073__, new_new_n25074__, new_new_n25075__, new_new_n25076__,
    new_new_n25077__, new_new_n25078__, new_new_n25079__, new_new_n25080__,
    new_new_n25081__, new_new_n25082__, new_new_n25083__, new_new_n25084__,
    new_new_n25085__, new_new_n25086__, new_new_n25087__, new_new_n25088__,
    new_new_n25089__, new_new_n25090__, new_new_n25091__, new_new_n25092__,
    new_new_n25093__, new_new_n25094__, new_new_n25095__, new_new_n25096__,
    new_new_n25097__, new_new_n25098__, new_new_n25099__, new_new_n25100__,
    new_new_n25101__, new_new_n25102__, new_new_n25103__, new_new_n25104__,
    new_new_n25105__, new_new_n25106__, new_new_n25107__, new_new_n25108__,
    new_new_n25109__, new_new_n25110__, new_new_n25111__, new_new_n25112__,
    new_new_n25113__, new_new_n25114__, new_new_n25115__, new_new_n25116__,
    new_new_n25117__, new_new_n25118__, new_new_n25119__, new_new_n25120__,
    new_new_n25121__, new_new_n25122__, new_new_n25123__, new_new_n25124__,
    new_new_n25125__, new_new_n25126__, new_new_n25127__, new_new_n25128__,
    new_new_n25129__, new_new_n25130__, new_new_n25131__, new_new_n25132__,
    new_new_n25133__, new_new_n25134__, new_new_n25135__, new_new_n25136__,
    new_new_n25137__, new_new_n25138__, new_new_n25139__, new_new_n25140__,
    new_new_n25141__, new_new_n25142__, new_new_n25143__, new_new_n25144__,
    new_new_n25145__, new_new_n25146__, new_new_n25147__, new_new_n25148__,
    new_new_n25149__, new_new_n25150__, new_new_n25151__, new_new_n25152__,
    new_new_n25153__, new_new_n25154__, new_new_n25155__, new_new_n25156__,
    new_new_n25157__, new_new_n25158__, new_new_n25159__, new_new_n25160__,
    new_new_n25161__, new_new_n25162__, new_new_n25163__, new_new_n25164__,
    new_new_n25165__, new_new_n25166__, new_new_n25167__, new_new_n25168__,
    new_new_n25169__, new_new_n25170__, new_new_n25171__, new_new_n25172__,
    new_new_n25173__, new_new_n25174__, new_new_n25175__, new_new_n25176__,
    new_new_n25177__, new_new_n25178__, new_new_n25179__, new_new_n25180__,
    new_new_n25181__, new_new_n25182__, new_new_n25183__, new_new_n25184__,
    new_new_n25185__, new_new_n25186__, new_new_n25187__, new_new_n25188__,
    new_new_n25189__, new_new_n25190__, new_new_n25191__, new_new_n25192__,
    new_new_n25193__, new_new_n25194__, new_new_n25195__, new_new_n25196__,
    new_new_n25197__, new_new_n25198__, new_new_n25199__, new_new_n25200__,
    new_new_n25201__, new_new_n25202__, new_new_n25203__, new_new_n25204__,
    new_new_n25205__, new_new_n25206__, new_new_n25207__, new_new_n25208__,
    new_new_n25209__, new_new_n25210__, new_new_n25211__, new_new_n25212__,
    new_new_n25213__, new_new_n25214__, new_new_n25215__, new_new_n25216__,
    new_new_n25217__, new_new_n25218__, new_new_n25219__, new_new_n25220__,
    new_new_n25221__, new_new_n25222__, new_new_n25223__, new_new_n25224__,
    new_new_n25225__, new_new_n25226__, new_new_n25227__, new_new_n25228__,
    new_new_n25229__, new_new_n25230__, new_new_n25231__, new_new_n25232__,
    new_new_n25233__, new_new_n25234__, new_new_n25235__, new_new_n25236__,
    new_new_n25237__, new_new_n25238__, new_new_n25239__, new_new_n25240__,
    new_new_n25241__, new_new_n25242__, new_new_n25243__, new_new_n25244__,
    new_new_n25245__, new_new_n25246__, new_new_n25247__, new_new_n25248__,
    new_new_n25249__, new_new_n25250__, new_new_n25251__, new_new_n25252__,
    new_new_n25253__, new_new_n25254__, new_new_n25255__, new_new_n25256__,
    new_new_n25257__, new_new_n25258__, new_new_n25259__, new_new_n25260__,
    new_new_n25261__, new_new_n25262__, new_new_n25263__, new_new_n25264__,
    new_new_n25265__, new_new_n25266__, new_new_n25267__, new_new_n25268__,
    new_new_n25269__, new_new_n25270__, new_new_n25271__, new_new_n25272__,
    new_new_n25273__, new_new_n25274__, new_new_n25275__, new_new_n25276__,
    new_new_n25277__, new_new_n25278__, new_new_n25279__, new_new_n25280__,
    new_new_n25281__, new_new_n25282__, new_new_n25283__, new_new_n25284__,
    new_new_n25285__, new_new_n25286__, new_new_n25287__, new_new_n25288__,
    new_new_n25289__, new_new_n25290__, new_new_n25291__, new_new_n25292__,
    new_new_n25293__, new_new_n25294__, new_new_n25295__, new_new_n25296__,
    new_new_n25297__, new_new_n25298__, new_new_n25299__, new_new_n25300__,
    new_new_n25301__, new_new_n25302__, new_new_n25303__, new_new_n25304__,
    new_new_n25305__, new_new_n25306__, new_new_n25307__, new_new_n25308__,
    new_new_n25309__, new_new_n25310__, new_new_n25311__, new_new_n25312__,
    new_new_n25313__, new_new_n25314__, new_new_n25315__, new_new_n25316__,
    new_new_n25317__, new_new_n25318__, new_new_n25319__, new_new_n25320__,
    new_new_n25321__, new_new_n25322__, new_new_n25323__, new_new_n25324__,
    new_new_n25325__, new_new_n25326__, new_new_n25327__, new_new_n25328__,
    new_new_n25329__, new_new_n25330__, new_new_n25331__, new_new_n25332__,
    new_new_n25333__, new_new_n25334__, new_new_n25335__, new_new_n25336__,
    new_new_n25337__, new_new_n25338__, new_new_n25339__, new_new_n25340__,
    new_new_n25341__, new_new_n25342__, new_new_n25343__, new_new_n25344__,
    new_new_n25345__, new_new_n25346__, new_new_n25347__, new_new_n25348__,
    new_new_n25349__, new_new_n25350__, new_new_n25351__, new_new_n25352__,
    new_new_n25353__, new_new_n25354__, new_new_n25355__, new_new_n25356__,
    new_new_n25357__, new_new_n25358__, new_new_n25359__, new_new_n25360__,
    new_new_n25361__, new_new_n25362__, new_new_n25363__, new_new_n25364__,
    new_new_n25365__, new_new_n25366__, new_new_n25367__, new_new_n25368__,
    new_new_n25369__, new_new_n25370__, new_new_n25371__, new_new_n25372__,
    new_new_n25373__, new_new_n25374__, new_new_n25375__, new_new_n25376__,
    new_new_n25377__, new_new_n25378__, new_new_n25379__, new_new_n25380__,
    new_new_n25381__, new_new_n25382__, new_new_n25383__, new_new_n25384__,
    new_new_n25385__, new_new_n25386__, new_new_n25387__, new_new_n25388__,
    new_new_n25389__, new_new_n25390__, new_new_n25391__, new_new_n25392__,
    new_new_n25393__, new_new_n25394__, new_new_n25395__, new_new_n25396__,
    new_new_n25397__, new_new_n25398__, new_new_n25399__, new_new_n25400__,
    new_new_n25401__, new_new_n25402__, new_new_n25403__, new_new_n25404__,
    new_new_n25405__, new_new_n25406__, new_new_n25407__, new_new_n25408__,
    new_new_n25409__, new_new_n25410__, new_new_n25411__, new_new_n25412__,
    new_new_n25413__, new_new_n25414__, new_new_n25415__, new_new_n25416__,
    new_new_n25417__, new_new_n25418__, new_new_n25419__, new_new_n25420__,
    new_new_n25421__, new_new_n25422__, new_new_n25423__, new_new_n25424__,
    new_new_n25425__, new_new_n25426__, new_new_n25427__, new_new_n25428__,
    new_new_n25429__, new_new_n25430__, new_new_n25431__, new_new_n25432__,
    new_new_n25433__, new_new_n25434__, new_new_n25435__, new_new_n25436__,
    new_new_n25437__, new_new_n25438__, new_new_n25439__, new_new_n25440__,
    new_new_n25441__, new_new_n25442__, new_new_n25443__, new_new_n25444__,
    new_new_n25445__, new_new_n25446__, new_new_n25447__, new_new_n25448__,
    new_new_n25449__, new_new_n25450__, new_new_n25451__, new_new_n25452__,
    new_new_n25453__, new_new_n25454__, new_new_n25455__, new_new_n25456__,
    new_new_n25457__, new_new_n25458__, new_new_n25459__, new_new_n25460__,
    new_new_n25461__, new_new_n25462__, new_new_n25463__, new_new_n25464__,
    new_new_n25465__, new_new_n25466__, new_new_n25467__, new_new_n25468__,
    new_new_n25469__, new_new_n25470__, new_new_n25471__, new_new_n25472__,
    new_new_n25473__, new_new_n25474__, new_new_n25475__, new_new_n25476__,
    new_new_n25477__, new_new_n25478__, new_new_n25479__, new_new_n25480__,
    new_new_n25481__, new_new_n25482__, new_new_n25483__, new_new_n25484__,
    new_new_n25485__, new_new_n25486__, new_new_n25487__, new_new_n25488__,
    new_new_n25489__, new_new_n25490__, new_new_n25491__, new_new_n25492__,
    new_new_n25493__, new_new_n25494__, new_new_n25495__, new_new_n25496__,
    new_new_n25497__, new_new_n25498__, new_new_n25499__, new_new_n25500__,
    new_new_n25501__, new_new_n25502__, new_new_n25503__, new_new_n25504__,
    new_new_n25505__, new_new_n25506__, new_new_n25507__, new_new_n25508__,
    new_new_n25509__, new_new_n25510__, new_new_n25511__, new_new_n25512__,
    new_new_n25513__, new_new_n25514__, new_new_n25515__, new_new_n25516__,
    new_new_n25517__, new_new_n25518__, new_new_n25519__, new_new_n25520__,
    new_new_n25521__, new_new_n25522__, new_new_n25523__, new_new_n25524__,
    new_new_n25525__, new_new_n25526__, new_new_n25527__, new_new_n25528__,
    new_new_n25529__, new_new_n25530__, new_new_n25531__, new_new_n25532__,
    new_new_n25533__, new_new_n25534__, new_new_n25535__, new_new_n25536__,
    new_new_n25537__, new_new_n25538__, new_new_n25539__, new_new_n25540__,
    new_new_n25541__, new_new_n25542__, new_new_n25543__, new_new_n25544__,
    new_new_n25545__, new_new_n25546__, new_new_n25547__, new_new_n25548__,
    new_new_n25549__, new_new_n25550__, new_new_n25551__, new_new_n25552__,
    new_new_n25553__, new_new_n25554__, new_new_n25555__, new_new_n25556__,
    new_new_n25557__, new_new_n25558__, new_new_n25559__, new_new_n25560__,
    new_new_n25561__, new_new_n25562__, new_new_n25563__, new_new_n25564__,
    new_new_n25565__, new_new_n25566__, new_new_n25567__, new_new_n25568__,
    new_new_n25569__, new_new_n25570__, new_new_n25571__, new_new_n25572__,
    new_new_n25573__, new_new_n25574__, new_new_n25575__, new_new_n25576__,
    new_new_n25577__, new_new_n25578__, new_new_n25579__, new_new_n25580__,
    new_new_n25581__, new_new_n25582__, new_new_n25583__, new_new_n25584__,
    new_new_n25585__, new_new_n25586__, new_new_n25587__, new_new_n25588__,
    new_new_n25589__, new_new_n25590__, new_new_n25591__, new_new_n25592__,
    new_new_n25593__, new_new_n25594__, new_new_n25595__, new_new_n25596__,
    new_new_n25597__, new_new_n25598__, new_new_n25599__, new_new_n25600__,
    new_new_n25601__, new_new_n25602__, new_new_n25603__, new_new_n25604__,
    new_new_n25605__, new_new_n25606__, new_new_n25607__, new_new_n25608__,
    new_new_n25609__, new_new_n25610__, new_new_n25611__, new_new_n25612__,
    new_new_n25613__, new_new_n25614__, new_new_n25615__, new_new_n25616__,
    new_new_n25617__, new_new_n25618__, new_new_n25619__, new_new_n25620__,
    new_new_n25621__, new_new_n25622__, new_new_n25623__, new_new_n25624__,
    new_new_n25625__, new_new_n25626__, new_new_n25627__, new_new_n25628__,
    new_new_n25629__, new_new_n25630__, new_new_n25631__, new_new_n25632__,
    new_new_n25633__, new_new_n25634__, new_new_n25635__, new_new_n25636__,
    new_new_n25637__, new_new_n25638__, new_new_n25639__, new_new_n25640__,
    new_new_n25641__, new_new_n25642__, new_new_n25643__, new_new_n25644__,
    new_new_n25645__, new_new_n25646__, new_new_n25647__, new_new_n25648__,
    new_new_n25649__, new_new_n25650__, new_new_n25651__, new_new_n25652__,
    new_new_n25653__, new_new_n25654__, new_new_n25655__, new_new_n25656__,
    new_new_n25657__, new_new_n25658__, new_new_n25659__, new_new_n25660__,
    new_new_n25661__, new_new_n25662__, new_new_n25663__, new_new_n25664__,
    new_new_n25665__, new_new_n25666__, new_new_n25667__, new_new_n25668__,
    new_new_n25669__, new_new_n25670__, new_new_n25671__, new_new_n25672__,
    new_new_n25673__, new_new_n25674__, new_new_n25675__, new_new_n25676__,
    new_new_n25677__, new_new_n25678__, new_new_n25679__, new_new_n25680__,
    new_new_n25681__, new_new_n25682__, new_new_n25683__, new_new_n25684__,
    new_new_n25685__, new_new_n25686__, new_new_n25687__, new_new_n25688__,
    new_new_n25689__, new_new_n25690__, new_new_n25691__, new_new_n25692__,
    new_new_n25693__, new_new_n25694__, new_new_n25695__, new_new_n25696__,
    new_new_n25697__, new_new_n25698__, new_new_n25699__, new_new_n25700__,
    new_new_n25701__, new_new_n25702__, new_new_n25703__, new_new_n25704__,
    new_new_n25705__, new_new_n25706__, new_new_n25707__, new_new_n25708__,
    new_new_n25709__, new_new_n25710__, new_new_n25711__, new_new_n25712__,
    new_new_n25713__, new_new_n25714__, new_new_n25715__, new_new_n25716__,
    new_new_n25717__, new_new_n25718__, new_new_n25719__, new_new_n25720__,
    new_new_n25721__, new_new_n25722__, new_new_n25723__, new_new_n25724__,
    new_new_n25725__, new_new_n25726__, new_new_n25727__, new_new_n25728__,
    new_new_n25729__, new_new_n25730__, new_new_n25731__, new_new_n25732__,
    new_new_n25733__, new_new_n25734__, new_new_n25735__, new_new_n25736__,
    new_new_n25737__, new_new_n25738__, new_new_n25739__, new_new_n25740__,
    new_new_n25741__, new_new_n25742__, new_new_n25743__, new_new_n25744__,
    new_new_n25745__, new_new_n25746__, new_new_n25747__, new_new_n25748__,
    new_new_n25749__, new_new_n25750__, new_new_n25751__, new_new_n25752__,
    new_new_n25753__, new_new_n25754__, new_new_n25755__, new_new_n25756__,
    new_new_n25757__, new_new_n25758__, new_new_n25759__, new_new_n25760__,
    new_new_n25761__, new_new_n25762__, new_new_n25763__, new_new_n25764__,
    new_new_n25765__, new_new_n25766__, new_new_n25767__, new_new_n25768__,
    new_new_n25769__, new_new_n25770__, new_new_n25771__, new_new_n25772__,
    new_new_n25773__, new_new_n25774__, new_new_n25775__, new_new_n25776__,
    new_new_n25777__, new_new_n25778__, new_new_n25779__, new_new_n25780__,
    new_new_n25781__, new_new_n25782__, new_new_n25783__, new_new_n25784__,
    new_new_n25785__, new_new_n25786__, new_new_n25787__, new_new_n25788__,
    new_new_n25789__, new_new_n25790__, new_new_n25791__, new_new_n25792__,
    new_new_n25793__, new_new_n25794__, new_new_n25795__, new_new_n25796__,
    new_new_n25797__, new_new_n25798__, new_new_n25799__, new_new_n25800__,
    new_new_n25801__, new_new_n25802__, new_new_n25803__, new_new_n25804__,
    new_new_n25805__, new_new_n25806__, new_new_n25807__, new_new_n25808__,
    new_new_n25809__, new_new_n25810__, new_new_n25811__, new_new_n25812__,
    new_new_n25813__, new_new_n25814__, new_new_n25815__, new_new_n25816__,
    new_new_n25817__, new_new_n25818__, new_new_n25819__, new_new_n25820__,
    new_new_n25821__, new_new_n25822__, new_new_n25823__, new_new_n25824__,
    new_new_n25825__, new_new_n25826__, new_new_n25827__, new_new_n25828__,
    new_new_n25829__, new_new_n25830__, new_new_n25831__, new_new_n25832__,
    new_new_n25833__, new_new_n25834__, new_new_n25835__, new_new_n25836__,
    new_new_n25837__, new_new_n25838__, new_new_n25839__, new_new_n25840__,
    new_new_n25841__, new_new_n25842__, new_new_n25843__, new_new_n25844__,
    new_new_n25845__, new_new_n25846__, new_new_n25847__, new_new_n25848__,
    new_new_n25849__, new_new_n25850__, new_new_n25851__, new_new_n25852__,
    new_new_n25853__, new_new_n25854__, new_new_n25855__, new_new_n25856__,
    new_new_n25857__, new_new_n25858__, new_new_n25859__, new_new_n25860__,
    new_new_n25861__, new_new_n25862__, new_new_n25863__, new_new_n25864__,
    new_new_n25865__, new_new_n25866__, new_new_n25867__, new_new_n25868__,
    new_new_n25869__, new_new_n25870__, new_new_n25871__, new_new_n25872__,
    new_new_n25873__, new_new_n25874__, new_new_n25875__, new_new_n25876__,
    new_new_n25877__, new_new_n25878__, new_new_n25879__, new_new_n25880__,
    new_new_n25881__, new_new_n25882__, new_new_n25883__, new_new_n25884__,
    new_new_n25885__, new_new_n25886__, new_new_n25887__, new_new_n25888__,
    new_new_n25889__, new_new_n25890__, new_new_n25891__, new_new_n25892__,
    new_new_n25893__, new_new_n25894__, new_new_n25895__, new_new_n25896__,
    new_new_n25897__, new_new_n25898__, new_new_n25899__, new_new_n25900__,
    new_new_n25901__, new_new_n25902__, new_new_n25903__, new_new_n25904__,
    new_new_n25905__, new_new_n25906__, new_new_n25907__, new_new_n25908__,
    new_new_n25909__, new_new_n25910__, new_new_n25911__, new_new_n25912__,
    new_new_n25913__, new_new_n25914__, new_new_n25915__, new_new_n25916__,
    new_new_n25917__, new_new_n25918__, new_new_n25919__, new_new_n25920__,
    new_new_n25921__, new_new_n25922__, new_new_n25923__, new_new_n25924__,
    new_new_n25925__, new_new_n25926__, new_new_n25927__, new_new_n25928__,
    new_new_n25929__, new_new_n25930__, new_new_n25931__, new_new_n25932__,
    new_new_n25933__, new_new_n25934__, new_new_n25935__, new_new_n25936__,
    new_new_n25937__, new_new_n25938__, new_new_n25939__, new_new_n25940__,
    new_new_n25941__, new_new_n25942__, new_new_n25943__, new_new_n25944__,
    new_new_n25945__, new_new_n25946__, new_new_n25947__, new_new_n25948__,
    new_new_n25949__, new_new_n25950__, new_new_n25951__, new_new_n25952__,
    new_new_n25953__, new_new_n25954__, new_new_n25955__, new_new_n25956__,
    new_new_n25957__, new_new_n25958__, new_new_n25959__, new_new_n25960__,
    new_new_n25961__, new_new_n25962__, new_new_n25963__, new_new_n25964__,
    new_new_n25965__, new_new_n25966__, new_new_n25967__, new_new_n25968__,
    new_new_n25969__, new_new_n25970__, new_new_n25971__, new_new_n25972__,
    new_new_n25973__, new_new_n25974__, new_new_n25975__, new_new_n25976__,
    new_new_n25977__, new_new_n25978__, new_new_n25979__, new_new_n25980__,
    new_new_n25981__, new_new_n25982__, new_new_n25983__, new_new_n25984__,
    new_new_n25985__, new_new_n25986__, new_new_n25987__, new_new_n25988__,
    new_new_n25989__, new_new_n25990__, new_new_n25991__, new_new_n25992__,
    new_new_n25993__, new_new_n25994__, new_new_n25995__, new_new_n25996__,
    new_new_n25997__, new_new_n25998__, new_new_n25999__, new_new_n26000__,
    new_new_n26001__, new_new_n26002__, new_new_n26003__, new_new_n26004__,
    new_new_n26005__, new_new_n26006__, new_new_n26007__, new_new_n26008__,
    new_new_n26009__, new_new_n26010__, new_new_n26011__, new_new_n26012__,
    new_new_n26013__, new_new_n26014__, new_new_n26015__, new_new_n26016__,
    new_new_n26017__, new_new_n26018__, new_new_n26019__, new_new_n26020__,
    new_new_n26021__, new_new_n26022__, new_new_n26023__, new_new_n26024__,
    new_new_n26025__, new_new_n26026__, new_new_n26027__, new_new_n26028__,
    new_new_n26029__, new_new_n26030__, new_new_n26031__, new_new_n26032__,
    new_new_n26033__, new_new_n26034__, new_new_n26035__, new_new_n26036__,
    new_new_n26037__, new_new_n26038__, new_new_n26039__, new_new_n26040__,
    new_new_n26041__, new_new_n26042__, new_new_n26043__, new_new_n26044__,
    new_new_n26045__, new_new_n26046__, new_new_n26047__, new_new_n26048__,
    new_new_n26049__, new_new_n26050__, new_new_n26051__, new_new_n26052__,
    new_new_n26053__, new_new_n26054__, new_new_n26055__, new_new_n26056__,
    new_new_n26057__, new_new_n26058__, new_new_n26059__, new_new_n26060__,
    new_new_n26061__, new_new_n26062__, new_new_n26063__, new_new_n26064__,
    new_new_n26065__, new_new_n26066__, new_new_n26067__, new_new_n26068__,
    new_new_n26069__, new_new_n26070__, new_new_n26071__, new_new_n26072__,
    new_new_n26073__, new_new_n26074__, new_new_n26075__, new_new_n26076__,
    new_new_n26077__, new_new_n26078__, new_new_n26079__, new_new_n26080__,
    new_new_n26081__, new_new_n26082__, new_new_n26083__, new_new_n26084__,
    new_new_n26085__, new_new_n26086__, new_new_n26087__, new_new_n26088__,
    new_new_n26089__, new_new_n26090__, new_new_n26091__, new_new_n26092__,
    new_new_n26093__, new_new_n26094__, new_new_n26095__, new_new_n26096__,
    new_new_n26097__, new_new_n26098__, new_new_n26099__, new_new_n26100__,
    new_new_n26101__, new_new_n26102__, new_new_n26103__, new_new_n26104__,
    new_new_n26105__, new_new_n26106__, new_new_n26107__, new_new_n26108__,
    new_new_n26109__, new_new_n26110__, new_new_n26111__, new_new_n26112__,
    new_new_n26113__, new_new_n26114__, new_new_n26115__, new_new_n26116__,
    new_new_n26117__, new_new_n26118__, new_new_n26119__, new_new_n26120__,
    new_new_n26121__, new_new_n26122__, new_new_n26123__, new_new_n26124__,
    new_new_n26125__, new_new_n26126__, new_new_n26127__, new_new_n26128__,
    new_new_n26129__, new_new_n26130__, new_new_n26131__, new_new_n26132__,
    new_new_n26133__, new_new_n26134__, new_new_n26135__, new_new_n26136__,
    new_new_n26137__, new_new_n26138__, new_new_n26139__, new_new_n26140__,
    new_new_n26141__, new_new_n26142__, new_new_n26143__, new_new_n26144__,
    new_new_n26145__, new_new_n26146__, new_new_n26147__, new_new_n26148__,
    new_new_n26149__, new_new_n26150__, new_new_n26151__, new_new_n26152__,
    new_new_n26153__, new_new_n26154__, new_new_n26155__, new_new_n26156__,
    new_new_n26157__, new_new_n26158__, new_new_n26159__, new_new_n26160__,
    new_new_n26161__, new_new_n26162__, new_new_n26163__, new_new_n26164__,
    new_new_n26165__, new_new_n26166__, new_new_n26167__, new_new_n26168__,
    new_new_n26169__, new_new_n26170__, new_new_n26171__, new_new_n26172__,
    new_new_n26173__, new_new_n26174__, new_new_n26175__, new_new_n26176__,
    new_new_n26177__, new_new_n26178__, new_new_n26179__, new_new_n26180__,
    new_new_n26181__, new_new_n26182__, new_new_n26183__, new_new_n26184__,
    new_new_n26185__, new_new_n26186__, new_new_n26187__, new_new_n26188__,
    new_new_n26189__, new_new_n26190__, new_new_n26191__, new_new_n26192__,
    new_new_n26193__, new_new_n26194__, new_new_n26195__, new_new_n26196__,
    new_new_n26197__, new_new_n26198__, new_new_n26199__, new_new_n26200__,
    new_new_n26201__, new_new_n26202__, new_new_n26203__, new_new_n26204__,
    new_new_n26205__, new_new_n26206__, new_new_n26207__, new_new_n26208__,
    new_new_n26209__, new_new_n26210__, new_new_n26211__, new_new_n26212__,
    new_new_n26213__, new_new_n26214__, new_new_n26215__, new_new_n26216__,
    new_new_n26217__, new_new_n26218__, new_new_n26219__, new_new_n26220__,
    new_new_n26221__, new_new_n26222__, new_new_n26223__, new_new_n26224__,
    new_new_n26225__, new_new_n26226__, new_new_n26227__, new_new_n26228__,
    new_new_n26229__, new_new_n26230__, new_new_n26231__, new_new_n26232__,
    new_new_n26233__, new_new_n26234__, new_new_n26235__, new_new_n26236__,
    new_new_n26237__, new_new_n26238__, new_new_n26239__, new_new_n26240__,
    new_new_n26241__, new_new_n26242__, new_new_n26243__, new_new_n26244__,
    new_new_n26245__, new_new_n26246__, new_new_n26247__, new_new_n26248__,
    new_new_n26249__, new_new_n26250__, new_new_n26251__, new_new_n26252__,
    new_new_n26253__, new_new_n26254__, new_new_n26255__, new_new_n26256__,
    new_new_n26257__, new_new_n26258__, new_new_n26259__, new_new_n26260__,
    new_new_n26261__, new_new_n26262__, new_new_n26263__, new_new_n26264__,
    new_new_n26265__, new_new_n26266__, new_new_n26267__, new_new_n26268__,
    new_new_n26269__, new_new_n26270__, new_new_n26271__, new_new_n26272__,
    new_new_n26273__, new_new_n26274__, new_new_n26275__, new_new_n26276__,
    new_new_n26277__, new_new_n26278__, new_new_n26279__, new_new_n26280__,
    new_new_n26281__, new_new_n26282__, new_new_n26283__, new_new_n26284__,
    new_new_n26285__, new_new_n26286__, new_new_n26287__, new_new_n26288__,
    new_new_n26289__, new_new_n26290__, new_new_n26291__, new_new_n26292__,
    new_new_n26293__, new_new_n26294__, new_new_n26295__, new_new_n26296__,
    new_new_n26297__, new_new_n26298__, new_new_n26299__, new_new_n26300__,
    new_new_n26301__, new_new_n26302__, new_new_n26303__, new_new_n26304__,
    new_new_n26305__, new_new_n26306__, new_new_n26307__, new_new_n26308__,
    new_new_n26309__, new_new_n26310__, new_new_n26311__, new_new_n26312__,
    new_new_n26313__, new_new_n26314__, new_new_n26315__, new_new_n26316__,
    new_new_n26317__, new_new_n26318__, new_new_n26319__, new_new_n26320__,
    new_new_n26321__, new_new_n26322__, new_new_n26323__, new_new_n26324__,
    new_new_n26325__, new_new_n26326__, new_new_n26327__, new_new_n26328__,
    new_new_n26329__, new_new_n26330__, new_new_n26331__, new_new_n26332__,
    new_new_n26333__, new_new_n26334__, new_new_n26335__, new_new_n26336__,
    new_new_n26337__, new_new_n26338__, new_new_n26339__, new_new_n26340__,
    new_new_n26341__, new_new_n26342__, new_new_n26343__, new_new_n26344__,
    new_new_n26345__, new_new_n26346__, new_new_n26347__, new_new_n26348__,
    new_new_n26349__, new_new_n26350__, new_new_n26351__, new_new_n26352__,
    new_new_n26353__, new_new_n26354__, new_new_n26355__, new_new_n26356__,
    new_new_n26357__, new_new_n26358__, new_new_n26359__, new_new_n26360__,
    new_new_n26361__, new_new_n26362__, new_new_n26363__, new_new_n26364__,
    new_new_n26365__, new_new_n26366__, new_new_n26367__, new_new_n26368__,
    new_new_n26369__, new_new_n26370__, new_new_n26371__, new_new_n26372__,
    new_new_n26373__, new_new_n26374__, new_new_n26375__, new_new_n26376__,
    new_new_n26377__, new_new_n26378__, new_new_n26379__, new_new_n26380__,
    new_new_n26381__, new_new_n26382__, new_new_n26383__, new_new_n26384__,
    new_new_n26385__, new_new_n26386__, new_new_n26387__, new_new_n26388__,
    new_new_n26389__, new_new_n26390__, new_new_n26391__, new_new_n26392__,
    new_new_n26393__, new_new_n26394__, new_new_n26395__, new_new_n26396__,
    new_new_n26397__, new_new_n26398__, new_new_n26399__, new_new_n26400__,
    new_new_n26401__, new_new_n26402__, new_new_n26403__, new_new_n26404__,
    new_new_n26405__, new_new_n26406__, new_new_n26407__, new_new_n26408__,
    new_new_n26409__, new_new_n26410__, new_new_n26411__, new_new_n26412__,
    new_new_n26413__, new_new_n26414__, new_new_n26415__, new_new_n26416__,
    new_new_n26417__, new_new_n26418__, new_new_n26419__, new_new_n26420__,
    new_new_n26421__, new_new_n26422__, new_new_n26423__, new_new_n26424__,
    new_new_n26425__, new_new_n26426__, new_new_n26427__, new_new_n26428__,
    new_new_n26429__, new_new_n26430__, new_new_n26431__, new_new_n26432__,
    new_new_n26433__, new_new_n26434__, new_new_n26435__, new_new_n26436__,
    new_new_n26437__, new_new_n26438__, new_new_n26439__, new_new_n26440__,
    new_new_n26441__, new_new_n26442__, new_new_n26443__, new_new_n26444__,
    new_new_n26445__, new_new_n26446__, new_new_n26447__, new_new_n26448__,
    new_new_n26449__, new_new_n26450__, new_new_n26451__, new_new_n26452__,
    new_new_n26453__, new_new_n26454__, new_new_n26455__, new_new_n26456__,
    new_new_n26457__, new_new_n26458__, new_new_n26459__, new_new_n26460__,
    new_new_n26461__, new_new_n26462__, new_new_n26463__, new_new_n26464__,
    new_new_n26465__, new_new_n26466__, new_new_n26467__, new_new_n26468__,
    new_new_n26469__, new_new_n26470__, new_new_n26471__, new_new_n26472__,
    new_new_n26473__, new_new_n26474__, new_new_n26475__, new_new_n26476__,
    new_new_n26477__, new_new_n26478__, new_new_n26479__, new_new_n26480__,
    new_new_n26481__, new_new_n26482__, new_new_n26483__, new_new_n26484__,
    new_new_n26485__, new_new_n26486__, new_new_n26487__, new_new_n26488__,
    new_new_n26489__, new_new_n26490__, new_new_n26491__, new_new_n26492__,
    new_new_n26493__, new_new_n26494__, new_new_n26495__, new_new_n26496__,
    new_new_n26497__, new_new_n26498__, new_new_n26499__, new_new_n26500__,
    new_new_n26501__, new_new_n26502__, new_new_n26503__, new_new_n26504__,
    new_new_n26505__, new_new_n26506__, new_new_n26507__, new_new_n26508__,
    new_new_n26509__, new_new_n26510__, new_new_n26511__, new_new_n26512__,
    new_new_n26513__, new_new_n26514__, new_new_n26515__, new_new_n26516__,
    new_new_n26517__, new_new_n26518__, new_new_n26519__, new_new_n26520__,
    new_new_n26521__, new_new_n26522__, new_new_n26523__, new_new_n26524__,
    new_new_n26525__, new_new_n26526__, new_new_n26527__, new_new_n26528__,
    new_new_n26529__, new_new_n26530__, new_new_n26531__, new_new_n26532__,
    new_new_n26533__, new_new_n26534__, new_new_n26535__, new_new_n26536__,
    new_new_n26537__, new_new_n26538__, new_new_n26539__, new_new_n26540__,
    new_new_n26541__, new_new_n26542__, new_new_n26543__, new_new_n26544__,
    new_new_n26545__, new_new_n26546__, new_new_n26547__, new_new_n26548__,
    new_new_n26549__, new_new_n26550__, new_new_n26551__, new_new_n26552__,
    new_new_n26553__, new_new_n26554__, new_new_n26555__, new_new_n26556__,
    new_new_n26557__, new_new_n26558__, new_new_n26559__, new_new_n26560__,
    new_new_n26561__, new_new_n26562__, new_new_n26563__, new_new_n26564__,
    new_new_n26565__, new_new_n26566__, new_new_n26567__, new_new_n26568__,
    new_new_n26569__, new_new_n26570__, new_new_n26571__, new_new_n26572__,
    new_new_n26573__, new_new_n26574__, new_new_n26575__, new_new_n26576__,
    new_new_n26577__, new_new_n26578__, new_new_n26579__, new_new_n26580__,
    new_new_n26581__, new_new_n26582__, new_new_n26583__, new_new_n26584__,
    new_new_n26585__, new_new_n26586__, new_new_n26587__, new_new_n26588__,
    new_new_n26589__, new_new_n26590__, new_new_n26591__, new_new_n26592__,
    new_new_n26593__, new_new_n26594__, new_new_n26595__, new_new_n26596__,
    new_new_n26597__, new_new_n26598__, new_new_n26599__, new_new_n26600__,
    new_new_n26601__, new_new_n26602__, new_new_n26603__, new_new_n26604__,
    new_new_n26605__, new_new_n26606__, new_new_n26607__, new_new_n26608__,
    new_new_n26609__, new_new_n26610__, new_new_n26611__, new_new_n26612__,
    new_new_n26613__, new_new_n26614__, new_new_n26615__, new_new_n26616__,
    new_new_n26617__, new_new_n26618__, new_new_n26619__, new_new_n26620__,
    new_new_n26621__, new_new_n26622__, new_new_n26623__, new_new_n26624__,
    new_new_n26625__, new_new_n26626__, new_new_n26627__, new_new_n26628__,
    new_new_n26629__, new_new_n26630__, new_new_n26631__, new_new_n26632__,
    new_new_n26633__, new_new_n26634__, new_new_n26635__, new_new_n26636__,
    new_new_n26637__, new_new_n26638__, new_new_n26639__, new_new_n26640__,
    new_new_n26641__, new_new_n26642__, new_new_n26643__, new_new_n26644__,
    new_new_n26645__, new_new_n26646__, new_new_n26647__, new_new_n26648__,
    new_new_n26649__, new_new_n26650__, new_new_n26651__, new_new_n26652__,
    new_new_n26653__, new_new_n26654__, new_new_n26655__, new_new_n26656__,
    new_new_n26657__, new_new_n26658__, new_new_n26659__, new_new_n26660__,
    new_new_n26661__, new_new_n26662__, new_new_n26663__, new_new_n26664__,
    new_new_n26665__, new_new_n26666__, new_new_n26667__, new_new_n26668__,
    new_new_n26669__, new_new_n26670__, new_new_n26671__, new_new_n26672__,
    new_new_n26673__, new_new_n26674__, new_new_n26675__, new_new_n26676__,
    new_new_n26677__, new_new_n26678__, new_new_n26679__, new_new_n26680__,
    new_new_n26681__, new_new_n26682__, new_new_n26683__, new_new_n26684__,
    new_new_n26685__, new_new_n26686__, new_new_n26687__, new_new_n26688__,
    new_new_n26689__, new_new_n26690__, new_new_n26691__, new_new_n26692__,
    new_new_n26693__, new_new_n26694__, new_new_n26695__, new_new_n26696__,
    new_new_n26697__, new_new_n26698__, new_new_n26699__, new_new_n26700__,
    new_new_n26701__, new_new_n26702__, new_new_n26703__, new_new_n26704__,
    new_new_n26705__, new_new_n26706__, new_new_n26707__, new_new_n26708__,
    new_new_n26709__, new_new_n26710__, new_new_n26711__, new_new_n26712__,
    new_new_n26713__, new_new_n26714__, new_new_n26715__, new_new_n26716__,
    new_new_n26717__, new_new_n26718__, new_new_n26719__, new_new_n26720__,
    new_new_n26721__, new_new_n26722__, new_new_n26723__, new_new_n26724__,
    new_new_n26725__, new_new_n26726__, new_new_n26727__, new_new_n26728__,
    new_new_n26729__, new_new_n26730__, new_new_n26731__, new_new_n26732__,
    new_new_n26733__, new_new_n26734__, new_new_n26735__, new_new_n26736__,
    new_new_n26737__, new_new_n26738__, new_new_n26739__, new_new_n26740__,
    new_new_n26741__, new_new_n26742__, new_new_n26743__, new_new_n26744__,
    new_new_n26745__, new_new_n26746__, new_new_n26747__, new_new_n26748__,
    new_new_n26749__, new_new_n26750__, new_new_n26751__, new_new_n26752__,
    new_new_n26753__, new_new_n26754__, new_new_n26755__, new_new_n26756__,
    new_new_n26757__, new_new_n26758__, new_new_n26759__, new_new_n26760__,
    new_new_n26761__, new_new_n26762__, new_new_n26763__, new_new_n26764__,
    new_new_n26765__, new_new_n26766__, new_new_n26767__, new_new_n26768__,
    new_new_n26769__, new_new_n26770__, new_new_n26771__, new_new_n26772__,
    new_new_n26773__, new_new_n26774__, new_new_n26775__, new_new_n26776__,
    new_new_n26777__, new_new_n26778__, new_new_n26779__, new_new_n26780__,
    new_new_n26781__, new_new_n26782__, new_new_n26783__, new_new_n26784__,
    new_new_n26785__, new_new_n26786__, new_new_n26787__, new_new_n26788__,
    new_new_n26789__, new_new_n26790__, new_new_n26791__, new_new_n26792__,
    new_new_n26793__, new_new_n26794__, new_new_n26795__, new_new_n26796__,
    new_new_n26797__, new_new_n26798__, new_new_n26799__, new_new_n26800__,
    new_new_n26801__, new_new_n26802__, new_new_n26803__, new_new_n26804__,
    new_new_n26805__, new_new_n26806__, new_new_n26807__, new_new_n26808__,
    new_new_n26809__, new_new_n26810__, new_new_n26811__, new_new_n26812__,
    new_new_n26813__, new_new_n26814__, new_new_n26815__, new_new_n26816__,
    new_new_n26817__, new_new_n26818__, new_new_n26819__, new_new_n26820__,
    new_new_n26821__, new_new_n26822__, new_new_n26823__, new_new_n26824__,
    new_new_n26825__, new_new_n26826__, new_new_n26827__, new_new_n26828__,
    new_new_n26829__, new_new_n26830__, new_new_n26831__, new_new_n26832__,
    new_new_n26833__, new_new_n26834__, new_new_n26835__, new_new_n26836__,
    new_new_n26837__, new_new_n26838__, new_new_n26839__, new_new_n26840__,
    new_new_n26841__, new_new_n26842__, new_new_n26843__, new_new_n26844__,
    new_new_n26845__, new_new_n26846__, new_new_n26847__, new_new_n26848__,
    new_new_n26849__, new_new_n26850__, new_new_n26851__, new_new_n26852__,
    new_new_n26853__, new_new_n26854__, new_new_n26855__, new_new_n26856__,
    new_new_n26857__, new_new_n26858__, new_new_n26859__, new_new_n26860__,
    new_new_n26861__, new_new_n26862__, new_new_n26863__, new_new_n26864__,
    new_new_n26865__, new_new_n26866__, new_new_n26867__, new_new_n26868__,
    new_new_n26869__, new_new_n26870__, new_new_n26871__, new_new_n26872__,
    new_new_n26873__, new_new_n26874__, new_new_n26875__, new_new_n26876__,
    new_new_n26877__, new_new_n26878__, new_new_n26879__, new_new_n26880__,
    new_new_n26881__, new_new_n26882__, new_new_n26883__, new_new_n26884__,
    new_new_n26885__, new_new_n26886__, new_new_n26887__, new_new_n26888__,
    new_new_n26889__, new_new_n26890__, new_new_n26891__, new_new_n26892__,
    new_new_n26893__, new_new_n26894__, new_new_n26895__, new_new_n26896__,
    new_new_n26897__, new_new_n26898__, new_new_n26899__, new_new_n26900__,
    new_new_n26901__, new_new_n26902__, new_new_n26903__, new_new_n26904__,
    new_new_n26905__, new_new_n26906__, new_new_n26907__, new_new_n26908__,
    new_new_n26909__, new_new_n26910__, new_new_n26911__, new_new_n26912__,
    new_new_n26913__, new_new_n26914__, new_new_n26915__, new_new_n26916__,
    new_new_n26917__, new_new_n26918__, new_new_n26919__, new_new_n26920__,
    new_new_n26921__, new_new_n26922__, new_new_n26923__, new_new_n26924__,
    new_new_n26925__, new_new_n26926__, new_new_n26927__, new_new_n26928__,
    new_new_n26929__, new_new_n26930__, new_new_n26931__, new_new_n26932__,
    new_new_n26933__, new_new_n26934__, new_new_n26935__, new_new_n26936__,
    new_new_n26937__, new_new_n26938__, new_new_n26939__, new_new_n26940__,
    new_new_n26941__, new_new_n26942__, new_new_n26943__, new_new_n26944__,
    new_new_n26945__, new_new_n26946__, new_new_n26947__, new_new_n26948__,
    new_new_n26949__, new_new_n26950__, new_new_n26951__, new_new_n26952__,
    new_new_n26953__, new_new_n26954__, new_new_n26955__, new_new_n26956__,
    new_new_n26957__, new_new_n26958__, new_new_n26959__, new_new_n26960__,
    new_new_n26961__, new_new_n26962__, new_new_n26963__, new_new_n26964__,
    new_new_n26965__, new_new_n26966__, new_new_n26967__, new_new_n26968__,
    new_new_n26969__, new_new_n26970__, new_new_n26971__, new_new_n26972__,
    new_new_n26973__, new_new_n26974__, new_new_n26975__, new_new_n26976__,
    new_new_n26977__, new_new_n26978__, new_new_n26979__, new_new_n26980__,
    new_new_n26981__, new_new_n26982__, new_new_n26983__, new_new_n26984__,
    new_new_n26985__, new_new_n26986__, new_new_n26987__, new_new_n26988__,
    new_new_n26989__, new_new_n26990__, new_new_n26991__, new_new_n26992__,
    new_new_n26993__, new_new_n26994__, new_new_n26995__, new_new_n26996__,
    new_new_n26997__, new_new_n26998__, new_new_n26999__, new_new_n27000__,
    new_new_n27001__, new_new_n27002__, new_new_n27003__, new_new_n27004__,
    new_new_n27005__, new_new_n27006__, new_new_n27007__, new_new_n27008__,
    new_new_n27009__, new_new_n27010__, new_new_n27011__, new_new_n27012__,
    new_new_n27013__, new_new_n27014__, new_new_n27015__, new_new_n27016__,
    new_new_n27017__, new_new_n27018__, new_new_n27019__, new_new_n27020__,
    new_new_n27021__, new_new_n27022__, new_new_n27023__, new_new_n27024__,
    new_new_n27025__, new_new_n27026__, new_new_n27027__, new_new_n27028__,
    new_new_n27029__, new_new_n27030__, new_new_n27031__, new_new_n27032__,
    new_new_n27033__, new_new_n27034__, new_new_n27035__, new_new_n27036__,
    new_new_n27037__, new_new_n27038__, new_new_n27039__, new_new_n27040__,
    new_new_n27041__, new_new_n27042__, new_new_n27043__, new_new_n27044__,
    new_new_n27045__, new_new_n27046__, new_new_n27047__, new_new_n27048__,
    new_new_n27049__, new_new_n27050__, new_new_n27051__, new_new_n27052__,
    new_new_n27053__, new_new_n27054__, new_new_n27055__, new_new_n27056__,
    new_new_n27057__, new_new_n27058__, new_new_n27059__, new_new_n27060__,
    new_new_n27061__, new_new_n27062__, new_new_n27063__, new_new_n27064__,
    new_new_n27065__, new_new_n27066__, new_new_n27067__, new_new_n27068__,
    new_new_n27069__, new_new_n27070__, new_new_n27071__, new_new_n27072__,
    new_new_n27073__, new_new_n27074__, new_new_n27075__, new_new_n27076__,
    new_new_n27077__, new_new_n27078__, new_new_n27079__, new_new_n27080__,
    new_new_n27081__, new_new_n27082__, new_new_n27083__, new_new_n27084__,
    new_new_n27085__, new_new_n27086__, new_new_n27087__, new_new_n27088__,
    new_new_n27089__, new_new_n27090__, new_new_n27091__, new_new_n27092__,
    new_new_n27093__, new_new_n27094__, new_new_n27095__, new_new_n27096__,
    new_new_n27097__, new_new_n27098__, new_new_n27099__, new_new_n27100__,
    new_new_n27101__, new_new_n27102__, new_new_n27103__, new_new_n27104__,
    new_new_n27105__, new_new_n27106__, new_new_n27107__, new_new_n27108__,
    new_new_n27109__, new_new_n27110__, new_new_n27111__, new_new_n27112__,
    new_new_n27113__, new_new_n27114__, new_new_n27115__, new_new_n27116__,
    new_new_n27117__, new_new_n27118__, new_new_n27119__, new_new_n27120__,
    new_new_n27121__, new_new_n27122__, new_new_n27123__, new_new_n27124__,
    new_new_n27125__, new_new_n27126__, new_new_n27127__, new_new_n27128__,
    new_new_n27129__, new_new_n27130__, new_new_n27131__, new_new_n27132__,
    new_new_n27133__, new_new_n27134__, new_new_n27135__, new_new_n27136__,
    new_new_n27137__, new_new_n27138__, new_new_n27139__, new_new_n27140__,
    new_new_n27141__, new_new_n27142__, new_new_n27143__, new_new_n27144__,
    new_new_n27145__, new_new_n27146__, new_new_n27147__, new_new_n27148__,
    new_new_n27149__, new_new_n27150__, new_new_n27151__, new_new_n27152__,
    new_new_n27153__, new_new_n27154__, new_new_n27155__, new_new_n27156__,
    new_new_n27157__, new_new_n27158__, new_new_n27159__, new_new_n27160__,
    new_new_n27161__, new_new_n27162__, new_new_n27163__, new_new_n27164__,
    new_new_n27165__, new_new_n27166__, new_new_n27167__, new_new_n27168__,
    new_new_n27169__, new_new_n27170__, new_new_n27171__, new_new_n27172__,
    new_new_n27173__, new_new_n27174__, new_new_n27175__, new_new_n27176__,
    new_new_n27177__, new_new_n27178__, new_new_n27179__, new_new_n27180__,
    new_new_n27181__, new_new_n27182__, new_new_n27183__, new_new_n27184__,
    new_new_n27185__, new_new_n27186__, new_new_n27187__, new_new_n27188__,
    new_new_n27189__, new_new_n27190__, new_new_n27191__, new_new_n27192__,
    new_new_n27193__, new_new_n27194__, new_new_n27195__, new_new_n27196__,
    new_new_n27197__, new_new_n27198__, new_new_n27199__, new_new_n27200__,
    new_new_n27201__, new_new_n27202__, new_new_n27203__, new_new_n27204__,
    new_new_n27205__, new_new_n27206__, new_new_n27207__, new_new_n27208__,
    new_new_n27209__, new_new_n27210__, new_new_n27211__, new_new_n27212__,
    new_new_n27213__, new_new_n27214__, new_new_n27215__, new_new_n27216__,
    new_new_n27217__, new_new_n27218__, new_new_n27219__, new_new_n27220__,
    new_new_n27221__, new_new_n27222__, new_new_n27223__, new_new_n27224__,
    new_new_n27225__, new_new_n27226__, new_new_n27227__, new_new_n27228__,
    new_new_n27229__, new_new_n27230__, new_new_n27231__, new_new_n27232__,
    new_new_n27233__, new_new_n27234__, new_new_n27235__, new_new_n27236__,
    new_new_n27237__, new_new_n27238__, new_new_n27239__, new_new_n27240__,
    new_new_n27241__, new_new_n27242__, new_new_n27243__, new_new_n27244__,
    new_new_n27245__, new_new_n27246__, new_new_n27247__, new_new_n27248__,
    new_new_n27249__, new_new_n27250__, new_new_n27251__, new_new_n27252__,
    new_new_n27253__, new_new_n27254__, new_new_n27255__, new_new_n27256__,
    new_new_n27257__, new_new_n27258__, new_new_n27259__, new_new_n27260__,
    new_new_n27261__, new_new_n27262__, new_new_n27263__, new_new_n27264__,
    new_new_n27265__, new_new_n27266__, new_new_n27267__, new_new_n27268__,
    new_new_n27269__, new_new_n27270__, new_new_n27271__, new_new_n27272__,
    new_new_n27273__, new_new_n27274__, new_new_n27275__, new_new_n27276__,
    new_new_n27277__, new_new_n27278__, new_new_n27279__, new_new_n27280__,
    new_new_n27281__, new_new_n27282__, new_new_n27283__, new_new_n27284__,
    new_new_n27285__, new_new_n27286__, new_new_n27287__, new_new_n27288__,
    new_new_n27289__, new_new_n27290__, new_new_n27291__, new_new_n27292__,
    new_new_n27293__, new_new_n27294__, new_new_n27295__, new_new_n27296__,
    new_new_n27297__, new_new_n27298__, new_new_n27299__, new_new_n27300__,
    new_new_n27301__, new_new_n27302__, new_new_n27303__, new_new_n27304__,
    new_new_n27305__, new_new_n27306__, new_new_n27307__, new_new_n27308__,
    new_new_n27309__, new_new_n27310__, new_new_n27311__, new_new_n27312__,
    new_new_n27313__, new_new_n27314__, new_new_n27315__, new_new_n27316__,
    new_new_n27317__, new_new_n27318__, new_new_n27319__, new_new_n27320__,
    new_new_n27321__, new_new_n27322__, new_new_n27323__, new_new_n27324__,
    new_new_n27325__, new_new_n27326__, new_new_n27327__, new_new_n27328__,
    new_new_n27329__, new_new_n27330__, new_new_n27331__, new_new_n27332__,
    new_new_n27333__, new_new_n27334__, new_new_n27335__, new_new_n27336__,
    new_new_n27337__, new_new_n27338__, new_new_n27339__, new_new_n27340__,
    new_new_n27341__, new_new_n27342__, new_new_n27343__, new_new_n27344__,
    new_new_n27345__, new_new_n27346__, new_new_n27347__, new_new_n27348__,
    new_new_n27349__, new_new_n27350__, new_new_n27351__, new_new_n27352__,
    new_new_n27353__, new_new_n27354__, new_new_n27355__, new_new_n27356__,
    new_new_n27357__, new_new_n27358__, new_new_n27359__, new_new_n27360__,
    new_new_n27361__, new_new_n27362__, new_new_n27363__, new_new_n27364__,
    new_new_n27365__, new_new_n27366__, new_new_n27367__, new_new_n27368__,
    new_new_n27369__, new_new_n27370__, new_new_n27371__, new_new_n27372__,
    new_new_n27373__, new_new_n27374__, new_new_n27375__, new_new_n27376__,
    new_new_n27377__, new_new_n27378__, new_new_n27379__, new_new_n27380__,
    new_new_n27381__, new_new_n27382__, new_new_n27383__, new_new_n27384__,
    new_new_n27385__, new_new_n27386__, new_new_n27387__, new_new_n27388__,
    new_new_n27389__, new_new_n27390__, new_new_n27391__, new_new_n27392__,
    new_new_n27393__, new_new_n27394__, new_new_n27395__, new_new_n27396__,
    new_new_n27397__, new_new_n27398__, new_new_n27399__, new_new_n27400__,
    new_new_n27401__, new_new_n27402__, new_new_n27403__, new_new_n27404__,
    new_new_n27405__, new_new_n27406__, new_new_n27407__, new_new_n27408__,
    new_new_n27409__, new_new_n27410__, new_new_n27411__, new_new_n27412__,
    new_new_n27413__, new_new_n27414__, new_new_n27415__, new_new_n27416__,
    new_new_n27417__, new_new_n27418__, new_new_n27419__, new_new_n27420__,
    new_new_n27421__, new_new_n27422__, new_new_n27423__, new_new_n27424__,
    new_new_n27425__, new_new_n27426__, new_new_n27427__, new_new_n27428__,
    new_new_n27429__, new_new_n27430__, new_new_n27431__, new_new_n27432__,
    new_new_n27433__, new_new_n27434__, new_new_n27435__, new_new_n27436__,
    new_new_n27437__, new_new_n27438__, new_new_n27439__, new_new_n27440__,
    new_new_n27441__, new_new_n27442__, new_new_n27443__, new_new_n27444__,
    new_new_n27445__, new_new_n27446__, new_new_n27447__, new_new_n27448__,
    new_new_n27449__, new_new_n27450__, new_new_n27451__, new_new_n27452__,
    new_new_n27453__, new_new_n27454__, new_new_n27455__, new_new_n27456__,
    new_new_n27457__, new_new_n27458__, new_new_n27459__, new_new_n27460__,
    new_new_n27461__, new_new_n27462__, new_new_n27463__, new_new_n27464__,
    new_new_n27465__, new_new_n27466__, new_new_n27467__, new_new_n27468__,
    new_new_n27469__, new_new_n27470__, new_new_n27471__, new_new_n27472__,
    new_new_n27473__, new_new_n27474__, new_new_n27475__, new_new_n27476__,
    new_new_n27477__, new_new_n27478__, new_new_n27479__, new_new_n27480__,
    new_new_n27481__, new_new_n27482__, new_new_n27483__, new_new_n27484__,
    new_new_n27485__, new_new_n27486__, new_new_n27487__, new_new_n27488__,
    new_new_n27489__, new_new_n27490__, new_new_n27491__, new_new_n27492__,
    new_new_n27493__, new_new_n27494__, new_new_n27495__, new_new_n27496__,
    new_new_n27497__, new_new_n27498__, new_new_n27499__, new_new_n27500__,
    new_new_n27501__, new_new_n27502__, new_new_n27503__, new_new_n27504__,
    new_new_n27505__, new_new_n27506__, new_new_n27507__, new_new_n27508__,
    new_new_n27509__, new_new_n27510__, new_new_n27511__, new_new_n27512__,
    new_new_n27513__, new_new_n27514__, new_new_n27515__, new_new_n27516__,
    new_new_n27517__, new_new_n27518__, new_new_n27519__, new_new_n27520__,
    new_new_n27521__, new_new_n27522__, new_new_n27523__, new_new_n27524__,
    new_new_n27525__, new_new_n27526__, new_new_n27527__, new_new_n27528__,
    new_new_n27529__, new_new_n27530__, new_new_n27531__, new_new_n27532__,
    new_new_n27533__, new_new_n27534__, new_new_n27535__, new_new_n27536__,
    new_new_n27537__, new_new_n27538__, new_new_n27539__, new_new_n27540__,
    new_new_n27541__, new_new_n27542__, new_new_n27543__, new_new_n27544__,
    new_new_n27545__, new_new_n27546__, new_new_n27547__, new_new_n27548__,
    new_new_n27549__, new_new_n27550__, new_new_n27551__, new_new_n27552__,
    new_new_n27553__, new_new_n27554__, new_new_n27555__, new_new_n27556__,
    new_new_n27557__, new_new_n27558__, new_new_n27559__, new_new_n27560__,
    new_new_n27561__, new_new_n27562__, new_new_n27563__, new_new_n27564__,
    new_new_n27565__, new_new_n27566__, new_new_n27567__, new_new_n27568__,
    new_new_n27569__, new_new_n27570__, new_new_n27571__, new_new_n27572__,
    new_new_n27573__, new_new_n27574__, new_new_n27575__, new_new_n27576__,
    new_new_n27577__, new_new_n27578__, new_new_n27579__, new_new_n27580__,
    new_new_n27581__, new_new_n27582__, new_new_n27583__, new_new_n27584__,
    new_new_n27585__, new_new_n27586__, new_new_n27587__, new_new_n27588__,
    new_new_n27589__, new_new_n27590__, new_new_n27591__, new_new_n27592__,
    new_new_n27593__, new_new_n27594__, new_new_n27595__, new_new_n27596__,
    new_new_n27597__, new_new_n27598__, new_new_n27599__, new_new_n27600__,
    new_new_n27601__, new_new_n27602__, new_new_n27603__, new_new_n27604__,
    new_new_n27605__, new_new_n27606__, new_new_n27607__, new_new_n27608__,
    new_new_n27609__, new_new_n27610__, new_new_n27611__, new_new_n27612__,
    new_new_n27613__, new_new_n27614__, new_new_n27615__, new_new_n27616__,
    new_new_n27617__, new_new_n27618__, new_new_n27619__, new_new_n27620__,
    new_new_n27621__, new_new_n27622__, new_new_n27623__, new_new_n27624__,
    new_new_n27625__, new_new_n27626__, new_new_n27627__, new_new_n27628__,
    new_new_n27629__, new_new_n27630__, new_new_n27631__, new_new_n27632__,
    new_new_n27633__, new_new_n27634__, new_new_n27635__, new_new_n27636__,
    new_new_n27637__, new_new_n27638__, new_new_n27639__, new_new_n27640__,
    new_new_n27641__, new_new_n27642__, new_new_n27643__, new_new_n27644__,
    new_new_n27645__, new_new_n27646__, new_new_n27647__, new_new_n27648__,
    new_new_n27649__, new_new_n27650__, new_new_n27651__, new_new_n27652__,
    new_new_n27653__, new_new_n27654__, new_new_n27655__, new_new_n27656__,
    new_new_n27657__, new_new_n27658__, new_new_n27659__, new_new_n27660__,
    new_new_n27661__, new_new_n27662__, new_new_n27663__, new_new_n27664__,
    new_new_n27665__, new_new_n27666__, new_new_n27667__, new_new_n27668__,
    new_new_n27669__, new_new_n27670__, new_new_n27671__, new_new_n27672__,
    new_new_n27673__, new_new_n27674__, new_new_n27675__, new_new_n27676__,
    new_new_n27677__, new_new_n27678__, new_new_n27679__, new_new_n27680__,
    new_new_n27681__, new_new_n27682__, new_new_n27683__, new_new_n27684__,
    new_new_n27685__, new_new_n27686__, new_new_n27687__, new_new_n27688__,
    new_new_n27689__, new_new_n27690__, new_new_n27691__, new_new_n27692__,
    new_new_n27693__, new_new_n27694__, new_new_n27695__, new_new_n27696__,
    new_new_n27697__, new_new_n27698__, new_new_n27699__, new_new_n27700__,
    new_new_n27701__, new_new_n27702__, new_new_n27703__, new_new_n27704__,
    new_new_n27705__, new_new_n27706__, new_new_n27707__, new_new_n27708__,
    new_new_n27709__, new_new_n27710__, new_new_n27711__, new_new_n27712__,
    new_new_n27713__, new_new_n27714__, new_new_n27715__, new_new_n27716__,
    new_new_n27717__, new_new_n27718__, new_new_n27719__, new_new_n27720__,
    new_new_n27721__, new_new_n27722__, new_new_n27723__, new_new_n27724__,
    new_new_n27725__, new_new_n27726__, new_new_n27727__, new_new_n27728__,
    new_new_n27729__, new_new_n27730__, new_new_n27731__, new_new_n27732__,
    new_new_n27733__, new_new_n27734__, new_new_n27735__, new_new_n27736__,
    new_new_n27737__, new_new_n27738__, new_new_n27739__, new_new_n27740__,
    new_new_n27741__, new_new_n27742__, new_new_n27743__, new_new_n27744__,
    new_new_n27745__, new_new_n27746__, new_new_n27747__, new_new_n27748__,
    new_new_n27749__, new_new_n27750__, new_new_n27751__, new_new_n27752__,
    new_new_n27753__, new_new_n27754__, new_new_n27755__, new_new_n27756__,
    new_new_n27757__, new_new_n27758__, new_new_n27759__, new_new_n27760__,
    new_new_n27761__, new_new_n27762__, new_new_n27763__, new_new_n27764__,
    new_new_n27765__, new_new_n27766__, new_new_n27767__, new_new_n27768__,
    new_new_n27769__, new_new_n27770__, new_new_n27771__, new_new_n27772__,
    new_new_n27773__, new_new_n27774__, new_new_n27775__, new_new_n27776__,
    new_new_n27777__, new_new_n27778__, new_new_n27779__, new_new_n27780__,
    new_new_n27781__, new_new_n27782__, new_new_n27783__, new_new_n27784__,
    new_new_n27785__, new_new_n27786__, new_new_n27787__, new_new_n27788__,
    new_new_n27789__, new_new_n27790__, new_new_n27791__, new_new_n27792__,
    new_new_n27793__, new_new_n27794__, new_new_n27795__, new_new_n27796__,
    new_new_n27797__, new_new_n27798__, new_new_n27799__, new_new_n27800__,
    new_new_n27801__, new_new_n27802__, new_new_n27803__, new_new_n27804__,
    new_new_n27805__, new_new_n27806__, new_new_n27807__, new_new_n27808__,
    new_new_n27809__, new_new_n27810__, new_new_n27811__, new_new_n27812__,
    new_new_n27813__, new_new_n27814__, new_new_n27815__, new_new_n27816__,
    new_new_n27817__, new_new_n27818__, new_new_n27819__, new_new_n27820__,
    new_new_n27821__, new_new_n27822__, new_new_n27823__, new_new_n27824__,
    new_new_n27825__, new_new_n27826__, new_new_n27827__, new_new_n27828__,
    new_new_n27829__, new_new_n27830__, new_new_n27831__, new_new_n27832__,
    new_new_n27833__, new_new_n27834__, new_new_n27835__, new_new_n27836__,
    new_new_n27837__, new_new_n27838__, new_new_n27839__, new_new_n27840__,
    new_new_n27841__, new_new_n27842__, new_new_n27843__, new_new_n27844__,
    new_new_n27845__, new_new_n27846__, new_new_n27847__, new_new_n27848__,
    new_new_n27849__, new_new_n27850__, new_new_n27851__, new_new_n27852__,
    new_new_n27853__, new_new_n27854__, new_new_n27855__, new_new_n27856__,
    new_new_n27857__, new_new_n27858__, new_new_n27859__, new_new_n27860__,
    new_new_n27861__, new_new_n27862__, new_new_n27863__, new_new_n27864__,
    new_new_n27865__, new_new_n27866__, new_new_n27867__, new_new_n27868__,
    new_new_n27869__, new_new_n27870__, new_new_n27871__, new_new_n27872__,
    new_new_n27873__, new_new_n27874__, new_new_n27875__, new_new_n27876__,
    new_new_n27877__, new_new_n27878__, new_new_n27879__, new_new_n27880__,
    new_new_n27881__, new_new_n27882__, new_new_n27883__, new_new_n27884__,
    new_new_n27885__, new_new_n27886__, new_new_n27887__, new_new_n27888__,
    new_new_n27889__, new_new_n27890__, new_new_n27891__, new_new_n27892__,
    new_new_n27893__, new_new_n27894__, new_new_n27895__, new_new_n27896__,
    new_new_n27897__, new_new_n27898__, new_new_n27899__, new_new_n27900__,
    new_new_n27901__, new_new_n27902__, new_new_n27903__, new_new_n27904__,
    new_new_n27905__, new_new_n27906__, new_new_n27907__, new_new_n27908__,
    new_new_n27909__, new_new_n27910__, new_new_n27911__, new_new_n27912__,
    new_new_n27913__, new_new_n27914__, new_new_n27915__, new_new_n27916__,
    new_new_n27917__, new_new_n27918__, new_new_n27919__, new_new_n27920__,
    new_new_n27921__, new_new_n27922__, new_new_n27923__, new_new_n27924__,
    new_new_n27925__, new_new_n27926__, new_new_n27927__, new_new_n27928__,
    new_new_n27929__, new_new_n27930__, new_new_n27931__, new_new_n27932__,
    new_new_n27933__, new_new_n27934__, new_new_n27935__, new_new_n27936__,
    new_new_n27937__, new_new_n27938__, new_new_n27939__, new_new_n27940__,
    new_new_n27941__, new_new_n27942__, new_new_n27943__, new_new_n27944__,
    new_new_n27945__, new_new_n27946__, new_new_n27947__, new_new_n27948__,
    new_new_n27949__, new_new_n27950__, new_new_n27951__, new_new_n27952__,
    new_new_n27953__, new_new_n27954__, new_new_n27955__, new_new_n27956__,
    new_new_n27957__, new_new_n27958__, new_new_n27959__, new_new_n27960__,
    new_new_n27961__, new_new_n27962__, new_new_n27963__, new_new_n27964__,
    new_new_n27965__, new_new_n27966__, new_new_n27967__, new_new_n27968__,
    new_new_n27969__, new_new_n27970__, new_new_n27971__, new_new_n27972__,
    new_new_n27973__, new_new_n27974__, new_new_n27975__, new_new_n27976__,
    new_new_n27977__, new_new_n27978__, new_new_n27979__, new_new_n27980__,
    new_new_n27981__, new_new_n27982__, new_new_n27983__, new_new_n27984__,
    new_new_n27985__, new_new_n27986__, new_new_n27987__, new_new_n27988__,
    new_new_n27989__, new_new_n27990__, new_new_n27991__, new_new_n27992__,
    new_new_n27993__, new_new_n27994__, new_new_n27995__, new_new_n27996__,
    new_new_n27997__, new_new_n27998__, new_new_n27999__, new_new_n28000__,
    new_new_n28001__, new_new_n28002__, new_new_n28003__, new_new_n28004__,
    new_new_n28005__, new_new_n28006__, new_new_n28007__, new_new_n28008__,
    new_new_n28009__, new_new_n28010__, new_new_n28011__, new_new_n28012__,
    new_new_n28013__, new_new_n28014__, new_new_n28015__, new_new_n28016__,
    new_new_n28017__, new_new_n28018__, new_new_n28019__, new_new_n28020__,
    new_new_n28021__, new_new_n28022__, new_new_n28023__, new_new_n28024__,
    new_new_n28025__, new_new_n28026__, new_new_n28027__, new_new_n28028__,
    new_new_n28029__, new_new_n28030__, new_new_n28031__, new_new_n28032__,
    new_new_n28033__, new_new_n28034__, new_new_n28035__, new_new_n28036__,
    new_new_n28037__, new_new_n28038__, new_new_n28039__, new_new_n28040__,
    new_new_n28041__, new_new_n28042__, new_new_n28043__, new_new_n28044__,
    new_new_n28045__, new_new_n28046__, new_new_n28047__, new_new_n28048__,
    new_new_n28049__, new_new_n28050__, new_new_n28051__, new_new_n28052__,
    new_new_n28053__, new_new_n28054__, new_new_n28055__, new_new_n28056__,
    new_new_n28057__, new_new_n28058__, new_new_n28059__, new_new_n28060__,
    new_new_n28061__, new_new_n28062__, new_new_n28063__, new_new_n28064__,
    new_new_n28065__, new_new_n28066__, new_new_n28067__, new_new_n28068__,
    new_new_n28069__, new_new_n28070__, new_new_n28071__, new_new_n28072__,
    new_new_n28073__, new_new_n28074__, new_new_n28075__, new_new_n28076__,
    new_new_n28077__, new_new_n28078__, new_new_n28079__, new_new_n28080__,
    new_new_n28081__, new_new_n28082__, new_new_n28083__, new_new_n28084__,
    new_new_n28085__, new_new_n28086__, new_new_n28087__, new_new_n28088__,
    new_new_n28089__, new_new_n28090__, new_new_n28091__, new_new_n28092__,
    new_new_n28093__, new_new_n28094__, new_new_n28095__, new_new_n28096__,
    new_new_n28097__, new_new_n28098__, new_new_n28099__, new_new_n28100__,
    new_new_n28101__, new_new_n28102__, new_new_n28103__, new_new_n28104__,
    new_new_n28105__, new_new_n28106__, new_new_n28107__, new_new_n28108__,
    new_new_n28109__, new_new_n28110__, new_new_n28111__, new_new_n28112__,
    new_new_n28113__, new_new_n28114__, new_new_n28115__, new_new_n28116__,
    new_new_n28117__, new_new_n28118__, new_new_n28119__, new_new_n28120__,
    new_new_n28121__, new_new_n28122__, new_new_n28123__, new_new_n28124__,
    new_new_n28125__, new_new_n28126__, new_new_n28127__, new_new_n28128__,
    new_new_n28129__, new_new_n28130__, new_new_n28131__, new_new_n28132__,
    new_new_n28133__, new_new_n28134__, new_new_n28135__, new_new_n28136__,
    new_new_n28137__, new_new_n28138__, new_new_n28139__, new_new_n28140__,
    new_new_n28141__, new_new_n28142__, new_new_n28143__, new_new_n28144__,
    new_new_n28145__, new_new_n28146__, new_new_n28147__, new_new_n28148__,
    new_new_n28149__, new_new_n28150__, new_new_n28151__, new_new_n28152__,
    new_new_n28153__, new_new_n28154__, new_new_n28155__, new_new_n28156__,
    new_new_n28157__, new_new_n28158__, new_new_n28159__, new_new_n28160__,
    new_new_n28161__, new_new_n28162__, new_new_n28163__, new_new_n28164__,
    new_new_n28165__, new_new_n28166__, new_new_n28167__, new_new_n28168__,
    new_new_n28169__, new_new_n28170__, new_new_n28171__, new_new_n28172__,
    new_new_n28173__, new_new_n28174__, new_new_n28175__, new_new_n28176__,
    new_new_n28177__, new_new_n28178__, new_new_n28179__, new_new_n28180__,
    new_new_n28181__, new_new_n28182__, new_new_n28183__, new_new_n28184__,
    new_new_n28185__, new_new_n28186__, new_new_n28187__, new_new_n28188__,
    new_new_n28189__, new_new_n28190__, new_new_n28191__, new_new_n28192__,
    new_new_n28193__, new_new_n28194__, new_new_n28195__, new_new_n28196__,
    new_new_n28197__, new_new_n28198__, new_new_n28199__, new_new_n28200__,
    new_new_n28201__, new_new_n28202__, new_new_n28203__, new_new_n28204__,
    new_new_n28205__, new_new_n28206__, new_new_n28207__, new_new_n28208__,
    new_new_n28209__, new_new_n28210__, new_new_n28211__, new_new_n28212__,
    new_new_n28213__, new_new_n28214__, new_new_n28215__, new_new_n28216__,
    new_new_n28217__, new_new_n28218__, new_new_n28219__, new_new_n28220__,
    new_new_n28221__, new_new_n28222__, new_new_n28223__, new_new_n28224__,
    new_new_n28225__, new_new_n28226__, new_new_n28227__, new_new_n28228__,
    new_new_n28229__, new_new_n28230__, new_new_n28231__, new_new_n28232__,
    new_new_n28233__, new_new_n28234__, new_new_n28235__, new_new_n28236__,
    new_new_n28237__, new_new_n28238__, new_new_n28239__, new_new_n28240__,
    new_new_n28241__, new_new_n28242__, new_new_n28243__, new_new_n28244__,
    new_new_n28245__, new_new_n28246__, new_new_n28247__, new_new_n28248__,
    new_new_n28249__, new_new_n28250__, new_new_n28251__, new_new_n28252__,
    new_new_n28253__, new_new_n28254__, new_new_n28255__, new_new_n28256__,
    new_new_n28257__, new_new_n28258__, new_new_n28259__, new_new_n28260__,
    new_new_n28261__, new_new_n28262__, new_new_n28263__, new_new_n28264__,
    new_new_n28265__, new_new_n28266__, new_new_n28267__, new_new_n28268__,
    new_new_n28269__, new_new_n28270__, new_new_n28271__, new_new_n28272__,
    new_new_n28273__, new_new_n28274__, new_new_n28275__, new_new_n28276__,
    new_new_n28277__, new_new_n28278__, new_new_n28279__, new_new_n28280__,
    new_new_n28281__, new_new_n28282__, new_new_n28283__, new_new_n28284__,
    new_new_n28285__, new_new_n28286__, new_new_n28287__, new_new_n28288__,
    new_new_n28289__, new_new_n28290__, new_new_n28291__, new_new_n28292__,
    new_new_n28293__, new_new_n28294__, new_new_n28295__, new_new_n28296__,
    new_new_n28297__, new_new_n28298__, new_new_n28299__, new_new_n28300__,
    new_new_n28301__, new_new_n28302__, new_new_n28303__, new_new_n28304__,
    new_new_n28305__, new_new_n28306__, new_new_n28307__, new_new_n28308__,
    new_new_n28309__, new_new_n28310__, new_new_n28311__, new_new_n28312__,
    new_new_n28313__, new_new_n28314__, new_new_n28315__, new_new_n28316__,
    new_new_n28317__, new_new_n28318__, new_new_n28319__, new_new_n28320__,
    new_new_n28321__, new_new_n28322__, new_new_n28323__, new_new_n28324__,
    new_new_n28325__, new_new_n28326__, new_new_n28327__, new_new_n28328__,
    new_new_n28329__, new_new_n28330__, new_new_n28331__, new_new_n28332__,
    new_new_n28333__, new_new_n28334__, new_new_n28335__, new_new_n28336__,
    new_new_n28337__, new_new_n28338__, new_new_n28339__, new_new_n28340__,
    new_new_n28341__, new_new_n28342__, new_new_n28343__, new_new_n28344__,
    new_new_n28345__, new_new_n28346__, new_new_n28347__, new_new_n28348__,
    new_new_n28349__, new_new_n28350__, new_new_n28351__, new_new_n28352__,
    new_new_n28353__, new_new_n28354__, new_new_n28355__, new_new_n28356__,
    new_new_n28357__, new_new_n28358__, new_new_n28359__, new_new_n28360__,
    new_new_n28361__, new_new_n28362__, new_new_n28363__, new_new_n28364__,
    new_new_n28365__, new_new_n28366__, new_new_n28367__, new_new_n28368__,
    new_new_n28369__, new_new_n28370__, new_new_n28371__, new_new_n28372__,
    new_new_n28373__, new_new_n28374__, new_new_n28375__, new_new_n28376__,
    new_new_n28377__, new_new_n28378__, new_new_n28379__, new_new_n28380__,
    new_new_n28381__, new_new_n28382__, new_new_n28383__, new_new_n28384__,
    new_new_n28385__, new_new_n28386__, new_new_n28387__, new_new_n28388__,
    new_new_n28389__, new_new_n28390__, new_new_n28391__, new_new_n28392__,
    new_new_n28393__, new_new_n28394__, new_new_n28395__, new_new_n28396__,
    new_new_n28397__, new_new_n28398__, new_new_n28399__, new_new_n28400__,
    new_new_n28401__, new_new_n28402__, new_new_n28403__, new_new_n28404__,
    new_new_n28405__, new_new_n28406__, new_new_n28407__, new_new_n28408__,
    new_new_n28409__, new_new_n28410__, new_new_n28411__, new_new_n28412__,
    new_new_n28413__, new_new_n28414__, new_new_n28415__, new_new_n28416__,
    new_new_n28417__, new_new_n28418__, new_new_n28419__, new_new_n28420__,
    new_new_n28421__, new_new_n28422__, new_new_n28423__, new_new_n28424__,
    new_new_n28425__, new_new_n28426__, new_new_n28427__, new_new_n28428__,
    new_new_n28429__, new_new_n28430__, new_new_n28431__, new_new_n28432__,
    new_new_n28433__, new_new_n28434__, new_new_n28435__, new_new_n28436__,
    new_new_n28437__, new_new_n28438__, new_new_n28439__, new_new_n28440__,
    new_new_n28441__, new_new_n28442__, new_new_n28443__, new_new_n28444__,
    new_new_n28445__, new_new_n28446__, new_new_n28447__, new_new_n28448__,
    new_new_n28449__, new_new_n28450__, new_new_n28451__, new_new_n28452__,
    new_new_n28453__, new_new_n28454__, new_new_n28455__, new_new_n28456__,
    new_new_n28457__, new_new_n28458__, new_new_n28459__, new_new_n28460__,
    new_new_n28461__, new_new_n28462__, new_new_n28463__, new_new_n28464__,
    new_new_n28465__, new_new_n28466__, new_new_n28467__, new_new_n28468__,
    new_new_n28469__, new_new_n28470__, new_new_n28471__, new_new_n28472__,
    new_new_n28473__, new_new_n28474__, new_new_n28475__, new_new_n28476__,
    new_new_n28477__, new_new_n28478__, new_new_n28479__, new_new_n28480__,
    new_new_n28481__, new_new_n28482__, new_new_n28483__, new_new_n28484__,
    new_new_n28485__, new_new_n28486__, new_new_n28487__, new_new_n28488__,
    new_new_n28489__, new_new_n28490__, new_new_n28491__, new_new_n28492__,
    new_new_n28493__, new_new_n28494__, new_new_n28495__, new_new_n28496__,
    new_new_n28497__, new_new_n28498__, new_new_n28499__, new_new_n28500__,
    new_new_n28501__, new_new_n28502__, new_new_n28503__, new_new_n28504__,
    new_new_n28505__, new_new_n28506__, new_new_n28507__, new_new_n28508__,
    new_new_n28509__, new_new_n28510__, new_new_n28511__, new_new_n28512__,
    new_new_n28513__, new_new_n28514__, new_new_n28515__, new_new_n28516__,
    new_new_n28517__, new_new_n28518__, new_new_n28519__, new_new_n28520__,
    new_new_n28521__, new_new_n28522__, new_new_n28523__, new_new_n28524__,
    new_new_n28525__, new_new_n28526__, new_new_n28527__, new_new_n28528__,
    new_new_n28529__, new_new_n28530__, new_new_n28531__, new_new_n28532__,
    new_new_n28533__, new_new_n28534__, new_new_n28535__, new_new_n28536__,
    new_new_n28537__, new_new_n28538__, new_new_n28539__, new_new_n28540__,
    new_new_n28541__, new_new_n28542__, new_new_n28543__, new_new_n28544__,
    new_new_n28545__, new_new_n28546__, new_new_n28547__, new_new_n28548__,
    new_new_n28549__, new_new_n28550__, new_new_n28551__, new_new_n28552__,
    new_new_n28553__, new_new_n28554__, new_new_n28555__, new_new_n28556__,
    new_new_n28557__, new_new_n28558__, new_new_n28559__, new_new_n28560__,
    new_new_n28561__, new_new_n28562__, new_new_n28563__, new_new_n28564__,
    new_new_n28565__, new_new_n28566__, new_new_n28567__, new_new_n28568__,
    new_new_n28569__, new_new_n28570__, new_new_n28571__, new_new_n28572__,
    new_new_n28573__, new_new_n28574__, new_new_n28575__, new_new_n28576__,
    new_new_n28577__, new_new_n28578__, new_new_n28579__, new_new_n28580__,
    new_new_n28581__, new_new_n28582__, new_new_n28583__, new_new_n28584__,
    new_new_n28585__, new_new_n28586__, new_new_n28587__, new_new_n28588__,
    new_new_n28589__, new_new_n28590__, new_new_n28591__, new_new_n28592__,
    new_new_n28593__, new_new_n28594__, new_new_n28595__, new_new_n28596__,
    new_new_n28597__, new_new_n28598__, new_new_n28599__, new_new_n28600__,
    new_new_n28601__, new_new_n28602__, new_new_n28603__, new_new_n28604__,
    new_new_n28605__, new_new_n28606__, new_new_n28607__, new_new_n28608__,
    new_new_n28609__, new_new_n28610__, new_new_n28611__, new_new_n28612__,
    new_new_n28613__, new_new_n28614__, new_new_n28615__, new_new_n28616__,
    new_new_n28617__, new_new_n28618__, new_new_n28619__, new_new_n28620__,
    new_new_n28621__, new_new_n28622__, new_new_n28623__, new_new_n28624__,
    new_new_n28625__, new_new_n28626__, new_new_n28627__, new_new_n28628__,
    new_new_n28629__, new_new_n28630__, new_new_n28631__, new_new_n28632__,
    new_new_n28633__, new_new_n28634__, new_new_n28635__, new_new_n28636__,
    new_new_n28637__, new_new_n28638__, new_new_n28639__, new_new_n28640__,
    new_new_n28641__, new_new_n28642__, new_new_n28643__, new_new_n28644__,
    new_new_n28645__, new_new_n28646__, new_new_n28647__, new_new_n28648__,
    new_new_n28649__, new_new_n28650__, new_new_n28651__, new_new_n28652__,
    new_new_n28653__, new_new_n28654__, new_new_n28655__, new_new_n28656__,
    new_new_n28657__, new_new_n28658__, new_new_n28659__, new_new_n28660__,
    new_new_n28661__, new_new_n28662__, new_new_n28663__, new_new_n28664__,
    new_new_n28665__, new_new_n28666__, new_new_n28667__, new_new_n28668__,
    new_new_n28669__, new_new_n28670__, new_new_n28671__, new_new_n28672__,
    new_new_n28673__, new_new_n28674__, new_new_n28675__, new_new_n28676__,
    new_new_n28677__, new_new_n28678__, new_new_n28679__, new_new_n28680__,
    new_new_n28681__, new_new_n28682__, new_new_n28683__, new_new_n28684__,
    new_new_n28685__, new_new_n28686__, new_new_n28687__, new_new_n28688__,
    new_new_n28689__, new_new_n28690__, new_new_n28691__, new_new_n28692__,
    new_new_n28693__, new_new_n28694__, new_new_n28695__, new_new_n28696__,
    new_new_n28697__, new_new_n28698__, new_new_n28699__, new_new_n28700__,
    new_new_n28701__, new_new_n28702__, new_new_n28703__, new_new_n28704__,
    new_new_n28705__, new_new_n28706__, new_new_n28707__, new_new_n28708__,
    new_new_n28709__, new_new_n28710__, new_new_n28711__, new_new_n28712__,
    new_new_n28713__, new_new_n28714__, new_new_n28715__, new_new_n28716__,
    new_new_n28717__, new_new_n28718__, new_new_n28719__, new_new_n28720__,
    new_new_n28721__, new_new_n28722__, new_new_n28723__, new_new_n28724__,
    new_new_n28725__, new_new_n28726__, new_new_n28727__, new_new_n28728__,
    new_new_n28729__, new_new_n28730__, new_new_n28731__, new_new_n28732__,
    new_new_n28733__, new_new_n28734__, new_new_n28735__, new_new_n28736__,
    new_new_n28737__, new_new_n28738__, new_new_n28739__, new_new_n28740__,
    new_new_n28741__, new_new_n28742__, new_new_n28743__, new_new_n28744__,
    new_new_n28745__, new_new_n28746__, new_new_n28747__, new_new_n28748__,
    new_new_n28749__, new_new_n28750__, new_new_n28751__, new_new_n28752__,
    new_new_n28753__, new_new_n28754__, new_new_n28755__, new_new_n28756__,
    new_new_n28757__, new_new_n28758__, new_new_n28759__, new_new_n28760__,
    new_new_n28761__, new_new_n28762__, new_new_n28763__, new_new_n28764__,
    new_new_n28765__, new_new_n28766__, new_new_n28767__, new_new_n28768__,
    new_new_n28769__, new_new_n28770__, new_new_n28771__, new_new_n28772__,
    new_new_n28773__, new_new_n28774__, new_new_n28775__, new_new_n28776__,
    new_new_n28777__, new_new_n28778__, new_new_n28779__, new_new_n28780__,
    new_new_n28781__, new_new_n28782__, new_new_n28783__, new_new_n28784__,
    new_new_n28785__, new_new_n28786__, new_new_n28787__, new_new_n28788__,
    new_new_n28789__, new_new_n28790__, new_new_n28791__, new_new_n28792__,
    new_new_n28793__, new_new_n28794__, new_new_n28795__, new_new_n28796__,
    new_new_n28797__, new_new_n28798__, new_new_n28799__, new_new_n28800__,
    new_new_n28801__, new_new_n28802__, new_new_n28803__, new_new_n28804__,
    new_new_n28805__, new_new_n28806__, new_new_n28807__, new_new_n28808__,
    new_new_n28809__, new_new_n28810__, new_new_n28811__, new_new_n28812__,
    new_new_n28813__, new_new_n28814__, new_new_n28815__, new_new_n28816__,
    new_new_n28817__, new_new_n28818__, new_new_n28819__, new_new_n28820__,
    new_new_n28821__, new_new_n28822__, new_new_n28823__, new_new_n28824__,
    new_new_n28825__, new_new_n28826__, new_new_n28827__, new_new_n28828__,
    new_new_n28829__, new_new_n28830__, new_new_n28831__, new_new_n28832__,
    new_new_n28833__, new_new_n28834__, new_new_n28835__, new_new_n28836__,
    new_new_n28837__, new_new_n28838__, new_new_n28839__, new_new_n28840__,
    new_new_n28841__, new_new_n28842__, new_new_n28843__, new_new_n28844__,
    new_new_n28845__, new_new_n28846__, new_new_n28847__, new_new_n28848__,
    new_new_n28849__, new_new_n28850__, new_new_n28851__, new_new_n28852__,
    new_new_n28853__, new_new_n28854__, new_new_n28855__, new_new_n28856__,
    new_new_n28857__, new_new_n28858__, new_new_n28859__, new_new_n28860__,
    new_new_n28861__, new_new_n28862__, new_new_n28863__, new_new_n28864__,
    new_new_n28865__, new_new_n28866__, new_new_n28867__, new_new_n28868__,
    new_new_n28869__, new_new_n28870__, new_new_n28871__, new_new_n28872__,
    new_new_n28873__, new_new_n28874__, new_new_n28875__, new_new_n28876__,
    new_new_n28877__, new_new_n28878__, new_new_n28879__, new_new_n28880__,
    new_new_n28881__, new_new_n28882__, new_new_n28883__, new_new_n28884__,
    new_new_n28885__, new_new_n28886__, new_new_n28887__, new_new_n28888__,
    new_new_n28889__, new_new_n28890__, new_new_n28891__, new_new_n28892__,
    new_new_n28893__, new_new_n28894__, new_new_n28895__, new_new_n28896__,
    new_new_n28897__, new_new_n28898__, new_new_n28899__, new_new_n28900__,
    new_new_n28901__, new_new_n28902__, new_new_n28903__, new_new_n28904__,
    new_new_n28905__, new_new_n28906__, new_new_n28907__, new_new_n28908__,
    new_new_n28909__, new_new_n28910__, new_new_n28911__, new_new_n28912__,
    new_new_n28913__, new_new_n28914__, new_new_n28915__, new_new_n28916__,
    new_new_n28917__, new_new_n28918__, new_new_n28919__, new_new_n28920__,
    new_new_n28921__, new_new_n28922__, new_new_n28923__, new_new_n28924__,
    new_new_n28925__, new_new_n28926__, new_new_n28927__, new_new_n28928__,
    new_new_n28929__, new_new_n28930__, new_new_n28931__, new_new_n28932__,
    new_new_n28933__, new_new_n28934__, new_new_n28935__, new_new_n28936__,
    new_new_n28937__, new_new_n28938__, new_new_n28939__, new_new_n28940__,
    new_new_n28941__, new_new_n28942__, new_new_n28943__, new_new_n28944__,
    new_new_n28945__, new_new_n28946__, new_new_n28947__, new_new_n28948__,
    new_new_n28949__, new_new_n28950__, new_new_n28951__, new_new_n28952__,
    new_new_n28953__, new_new_n28954__, new_new_n28955__, new_new_n28956__,
    new_new_n28957__, new_new_n28958__, new_new_n28959__, new_new_n28960__,
    new_new_n28961__, new_new_n28962__, new_new_n28963__, new_new_n28964__,
    new_new_n28965__, new_new_n28966__, new_new_n28967__, new_new_n28968__,
    new_new_n28969__, new_new_n28970__, new_new_n28971__, new_new_n28972__,
    new_new_n28973__, new_new_n28974__, new_new_n28975__, new_new_n28976__,
    new_new_n28977__, new_new_n28978__, new_new_n28979__, new_new_n28980__,
    new_new_n28981__, new_new_n28982__, new_new_n28983__, new_new_n28984__,
    new_new_n28985__, new_new_n28986__, new_new_n28987__, new_new_n28988__,
    new_new_n28989__, new_new_n28990__, new_new_n28991__, new_new_n28992__,
    new_new_n28993__, new_new_n28994__, new_new_n28995__, new_new_n28996__,
    new_new_n28997__, new_new_n28998__, new_new_n28999__, new_new_n29000__,
    new_new_n29001__, new_new_n29002__, new_new_n29003__, new_new_n29004__,
    new_new_n29005__, new_new_n29006__, new_new_n29007__, new_new_n29008__,
    new_new_n29009__, new_new_n29010__, new_new_n29011__, new_new_n29012__,
    new_new_n29013__, new_new_n29014__, new_new_n29015__, new_new_n29016__,
    new_new_n29017__, new_new_n29018__, new_new_n29019__, new_new_n29020__,
    new_new_n29021__, new_new_n29022__, new_new_n29023__, new_new_n29024__,
    new_new_n29025__, new_new_n29026__, new_new_n29027__, new_new_n29028__,
    new_new_n29029__, new_new_n29030__, new_new_n29031__, new_new_n29032__,
    new_new_n29033__, new_new_n29034__, new_new_n29035__, new_new_n29036__,
    new_new_n29037__, new_new_n29038__, new_new_n29039__, new_new_n29040__,
    new_new_n29041__, new_new_n29042__, new_new_n29043__, new_new_n29044__,
    new_new_n29045__, new_new_n29046__, new_new_n29047__, new_new_n29048__,
    new_new_n29049__, new_new_n29050__, new_new_n29051__, new_new_n29052__,
    new_new_n29053__, new_new_n29054__, new_new_n29055__, new_new_n29056__,
    new_new_n29057__, new_new_n29058__, new_new_n29059__, new_new_n29060__,
    new_new_n29061__, new_new_n29062__, new_new_n29063__, new_new_n29064__,
    new_new_n29065__, new_new_n29066__, new_new_n29067__, new_new_n29068__,
    new_new_n29069__, new_new_n29070__, new_new_n29071__, new_new_n29072__,
    new_new_n29073__, new_new_n29074__, new_new_n29075__, new_new_n29076__,
    new_new_n29077__, new_new_n29078__, new_new_n29079__, new_new_n29080__,
    new_new_n29081__, new_new_n29082__, new_new_n29083__, new_new_n29084__,
    new_new_n29085__, new_new_n29086__, new_new_n29087__, new_new_n29088__,
    new_new_n29089__, new_new_n29090__, new_new_n29091__, new_new_n29092__,
    new_new_n29093__, new_new_n29094__, new_new_n29095__, new_new_n29096__,
    new_new_n29097__, new_new_n29098__, new_new_n29099__, new_new_n29100__,
    new_new_n29101__, new_new_n29102__, new_new_n29103__, new_new_n29104__,
    new_new_n29105__, new_new_n29106__, new_new_n29107__, new_new_n29108__,
    new_new_n29109__, new_new_n29110__, new_new_n29111__, new_new_n29112__,
    new_new_n29113__, new_new_n29114__, new_new_n29115__, new_new_n29116__,
    new_new_n29117__, new_new_n29118__, new_new_n29119__, new_new_n29120__,
    new_new_n29121__, new_new_n29122__, new_new_n29123__, new_new_n29124__,
    new_new_n29125__, new_new_n29126__, new_new_n29127__, new_new_n29128__,
    new_new_n29129__, new_new_n29130__, new_new_n29131__, new_new_n29132__,
    new_new_n29133__, new_new_n29134__, new_new_n29135__, new_new_n29136__,
    new_new_n29137__, new_new_n29138__, new_new_n29139__, new_new_n29140__,
    new_new_n29141__, new_new_n29142__, new_new_n29143__, new_new_n29144__,
    new_new_n29145__, new_new_n29146__, new_new_n29147__, new_new_n29148__,
    new_new_n29149__, new_new_n29150__, new_new_n29151__, new_new_n29152__,
    new_new_n29153__, new_new_n29154__, new_new_n29155__, new_new_n29156__,
    new_new_n29157__, new_new_n29158__, new_new_n29159__, new_new_n29160__,
    new_new_n29161__, new_new_n29162__, new_new_n29163__, new_new_n29164__,
    new_new_n29165__, new_new_n29166__, new_new_n29167__, new_new_n29168__,
    new_new_n29169__, new_new_n29170__, new_new_n29171__, new_new_n29172__,
    new_new_n29173__, new_new_n29174__, new_new_n29175__, new_new_n29176__,
    new_new_n29177__, new_new_n29178__, new_new_n29179__, new_new_n29180__,
    new_new_n29181__, new_new_n29182__, new_new_n29183__, new_new_n29184__,
    new_new_n29185__, new_new_n29186__, new_new_n29187__, new_new_n29188__,
    new_new_n29189__, new_new_n29190__, new_new_n29191__, new_new_n29192__,
    new_new_n29193__, new_new_n29194__, new_new_n29195__, new_new_n29196__,
    new_new_n29197__, new_new_n29198__, new_new_n29199__, new_new_n29200__,
    new_new_n29201__, new_new_n29202__, new_new_n29203__, new_new_n29204__,
    new_new_n29205__, new_new_n29206__, new_new_n29207__, new_new_n29208__,
    new_new_n29209__, new_new_n29210__, new_new_n29211__, new_new_n29212__,
    new_new_n29213__, new_new_n29214__, new_new_n29215__, new_new_n29216__,
    new_new_n29217__, new_new_n29218__, new_new_n29219__, new_new_n29220__,
    new_new_n29221__, new_new_n29222__, new_new_n29223__, new_new_n29224__,
    new_new_n29225__, new_new_n29226__, new_new_n29227__, new_new_n29228__,
    new_new_n29229__, new_new_n29230__, new_new_n29231__, new_new_n29232__,
    new_new_n29233__, new_new_n29234__, new_new_n29235__, new_new_n29236__,
    new_new_n29237__, new_new_n29238__, new_new_n29239__, new_new_n29240__,
    new_new_n29241__, new_new_n29242__, new_new_n29243__, new_new_n29244__,
    new_new_n29245__, new_new_n29246__, new_new_n29247__, new_new_n29248__,
    new_new_n29249__, new_new_n29250__, new_new_n29251__, new_new_n29252__,
    new_new_n29253__, new_new_n29254__, new_new_n29255__, new_new_n29256__,
    new_new_n29257__, new_new_n29258__, new_new_n29259__, new_new_n29260__,
    new_new_n29261__, new_new_n29262__, new_new_n29263__, new_new_n29264__,
    new_new_n29265__, new_new_n29266__, new_new_n29267__, new_new_n29268__,
    new_new_n29269__, new_new_n29270__, new_new_n29271__, new_new_n29272__,
    new_new_n29273__, new_new_n29274__, new_new_n29275__, new_new_n29276__,
    new_new_n29277__, new_new_n29278__, new_new_n29279__, new_new_n29280__,
    new_new_n29281__, new_new_n29282__, new_new_n29283__, new_new_n29284__,
    new_new_n29285__, new_new_n29286__, new_new_n29287__, new_new_n29288__,
    new_new_n29289__, new_new_n29290__, new_new_n29291__, new_new_n29292__,
    new_new_n29293__, new_new_n29294__, new_new_n29295__, new_new_n29296__,
    new_new_n29297__, new_new_n29298__, new_new_n29299__, new_new_n29300__,
    new_new_n29301__, new_new_n29302__, new_new_n29303__, new_new_n29304__,
    new_new_n29305__, new_new_n29306__, new_new_n29307__, new_new_n29308__,
    new_new_n29309__, new_new_n29310__, new_new_n29311__, new_new_n29312__,
    new_new_n29313__, new_new_n29314__, new_new_n29315__, new_new_n29316__,
    new_new_n29317__, new_new_n29318__, new_new_n29319__, new_new_n29320__,
    new_new_n29321__, new_new_n29322__, new_new_n29323__, new_new_n29324__,
    new_new_n29325__, new_new_n29326__, new_new_n29327__, new_new_n29328__,
    new_new_n29329__, new_new_n29330__, new_new_n29331__, new_new_n29332__,
    new_new_n29333__, new_new_n29334__, new_new_n29335__, new_new_n29336__,
    new_new_n29337__, new_new_n29338__, new_new_n29339__, new_new_n29340__,
    new_new_n29341__, new_new_n29342__, new_new_n29343__, new_new_n29344__,
    new_new_n29345__, new_new_n29346__, new_new_n29347__, new_new_n29348__,
    new_new_n29349__, new_new_n29350__, new_new_n29351__, new_new_n29352__,
    new_new_n29353__, new_new_n29354__, new_new_n29355__, new_new_n29356__,
    new_new_n29357__, new_new_n29358__, new_new_n29359__, new_new_n29360__,
    new_new_n29361__, new_new_n29362__, new_new_n29363__, new_new_n29364__,
    new_new_n29365__, new_new_n29366__, new_new_n29367__, new_new_n29368__,
    new_new_n29369__, new_new_n29370__, new_new_n29371__, new_new_n29372__,
    new_new_n29373__, new_new_n29374__, new_new_n29375__, new_new_n29376__,
    new_new_n29377__, new_new_n29378__, new_new_n29379__, new_new_n29380__,
    new_new_n29381__, new_new_n29382__, new_new_n29383__, new_new_n29384__,
    new_new_n29385__, new_new_n29386__, new_new_n29387__, new_new_n29388__,
    new_new_n29389__, new_new_n29390__, new_new_n29391__, new_new_n29392__,
    new_new_n29393__, new_new_n29394__, new_new_n29395__, new_new_n29396__,
    new_new_n29397__, new_new_n29398__, new_new_n29399__, new_new_n29400__,
    new_new_n29401__, new_new_n29402__, new_new_n29403__, new_new_n29404__,
    new_new_n29405__, new_new_n29406__, new_new_n29407__, new_new_n29408__,
    new_new_n29409__, new_new_n29410__, new_new_n29411__, new_new_n29412__,
    new_new_n29413__, new_new_n29414__, new_new_n29415__, new_new_n29416__,
    new_new_n29417__, new_new_n29418__, new_new_n29419__, new_new_n29420__,
    new_new_n29421__, new_new_n29422__, new_new_n29423__, new_new_n29424__,
    new_new_n29425__, new_new_n29426__, new_new_n29427__, new_new_n29428__,
    new_new_n29429__, new_new_n29430__, new_new_n29431__, new_new_n29432__,
    new_new_n29433__, new_new_n29434__, new_new_n29435__, new_new_n29436__,
    new_new_n29437__, new_new_n29438__, new_new_n29439__, new_new_n29440__,
    new_new_n29441__, new_new_n29442__, new_new_n29443__, new_new_n29444__,
    new_new_n29445__, new_new_n29446__, new_new_n29447__, new_new_n29448__,
    new_new_n29449__, new_new_n29450__, new_new_n29451__, new_new_n29452__,
    new_new_n29453__, new_new_n29454__, new_new_n29455__, new_new_n29456__,
    new_new_n29457__, new_new_n29458__, new_new_n29459__, new_new_n29460__,
    new_new_n29461__, new_new_n29462__, new_new_n29463__, new_new_n29464__,
    new_new_n29465__, new_new_n29466__, new_new_n29467__, new_new_n29468__,
    new_new_n29469__, new_new_n29470__, new_new_n29471__, new_new_n29472__,
    new_new_n29473__, new_new_n29474__, new_new_n29475__, new_new_n29476__,
    new_new_n29477__, new_new_n29478__, new_new_n29479__, new_new_n29480__,
    new_new_n29481__, new_new_n29482__, new_new_n29483__, new_new_n29484__,
    new_new_n29485__, new_new_n29486__, new_new_n29487__, new_new_n29488__,
    new_new_n29489__, new_new_n29490__, new_new_n29491__, new_new_n29492__,
    new_new_n29493__, new_new_n29494__, new_new_n29495__, new_new_n29496__,
    new_new_n29497__, new_new_n29498__, new_new_n29499__, new_new_n29500__,
    new_new_n29501__, new_new_n29502__, new_new_n29503__, new_new_n29504__,
    new_new_n29505__, new_new_n29506__, new_new_n29507__, new_new_n29508__,
    new_new_n29509__, new_new_n29510__, new_new_n29511__, new_new_n29512__,
    new_new_n29513__, new_new_n29514__, new_new_n29515__, new_new_n29516__,
    new_new_n29517__, new_new_n29518__, new_new_n29519__, new_new_n29520__,
    new_new_n29521__, new_new_n29522__, new_new_n29523__, new_new_n29524__,
    new_new_n29525__, new_new_n29526__, new_new_n29527__, new_new_n29528__,
    new_new_n29529__, new_new_n29530__, new_new_n29531__, new_new_n29532__,
    new_new_n29533__, new_new_n29534__, new_new_n29535__, new_new_n29536__,
    new_new_n29537__, new_new_n29538__, new_new_n29539__, new_new_n29540__,
    new_new_n29541__, new_new_n29542__, new_new_n29543__, new_new_n29544__,
    new_new_n29545__, new_new_n29546__, new_new_n29547__, new_new_n29548__,
    new_new_n29549__, new_new_n29550__, new_new_n29551__, new_new_n29552__,
    new_new_n29553__, new_new_n29554__, new_new_n29555__, new_new_n29556__,
    new_new_n29557__, new_new_n29558__, new_new_n29559__, new_new_n29560__,
    new_new_n29561__, new_new_n29562__, new_new_n29563__, new_new_n29564__,
    new_new_n29565__, new_new_n29566__, new_new_n29567__, new_new_n29568__,
    new_new_n29569__, new_new_n29570__, new_new_n29571__, new_new_n29572__,
    new_new_n29573__, new_new_n29574__, new_new_n29575__, new_new_n29576__,
    new_new_n29577__, new_new_n29578__, new_new_n29579__, new_new_n29580__,
    new_new_n29581__, new_new_n29582__, new_new_n29583__, new_new_n29584__,
    new_new_n29585__, new_new_n29586__, new_new_n29587__, new_new_n29588__,
    new_new_n29589__, new_new_n29590__, new_new_n29591__, new_new_n29592__,
    new_new_n29593__, new_new_n29594__, new_new_n29595__, new_new_n29596__,
    new_new_n29597__, new_new_n29598__, new_new_n29599__, new_new_n29600__,
    new_new_n29601__, new_new_n29602__, new_new_n29603__, new_new_n29604__,
    new_new_n29605__, new_new_n29606__, new_new_n29607__, new_new_n29608__,
    new_new_n29609__, new_new_n29610__, new_new_n29611__, new_new_n29612__,
    new_new_n29613__, new_new_n29614__, new_new_n29615__, new_new_n29616__,
    new_new_n29617__, new_new_n29618__, new_new_n29619__, new_new_n29620__,
    new_new_n29621__, new_new_n29622__, new_new_n29623__, new_new_n29624__,
    new_new_n29625__, new_new_n29626__, new_new_n29627__, new_new_n29628__,
    new_new_n29629__, new_new_n29630__, new_new_n29631__, new_new_n29632__,
    new_new_n29633__, new_new_n29634__, new_new_n29635__, new_new_n29636__,
    new_new_n29637__, new_new_n29638__, new_new_n29639__, new_new_n29640__,
    new_new_n29641__, new_new_n29642__, new_new_n29643__, new_new_n29644__,
    new_new_n29645__, new_new_n29646__, new_new_n29647__, new_new_n29648__,
    new_new_n29649__, new_new_n29650__, new_new_n29651__, new_new_n29652__,
    new_new_n29653__, new_new_n29654__, new_new_n29655__, new_new_n29656__,
    new_new_n29657__, new_new_n29658__, new_new_n29659__, new_new_n29660__,
    new_new_n29661__, new_new_n29662__, new_new_n29663__, new_new_n29664__,
    new_new_n29665__, new_new_n29666__, new_new_n29667__, new_new_n29668__,
    new_new_n29669__, new_new_n29670__, new_new_n29671__, new_new_n29672__,
    new_new_n29673__, new_new_n29674__, new_new_n29675__, new_new_n29676__,
    new_new_n29677__, new_new_n29678__, new_new_n29679__, new_new_n29680__,
    new_new_n29681__, new_new_n29682__, new_new_n29683__, new_new_n29684__,
    new_new_n29685__, new_new_n29686__, new_new_n29687__, new_new_n29688__,
    new_new_n29689__, new_new_n29690__, new_new_n29691__, new_new_n29692__,
    new_new_n29693__, new_new_n29694__, new_new_n29695__, new_new_n29696__,
    new_new_n29697__, new_new_n29698__, new_new_n29699__, new_new_n29700__,
    new_new_n29701__, new_new_n29702__, new_new_n29703__, new_new_n29704__,
    new_new_n29705__, new_new_n29706__, new_new_n29707__, new_new_n29708__,
    new_new_n29709__, new_new_n29710__, new_new_n29711__, new_new_n29712__,
    new_new_n29713__, new_new_n29714__, new_new_n29715__, new_new_n29716__,
    new_new_n29717__, new_new_n29718__, new_new_n29719__, new_new_n29720__,
    new_new_n29721__, new_new_n29722__, new_new_n29723__, new_new_n29724__,
    new_new_n29725__, new_new_n29726__, new_new_n29727__, new_new_n29728__,
    new_new_n29729__, new_new_n29730__, new_new_n29731__, new_new_n29732__,
    new_new_n29733__, new_new_n29734__, new_new_n29735__, new_new_n29736__,
    new_new_n29737__, new_new_n29738__, new_new_n29739__, new_new_n29740__,
    new_new_n29741__, new_new_n29742__, new_new_n29743__, new_new_n29744__,
    new_new_n29745__, new_new_n29746__, new_new_n29747__, new_new_n29748__,
    new_new_n29749__, new_new_n29750__, new_new_n29751__, new_new_n29752__,
    new_new_n29753__, new_new_n29754__, new_new_n29755__, new_new_n29756__,
    new_new_n29757__, new_new_n29758__, new_new_n29759__, new_new_n29760__,
    new_new_n29761__, new_new_n29762__, new_new_n29763__, new_new_n29764__,
    new_new_n29765__, new_new_n29766__, new_new_n29767__, new_new_n29768__,
    new_new_n29769__, new_new_n29770__, new_new_n29771__, new_new_n29772__,
    new_new_n29773__, new_new_n29774__, new_new_n29775__, new_new_n29776__,
    new_new_n29777__, new_new_n29778__, new_new_n29779__, new_new_n29780__,
    new_new_n29781__, new_new_n29782__, new_new_n29783__, new_new_n29784__,
    new_new_n29785__, new_new_n29786__, new_new_n29787__, new_new_n29788__,
    new_new_n29789__, new_new_n29790__, new_new_n29791__, new_new_n29792__,
    new_new_n29793__, new_new_n29794__, new_new_n29795__, new_new_n29796__,
    new_new_n29797__, new_new_n29798__, new_new_n29799__, new_new_n29800__,
    new_new_n29801__, new_new_n29802__, new_new_n29803__, new_new_n29804__,
    new_new_n29805__, new_new_n29806__, new_new_n29807__, new_new_n29808__,
    new_new_n29809__, new_new_n29810__, new_new_n29811__, new_new_n29812__,
    new_new_n29813__, new_new_n29814__, new_new_n29815__, new_new_n29816__,
    new_new_n29817__, new_new_n29818__, new_new_n29819__, new_new_n29820__,
    new_new_n29821__, new_new_n29822__, new_new_n29823__, new_new_n29824__,
    new_new_n29825__, new_new_n29826__, new_new_n29827__, new_new_n29828__,
    new_new_n29829__, new_new_n29830__, new_new_n29831__, new_new_n29832__,
    new_new_n29833__, new_new_n29834__, new_new_n29835__, new_new_n29836__,
    new_new_n29837__, new_new_n29838__, new_new_n29839__, new_new_n29840__,
    new_new_n29841__, new_new_n29842__, new_new_n29843__, new_new_n29844__,
    new_new_n29845__, new_new_n29846__, new_new_n29847__, new_new_n29848__,
    new_new_n29849__, new_new_n29850__, new_new_n29851__, new_new_n29852__,
    new_new_n29853__, new_new_n29854__, new_new_n29855__, new_new_n29856__,
    new_new_n29857__, new_new_n29858__, new_new_n29859__, new_new_n29860__,
    new_new_n29861__, new_new_n29862__, new_new_n29863__, new_new_n29864__,
    new_new_n29865__, new_new_n29866__, new_new_n29867__, new_new_n29868__,
    new_new_n29869__, new_new_n29870__, new_new_n29871__, new_new_n29872__,
    new_new_n29873__, new_new_n29874__, new_new_n29875__, new_new_n29876__,
    new_new_n29877__, new_new_n29878__, new_new_n29879__, new_new_n29880__,
    new_new_n29881__, new_new_n29882__, new_new_n29883__, new_new_n29884__,
    new_new_n29885__, new_new_n29886__, new_new_n29887__, new_new_n29888__,
    new_new_n29889__, new_new_n29890__, new_new_n29891__, new_new_n29892__,
    new_new_n29893__, new_new_n29894__, new_new_n29895__, new_new_n29896__,
    new_new_n29897__, new_new_n29898__, new_new_n29899__, new_new_n29900__,
    new_new_n29901__, new_new_n29902__, new_new_n29903__, new_new_n29904__,
    new_new_n29905__, new_new_n29906__, new_new_n29907__, new_new_n29908__,
    new_new_n29909__, new_new_n29910__, new_new_n29911__, new_new_n29912__,
    new_new_n29913__, new_new_n29914__, new_new_n29915__, new_new_n29916__,
    new_new_n29917__, new_new_n29918__, new_new_n29919__, new_new_n29920__,
    new_new_n29921__, new_new_n29922__, new_new_n29923__, new_new_n29924__,
    new_new_n29925__, new_new_n29926__, new_new_n29927__, new_new_n29928__,
    new_new_n29929__, new_new_n29930__, new_new_n29931__, new_new_n29932__,
    new_new_n29933__, new_new_n29934__, new_new_n29935__, new_new_n29936__,
    new_new_n29937__, new_new_n29938__, new_new_n29939__, new_new_n29940__,
    new_new_n29941__, new_new_n29942__, new_new_n29943__, new_new_n29944__,
    new_new_n29945__, new_new_n29946__, new_new_n29947__, new_new_n29948__,
    new_new_n29949__, new_new_n29950__, new_new_n29951__, new_new_n29952__,
    new_new_n29953__, new_new_n29954__, new_new_n29955__, new_new_n29956__,
    new_new_n29957__, new_new_n29958__, new_new_n29959__, new_new_n29960__,
    new_new_n29961__, new_new_n29962__, new_new_n29963__, new_new_n29964__,
    new_new_n29965__, new_new_n29966__, new_new_n29967__, new_new_n29968__,
    new_new_n29969__, new_new_n29970__, new_new_n29971__, new_new_n29972__,
    new_new_n29973__, new_new_n29974__, new_new_n29975__, new_new_n29976__,
    new_new_n29977__, new_new_n29978__, new_new_n29979__, new_new_n29980__,
    new_new_n29981__, new_new_n29982__, new_new_n29983__, new_new_n29984__,
    new_new_n29985__, new_new_n29986__, new_new_n29987__, new_new_n29988__,
    new_new_n29989__, new_new_n29990__, new_new_n29991__, new_new_n29992__,
    new_new_n29993__, new_new_n29994__, new_new_n29995__, new_new_n29996__,
    new_new_n29997__, new_new_n29998__, new_new_n29999__, new_new_n30000__,
    new_new_n30001__, new_new_n30002__, new_new_n30003__, new_new_n30004__,
    new_new_n30005__, new_new_n30006__, new_new_n30007__, new_new_n30008__,
    new_new_n30009__, new_new_n30010__, new_new_n30011__, new_new_n30012__,
    new_new_n30013__, new_new_n30014__, new_new_n30015__, new_new_n30016__,
    new_new_n30017__, new_new_n30018__, new_new_n30019__, new_new_n30020__,
    new_new_n30021__, new_new_n30022__, new_new_n30023__, new_new_n30024__,
    new_new_n30025__, new_new_n30026__, new_new_n30027__, new_new_n30028__,
    new_new_n30029__, new_new_n30030__, new_new_n30031__, new_new_n30032__,
    new_new_n30033__, new_new_n30034__, new_new_n30035__, new_new_n30036__,
    new_new_n30037__, new_new_n30038__, new_new_n30039__, new_new_n30040__,
    new_new_n30041__, new_new_n30042__, new_new_n30043__, new_new_n30044__,
    new_new_n30045__, new_new_n30046__, new_new_n30047__, new_new_n30048__,
    new_new_n30049__, new_new_n30050__, new_new_n30051__, new_new_n30052__,
    new_new_n30053__, new_new_n30054__, new_new_n30055__, new_new_n30056__,
    new_new_n30057__, new_new_n30058__, new_new_n30059__, new_new_n30060__,
    new_new_n30061__, new_new_n30062__, new_new_n30063__, new_new_n30064__,
    new_new_n30065__, new_new_n30066__, new_new_n30067__, new_new_n30068__,
    new_new_n30069__, new_new_n30070__, new_new_n30071__, new_new_n30072__,
    new_new_n30073__, new_new_n30074__, new_new_n30075__, new_new_n30076__,
    new_new_n30077__, new_new_n30078__, new_new_n30079__, new_new_n30080__,
    new_new_n30081__, new_new_n30082__, new_new_n30083__, new_new_n30084__,
    new_new_n30085__, new_new_n30086__, new_new_n30087__, new_new_n30088__,
    new_new_n30089__, new_new_n30090__, new_new_n30091__, new_new_n30092__,
    new_new_n30093__, new_new_n30094__, new_new_n30095__, new_new_n30096__,
    new_new_n30097__, new_new_n30098__, new_new_n30099__, new_new_n30100__,
    new_new_n30101__, new_new_n30102__, new_new_n30103__, new_new_n30104__,
    new_new_n30105__, new_new_n30106__, new_new_n30107__, new_new_n30108__,
    new_new_n30109__, new_new_n30110__, new_new_n30111__, new_new_n30112__,
    new_new_n30113__, new_new_n30114__, new_new_n30115__, new_new_n30116__,
    new_new_n30117__, new_new_n30118__, new_new_n30119__, new_new_n30120__,
    new_new_n30121__, new_new_n30122__, new_new_n30123__, new_new_n30124__,
    new_new_n30125__, new_new_n30126__, new_new_n30127__, new_new_n30128__,
    new_new_n30129__, new_new_n30130__, new_new_n30131__, new_new_n30132__,
    new_new_n30133__, new_new_n30134__, new_new_n30135__, new_new_n30136__,
    new_new_n30137__, new_new_n30138__, new_new_n30139__, new_new_n30140__,
    new_new_n30141__, new_new_n30142__, new_new_n30143__, new_new_n30144__,
    new_new_n30145__, new_new_n30146__, new_new_n30147__, new_new_n30148__,
    new_new_n30149__, new_new_n30150__, new_new_n30151__, new_new_n30152__,
    new_new_n30153__, new_new_n30154__, new_new_n30155__, new_new_n30156__,
    new_new_n30157__, new_new_n30158__, new_new_n30159__, new_new_n30160__,
    new_new_n30161__, new_new_n30162__, new_new_n30163__, new_new_n30164__,
    new_new_n30165__, new_new_n30166__, new_new_n30167__, new_new_n30168__,
    new_new_n30169__, new_new_n30170__, new_new_n30171__, new_new_n30172__,
    new_new_n30173__, new_new_n30174__, new_new_n30175__, new_new_n30176__,
    new_new_n30177__, new_new_n30178__, new_new_n30179__, new_new_n30180__,
    new_new_n30181__, new_new_n30182__, new_new_n30183__, new_new_n30184__,
    new_new_n30185__, new_new_n30186__, new_new_n30187__, new_new_n30188__,
    new_new_n30189__, new_new_n30190__, new_new_n30191__, new_new_n30192__,
    new_new_n30193__, new_new_n30194__, new_new_n30195__, new_new_n30196__,
    new_new_n30197__, new_new_n30198__, new_new_n30199__, new_new_n30200__,
    new_new_n30201__, new_new_n30202__, new_new_n30203__, new_new_n30204__,
    new_new_n30205__, new_new_n30206__, new_new_n30207__, new_new_n30208__,
    new_new_n30209__, new_new_n30210__, new_new_n30211__, new_new_n30212__,
    new_new_n30213__, new_new_n30214__, new_new_n30215__, new_new_n30216__,
    new_new_n30217__, new_new_n30218__, new_new_n30219__, new_new_n30220__,
    new_new_n30221__, new_new_n30222__, new_new_n30223__, new_new_n30224__,
    new_new_n30225__, new_new_n30226__, new_new_n30227__, new_new_n30228__,
    new_new_n30229__, new_new_n30230__, new_new_n30231__, new_new_n30232__,
    new_new_n30233__, new_new_n30234__, new_new_n30235__, new_new_n30236__,
    new_new_n30237__, new_new_n30238__, new_new_n30239__, new_new_n30240__,
    new_new_n30241__, new_new_n30242__, new_new_n30243__, new_new_n30244__,
    new_new_n30245__, new_new_n30246__, new_new_n30247__, new_new_n30248__,
    new_new_n30249__, new_new_n30250__, new_new_n30251__, new_new_n30252__,
    new_new_n30253__, new_new_n30254__, new_new_n30255__, new_new_n30256__,
    new_new_n30257__, new_new_n30258__, new_new_n30259__, new_new_n30260__,
    new_new_n30261__, new_new_n30262__, new_new_n30263__, new_new_n30264__,
    new_new_n30265__, new_new_n30266__, new_new_n30267__, new_new_n30268__,
    new_new_n30269__, new_new_n30270__, new_new_n30271__, new_new_n30272__,
    new_new_n30273__, new_new_n30274__, new_new_n30275__, new_new_n30276__,
    new_new_n30277__, new_new_n30278__, new_new_n30279__, new_new_n30280__,
    new_new_n30281__, new_new_n30282__, new_new_n30283__, new_new_n30284__,
    new_new_n30285__, new_new_n30286__, new_new_n30287__, new_new_n30288__,
    new_new_n30289__, new_new_n30290__, new_new_n30291__, new_new_n30292__,
    new_new_n30293__, new_new_n30294__, new_new_n30295__, new_new_n30296__,
    new_new_n30297__, new_new_n30298__, new_new_n30299__, new_new_n30300__,
    new_new_n30301__, new_new_n30302__, new_new_n30303__, new_new_n30304__,
    new_new_n30305__, new_new_n30306__, new_new_n30307__, new_new_n30308__,
    new_new_n30309__, new_new_n30310__, new_new_n30311__, new_new_n30312__,
    new_new_n30313__, new_new_n30314__, new_new_n30315__, new_new_n30316__,
    new_new_n30317__, new_new_n30318__, new_new_n30319__, new_new_n30320__,
    new_new_n30321__, new_new_n30322__, new_new_n30323__, new_new_n30324__,
    new_new_n30325__, new_new_n30326__, new_new_n30327__, new_new_n30328__,
    new_new_n30329__, new_new_n30330__, new_new_n30331__, new_new_n30332__,
    new_new_n30333__, new_new_n30334__, new_new_n30335__, new_new_n30336__,
    new_new_n30337__, new_new_n30338__, new_new_n30339__, new_new_n30340__,
    new_new_n30341__, new_new_n30342__, new_new_n30343__, new_new_n30344__,
    new_new_n30345__, new_new_n30346__, new_new_n30347__, new_new_n30348__,
    new_new_n30349__, new_new_n30350__, new_new_n30351__, new_new_n30352__,
    new_new_n30353__, new_new_n30354__, new_new_n30355__, new_new_n30356__,
    new_new_n30357__, new_new_n30358__, new_new_n30359__, new_new_n30360__,
    new_new_n30361__, new_new_n30362__, new_new_n30363__, new_new_n30364__,
    new_new_n30365__, new_new_n30366__, new_new_n30367__, new_new_n30368__,
    new_new_n30369__, new_new_n30370__, new_new_n30371__, new_new_n30372__,
    new_new_n30373__, new_new_n30374__, new_new_n30375__, new_new_n30376__,
    new_new_n30377__, new_new_n30378__, new_new_n30379__, new_new_n30380__,
    new_new_n30381__, new_new_n30382__, new_new_n30383__, new_new_n30384__,
    new_new_n30385__, new_new_n30386__, new_new_n30387__, new_new_n30388__,
    new_new_n30389__, new_new_n30390__, new_new_n30391__, new_new_n30392__,
    new_new_n30393__, new_new_n30394__, new_new_n30395__, new_new_n30396__,
    new_new_n30397__, new_new_n30398__, new_new_n30399__, new_new_n30400__,
    new_new_n30401__, new_new_n30402__, new_new_n30403__, new_new_n30404__,
    new_new_n30405__, new_new_n30406__, new_new_n30407__, new_new_n30408__,
    new_new_n30409__, new_new_n30410__, new_new_n30411__, new_new_n30412__,
    new_new_n30413__, new_new_n30414__, new_new_n30415__, new_new_n30416__,
    new_new_n30417__, new_new_n30418__, new_new_n30419__, new_new_n30420__,
    new_new_n30421__, new_new_n30422__, new_new_n30423__, new_new_n30424__,
    new_new_n30425__, new_new_n30426__, new_new_n30427__, new_new_n30428__,
    new_new_n30429__, new_new_n30430__, new_new_n30431__, new_new_n30432__,
    new_new_n30433__, new_new_n30434__, new_new_n30435__, new_new_n30436__,
    new_new_n30437__, new_new_n30438__, new_new_n30439__, new_new_n30440__,
    new_new_n30441__, new_new_n30442__, new_new_n30443__, new_new_n30444__,
    new_new_n30445__, new_new_n30446__, new_new_n30447__, new_new_n30448__,
    new_new_n30449__, new_new_n30450__, new_new_n30451__, new_new_n30452__,
    new_new_n30453__, new_new_n30454__, new_new_n30455__, new_new_n30456__,
    new_new_n30457__, new_new_n30458__, new_new_n30459__, new_new_n30460__,
    new_new_n30461__, new_new_n30462__, new_new_n30463__, new_new_n30464__,
    new_new_n30465__, new_new_n30466__, new_new_n30467__, new_new_n30468__,
    new_new_n30469__, new_new_n30470__, new_new_n30471__, new_new_n30472__,
    new_new_n30473__, new_new_n30474__, new_new_n30475__, new_new_n30476__,
    new_new_n30477__, new_new_n30478__, new_new_n30479__, new_new_n30480__,
    new_new_n30481__, new_new_n30482__, new_new_n30483__, new_new_n30484__,
    new_new_n30485__, new_new_n30486__, new_new_n30487__, new_new_n30488__,
    new_new_n30489__, new_new_n30490__, new_new_n30491__, new_new_n30492__,
    new_new_n30493__, new_new_n30494__, new_new_n30495__, new_new_n30496__,
    new_new_n30497__, new_new_n30498__, new_new_n30499__, new_new_n30500__,
    new_new_n30501__, new_new_n30502__, new_new_n30503__, new_new_n30504__,
    new_new_n30505__, new_new_n30506__, new_new_n30507__, new_new_n30508__,
    new_new_n30509__, new_new_n30510__, new_new_n30511__, new_new_n30512__,
    new_new_n30513__, new_new_n30514__, new_new_n30515__, new_new_n30516__,
    new_new_n30517__, new_new_n30518__, new_new_n30519__, new_new_n30520__,
    new_new_n30521__, new_new_n30522__, new_new_n30523__, new_new_n30524__,
    new_new_n30525__, new_new_n30526__, new_new_n30527__, new_new_n30528__,
    new_new_n30529__, new_new_n30530__, new_new_n30531__, new_new_n30532__,
    new_new_n30533__, new_new_n30534__, new_new_n30535__, new_new_n30536__,
    new_new_n30537__, new_new_n30538__, new_new_n30539__, new_new_n30540__,
    new_new_n30541__, new_new_n30542__, new_new_n30543__, new_new_n30544__,
    new_new_n30545__, new_new_n30546__, new_new_n30547__, new_new_n30548__,
    new_new_n30549__, new_new_n30550__, new_new_n30551__, new_new_n30552__,
    new_new_n30553__, new_new_n30554__, new_new_n30555__, new_new_n30556__,
    new_new_n30557__, new_new_n30558__, new_new_n30559__, new_new_n30560__,
    new_new_n30561__, new_new_n30562__, new_new_n30563__, new_new_n30564__,
    new_new_n30565__, new_new_n30566__, new_new_n30567__, new_new_n30568__,
    new_new_n30569__, new_new_n30570__, new_new_n30571__, new_new_n30572__,
    new_new_n30573__, new_new_n30574__, new_new_n30575__, new_new_n30576__,
    new_new_n30577__, new_new_n30578__, new_new_n30579__, new_new_n30580__,
    new_new_n30581__, new_new_n30582__, new_new_n30583__, new_new_n30584__,
    new_new_n30585__, new_new_n30586__, new_new_n30587__, new_new_n30588__,
    new_new_n30589__, new_new_n30590__, new_new_n30591__, new_new_n30592__,
    new_new_n30593__, new_new_n30594__, new_new_n30595__, new_new_n30596__,
    new_new_n30597__, new_new_n30598__, new_new_n30599__, new_new_n30600__,
    new_new_n30601__, new_new_n30602__, new_new_n30603__, new_new_n30604__,
    new_new_n30605__, new_new_n30606__, new_new_n30607__, new_new_n30608__,
    new_new_n30609__, new_new_n30610__, new_new_n30611__, new_new_n30612__,
    new_new_n30613__, new_new_n30614__, new_new_n30615__, new_new_n30616__,
    new_new_n30617__, new_new_n30618__, new_new_n30619__, new_new_n30620__,
    new_new_n30621__, new_new_n30622__, new_new_n30623__, new_new_n30624__,
    new_new_n30625__, new_new_n30626__, new_new_n30627__, new_new_n30628__,
    new_new_n30629__, new_new_n30630__, new_new_n30631__, new_new_n30632__,
    new_new_n30633__, new_new_n30634__, new_new_n30635__, new_new_n30636__,
    new_new_n30637__, new_new_n30638__, new_new_n30639__, new_new_n30640__,
    new_new_n30641__, new_new_n30642__, new_new_n30643__, new_new_n30644__,
    new_new_n30645__, new_new_n30646__, new_new_n30647__, new_new_n30648__,
    new_new_n30649__, new_new_n30650__, new_new_n30651__, new_new_n30652__,
    new_new_n30653__, new_new_n30654__, new_new_n30655__, new_new_n30656__,
    new_new_n30657__, new_new_n30658__, new_new_n30659__, new_new_n30660__,
    new_new_n30661__, new_new_n30662__, new_new_n30663__, new_new_n30664__,
    new_new_n30665__, new_new_n30666__, new_new_n30667__, new_new_n30668__,
    new_new_n30669__, new_new_n30670__, new_new_n30671__, new_new_n30672__,
    new_new_n30673__, new_new_n30674__, new_new_n30675__, new_new_n30676__,
    new_new_n30677__, new_new_n30678__, new_new_n30679__, new_new_n30680__,
    new_new_n30681__, new_new_n30682__, new_new_n30683__, new_new_n30684__,
    new_new_n30685__, new_new_n30686__, new_new_n30687__, new_new_n30688__,
    new_new_n30689__, new_new_n30690__, new_new_n30691__, new_new_n30692__,
    new_new_n30693__, new_new_n30694__, new_new_n30695__, new_new_n30696__,
    new_new_n30697__, new_new_n30698__, new_new_n30699__, new_new_n30700__,
    new_new_n30701__, new_new_n30702__, new_new_n30703__, new_new_n30704__,
    new_new_n30705__, new_new_n30706__, new_new_n30707__, new_new_n30708__,
    new_new_n30709__, new_new_n30710__, new_new_n30711__, new_new_n30712__,
    new_new_n30713__, new_new_n30714__, new_new_n30715__, new_new_n30716__,
    new_new_n30717__, new_new_n30718__, new_new_n30719__, new_new_n30720__,
    new_new_n30721__, new_new_n30722__, new_new_n30723__, new_new_n30724__,
    new_new_n30725__, new_new_n30726__, new_new_n30727__, new_new_n30728__,
    new_new_n30729__, new_new_n30730__, new_new_n30731__, new_new_n30732__,
    new_new_n30733__, new_new_n30734__, new_new_n30735__, new_new_n30736__,
    new_new_n30737__, new_new_n30738__, new_new_n30739__, new_new_n30740__,
    new_new_n30741__, new_new_n30742__, new_new_n30743__, new_new_n30744__,
    new_new_n30745__, new_new_n30746__, new_new_n30747__, new_new_n30748__,
    new_new_n30749__, new_new_n30750__, new_new_n30751__, new_new_n30752__,
    new_new_n30753__, new_new_n30754__, new_new_n30755__, new_new_n30756__,
    new_new_n30757__, new_new_n30758__, new_new_n30759__, new_new_n30760__,
    new_new_n30761__, new_new_n30762__, new_new_n30763__, new_new_n30764__,
    new_new_n30765__, new_new_n30766__, new_new_n30767__, new_new_n30768__,
    new_new_n30769__, new_new_n30770__, new_new_n30771__, new_new_n30772__,
    new_new_n30773__, new_new_n30774__, new_new_n30775__, new_new_n30776__,
    new_new_n30777__, new_new_n30778__, new_new_n30779__, new_new_n30780__,
    new_new_n30781__, new_new_n30782__, new_new_n30783__, new_new_n30784__,
    new_new_n30785__, new_new_n30786__, new_new_n30787__, new_new_n30788__,
    new_new_n30789__, new_new_n30790__, new_new_n30791__, new_new_n30792__,
    new_new_n30793__, new_new_n30794__, new_new_n30795__, new_new_n30796__,
    new_new_n30797__, new_new_n30798__, new_new_n30799__, new_new_n30800__,
    new_new_n30801__, new_new_n30802__, new_new_n30803__, new_new_n30804__,
    new_new_n30805__, new_new_n30806__, new_new_n30807__, new_new_n30808__,
    new_new_n30809__, new_new_n30810__, new_new_n30811__, new_new_n30812__,
    new_new_n30813__, new_new_n30814__, new_new_n30815__, new_new_n30816__,
    new_new_n30817__, new_new_n30818__, new_new_n30819__, new_new_n30820__,
    new_new_n30821__, new_new_n30822__, new_new_n30823__, new_new_n30824__,
    new_new_n30825__, new_new_n30826__, new_new_n30827__, new_new_n30828__,
    new_new_n30829__, new_new_n30830__, new_new_n30831__, new_new_n30832__,
    new_new_n30833__, new_new_n30834__, new_new_n30835__, new_new_n30836__,
    new_new_n30837__, new_new_n30838__, new_new_n30839__, new_new_n30840__,
    new_new_n30841__, new_new_n30842__, new_new_n30843__, new_new_n30844__,
    new_new_n30845__, new_new_n30846__, new_new_n30847__, new_new_n30848__,
    new_new_n30849__, new_new_n30850__, new_new_n30851__, new_new_n30852__,
    new_new_n30853__, new_new_n30854__, new_new_n30855__, new_new_n30856__,
    new_new_n30857__, new_new_n30858__, new_new_n30859__, new_new_n30860__,
    new_new_n30861__, new_new_n30862__, new_new_n30863__, new_new_n30864__,
    new_new_n30865__, new_new_n30866__, new_new_n30867__, new_new_n30868__,
    new_new_n30869__, new_new_n30870__, new_new_n30871__, new_new_n30872__,
    new_new_n30873__, new_new_n30874__, new_new_n30875__, new_new_n30876__,
    new_new_n30877__, new_new_n30878__, new_new_n30879__, new_new_n30880__,
    new_new_n30881__, new_new_n30882__, new_new_n30883__, new_new_n30884__,
    new_new_n30885__, new_new_n30886__, new_new_n30887__, new_new_n30888__,
    new_new_n30889__, new_new_n30890__, new_new_n30891__, new_new_n30892__,
    new_new_n30893__, new_new_n30894__, new_new_n30895__, new_new_n30896__,
    new_new_n30897__, new_new_n30898__, new_new_n30899__, new_new_n30900__,
    new_new_n30901__, new_new_n30902__, new_new_n30903__, new_new_n30904__,
    new_new_n30905__, new_new_n30906__, new_new_n30907__, new_new_n30908__,
    new_new_n30909__, new_new_n30910__, new_new_n30911__, new_new_n30912__,
    new_new_n30913__, new_new_n30914__, new_new_n30915__, new_new_n30916__,
    new_new_n30917__, new_new_n30918__, new_new_n30919__, new_new_n30920__,
    new_new_n30921__, new_new_n30922__, new_new_n30923__, new_new_n30924__,
    new_new_n30925__, new_new_n30926__, new_new_n30927__, new_new_n30928__,
    new_new_n30929__, new_new_n30930__, new_new_n30931__, new_new_n30932__,
    new_new_n30933__, new_new_n30934__, new_new_n30935__, new_new_n30936__,
    new_new_n30937__, new_new_n30938__, new_new_n30939__, new_new_n30940__,
    new_new_n30941__, new_new_n30942__, new_new_n30943__, new_new_n30944__,
    new_new_n30945__, new_new_n30946__, new_new_n30947__, new_new_n30948__,
    new_new_n30949__, new_new_n30950__, new_new_n30951__, new_new_n30952__,
    new_new_n30953__, new_new_n30954__, new_new_n30955__, new_new_n30956__,
    new_new_n30957__, new_new_n30958__, new_new_n30959__, new_new_n30960__,
    new_new_n30961__, new_new_n30962__, new_new_n30963__, new_new_n30964__,
    new_new_n30965__, new_new_n30966__, new_new_n30967__, new_new_n30968__,
    new_new_n30969__, new_new_n30970__, new_new_n30971__, new_new_n30972__,
    new_new_n30973__, new_new_n30974__, new_new_n30975__, new_new_n30976__,
    new_new_n30977__, new_new_n30978__, new_new_n30979__, new_new_n30980__,
    new_new_n30981__, new_new_n30982__, new_new_n30983__, new_new_n30984__,
    new_new_n30985__, new_new_n30986__, new_new_n30987__, new_new_n30988__,
    new_new_n30989__, new_new_n30990__, new_new_n30991__, new_new_n30992__,
    new_new_n30993__, new_new_n30994__, new_new_n30995__, new_new_n30996__,
    new_new_n30997__, new_new_n30998__, new_new_n30999__, new_new_n31000__,
    new_new_n31001__, new_new_n31002__, new_new_n31003__, new_new_n31004__,
    new_new_n31005__, new_new_n31006__, new_new_n31007__, new_new_n31008__,
    new_new_n31009__, new_new_n31010__, new_new_n31011__, new_new_n31012__,
    new_new_n31013__, new_new_n31014__, new_new_n31015__, new_new_n31016__,
    new_new_n31017__, new_new_n31018__, new_new_n31019__, new_new_n31020__,
    new_new_n31021__, new_new_n31022__, new_new_n31023__, new_new_n31024__,
    new_new_n31025__, new_new_n31026__, new_new_n31027__, new_new_n31028__,
    new_new_n31029__, new_new_n31030__, new_new_n31031__, new_new_n31032__,
    new_new_n31033__, new_new_n31034__, new_new_n31035__, new_new_n31036__,
    new_new_n31037__, new_new_n31038__, new_new_n31039__, new_new_n31040__,
    new_new_n31041__, new_new_n31042__, new_new_n31043__, new_new_n31044__,
    new_new_n31045__, new_new_n31046__, new_new_n31047__, new_new_n31048__,
    new_new_n31049__, new_new_n31050__, new_new_n31051__, new_new_n31052__,
    new_new_n31053__, new_new_n31054__, new_new_n31055__, new_new_n31056__,
    new_new_n31057__, new_new_n31058__, new_new_n31059__, new_new_n31060__,
    new_new_n31061__, new_new_n31062__, new_new_n31063__, new_new_n31064__,
    new_new_n31065__, new_new_n31066__, new_new_n31067__, new_new_n31068__,
    new_new_n31069__, new_new_n31070__, new_new_n31071__, new_new_n31072__,
    new_new_n31073__, new_new_n31074__, new_new_n31075__, new_new_n31076__,
    new_new_n31077__, new_new_n31078__, new_new_n31079__, new_new_n31080__,
    new_new_n31081__, new_new_n31082__, new_new_n31083__, new_new_n31084__,
    new_new_n31085__, new_new_n31086__, new_new_n31087__, new_new_n31088__,
    new_new_n31089__, new_new_n31090__, new_new_n31091__, new_new_n31092__,
    new_new_n31093__, new_new_n31094__, new_new_n31095__, new_new_n31096__,
    new_new_n31097__, new_new_n31098__, new_new_n31099__, new_new_n31100__,
    new_new_n31101__, new_new_n31102__, new_new_n31103__, new_new_n31104__,
    new_new_n31105__, new_new_n31106__, new_new_n31107__, new_new_n31108__,
    new_new_n31109__, new_new_n31110__, new_new_n31111__, new_new_n31112__,
    new_new_n31113__, new_new_n31114__, new_new_n31115__, new_new_n31116__,
    new_new_n31117__, new_new_n31118__, new_new_n31119__, new_new_n31120__,
    new_new_n31121__, new_new_n31122__, new_new_n31123__, new_new_n31124__,
    new_new_n31125__, new_new_n31126__, new_new_n31127__, new_new_n31128__,
    new_new_n31129__, new_new_n31130__, new_new_n31131__, new_new_n31132__,
    new_new_n31133__, new_new_n31134__, new_new_n31135__, new_new_n31136__,
    new_new_n31137__, new_new_n31138__, new_new_n31139__, new_new_n31140__,
    new_new_n31141__, new_new_n31142__, new_new_n31143__, new_new_n31144__,
    new_new_n31145__, new_new_n31146__, new_new_n31147__, new_new_n31148__,
    new_new_n31149__, new_new_n31150__, new_new_n31151__, new_new_n31152__,
    new_new_n31153__, new_new_n31154__, new_new_n31155__, new_new_n31156__,
    new_new_n31157__, new_new_n31158__, new_new_n31159__, new_new_n31160__,
    new_new_n31161__, new_new_n31162__, new_new_n31163__, new_new_n31164__,
    new_new_n31165__, new_new_n31166__, new_new_n31167__, new_new_n31168__,
    new_new_n31169__, new_new_n31170__, new_new_n31171__, new_new_n31172__,
    new_new_n31173__, new_new_n31174__, new_new_n31175__, new_new_n31176__,
    new_new_n31177__, new_new_n31178__, new_new_n31179__, new_new_n31180__,
    new_new_n31181__, new_new_n31182__, new_new_n31183__, new_new_n31184__,
    new_new_n31185__, new_new_n31186__, new_new_n31187__, new_new_n31188__,
    new_new_n31189__, new_new_n31190__, new_new_n31191__, new_new_n31192__,
    new_new_n31193__, new_new_n31194__, new_new_n31195__, new_new_n31196__,
    new_new_n31197__, new_new_n31198__, new_new_n31199__, new_new_n31200__,
    new_new_n31201__, new_new_n31202__, new_new_n31203__, new_new_n31204__,
    new_new_n31205__, new_new_n31206__, new_new_n31207__, new_new_n31208__,
    new_new_n31209__, new_new_n31210__, new_new_n31211__, new_new_n31212__,
    new_new_n31213__, new_new_n31214__, new_new_n31215__, new_new_n31216__,
    new_new_n31217__, new_new_n31218__, new_new_n31219__, new_new_n31220__,
    new_new_n31221__, new_new_n31222__, new_new_n31223__, new_new_n31224__,
    new_new_n31225__, new_new_n31226__, new_new_n31227__, new_new_n31228__,
    new_new_n31229__, new_new_n31230__, new_new_n31231__, new_new_n31232__,
    new_new_n31233__, new_new_n31234__, new_new_n31235__, new_new_n31236__,
    new_new_n31237__, new_new_n31238__, new_new_n31239__, new_new_n31240__,
    new_new_n31241__, new_new_n31242__, new_new_n31243__, new_new_n31244__,
    new_new_n31245__, new_new_n31246__, new_new_n31247__, new_new_n31248__,
    new_new_n31249__, new_new_n31250__, new_new_n31251__, new_new_n31252__,
    new_new_n31253__, new_new_n31254__, new_new_n31255__, new_new_n31256__,
    new_new_n31257__, new_new_n31258__, new_new_n31259__, new_new_n31260__,
    new_new_n31261__, new_new_n31262__, new_new_n31263__, new_new_n31264__,
    new_new_n31265__, new_new_n31266__, new_new_n31267__, new_new_n31268__,
    new_new_n31269__, new_new_n31270__, new_new_n31271__, new_new_n31272__,
    new_new_n31273__, new_new_n31274__, new_new_n31275__, new_new_n31276__,
    new_new_n31277__, new_new_n31278__, new_new_n31279__, new_new_n31280__,
    new_new_n31281__, new_new_n31282__, new_new_n31283__, new_new_n31284__,
    new_new_n31285__, new_new_n31286__, new_new_n31287__, new_new_n31288__,
    new_new_n31289__, new_new_n31290__, new_new_n31291__, new_new_n31292__,
    new_new_n31293__, new_new_n31294__, new_new_n31295__, new_new_n31296__,
    new_new_n31297__, new_new_n31298__, new_new_n31299__, new_new_n31300__,
    new_new_n31301__, new_new_n31302__, new_new_n31303__, new_new_n31304__,
    new_new_n31305__, new_new_n31306__, new_new_n31307__, new_new_n31308__,
    new_new_n31309__, new_new_n31310__, new_new_n31311__, new_new_n31312__,
    new_new_n31313__, new_new_n31314__, new_new_n31315__, new_new_n31316__,
    new_new_n31317__, new_new_n31318__, new_new_n31319__, new_new_n31320__,
    new_new_n31321__, new_new_n31322__, new_new_n31323__, new_new_n31324__,
    new_new_n31325__, new_new_n31326__, new_new_n31327__, new_new_n31328__,
    new_new_n31329__, new_new_n31330__, new_new_n31331__, new_new_n31332__,
    new_new_n31333__, new_new_n31334__, new_new_n31335__, new_new_n31336__,
    new_new_n31337__, new_new_n31338__, new_new_n31339__, new_new_n31340__,
    new_new_n31341__, new_new_n31342__, new_new_n31343__, new_new_n31344__,
    new_new_n31345__, new_new_n31346__, new_new_n31347__, new_new_n31348__,
    new_new_n31349__, new_new_n31350__, new_new_n31351__, new_new_n31352__,
    new_new_n31353__, new_new_n31354__, new_new_n31355__, new_new_n31356__,
    new_new_n31357__, new_new_n31358__, new_new_n31359__, new_new_n31360__,
    new_new_n31361__, new_new_n31362__, new_new_n31363__, new_new_n31364__,
    new_new_n31365__, new_new_n31366__, new_new_n31367__, new_new_n31368__,
    new_new_n31369__, new_new_n31370__, new_new_n31371__, new_new_n31372__,
    new_new_n31373__, new_new_n31374__, new_new_n31375__, new_new_n31376__,
    new_new_n31377__, new_new_n31378__, new_new_n31379__, new_new_n31380__,
    new_new_n31381__, new_new_n31382__, new_new_n31383__, new_new_n31384__,
    new_new_n31385__, new_new_n31386__, new_new_n31387__, new_new_n31388__,
    new_new_n31389__, new_new_n31390__, new_new_n31391__, new_new_n31392__,
    new_new_n31393__, new_new_n31394__, new_new_n31395__, new_new_n31396__,
    new_new_n31397__, new_new_n31398__, new_new_n31399__, new_new_n31400__,
    new_new_n31401__, new_new_n31402__, new_new_n31403__, new_new_n31404__,
    new_new_n31405__, new_new_n31406__, new_new_n31407__, new_new_n31408__,
    new_new_n31409__, new_new_n31410__, new_new_n31411__, new_new_n31412__,
    new_new_n31413__, new_new_n31414__, new_new_n31415__, new_new_n31416__,
    new_new_n31417__, new_new_n31418__, new_new_n31419__, new_new_n31420__,
    new_new_n31421__, new_new_n31422__, new_new_n31423__, new_new_n31424__,
    new_new_n31425__, new_new_n31426__, new_new_n31427__, new_new_n31428__,
    new_new_n31429__, new_new_n31430__, new_new_n31431__, new_new_n31432__,
    new_new_n31433__, new_new_n31434__, new_new_n31435__, new_new_n31436__,
    new_new_n31437__, new_new_n31438__, new_new_n31439__, new_new_n31440__,
    new_new_n31441__, new_new_n31442__, new_new_n31443__, new_new_n31444__,
    new_new_n31445__, new_new_n31446__, new_new_n31447__, new_new_n31448__,
    new_new_n31449__, new_new_n31450__, new_new_n31451__, new_new_n31452__,
    new_new_n31453__, new_new_n31454__, new_new_n31455__, new_new_n31456__,
    new_new_n31457__, new_new_n31458__, new_new_n31459__, new_new_n31460__,
    new_new_n31461__, new_new_n31462__, new_new_n31463__, new_new_n31464__,
    new_new_n31465__, new_new_n31466__, new_new_n31467__, new_new_n31468__,
    new_new_n31469__, new_new_n31470__, new_new_n31471__, new_new_n31472__,
    new_new_n31473__, new_new_n31474__, new_new_n31475__, new_new_n31476__,
    new_new_n31477__, new_new_n31478__, new_new_n31479__, new_new_n31480__,
    new_new_n31481__, new_new_n31482__, new_new_n31483__, new_new_n31484__,
    new_new_n31485__, new_new_n31486__, new_new_n31487__, new_new_n31488__,
    new_new_n31489__, new_new_n31490__, new_new_n31491__, new_new_n31492__,
    new_new_n31493__, new_new_n31494__, new_new_n31495__, new_new_n31496__,
    new_new_n31497__, new_new_n31498__, new_new_n31499__, new_new_n31500__,
    new_new_n31501__, new_new_n31502__, new_new_n31503__, new_new_n31504__,
    new_new_n31505__, new_new_n31506__, new_new_n31507__, new_new_n31508__,
    new_new_n31509__, new_new_n31510__, new_new_n31511__, new_new_n31512__,
    new_new_n31513__, new_new_n31514__, new_new_n31515__, new_new_n31516__,
    new_new_n31517__, new_new_n31518__, new_new_n31519__, new_new_n31520__,
    new_new_n31521__, new_new_n31522__, new_new_n31523__, new_new_n31524__,
    new_new_n31525__, new_new_n31526__, new_new_n31527__, new_new_n31528__,
    new_new_n31529__, new_new_n31530__, new_new_n31531__, new_new_n31532__,
    new_new_n31533__, new_new_n31534__, new_new_n31535__, new_new_n31536__,
    new_new_n31537__, new_new_n31538__, new_new_n31539__, new_new_n31540__,
    new_new_n31541__, new_new_n31542__, new_new_n31543__, new_new_n31544__,
    new_new_n31545__, new_new_n31546__, new_new_n31547__, new_new_n31548__,
    new_new_n31549__, new_new_n31550__, new_new_n31551__, new_new_n31552__,
    new_new_n31553__, new_new_n31554__, new_new_n31555__, new_new_n31556__,
    new_new_n31557__, new_new_n31558__, new_new_n31559__, new_new_n31560__,
    new_new_n31561__, new_new_n31562__, new_new_n31563__, new_new_n31564__,
    new_new_n31565__, new_new_n31566__, new_new_n31567__, new_new_n31568__,
    new_new_n31569__, new_new_n31570__, new_new_n31571__, new_new_n31572__,
    new_new_n31573__, new_new_n31574__, new_new_n31575__, new_new_n31576__,
    new_new_n31577__, new_new_n31578__, new_new_n31579__, new_new_n31580__,
    new_new_n31581__, new_new_n31582__, new_new_n31583__, new_new_n31584__,
    new_new_n31585__, new_new_n31586__, new_new_n31587__, new_new_n31588__,
    new_new_n31589__, new_new_n31590__, new_new_n31591__, new_new_n31592__,
    new_new_n31593__, new_new_n31594__, new_new_n31595__, new_new_n31596__,
    new_new_n31597__, new_new_n31598__, new_new_n31599__, new_new_n31600__,
    new_new_n31601__, new_new_n31602__, new_new_n31603__, new_new_n31604__,
    new_new_n31605__, new_new_n31606__, new_new_n31607__, new_new_n31608__,
    new_new_n31609__, new_new_n31610__, new_new_n31611__, new_new_n31612__,
    new_new_n31613__, new_new_n31614__, new_new_n31615__, new_new_n31616__,
    new_new_n31617__, new_new_n31618__, new_new_n31619__, new_new_n31620__,
    new_new_n31621__, new_new_n31622__, new_new_n31623__, new_new_n31624__,
    new_new_n31625__, new_new_n31626__, new_new_n31627__, new_new_n31628__,
    new_new_n31629__, new_new_n31630__, new_new_n31631__, new_new_n31632__,
    new_new_n31633__, new_new_n31634__, new_new_n31635__, new_new_n31636__,
    new_new_n31637__, new_new_n31638__, new_new_n31639__, new_new_n31640__,
    new_new_n31641__, new_new_n31642__, new_new_n31643__, new_new_n31644__,
    new_new_n31645__, new_new_n31646__, new_new_n31647__, new_new_n31648__,
    new_new_n31649__, new_new_n31650__, new_new_n31651__, new_new_n31652__,
    new_new_n31653__, new_new_n31654__, new_new_n31655__, new_new_n31656__,
    new_new_n31657__, new_new_n31658__, new_new_n31659__, new_new_n31660__,
    new_new_n31661__, new_new_n31662__, new_new_n31663__, new_new_n31664__,
    new_new_n31665__, new_new_n31666__, new_new_n31667__, new_new_n31668__,
    new_new_n31669__, new_new_n31670__, new_new_n31671__, new_new_n31672__,
    new_new_n31673__, new_new_n31674__, new_new_n31675__, new_new_n31676__,
    new_new_n31677__, new_new_n31678__, new_new_n31679__, new_new_n31680__,
    new_new_n31681__, new_new_n31682__, new_new_n31683__, new_new_n31684__,
    new_new_n31685__, new_new_n31686__, new_new_n31687__, new_new_n31688__,
    new_new_n31689__, new_new_n31690__, new_new_n31691__, new_new_n31692__,
    new_new_n31693__, new_new_n31694__, new_new_n31695__, new_new_n31696__,
    new_new_n31697__, new_new_n31698__, new_new_n31699__, new_new_n31700__,
    new_new_n31701__, new_new_n31702__, new_new_n31703__, new_new_n31704__,
    new_new_n31705__, new_new_n31706__, new_new_n31707__, new_new_n31708__,
    new_new_n31709__, new_new_n31710__, new_new_n31711__, new_new_n31712__,
    new_new_n31713__, new_new_n31714__, new_new_n31715__, new_new_n31716__,
    new_new_n31717__, new_new_n31718__, new_new_n31719__, new_new_n31720__,
    new_new_n31721__, new_new_n31722__, new_new_n31723__, new_new_n31724__,
    new_new_n31725__, new_new_n31726__, new_new_n31727__, new_new_n31728__,
    new_new_n31729__, new_new_n31730__, new_new_n31731__, new_new_n31732__,
    new_new_n31733__, new_new_n31734__, new_new_n31735__, new_new_n31736__,
    new_new_n31737__, new_new_n31738__, new_new_n31739__, new_new_n31740__,
    new_new_n31741__, new_new_n31742__, new_new_n31743__, new_new_n31744__,
    new_new_n31745__, new_new_n31746__, new_new_n31747__, new_new_n31748__,
    new_new_n31749__, new_new_n31750__, new_new_n31751__, new_new_n31752__,
    new_new_n31753__, new_new_n31754__, new_new_n31755__, new_new_n31756__,
    new_new_n31757__, new_new_n31758__, new_new_n31759__, new_new_n31760__,
    new_new_n31761__, new_new_n31762__, new_new_n31763__, new_new_n31764__,
    new_new_n31765__, new_new_n31766__, new_new_n31767__, new_new_n31768__,
    new_new_n31769__, new_new_n31770__, new_new_n31771__, new_new_n31772__,
    new_new_n31773__, new_new_n31774__, new_new_n31775__, new_new_n31776__,
    new_new_n31777__, new_new_n31778__, new_new_n31779__, new_new_n31780__,
    new_new_n31781__, new_new_n31782__, new_new_n31783__, new_new_n31784__,
    new_new_n31785__, new_new_n31786__, new_new_n31787__, new_new_n31788__,
    new_new_n31789__, new_new_n31790__, new_new_n31791__, new_new_n31792__,
    new_new_n31793__, new_new_n31794__, new_new_n31795__, new_new_n31796__,
    new_new_n31797__, new_new_n31798__, new_new_n31799__, new_new_n31800__,
    new_new_n31801__, new_new_n31802__, new_new_n31803__, new_new_n31804__,
    new_new_n31805__, new_new_n31806__, new_new_n31807__, new_new_n31808__,
    new_new_n31809__, new_new_n31810__, new_new_n31811__, new_new_n31812__,
    new_new_n31813__, new_new_n31814__, new_new_n31815__, new_new_n31816__,
    new_new_n31817__, new_new_n31818__, new_new_n31819__, new_new_n31820__,
    new_new_n31821__, new_new_n31822__, new_new_n31823__, new_new_n31824__,
    new_new_n31825__, new_new_n31826__, new_new_n31827__, new_new_n31828__,
    new_new_n31829__, new_new_n31830__, new_new_n31831__, new_new_n31832__,
    new_new_n31833__, new_new_n31834__, new_new_n31835__, new_new_n31836__,
    new_new_n31837__, new_new_n31838__, new_new_n31839__, new_new_n31840__,
    new_new_n31841__, new_new_n31842__, new_new_n31843__, new_new_n31844__,
    new_new_n31845__, new_new_n31846__, new_new_n31847__, new_new_n31848__,
    new_new_n31849__, new_new_n31850__, new_new_n31851__, new_new_n31852__,
    new_new_n31853__, new_new_n31854__, new_new_n31855__, new_new_n31856__,
    new_new_n31857__, new_new_n31858__, new_new_n31859__, new_new_n31860__,
    new_new_n31861__, new_new_n31862__, new_new_n31863__, new_new_n31864__,
    new_new_n31865__, new_new_n31866__, new_new_n31867__, new_new_n31868__,
    new_new_n31869__, new_new_n31870__, new_new_n31871__, new_new_n31872__,
    new_new_n31873__, new_new_n31874__, new_new_n31875__, new_new_n31876__,
    new_new_n31877__, new_new_n31878__, new_new_n31879__, new_new_n31880__,
    new_new_n31881__, new_new_n31882__, new_new_n31883__, new_new_n31884__,
    new_new_n31885__, new_new_n31886__, new_new_n31887__, new_new_n31888__,
    new_new_n31889__, new_new_n31890__, new_new_n31891__, new_new_n31892__,
    new_new_n31893__, new_new_n31894__, new_new_n31895__, new_new_n31896__,
    new_new_n31897__, new_new_n31898__, new_new_n31899__, new_new_n31900__,
    new_new_n31901__, new_new_n31902__, new_new_n31903__, new_new_n31904__,
    new_new_n31905__, new_new_n31906__, new_new_n31907__, new_new_n31908__,
    new_new_n31909__, new_new_n31910__, new_new_n31911__, new_new_n31912__,
    new_new_n31913__, new_new_n31914__, new_new_n31915__, new_new_n31916__,
    new_new_n31917__, new_new_n31918__, new_new_n31919__, new_new_n31920__,
    new_new_n31921__, new_new_n31922__, new_new_n31923__, new_new_n31924__,
    new_new_n31925__, new_new_n31926__, new_new_n31927__, new_new_n31928__,
    new_new_n31929__, new_new_n31930__, new_new_n31931__, new_new_n31932__,
    new_new_n31933__, new_new_n31934__, new_new_n31935__, new_new_n31936__,
    new_new_n31937__, new_new_n31938__, new_new_n31939__, new_new_n31940__,
    new_new_n31941__, new_new_n31942__, new_new_n31943__, new_new_n31944__,
    new_new_n31945__, new_new_n31946__, new_new_n31947__, new_new_n31948__,
    new_new_n31949__, new_new_n31950__, new_new_n31951__, new_new_n31952__,
    new_new_n31953__, new_new_n31954__, new_new_n31955__, new_new_n31956__,
    new_new_n31957__, new_new_n31958__, new_new_n31959__, new_new_n31960__,
    new_new_n31961__, new_new_n31962__, new_new_n31963__, new_new_n31964__,
    new_new_n31965__, new_new_n31966__, new_new_n31967__, new_new_n31968__,
    new_new_n31969__, new_new_n31970__, new_new_n31971__, new_new_n31972__,
    new_new_n31973__, new_new_n31974__, new_new_n31975__, new_new_n31976__,
    new_new_n31977__, new_new_n31978__, new_new_n31979__, new_new_n31980__,
    new_new_n31981__, new_new_n31982__, new_new_n31983__, new_new_n31984__,
    new_new_n31985__, new_new_n31986__, new_new_n31987__, new_new_n31988__,
    new_new_n31989__, new_new_n31990__, new_new_n31991__, new_new_n31992__,
    new_new_n31993__, new_new_n31994__, new_new_n31995__, new_new_n31996__,
    new_new_n31997__, new_new_n31998__, new_new_n31999__, new_new_n32000__,
    new_new_n32001__, new_new_n32002__, new_new_n32003__, new_new_n32004__,
    new_new_n32005__, new_new_n32006__, new_new_n32007__, new_new_n32008__,
    new_new_n32009__, new_new_n32010__, new_new_n32011__, new_new_n32012__,
    new_new_n32013__, new_new_n32014__, new_new_n32015__, new_new_n32016__,
    new_new_n32017__, new_new_n32018__, new_new_n32019__, new_new_n32020__,
    new_new_n32021__, new_new_n32022__, new_new_n32023__, new_new_n32024__,
    new_new_n32025__, new_new_n32026__, new_new_n32027__, new_new_n32028__,
    new_new_n32029__, new_new_n32030__, new_new_n32031__, new_new_n32032__,
    new_new_n32033__, new_new_n32034__, new_new_n32035__, new_new_n32036__,
    new_new_n32037__, new_new_n32038__, new_new_n32039__, new_new_n32040__,
    new_new_n32041__, new_new_n32042__, new_new_n32043__, new_new_n32044__,
    new_new_n32045__, new_new_n32046__, new_new_n32047__, new_new_n32048__,
    new_new_n32049__, new_new_n32050__, new_new_n32051__, new_new_n32052__,
    new_new_n32053__, new_new_n32054__, new_new_n32055__, new_new_n32056__,
    new_new_n32057__, new_new_n32058__, new_new_n32059__, new_new_n32060__,
    new_new_n32061__, new_new_n32062__, new_new_n32063__, new_new_n32064__,
    new_new_n32065__, new_new_n32066__, new_new_n32067__, new_new_n32068__,
    new_new_n32069__, new_new_n32070__, new_new_n32071__, new_new_n32072__,
    new_new_n32073__, new_new_n32074__, new_new_n32075__, new_new_n32076__,
    new_new_n32077__, new_new_n32078__, new_new_n32079__, new_new_n32080__,
    new_new_n32081__, new_new_n32082__, new_new_n32083__, new_new_n32084__,
    new_new_n32085__, new_new_n32086__, new_new_n32087__, new_new_n32088__,
    new_new_n32089__, new_new_n32090__, new_new_n32091__, new_new_n32092__,
    new_new_n32093__, new_new_n32094__, new_new_n32095__, new_new_n32096__,
    new_new_n32097__, new_new_n32098__, new_new_n32099__, new_new_n32100__,
    new_new_n32101__, new_new_n32102__, new_new_n32103__, new_new_n32104__,
    new_new_n32105__, new_new_n32106__, new_new_n32107__, new_new_n32108__,
    new_new_n32109__, new_new_n32110__, new_new_n32111__, new_new_n32112__,
    new_new_n32113__, new_new_n32114__, new_new_n32115__, new_new_n32116__,
    new_new_n32117__, new_new_n32118__, new_new_n32119__, new_new_n32120__,
    new_new_n32121__, new_new_n32122__, new_new_n32123__, new_new_n32124__,
    new_new_n32125__, new_new_n32126__, new_new_n32127__, new_new_n32128__,
    new_new_n32129__, new_new_n32130__, new_new_n32131__, new_new_n32132__,
    new_new_n32133__, new_new_n32134__, new_new_n32135__, new_new_n32136__,
    new_new_n32137__, new_new_n32138__, new_new_n32139__, new_new_n32140__,
    new_new_n32141__, new_new_n32142__, new_new_n32143__, new_new_n32144__,
    new_new_n32145__, new_new_n32146__, new_new_n32147__, new_new_n32148__,
    new_new_n32149__, new_new_n32150__, new_new_n32151__, new_new_n32152__,
    new_new_n32153__, new_new_n32154__, new_new_n32155__, new_new_n32156__,
    new_new_n32157__, new_new_n32158__, new_new_n32159__, new_new_n32160__,
    new_new_n32161__, new_new_n32162__, new_new_n32163__, new_new_n32164__,
    new_new_n32165__, new_new_n32166__, new_new_n32167__, new_new_n32168__,
    new_new_n32169__, new_new_n32170__, new_new_n32171__, new_new_n32172__,
    new_new_n32173__, new_new_n32174__, new_new_n32175__, new_new_n32176__,
    new_new_n32177__, new_new_n32178__, new_new_n32179__, new_new_n32180__,
    new_new_n32181__, new_new_n32182__, new_new_n32183__, new_new_n32184__,
    new_new_n32185__, new_new_n32186__, new_new_n32187__, new_new_n32188__,
    new_new_n32189__, new_new_n32190__, new_new_n32191__, new_new_n32192__,
    new_new_n32193__, new_new_n32194__, new_new_n32195__, new_new_n32196__,
    new_new_n32197__, new_new_n32198__, new_new_n32199__, new_new_n32200__,
    new_new_n32201__, new_new_n32202__, new_new_n32203__, new_new_n32204__,
    new_new_n32205__, new_new_n32206__, new_new_n32207__, new_new_n32208__,
    new_new_n32209__, new_new_n32210__, new_new_n32211__, new_new_n32212__,
    new_new_n32213__, new_new_n32214__, new_new_n32215__, new_new_n32216__,
    new_new_n32217__, new_new_n32218__, new_new_n32219__, new_new_n32220__,
    new_new_n32221__, new_new_n32222__, new_new_n32223__, new_new_n32224__,
    new_new_n32225__, new_new_n32226__, new_new_n32227__, new_new_n32228__,
    new_new_n32229__, new_new_n32230__, new_new_n32231__, new_new_n32232__,
    new_new_n32233__, new_new_n32234__, new_new_n32235__, new_new_n32236__,
    new_new_n32237__, new_new_n32238__, new_new_n32239__, new_new_n32240__,
    new_new_n32241__, new_new_n32242__, new_new_n32243__, new_new_n32244__,
    new_new_n32245__, new_new_n32246__, new_new_n32247__, new_new_n32248__,
    new_new_n32249__, new_new_n32250__, new_new_n32251__, new_new_n32252__,
    new_new_n32253__, new_new_n32254__, new_new_n32255__, new_new_n32256__,
    new_new_n32257__, new_new_n32258__, new_new_n32259__, new_new_n32260__,
    new_new_n32261__, new_new_n32262__, new_new_n32263__, new_new_n32264__,
    new_new_n32265__, new_new_n32266__, new_new_n32267__, new_new_n32268__,
    new_new_n32269__, new_new_n32270__, new_new_n32271__, new_new_n32272__,
    new_new_n32273__, new_new_n32274__, new_new_n32275__, new_new_n32276__,
    new_new_n32277__, new_new_n32278__, new_new_n32279__, new_new_n32280__,
    new_new_n32281__, new_new_n32282__, new_new_n32283__, new_new_n32284__,
    new_new_n32285__, new_new_n32286__, new_new_n32287__, new_new_n32288__,
    new_new_n32289__, new_new_n32290__, new_new_n32291__, new_new_n32292__,
    new_new_n32293__, new_new_n32294__, new_new_n32295__, new_new_n32296__,
    new_new_n32297__, new_new_n32298__, new_new_n32299__, new_new_n32300__,
    new_new_n32301__, new_new_n32302__, new_new_n32303__, new_new_n32304__,
    new_new_n32305__, new_new_n32306__, new_new_n32307__, new_new_n32308__,
    new_new_n32309__, new_new_n32310__, new_new_n32311__, new_new_n32312__,
    new_new_n32313__, new_new_n32314__, new_new_n32315__, new_new_n32316__,
    new_new_n32317__, new_new_n32318__, new_new_n32319__, new_new_n32320__,
    new_new_n32321__, new_new_n32322__, new_new_n32323__, new_new_n32324__,
    new_new_n32325__, new_new_n32326__, new_new_n32328__, new_new_n32329__,
    new_new_n32330__, new_new_n32331__, new_new_n32332__, new_new_n32333__,
    new_new_n32334__, new_new_n32335__, new_new_n32336__, new_new_n32337__,
    new_new_n32338__, new_new_n32339__, new_new_n32340__, new_new_n32341__,
    new_new_n32342__, new_new_n32343__, new_new_n32344__, new_new_n32345__,
    new_new_n32346__, new_new_n32347__, new_new_n32348__, new_new_n32349__,
    new_new_n32350__, new_new_n32351__, new_new_n32352__, new_new_n32353__,
    new_new_n32354__, new_new_n32355__, new_new_n32356__, new_new_n32357__,
    new_new_n32358__, new_new_n32359__, new_new_n32360__, new_new_n32361__,
    new_new_n32362__, new_new_n32363__, new_new_n32364__, new_new_n32365__,
    new_new_n32366__, new_new_n32367__, new_new_n32368__, new_new_n32369__,
    new_new_n32370__, new_new_n32371__, new_new_n32372__, new_new_n32373__,
    new_new_n32374__, new_new_n32375__, new_new_n32376__, new_new_n32377__,
    new_new_n32378__, new_new_n32379__, new_new_n32380__, new_new_n32381__,
    new_new_n32382__, new_new_n32383__, new_new_n32384__, new_new_n32385__,
    new_new_n32386__, new_new_n32387__, new_new_n32388__, new_new_n32389__,
    new_new_n32390__, new_new_n32391__, new_new_n32392__, new_new_n32393__,
    new_new_n32394__, new_new_n32395__, new_new_n32396__, new_new_n32397__,
    new_new_n32398__, new_new_n32399__, new_new_n32400__, new_new_n32401__,
    new_new_n32402__, new_new_n32403__, new_new_n32404__, new_new_n32405__,
    new_new_n32406__, new_new_n32407__, new_new_n32408__, new_new_n32409__,
    new_new_n32410__, new_new_n32411__, new_new_n32412__, new_new_n32413__,
    new_new_n32414__, new_new_n32415__, new_new_n32416__, new_new_n32417__,
    new_new_n32418__, new_new_n32419__, new_new_n32420__, new_new_n32421__,
    new_new_n32422__, new_new_n32423__, new_new_n32424__, new_new_n32425__,
    new_new_n32426__, new_new_n32427__, new_new_n32428__, new_new_n32429__,
    new_new_n32430__, new_new_n32431__, new_new_n32432__, new_new_n32433__,
    new_new_n32434__, new_new_n32435__, new_new_n32436__, new_new_n32437__,
    new_new_n32438__, new_new_n32439__, new_new_n32440__, new_new_n32441__,
    new_new_n32442__, new_new_n32443__, new_new_n32444__, new_new_n32445__,
    new_new_n32446__, new_new_n32447__, new_new_n32448__, new_new_n32449__,
    new_new_n32450__, new_new_n32451__, new_new_n32452__, new_new_n32453__,
    new_new_n32454__, new_new_n32455__, new_new_n32456__, new_new_n32457__,
    new_new_n32458__, new_new_n32459__, new_new_n32460__, new_new_n32461__,
    new_new_n32462__, new_new_n32463__, new_new_n32464__, new_new_n32465__,
    new_new_n32466__, new_new_n32467__, new_new_n32468__, new_new_n32469__,
    new_new_n32470__, new_new_n32471__, new_new_n32472__, new_new_n32473__,
    new_new_n32474__, new_new_n32475__, new_new_n32476__, new_new_n32477__,
    new_new_n32478__, new_new_n32479__, new_new_n32480__, new_new_n32481__,
    new_new_n32482__, new_new_n32483__, new_new_n32484__, new_new_n32485__,
    new_new_n32486__, new_new_n32487__, new_new_n32488__, new_new_n32489__,
    new_new_n32490__, new_new_n32491__, new_new_n32492__, new_new_n32493__,
    new_new_n32494__, new_new_n32495__, new_new_n32496__, new_new_n32497__,
    new_new_n32498__, new_new_n32499__, new_new_n32500__, new_new_n32501__,
    new_new_n32502__, new_new_n32503__, new_new_n32504__, new_new_n32505__,
    new_new_n32506__, new_new_n32507__, new_new_n32508__, new_new_n32509__,
    new_new_n32510__, new_new_n32511__, new_new_n32512__, new_new_n32513__,
    new_new_n32514__, new_new_n32515__, new_new_n32516__, new_new_n32517__,
    new_new_n32518__, new_new_n32519__, new_new_n32520__, new_new_n32521__,
    new_new_n32522__, new_new_n32523__, new_new_n32524__, new_new_n32525__,
    new_new_n32526__, new_new_n32527__, new_new_n32528__, new_new_n32529__,
    new_new_n32530__, new_new_n32531__, new_new_n32532__, new_new_n32533__,
    new_new_n32534__, new_new_n32535__, new_new_n32536__, new_new_n32537__,
    new_new_n32538__, new_new_n32539__, new_new_n32540__, new_new_n32541__,
    new_new_n32542__, new_new_n32543__, new_new_n32544__, new_new_n32545__,
    new_new_n32546__, new_new_n32547__, new_new_n32548__, new_new_n32549__,
    new_new_n32550__, new_new_n32551__, new_new_n32552__, new_new_n32553__,
    new_new_n32554__, new_new_n32555__, new_new_n32556__, new_new_n32557__,
    new_new_n32558__, new_new_n32559__, new_new_n32560__, new_new_n32561__,
    new_new_n32562__, new_new_n32563__, new_new_n32564__, new_new_n32565__,
    new_new_n32566__, new_new_n32567__, new_new_n32568__, new_new_n32569__,
    new_new_n32570__, new_new_n32571__, new_new_n32572__, new_new_n32573__,
    new_new_n32574__, new_new_n32575__, new_new_n32576__, new_new_n32577__,
    new_new_n32578__, new_new_n32579__, new_new_n32580__, new_new_n32581__,
    new_new_n32582__, new_new_n32583__, new_new_n32584__, new_new_n32585__,
    new_new_n32586__, new_new_n32587__, new_new_n32588__, new_new_n32589__,
    new_new_n32590__, new_new_n32591__, new_new_n32592__, new_new_n32593__,
    new_new_n32594__, new_new_n32595__, new_new_n32596__, new_new_n32597__,
    new_new_n32598__, new_new_n32599__, new_new_n32600__, new_new_n32601__,
    new_new_n32602__, new_new_n32603__, new_new_n32604__, new_new_n32605__,
    new_new_n32606__, new_new_n32607__, new_new_n32608__, new_new_n32609__,
    new_new_n32610__, new_new_n32611__, new_new_n32612__, new_new_n32613__,
    new_new_n32614__, new_new_n32615__, new_new_n32616__, new_new_n32617__,
    new_new_n32618__, new_new_n32619__, new_new_n32620__, new_new_n32621__,
    new_new_n32622__, new_new_n32623__, new_new_n32624__, new_new_n32625__,
    new_new_n32626__, new_new_n32627__, new_new_n32628__, new_new_n32629__,
    new_new_n32630__, new_new_n32631__, new_new_n32632__, new_new_n32633__,
    new_new_n32634__, new_new_n32635__, new_new_n32636__, new_new_n32637__,
    new_new_n32638__, new_new_n32639__, new_new_n32640__, new_new_n32641__,
    new_new_n32642__, new_new_n32643__, new_new_n32644__, new_new_n32645__,
    new_new_n32646__, new_new_n32647__, new_new_n32648__, new_new_n32649__,
    new_new_n32650__, new_new_n32651__, new_new_n32652__, new_new_n32653__,
    new_new_n32654__, new_new_n32655__, new_new_n32656__, new_new_n32657__,
    new_new_n32658__, new_new_n32659__, new_new_n32660__, new_new_n32661__,
    new_new_n32662__, new_new_n32663__, new_new_n32664__, new_new_n32665__,
    new_new_n32666__, new_new_n32667__, new_new_n32668__, new_new_n32669__,
    new_new_n32670__, new_new_n32671__, new_new_n32672__, new_new_n32673__,
    new_new_n32674__, new_new_n32675__, new_new_n32676__, new_new_n32678__,
    new_new_n32679__, new_new_n32680__, new_new_n32681__, new_new_n32682__,
    new_new_n32683__, new_new_n32684__, new_new_n32685__, new_new_n32686__,
    new_new_n32687__, new_new_n32688__, new_new_n32689__, new_new_n32690__,
    new_new_n32691__, new_new_n32692__, new_new_n32693__, new_new_n32694__,
    new_new_n32695__, new_new_n32696__, new_new_n32697__, new_new_n32698__,
    new_new_n32699__, new_new_n32700__, new_new_n32701__, new_new_n32702__,
    new_new_n32703__, new_new_n32704__, new_new_n32705__, new_new_n32706__,
    new_new_n32707__, new_new_n32708__, new_new_n32709__, new_new_n32710__,
    new_new_n32711__, new_new_n32712__, new_new_n32713__, new_new_n32714__,
    new_new_n32715__, new_new_n32716__, new_new_n32717__, new_new_n32718__,
    new_new_n32719__, new_new_n32720__, new_new_n32721__, new_new_n32722__,
    new_new_n32723__, new_new_n32724__, new_new_n32725__, new_new_n32726__,
    new_new_n32727__, new_new_n32728__, new_new_n32729__, new_new_n32730__,
    new_new_n32731__, new_new_n32732__, new_new_n32733__, new_new_n32734__,
    new_new_n32735__, new_new_n32736__, new_new_n32737__, new_new_n32738__,
    new_new_n32739__, new_new_n32740__, new_new_n32741__, new_new_n32742__,
    new_new_n32743__, new_new_n32744__, new_new_n32745__, new_new_n32746__,
    new_new_n32747__, new_new_n32748__, new_new_n32749__, new_new_n32750__,
    new_new_n32751__, new_new_n32752__, new_new_n32753__, new_new_n32754__,
    new_new_n32755__, new_new_n32756__, new_new_n32757__, new_new_n32758__,
    new_new_n32759__, new_new_n32760__, new_new_n32761__, new_new_n32762__,
    new_new_n32763__, new_new_n32764__, new_new_n32765__, new_new_n32766__,
    new_new_n32767__, new_new_n32768__, new_new_n32769__, new_new_n32770__,
    new_new_n32771__, new_new_n32772__, new_new_n32773__, new_new_n32774__,
    new_new_n32775__, new_new_n32776__, new_new_n32777__, new_new_n32778__,
    new_new_n32779__, new_new_n32780__, new_new_n32781__, new_new_n32782__,
    new_new_n32783__, new_new_n32784__, new_new_n32785__, new_new_n32786__,
    new_new_n32787__, new_new_n32788__, new_new_n32789__, new_new_n32790__,
    new_new_n32791__, new_new_n32792__, new_new_n32793__, new_new_n32794__,
    new_new_n32795__, new_new_n32796__, new_new_n32797__, new_new_n32798__,
    new_new_n32799__, new_new_n32800__, new_new_n32801__, new_new_n32802__,
    new_new_n32803__, new_new_n32804__, new_new_n32805__, new_new_n32806__,
    new_new_n32807__, new_new_n32808__, new_new_n32809__, new_new_n32810__,
    new_new_n32811__, new_new_n32812__, new_new_n32813__, new_new_n32814__,
    new_new_n32815__, new_new_n32816__, new_new_n32817__, new_new_n32818__,
    new_new_n32819__, new_new_n32820__, new_new_n32821__, new_new_n32822__,
    new_new_n32823__, new_new_n32824__, new_new_n32825__, new_new_n32826__,
    new_new_n32827__, new_new_n32828__, new_new_n32829__, new_new_n32830__,
    new_new_n32831__, new_new_n32832__, new_new_n32833__, new_new_n32834__,
    new_new_n32835__, new_new_n32836__, new_new_n32837__, new_new_n32838__,
    new_new_n32839__, new_new_n32840__, new_new_n32841__, new_new_n32842__,
    new_new_n32843__, new_new_n32844__, new_new_n32845__, new_new_n32846__,
    new_new_n32847__, new_new_n32848__, new_new_n32849__, new_new_n32850__,
    new_new_n32851__, new_new_n32852__, new_new_n32853__, new_new_n32854__,
    new_new_n32855__, new_new_n32856__, new_new_n32857__, new_new_n32858__,
    new_new_n32859__, new_new_n32860__, new_new_n32861__, new_new_n32862__,
    new_new_n32863__, new_new_n32864__, new_new_n32865__, new_new_n32866__,
    new_new_n32867__, new_new_n32868__, new_new_n32869__, new_new_n32870__,
    new_new_n32871__, new_new_n32872__, new_new_n32873__, new_new_n32874__,
    new_new_n32875__, new_new_n32876__, new_new_n32877__, new_new_n32878__,
    new_new_n32879__, new_new_n32880__, new_new_n32881__, new_new_n32882__,
    new_new_n32883__, new_new_n32884__, new_new_n32885__, new_new_n32886__,
    new_new_n32887__, new_new_n32888__, new_new_n32889__, new_new_n32890__,
    new_new_n32891__, new_new_n32892__, new_new_n32893__, new_new_n32894__,
    new_new_n32895__, new_new_n32896__, new_new_n32897__, new_new_n32898__,
    new_new_n32899__, new_new_n32900__, new_new_n32901__, new_new_n32902__,
    new_new_n32903__, new_new_n32904__, new_new_n32905__, new_new_n32906__,
    new_new_n32907__, new_new_n32908__, new_new_n32909__, new_new_n32910__,
    new_new_n32911__, new_new_n32912__, new_new_n32913__, new_new_n32914__,
    new_new_n32915__, new_new_n32916__, new_new_n32917__, new_new_n32918__,
    new_new_n32919__, new_new_n32920__, new_new_n32921__, new_new_n32922__,
    new_new_n32923__, new_new_n32924__, new_new_n32925__, new_new_n32926__,
    new_new_n32927__, new_new_n32928__, new_new_n32929__, new_new_n32930__,
    new_new_n32931__, new_new_n32932__, new_new_n32933__, new_new_n32934__,
    new_new_n32935__, new_new_n32936__, new_new_n32937__, new_new_n32938__,
    new_new_n32939__, new_new_n32940__, new_new_n32941__, new_new_n32942__,
    new_new_n32943__, new_new_n32944__, new_new_n32945__, new_new_n32946__,
    new_new_n32947__, new_new_n32948__, new_new_n32949__, new_new_n32950__,
    new_new_n32951__, new_new_n32952__, new_new_n32953__, new_new_n32954__,
    new_new_n32955__, new_new_n32956__, new_new_n32957__, new_new_n32958__,
    new_new_n32959__, new_new_n32960__, new_new_n32961__, new_new_n32962__,
    new_new_n32963__, new_new_n32964__, new_new_n32965__, new_new_n32966__,
    new_new_n32967__, new_new_n32968__, new_new_n32969__, new_new_n32970__,
    new_new_n32971__, new_new_n32972__, new_new_n32973__, new_new_n32974__,
    new_new_n32975__, new_new_n32976__, new_new_n32977__, new_new_n32978__,
    new_new_n32979__, new_new_n32980__, new_new_n32981__, new_new_n32982__,
    new_new_n32983__, new_new_n32984__, new_new_n32985__, new_new_n32986__,
    new_new_n32987__, new_new_n32988__, new_new_n32989__, new_new_n32990__,
    new_new_n32991__, new_new_n32992__, new_new_n32993__, new_new_n32994__,
    new_new_n32995__, new_new_n32996__, new_new_n32997__, new_new_n32998__,
    new_new_n32999__, new_new_n33000__, new_new_n33001__, new_new_n33002__,
    new_new_n33003__, new_new_n33004__, new_new_n33005__, new_new_n33006__,
    new_new_n33007__, new_new_n33008__, new_new_n33009__, new_new_n33010__,
    new_new_n33011__, new_new_n33012__, new_new_n33013__, new_new_n33014__,
    new_new_n33015__, new_new_n33016__, new_new_n33017__, new_new_n33018__,
    new_new_n33019__, new_new_n33020__, new_new_n33021__, new_new_n33022__,
    new_new_n33023__, new_new_n33024__, new_new_n33025__, new_new_n33026__,
    new_new_n33027__, new_new_n33028__, new_new_n33029__, new_new_n33030__,
    new_new_n33031__, new_new_n33032__, new_new_n33033__, new_new_n33034__,
    new_new_n33035__, new_new_n33036__, new_new_n33037__, new_new_n33038__,
    new_new_n33039__, new_new_n33040__, new_new_n33042__, new_new_n33043__,
    new_new_n33044__, new_new_n33045__, new_new_n33046__, new_new_n33047__,
    new_new_n33048__, new_new_n33049__, new_new_n33050__, new_new_n33051__,
    new_new_n33052__, new_new_n33053__, new_new_n33054__, new_new_n33055__,
    new_new_n33056__, new_new_n33057__, new_new_n33058__, new_new_n33059__,
    new_new_n33060__, new_new_n33061__, new_new_n33062__, new_new_n33063__,
    new_new_n33064__, new_new_n33065__, new_new_n33066__, new_new_n33067__,
    new_new_n33068__, new_new_n33069__, new_new_n33070__, new_new_n33071__,
    new_new_n33072__, new_new_n33073__, new_new_n33074__, new_new_n33075__,
    new_new_n33076__, new_new_n33077__, new_new_n33078__, new_new_n33079__,
    new_new_n33080__, new_new_n33081__, new_new_n33082__, new_new_n33083__,
    new_new_n33084__, new_new_n33085__, new_new_n33086__, new_new_n33087__,
    new_new_n33088__, new_new_n33089__, new_new_n33090__, new_new_n33091__,
    new_new_n33092__, new_new_n33093__, new_new_n33094__, new_new_n33095__,
    new_new_n33096__, new_new_n33097__, new_new_n33098__, new_new_n33099__,
    new_new_n33100__, new_new_n33101__, new_new_n33102__, new_new_n33103__,
    new_new_n33104__, new_new_n33105__, new_new_n33106__, new_new_n33107__,
    new_new_n33108__, new_new_n33109__, new_new_n33110__, new_new_n33111__,
    new_new_n33112__, new_new_n33113__, new_new_n33114__, new_new_n33115__,
    new_new_n33116__, new_new_n33117__, new_new_n33118__, new_new_n33119__,
    new_new_n33120__, new_new_n33121__, new_new_n33122__, new_new_n33123__,
    new_new_n33124__, new_new_n33125__, new_new_n33126__, new_new_n33127__,
    new_new_n33128__, new_new_n33129__, new_new_n33130__, new_new_n33131__,
    new_new_n33132__, new_new_n33133__, new_new_n33134__, new_new_n33135__,
    new_new_n33136__, new_new_n33137__, new_new_n33138__, new_new_n33139__,
    new_new_n33140__, new_new_n33141__, new_new_n33142__, new_new_n33143__,
    new_new_n33144__, new_new_n33145__, new_new_n33146__, new_new_n33147__,
    new_new_n33148__, new_new_n33149__, new_new_n33150__, new_new_n33151__,
    new_new_n33152__, new_new_n33153__, new_new_n33154__, new_new_n33155__,
    new_new_n33156__, new_new_n33157__, new_new_n33158__, new_new_n33159__,
    new_new_n33160__, new_new_n33161__, new_new_n33162__, new_new_n33163__,
    new_new_n33164__, new_new_n33165__, new_new_n33166__, new_new_n33167__,
    new_new_n33168__, new_new_n33169__, new_new_n33170__, new_new_n33171__,
    new_new_n33172__, new_new_n33173__, new_new_n33174__, new_new_n33175__,
    new_new_n33176__, new_new_n33177__, new_new_n33178__, new_new_n33179__,
    new_new_n33180__, new_new_n33181__, new_new_n33182__, new_new_n33183__,
    new_new_n33184__, new_new_n33185__, new_new_n33186__, new_new_n33187__,
    new_new_n33188__, new_new_n33189__, new_new_n33190__, new_new_n33191__,
    new_new_n33192__, new_new_n33193__, new_new_n33194__, new_new_n33195__,
    new_new_n33196__, new_new_n33197__, new_new_n33198__, new_new_n33199__,
    new_new_n33200__, new_new_n33201__, new_new_n33202__, new_new_n33203__,
    new_new_n33204__, new_new_n33205__, new_new_n33206__, new_new_n33207__,
    new_new_n33208__, new_new_n33209__, new_new_n33210__, new_new_n33211__,
    new_new_n33212__, new_new_n33213__, new_new_n33214__, new_new_n33215__,
    new_new_n33216__, new_new_n33217__, new_new_n33218__, new_new_n33219__,
    new_new_n33220__, new_new_n33221__, new_new_n33222__, new_new_n33223__,
    new_new_n33224__, new_new_n33225__, new_new_n33226__, new_new_n33227__,
    new_new_n33228__, new_new_n33229__, new_new_n33230__, new_new_n33231__,
    new_new_n33232__, new_new_n33233__, new_new_n33234__, new_new_n33235__,
    new_new_n33236__, new_new_n33237__, new_new_n33238__, new_new_n33239__,
    new_new_n33240__, new_new_n33241__, new_new_n33242__, new_new_n33243__,
    new_new_n33244__, new_new_n33245__, new_new_n33246__, new_new_n33247__,
    new_new_n33248__, new_new_n33249__, new_new_n33250__, new_new_n33251__,
    new_new_n33252__, new_new_n33253__, new_new_n33254__, new_new_n33255__,
    new_new_n33256__, new_new_n33257__, new_new_n33258__, new_new_n33259__,
    new_new_n33260__, new_new_n33261__, new_new_n33262__, new_new_n33263__,
    new_new_n33264__, new_new_n33265__, new_new_n33266__, new_new_n33267__,
    new_new_n33268__, new_new_n33269__, new_new_n33270__, new_new_n33271__,
    new_new_n33272__, new_new_n33273__, new_new_n33274__, new_new_n33275__,
    new_new_n33276__, new_new_n33277__, new_new_n33278__, new_new_n33279__,
    new_new_n33280__, new_new_n33281__, new_new_n33282__, new_new_n33283__,
    new_new_n33284__, new_new_n33285__, new_new_n33286__, new_new_n33287__,
    new_new_n33288__, new_new_n33289__, new_new_n33290__, new_new_n33291__,
    new_new_n33292__, new_new_n33293__, new_new_n33294__, new_new_n33295__,
    new_new_n33296__, new_new_n33297__, new_new_n33298__, new_new_n33299__,
    new_new_n33300__, new_new_n33301__, new_new_n33302__, new_new_n33303__,
    new_new_n33304__, new_new_n33305__, new_new_n33306__, new_new_n33307__,
    new_new_n33308__, new_new_n33309__, new_new_n33311__, new_new_n33312__,
    new_new_n33313__, new_new_n33314__, new_new_n33315__, new_new_n33316__,
    new_new_n33317__, new_new_n33318__, new_new_n33319__, new_new_n33320__,
    new_new_n33321__, new_new_n33322__, new_new_n33323__, new_new_n33324__,
    new_new_n33325__, new_new_n33326__, new_new_n33327__, new_new_n33328__,
    new_new_n33329__, new_new_n33330__, new_new_n33331__, new_new_n33332__,
    new_new_n33333__, new_new_n33334__, new_new_n33335__, new_new_n33336__,
    new_new_n33337__, new_new_n33338__, new_new_n33339__, new_new_n33340__,
    new_new_n33341__, new_new_n33342__, new_new_n33343__, new_new_n33344__,
    new_new_n33345__, new_new_n33346__, new_new_n33347__, new_new_n33348__,
    new_new_n33349__, new_new_n33350__, new_new_n33351__, new_new_n33352__,
    new_new_n33353__, new_new_n33354__, new_new_n33355__, new_new_n33356__,
    new_new_n33357__, new_new_n33358__, new_new_n33359__, new_new_n33360__,
    new_new_n33361__, new_new_n33362__, new_new_n33363__, new_new_n33364__,
    new_new_n33365__, new_new_n33366__, new_new_n33367__, new_new_n33368__,
    new_new_n33369__, new_new_n33370__, new_new_n33371__, new_new_n33372__,
    new_new_n33373__, new_new_n33374__, new_new_n33375__, new_new_n33376__,
    new_new_n33377__, new_new_n33378__, new_new_n33379__, new_new_n33380__,
    new_new_n33381__, new_new_n33382__, new_new_n33383__, new_new_n33384__,
    new_new_n33385__, new_new_n33386__, new_new_n33387__, new_new_n33388__,
    new_new_n33389__, new_new_n33390__, new_new_n33391__, new_new_n33392__,
    new_new_n33393__, new_new_n33394__, new_new_n33395__, new_new_n33396__,
    new_new_n33397__, new_new_n33398__, new_new_n33399__, new_new_n33400__,
    new_new_n33401__, new_new_n33402__, new_new_n33403__, new_new_n33404__,
    new_new_n33405__, new_new_n33406__, new_new_n33407__, new_new_n33408__,
    new_new_n33409__, new_new_n33410__, new_new_n33411__, new_new_n33412__,
    new_new_n33413__, new_new_n33414__, new_new_n33415__, new_new_n33416__,
    new_new_n33417__, new_new_n33418__, new_new_n33419__, new_new_n33420__,
    new_new_n33421__, new_new_n33422__, new_new_n33423__, new_new_n33424__,
    new_new_n33425__, new_new_n33426__, new_new_n33427__, new_new_n33428__,
    new_new_n33429__, new_new_n33430__, new_new_n33431__, new_new_n33432__,
    new_new_n33433__, new_new_n33434__, new_new_n33435__, new_new_n33436__,
    new_new_n33437__, new_new_n33438__, new_new_n33439__, new_new_n33440__,
    new_new_n33441__, new_new_n33442__, new_new_n33443__, new_new_n33444__,
    new_new_n33445__, new_new_n33446__, new_new_n33447__, new_new_n33448__,
    new_new_n33449__, new_new_n33450__, new_new_n33451__, new_new_n33452__,
    new_new_n33453__, new_new_n33454__, new_new_n33455__, new_new_n33456__,
    new_new_n33457__, new_new_n33458__, new_new_n33459__, new_new_n33460__,
    new_new_n33461__, new_new_n33462__, new_new_n33463__, new_new_n33464__,
    new_new_n33465__, new_new_n33466__, new_new_n33467__, new_new_n33468__,
    new_new_n33469__, new_new_n33470__, new_new_n33471__, new_new_n33472__,
    new_new_n33473__, new_new_n33474__, new_new_n33475__, new_new_n33476__,
    new_new_n33477__, new_new_n33478__, new_new_n33479__, new_new_n33480__,
    new_new_n33481__, new_new_n33482__, new_new_n33483__, new_new_n33484__,
    new_new_n33485__, new_new_n33486__, new_new_n33487__, new_new_n33488__,
    new_new_n33489__, new_new_n33490__, new_new_n33491__, new_new_n33492__,
    new_new_n33493__, new_new_n33494__, new_new_n33495__, new_new_n33496__,
    new_new_n33497__, new_new_n33498__, new_new_n33499__, new_new_n33500__,
    new_new_n33501__, new_new_n33502__, new_new_n33503__, new_new_n33504__,
    new_new_n33505__, new_new_n33506__, new_new_n33507__, new_new_n33508__,
    new_new_n33509__, new_new_n33510__, new_new_n33511__, new_new_n33512__,
    new_new_n33513__, new_new_n33514__, new_new_n33515__, new_new_n33516__,
    new_new_n33517__, new_new_n33518__, new_new_n33519__, new_new_n33520__,
    new_new_n33521__, new_new_n33522__, new_new_n33523__, new_new_n33524__,
    new_new_n33525__, new_new_n33526__, new_new_n33527__, new_new_n33528__,
    new_new_n33529__, new_new_n33530__, new_new_n33531__, new_new_n33532__,
    new_new_n33533__, new_new_n33534__, new_new_n33535__, new_new_n33536__,
    new_new_n33537__, new_new_n33538__, new_new_n33539__, new_new_n33540__,
    new_new_n33541__, new_new_n33542__, new_new_n33543__, new_new_n33544__,
    new_new_n33545__, new_new_n33546__, new_new_n33547__, new_new_n33548__,
    new_new_n33549__, new_new_n33550__, new_new_n33551__, new_new_n33552__,
    new_new_n33553__, new_new_n33554__, new_new_n33555__, new_new_n33556__,
    new_new_n33557__, new_new_n33558__, new_new_n33559__, new_new_n33560__,
    new_new_n33561__, new_new_n33562__, new_new_n33563__, new_new_n33564__,
    new_new_n33565__, new_new_n33566__, new_new_n33567__, new_new_n33568__,
    new_new_n33569__, new_new_n33570__, new_new_n33571__, new_new_n33572__,
    new_new_n33573__, new_new_n33574__, new_new_n33575__, new_new_n33576__,
    new_new_n33577__, new_new_n33578__, new_new_n33579__, new_new_n33580__,
    new_new_n33581__, new_new_n33582__, new_new_n33583__, new_new_n33584__,
    new_new_n33585__, new_new_n33586__, new_new_n33587__, new_new_n33588__,
    new_new_n33589__, new_new_n33590__, new_new_n33591__, new_new_n33592__,
    new_new_n33593__, new_new_n33594__, new_new_n33595__, new_new_n33597__,
    new_new_n33598__, new_new_n33599__, new_new_n33600__, new_new_n33601__,
    new_new_n33602__, new_new_n33603__, new_new_n33604__, new_new_n33605__,
    new_new_n33606__, new_new_n33607__, new_new_n33608__, new_new_n33609__,
    new_new_n33610__, new_new_n33611__, new_new_n33612__, new_new_n33613__,
    new_new_n33614__, new_new_n33615__, new_new_n33616__, new_new_n33617__,
    new_new_n33618__, new_new_n33619__, new_new_n33620__, new_new_n33621__,
    new_new_n33622__, new_new_n33623__, new_new_n33624__, new_new_n33625__,
    new_new_n33626__, new_new_n33627__, new_new_n33628__, new_new_n33629__,
    new_new_n33630__, new_new_n33631__, new_new_n33632__, new_new_n33633__,
    new_new_n33634__, new_new_n33635__, new_new_n33636__, new_new_n33637__,
    new_new_n33638__, new_new_n33639__, new_new_n33640__, new_new_n33641__,
    new_new_n33642__, new_new_n33643__, new_new_n33644__, new_new_n33645__,
    new_new_n33646__, new_new_n33647__, new_new_n33648__, new_new_n33649__,
    new_new_n33650__, new_new_n33651__, new_new_n33652__, new_new_n33653__,
    new_new_n33654__, new_new_n33655__, new_new_n33656__, new_new_n33657__,
    new_new_n33658__, new_new_n33659__, new_new_n33660__, new_new_n33661__,
    new_new_n33662__, new_new_n33663__, new_new_n33664__, new_new_n33665__,
    new_new_n33666__, new_new_n33667__, new_new_n33668__, new_new_n33669__,
    new_new_n33670__, new_new_n33671__, new_new_n33672__, new_new_n33673__,
    new_new_n33674__, new_new_n33675__, new_new_n33676__, new_new_n33677__,
    new_new_n33678__, new_new_n33679__, new_new_n33680__, new_new_n33681__,
    new_new_n33682__, new_new_n33683__, new_new_n33684__, new_new_n33685__,
    new_new_n33686__, new_new_n33687__, new_new_n33688__, new_new_n33689__,
    new_new_n33690__, new_new_n33691__, new_new_n33692__, new_new_n33693__,
    new_new_n33694__, new_new_n33695__, new_new_n33696__, new_new_n33697__,
    new_new_n33698__, new_new_n33699__, new_new_n33700__, new_new_n33701__,
    new_new_n33702__, new_new_n33703__, new_new_n33704__, new_new_n33705__,
    new_new_n33706__, new_new_n33707__, new_new_n33708__, new_new_n33709__,
    new_new_n33710__, new_new_n33711__, new_new_n33712__, new_new_n33713__,
    new_new_n33714__, new_new_n33715__, new_new_n33716__, new_new_n33717__,
    new_new_n33718__, new_new_n33719__, new_new_n33720__, new_new_n33721__,
    new_new_n33722__, new_new_n33723__, new_new_n33724__, new_new_n33725__,
    new_new_n33726__, new_new_n33727__, new_new_n33728__, new_new_n33729__,
    new_new_n33730__, new_new_n33731__, new_new_n33732__, new_new_n33733__,
    new_new_n33734__, new_new_n33735__, new_new_n33736__, new_new_n33737__,
    new_new_n33738__, new_new_n33739__, new_new_n33740__, new_new_n33741__,
    new_new_n33742__, new_new_n33743__, new_new_n33744__, new_new_n33745__,
    new_new_n33746__, new_new_n33747__, new_new_n33748__, new_new_n33749__,
    new_new_n33750__, new_new_n33751__, new_new_n33752__, new_new_n33753__,
    new_new_n33754__, new_new_n33755__, new_new_n33756__, new_new_n33757__,
    new_new_n33758__, new_new_n33759__, new_new_n33760__, new_new_n33761__,
    new_new_n33762__, new_new_n33763__, new_new_n33764__, new_new_n33765__,
    new_new_n33766__, new_new_n33767__, new_new_n33768__, new_new_n33769__,
    new_new_n33770__, new_new_n33771__, new_new_n33772__, new_new_n33773__,
    new_new_n33774__, new_new_n33775__, new_new_n33776__, new_new_n33777__,
    new_new_n33778__, new_new_n33779__, new_new_n33780__, new_new_n33781__,
    new_new_n33782__, new_new_n33783__, new_new_n33784__, new_new_n33785__,
    new_new_n33786__, new_new_n33787__, new_new_n33788__, new_new_n33789__,
    new_new_n33790__, new_new_n33791__, new_new_n33792__, new_new_n33793__,
    new_new_n33794__, new_new_n33795__, new_new_n33796__, new_new_n33797__,
    new_new_n33798__, new_new_n33799__, new_new_n33800__, new_new_n33801__,
    new_new_n33802__, new_new_n33803__, new_new_n33804__, new_new_n33805__,
    new_new_n33806__, new_new_n33807__, new_new_n33808__, new_new_n33809__,
    new_new_n33810__, new_new_n33811__, new_new_n33812__, new_new_n33813__,
    new_new_n33814__, new_new_n33815__, new_new_n33816__, new_new_n33817__,
    new_new_n33818__, new_new_n33819__, new_new_n33820__, new_new_n33821__,
    new_new_n33822__, new_new_n33823__, new_new_n33824__, new_new_n33825__,
    new_new_n33826__, new_new_n33827__, new_new_n33828__, new_new_n33829__,
    new_new_n33830__, new_new_n33831__, new_new_n33832__, new_new_n33833__,
    new_new_n33834__, new_new_n33835__, new_new_n33836__, new_new_n33837__,
    new_new_n33838__, new_new_n33839__, new_new_n33840__, new_new_n33841__,
    new_new_n33842__, new_new_n33843__, new_new_n33844__, new_new_n33845__,
    new_new_n33846__, new_new_n33847__, new_new_n33848__, new_new_n33849__,
    new_new_n33850__, new_new_n33851__, new_new_n33852__, new_new_n33853__,
    new_new_n33854__, new_new_n33855__, new_new_n33856__, new_new_n33857__,
    new_new_n33858__, new_new_n33859__, new_new_n33860__, new_new_n33861__,
    new_new_n33862__, new_new_n33863__, new_new_n33864__, new_new_n33865__,
    new_new_n33866__, new_new_n33867__, new_new_n33868__, new_new_n33869__,
    new_new_n33870__, new_new_n33871__, new_new_n33872__, new_new_n33873__,
    new_new_n33874__, new_new_n33875__, new_new_n33876__, new_new_n33877__,
    new_new_n33879__, new_new_n33880__, new_new_n33881__, new_new_n33882__,
    new_new_n33883__, new_new_n33884__, new_new_n33885__, new_new_n33886__,
    new_new_n33887__, new_new_n33888__, new_new_n33889__, new_new_n33890__,
    new_new_n33891__, new_new_n33892__, new_new_n33893__, new_new_n33894__,
    new_new_n33895__, new_new_n33896__, new_new_n33897__, new_new_n33898__,
    new_new_n33899__, new_new_n33900__, new_new_n33901__, new_new_n33902__,
    new_new_n33903__, new_new_n33904__, new_new_n33905__, new_new_n33906__,
    new_new_n33907__, new_new_n33908__, new_new_n33909__, new_new_n33910__,
    new_new_n33911__, new_new_n33912__, new_new_n33913__, new_new_n33914__,
    new_new_n33915__, new_new_n33916__, new_new_n33917__, new_new_n33918__,
    new_new_n33919__, new_new_n33920__, new_new_n33921__, new_new_n33922__,
    new_new_n33923__, new_new_n33924__, new_new_n33925__, new_new_n33926__,
    new_new_n33927__, new_new_n33928__, new_new_n33929__, new_new_n33930__,
    new_new_n33931__, new_new_n33932__, new_new_n33933__, new_new_n33934__,
    new_new_n33935__, new_new_n33936__, new_new_n33937__, new_new_n33938__,
    new_new_n33939__, new_new_n33940__, new_new_n33941__, new_new_n33942__,
    new_new_n33943__, new_new_n33944__, new_new_n33945__, new_new_n33946__,
    new_new_n33947__, new_new_n33948__, new_new_n33949__, new_new_n33950__,
    new_new_n33951__, new_new_n33952__, new_new_n33953__, new_new_n33954__,
    new_new_n33955__, new_new_n33956__, new_new_n33957__, new_new_n33958__,
    new_new_n33959__, new_new_n33960__, new_new_n33961__, new_new_n33962__,
    new_new_n33963__, new_new_n33964__, new_new_n33965__, new_new_n33966__,
    new_new_n33967__, new_new_n33968__, new_new_n33969__, new_new_n33970__,
    new_new_n33971__, new_new_n33972__, new_new_n33973__, new_new_n33974__,
    new_new_n33975__, new_new_n33976__, new_new_n33977__, new_new_n33978__,
    new_new_n33979__, new_new_n33980__, new_new_n33981__, new_new_n33982__,
    new_new_n33983__, new_new_n33984__, new_new_n33985__, new_new_n33986__,
    new_new_n33987__, new_new_n33988__, new_new_n33989__, new_new_n33990__,
    new_new_n33991__, new_new_n33992__, new_new_n33993__, new_new_n33994__,
    new_new_n33995__, new_new_n33996__, new_new_n33997__, new_new_n33998__,
    new_new_n33999__, new_new_n34000__, new_new_n34001__, new_new_n34002__,
    new_new_n34003__, new_new_n34004__, new_new_n34005__, new_new_n34006__,
    new_new_n34007__, new_new_n34008__, new_new_n34009__, new_new_n34010__,
    new_new_n34011__, new_new_n34012__, new_new_n34013__, new_new_n34014__,
    new_new_n34015__, new_new_n34016__, new_new_n34017__, new_new_n34018__,
    new_new_n34019__, new_new_n34020__, new_new_n34021__, new_new_n34022__,
    new_new_n34023__, new_new_n34024__, new_new_n34025__, new_new_n34026__,
    new_new_n34027__, new_new_n34028__, new_new_n34029__, new_new_n34030__,
    new_new_n34031__, new_new_n34032__, new_new_n34033__, new_new_n34034__,
    new_new_n34035__, new_new_n34036__, new_new_n34037__, new_new_n34038__,
    new_new_n34039__, new_new_n34040__, new_new_n34041__, new_new_n34042__,
    new_new_n34043__, new_new_n34044__, new_new_n34045__, new_new_n34046__,
    new_new_n34047__, new_new_n34048__, new_new_n34049__, new_new_n34050__,
    new_new_n34051__, new_new_n34052__, new_new_n34053__, new_new_n34054__,
    new_new_n34055__, new_new_n34056__, new_new_n34057__, new_new_n34058__,
    new_new_n34059__, new_new_n34060__, new_new_n34061__, new_new_n34062__,
    new_new_n34063__, new_new_n34064__, new_new_n34065__, new_new_n34066__,
    new_new_n34067__, new_new_n34068__, new_new_n34069__, new_new_n34070__,
    new_new_n34071__, new_new_n34072__, new_new_n34073__, new_new_n34074__,
    new_new_n34075__, new_new_n34076__, new_new_n34077__, new_new_n34078__,
    new_new_n34079__, new_new_n34080__, new_new_n34081__, new_new_n34082__,
    new_new_n34083__, new_new_n34084__, new_new_n34085__, new_new_n34086__,
    new_new_n34087__, new_new_n34088__, new_new_n34089__, new_new_n34090__,
    new_new_n34091__, new_new_n34092__, new_new_n34093__, new_new_n34094__,
    new_new_n34095__, new_new_n34096__, new_new_n34097__, new_new_n34098__,
    new_new_n34099__, new_new_n34100__, new_new_n34101__, new_new_n34102__,
    new_new_n34103__, new_new_n34104__, new_new_n34105__, new_new_n34106__,
    new_new_n34107__, new_new_n34108__, new_new_n34109__, new_new_n34110__,
    new_new_n34111__, new_new_n34112__, new_new_n34113__, new_new_n34114__,
    new_new_n34115__, new_new_n34116__, new_new_n34117__, new_new_n34118__,
    new_new_n34119__, new_new_n34120__, new_new_n34121__, new_new_n34122__,
    new_new_n34123__, new_new_n34124__, new_new_n34125__, new_new_n34126__,
    new_new_n34127__, new_new_n34128__, new_new_n34129__, new_new_n34130__,
    new_new_n34131__, new_new_n34132__, new_new_n34133__, new_new_n34134__,
    new_new_n34135__, new_new_n34136__, new_new_n34137__, new_new_n34138__,
    new_new_n34139__, new_new_n34140__, new_new_n34141__, new_new_n34142__,
    new_new_n34143__, new_new_n34145__, new_new_n34146__, new_new_n34147__,
    new_new_n34148__, new_new_n34149__, new_new_n34150__, new_new_n34151__,
    new_new_n34152__, new_new_n34153__, new_new_n34154__, new_new_n34155__,
    new_new_n34156__, new_new_n34157__, new_new_n34158__, new_new_n34159__,
    new_new_n34160__, new_new_n34161__, new_new_n34162__, new_new_n34163__,
    new_new_n34164__, new_new_n34165__, new_new_n34166__, new_new_n34167__,
    new_new_n34168__, new_new_n34169__, new_new_n34170__, new_new_n34171__,
    new_new_n34172__, new_new_n34173__, new_new_n34174__, new_new_n34175__,
    new_new_n34176__, new_new_n34177__, new_new_n34178__, new_new_n34179__,
    new_new_n34180__, new_new_n34181__, new_new_n34182__, new_new_n34183__,
    new_new_n34184__, new_new_n34185__, new_new_n34186__, new_new_n34187__,
    new_new_n34188__, new_new_n34189__, new_new_n34190__, new_new_n34191__,
    new_new_n34192__, new_new_n34193__, new_new_n34194__, new_new_n34195__,
    new_new_n34196__, new_new_n34197__, new_new_n34198__, new_new_n34199__,
    new_new_n34200__, new_new_n34201__, new_new_n34202__, new_new_n34203__,
    new_new_n34204__, new_new_n34205__, new_new_n34206__, new_new_n34207__,
    new_new_n34208__, new_new_n34209__, new_new_n34210__, new_new_n34211__,
    new_new_n34212__, new_new_n34213__, new_new_n34214__, new_new_n34215__,
    new_new_n34216__, new_new_n34217__, new_new_n34218__, new_new_n34219__,
    new_new_n34220__, new_new_n34221__, new_new_n34222__, new_new_n34223__,
    new_new_n34224__, new_new_n34225__, new_new_n34226__, new_new_n34227__,
    new_new_n34228__, new_new_n34229__, new_new_n34230__, new_new_n34231__,
    new_new_n34232__, new_new_n34233__, new_new_n34234__, new_new_n34235__,
    new_new_n34236__, new_new_n34237__, new_new_n34238__, new_new_n34239__,
    new_new_n34240__, new_new_n34241__, new_new_n34242__, new_new_n34243__,
    new_new_n34244__, new_new_n34245__, new_new_n34246__, new_new_n34247__,
    new_new_n34248__, new_new_n34249__, new_new_n34250__, new_new_n34251__,
    new_new_n34252__, new_new_n34253__, new_new_n34254__, new_new_n34255__,
    new_new_n34256__, new_new_n34257__, new_new_n34258__, new_new_n34259__,
    new_new_n34260__, new_new_n34261__, new_new_n34262__, new_new_n34263__,
    new_new_n34264__, new_new_n34265__, new_new_n34266__, new_new_n34267__,
    new_new_n34268__, new_new_n34269__, new_new_n34270__, new_new_n34271__,
    new_new_n34272__, new_new_n34273__, new_new_n34274__, new_new_n34275__,
    new_new_n34276__, new_new_n34277__, new_new_n34278__, new_new_n34279__,
    new_new_n34280__, new_new_n34281__, new_new_n34282__, new_new_n34283__,
    new_new_n34284__, new_new_n34285__, new_new_n34286__, new_new_n34287__,
    new_new_n34288__, new_new_n34289__, new_new_n34290__, new_new_n34291__,
    new_new_n34292__, new_new_n34293__, new_new_n34294__, new_new_n34295__,
    new_new_n34296__, new_new_n34297__, new_new_n34298__, new_new_n34299__,
    new_new_n34300__, new_new_n34301__, new_new_n34302__, new_new_n34303__,
    new_new_n34304__, new_new_n34305__, new_new_n34306__, new_new_n34307__,
    new_new_n34308__, new_new_n34309__, new_new_n34310__, new_new_n34311__,
    new_new_n34312__, new_new_n34313__, new_new_n34314__, new_new_n34315__,
    new_new_n34316__, new_new_n34317__, new_new_n34318__, new_new_n34319__,
    new_new_n34320__, new_new_n34321__, new_new_n34322__, new_new_n34323__,
    new_new_n34324__, new_new_n34325__, new_new_n34326__, new_new_n34327__,
    new_new_n34328__, new_new_n34329__, new_new_n34330__, new_new_n34331__,
    new_new_n34332__, new_new_n34333__, new_new_n34334__, new_new_n34335__,
    new_new_n34336__, new_new_n34337__, new_new_n34338__, new_new_n34339__,
    new_new_n34340__, new_new_n34341__, new_new_n34342__, new_new_n34343__,
    new_new_n34344__, new_new_n34345__, new_new_n34346__, new_new_n34347__,
    new_new_n34348__, new_new_n34349__, new_new_n34350__, new_new_n34351__,
    new_new_n34352__, new_new_n34353__, new_new_n34354__, new_new_n34355__,
    new_new_n34356__, new_new_n34357__, new_new_n34358__, new_new_n34359__,
    new_new_n34360__, new_new_n34361__, new_new_n34362__, new_new_n34363__,
    new_new_n34364__, new_new_n34365__, new_new_n34366__, new_new_n34367__,
    new_new_n34368__, new_new_n34369__, new_new_n34370__, new_new_n34371__,
    new_new_n34372__, new_new_n34373__, new_new_n34374__, new_new_n34375__,
    new_new_n34376__, new_new_n34377__, new_new_n34378__, new_new_n34379__,
    new_new_n34380__, new_new_n34381__, new_new_n34382__, new_new_n34383__,
    new_new_n34384__, new_new_n34385__, new_new_n34386__, new_new_n34387__,
    new_new_n34388__, new_new_n34389__, new_new_n34390__, new_new_n34391__,
    new_new_n34392__, new_new_n34393__, new_new_n34394__, new_new_n34395__,
    new_new_n34396__, new_new_n34397__, new_new_n34398__, new_new_n34399__,
    new_new_n34400__, new_new_n34401__, new_new_n34402__, new_new_n34403__,
    new_new_n34404__, new_new_n34405__, new_new_n34406__, new_new_n34407__,
    new_new_n34408__, new_new_n34409__, new_new_n34410__, new_new_n34411__,
    new_new_n34412__, new_new_n34413__, new_new_n34414__, new_new_n34415__,
    new_new_n34416__, new_new_n34417__, new_new_n34418__, new_new_n34419__,
    new_new_n34420__, new_new_n34421__, new_new_n34422__, new_new_n34423__,
    new_new_n34424__, new_new_n34425__, new_new_n34426__, new_new_n34427__,
    new_new_n34428__, new_new_n34429__, new_new_n34430__, new_new_n34431__,
    new_new_n34432__, new_new_n34433__, new_new_n34434__, new_new_n34435__,
    new_new_n34436__, new_new_n34437__, new_new_n34438__, new_new_n34439__,
    new_new_n34440__, new_new_n34441__, new_new_n34442__, new_new_n34443__,
    new_new_n34444__, new_new_n34445__, new_new_n34446__, new_new_n34447__,
    new_new_n34448__, new_new_n34449__, new_new_n34450__, new_new_n34451__,
    new_new_n34452__, new_new_n34453__, new_new_n34454__, new_new_n34456__,
    new_new_n34457__, new_new_n34458__, new_new_n34459__, new_new_n34460__,
    new_new_n34461__, new_new_n34462__, new_new_n34463__, new_new_n34464__,
    new_new_n34465__, new_new_n34466__, new_new_n34467__, new_new_n34468__,
    new_new_n34469__, new_new_n34470__, new_new_n34471__, new_new_n34472__,
    new_new_n34473__, new_new_n34474__, new_new_n34475__, new_new_n34476__,
    new_new_n34477__, new_new_n34478__, new_new_n34479__, new_new_n34480__,
    new_new_n34481__, new_new_n34482__, new_new_n34483__, new_new_n34484__,
    new_new_n34485__, new_new_n34486__, new_new_n34487__, new_new_n34488__,
    new_new_n34489__, new_new_n34490__, new_new_n34491__, new_new_n34492__,
    new_new_n34493__, new_new_n34494__, new_new_n34495__, new_new_n34496__,
    new_new_n34497__, new_new_n34498__, new_new_n34499__, new_new_n34500__,
    new_new_n34501__, new_new_n34502__, new_new_n34503__, new_new_n34504__,
    new_new_n34505__, new_new_n34506__, new_new_n34507__, new_new_n34508__,
    new_new_n34509__, new_new_n34510__, new_new_n34511__, new_new_n34512__,
    new_new_n34513__, new_new_n34514__, new_new_n34515__, new_new_n34516__,
    new_new_n34517__, new_new_n34518__, new_new_n34519__, new_new_n34520__,
    new_new_n34521__, new_new_n34522__, new_new_n34523__, new_new_n34524__,
    new_new_n34525__, new_new_n34526__, new_new_n34527__, new_new_n34528__,
    new_new_n34529__, new_new_n34530__, new_new_n34531__, new_new_n34532__,
    new_new_n34533__, new_new_n34534__, new_new_n34535__, new_new_n34536__,
    new_new_n34537__, new_new_n34538__, new_new_n34539__, new_new_n34540__,
    new_new_n34541__, new_new_n34542__, new_new_n34543__, new_new_n34544__,
    new_new_n34545__, new_new_n34546__, new_new_n34547__, new_new_n34548__,
    new_new_n34549__, new_new_n34550__, new_new_n34551__, new_new_n34552__,
    new_new_n34553__, new_new_n34554__, new_new_n34555__, new_new_n34556__,
    new_new_n34557__, new_new_n34558__, new_new_n34559__, new_new_n34560__,
    new_new_n34561__, new_new_n34562__, new_new_n34563__, new_new_n34564__,
    new_new_n34565__, new_new_n34566__, new_new_n34567__, new_new_n34568__,
    new_new_n34569__, new_new_n34570__, new_new_n34571__, new_new_n34572__,
    new_new_n34573__, new_new_n34574__, new_new_n34575__, new_new_n34576__,
    new_new_n34577__, new_new_n34578__, new_new_n34579__, new_new_n34580__,
    new_new_n34581__, new_new_n34582__, new_new_n34583__, new_new_n34584__,
    new_new_n34585__, new_new_n34586__, new_new_n34587__, new_new_n34588__,
    new_new_n34589__, new_new_n34590__, new_new_n34591__, new_new_n34592__,
    new_new_n34593__, new_new_n34594__, new_new_n34595__, new_new_n34596__,
    new_new_n34597__, new_new_n34598__, new_new_n34599__, new_new_n34600__,
    new_new_n34601__, new_new_n34602__, new_new_n34603__, new_new_n34604__,
    new_new_n34605__, new_new_n34606__, new_new_n34607__, new_new_n34608__,
    new_new_n34609__, new_new_n34610__, new_new_n34611__, new_new_n34612__,
    new_new_n34613__, new_new_n34614__, new_new_n34615__, new_new_n34616__,
    new_new_n34617__, new_new_n34618__, new_new_n34619__, new_new_n34620__,
    new_new_n34621__, new_new_n34622__, new_new_n34623__, new_new_n34624__,
    new_new_n34625__, new_new_n34626__, new_new_n34627__, new_new_n34628__,
    new_new_n34629__, new_new_n34630__, new_new_n34631__, new_new_n34632__,
    new_new_n34633__, new_new_n34634__, new_new_n34635__, new_new_n34636__,
    new_new_n34637__, new_new_n34638__, new_new_n34639__, new_new_n34640__,
    new_new_n34641__, new_new_n34642__, new_new_n34643__, new_new_n34644__,
    new_new_n34645__, new_new_n34646__, new_new_n34647__, new_new_n34648__,
    new_new_n34649__, new_new_n34650__, new_new_n34651__, new_new_n34652__,
    new_new_n34653__, new_new_n34654__, new_new_n34655__, new_new_n34656__,
    new_new_n34657__, new_new_n34658__, new_new_n34659__, new_new_n34660__,
    new_new_n34661__, new_new_n34662__, new_new_n34663__, new_new_n34664__,
    new_new_n34665__, new_new_n34666__, new_new_n34667__, new_new_n34668__,
    new_new_n34669__, new_new_n34670__, new_new_n34671__, new_new_n34672__,
    new_new_n34673__, new_new_n34674__, new_new_n34675__, new_new_n34676__,
    new_new_n34677__, new_new_n34678__, new_new_n34679__, new_new_n34680__,
    new_new_n34681__, new_new_n34682__, new_new_n34683__, new_new_n34684__,
    new_new_n34685__, new_new_n34686__, new_new_n34687__, new_new_n34688__,
    new_new_n34689__, new_new_n34690__, new_new_n34691__, new_new_n34692__,
    new_new_n34693__, new_new_n34694__, new_new_n34695__, new_new_n34696__,
    new_new_n34697__, new_new_n34698__, new_new_n34699__, new_new_n34700__,
    new_new_n34701__, new_new_n34703__, new_new_n34704__, new_new_n34705__,
    new_new_n34706__, new_new_n34707__, new_new_n34708__, new_new_n34709__,
    new_new_n34710__, new_new_n34711__, new_new_n34712__, new_new_n34713__,
    new_new_n34714__, new_new_n34715__, new_new_n34716__, new_new_n34717__,
    new_new_n34718__, new_new_n34719__, new_new_n34720__, new_new_n34721__,
    new_new_n34722__, new_new_n34723__, new_new_n34724__, new_new_n34725__,
    new_new_n34726__, new_new_n34727__, new_new_n34728__, new_new_n34729__,
    new_new_n34730__, new_new_n34731__, new_new_n34732__, new_new_n34733__,
    new_new_n34734__, new_new_n34735__, new_new_n34736__, new_new_n34737__,
    new_new_n34738__, new_new_n34739__, new_new_n34740__, new_new_n34741__,
    new_new_n34742__, new_new_n34743__, new_new_n34744__, new_new_n34745__,
    new_new_n34746__, new_new_n34747__, new_new_n34748__, new_new_n34749__,
    new_new_n34750__, new_new_n34751__, new_new_n34752__, new_new_n34753__,
    new_new_n34754__, new_new_n34755__, new_new_n34756__, new_new_n34757__,
    new_new_n34758__, new_new_n34759__, new_new_n34760__, new_new_n34761__,
    new_new_n34762__, new_new_n34763__, new_new_n34764__, new_new_n34765__,
    new_new_n34766__, new_new_n34767__, new_new_n34768__, new_new_n34769__,
    new_new_n34770__, new_new_n34771__, new_new_n34772__, new_new_n34773__,
    new_new_n34774__, new_new_n34775__, new_new_n34776__, new_new_n34777__,
    new_new_n34778__, new_new_n34779__, new_new_n34780__, new_new_n34781__,
    new_new_n34782__, new_new_n34783__, new_new_n34784__, new_new_n34785__,
    new_new_n34786__, new_new_n34787__, new_new_n34788__, new_new_n34789__,
    new_new_n34790__, new_new_n34791__, new_new_n34792__, new_new_n34793__,
    new_new_n34794__, new_new_n34795__, new_new_n34796__, new_new_n34797__,
    new_new_n34798__, new_new_n34799__, new_new_n34800__, new_new_n34801__,
    new_new_n34802__, new_new_n34803__, new_new_n34804__, new_new_n34805__,
    new_new_n34806__, new_new_n34807__, new_new_n34808__, new_new_n34809__,
    new_new_n34810__, new_new_n34811__, new_new_n34812__, new_new_n34813__,
    new_new_n34814__, new_new_n34815__, new_new_n34816__, new_new_n34817__,
    new_new_n34818__, new_new_n34819__, new_new_n34820__, new_new_n34821__,
    new_new_n34822__, new_new_n34823__, new_new_n34824__, new_new_n34825__,
    new_new_n34826__, new_new_n34827__, new_new_n34828__, new_new_n34829__,
    new_new_n34830__, new_new_n34831__, new_new_n34832__, new_new_n34833__,
    new_new_n34834__, new_new_n34835__, new_new_n34836__, new_new_n34837__,
    new_new_n34838__, new_new_n34839__, new_new_n34840__, new_new_n34841__,
    new_new_n34842__, new_new_n34843__, new_new_n34844__, new_new_n34845__,
    new_new_n34846__, new_new_n34847__, new_new_n34848__, new_new_n34849__,
    new_new_n34850__, new_new_n34851__, new_new_n34852__, new_new_n34853__,
    new_new_n34854__, new_new_n34855__, new_new_n34856__, new_new_n34857__,
    new_new_n34858__, new_new_n34859__, new_new_n34860__, new_new_n34861__,
    new_new_n34862__, new_new_n34863__, new_new_n34864__, new_new_n34865__,
    new_new_n34866__, new_new_n34867__, new_new_n34868__, new_new_n34869__,
    new_new_n34870__, new_new_n34871__, new_new_n34872__, new_new_n34873__,
    new_new_n34874__, new_new_n34875__, new_new_n34876__, new_new_n34877__,
    new_new_n34878__, new_new_n34879__, new_new_n34880__, new_new_n34881__,
    new_new_n34882__, new_new_n34883__, new_new_n34884__, new_new_n34885__,
    new_new_n34886__, new_new_n34887__, new_new_n34888__, new_new_n34889__,
    new_new_n34890__, new_new_n34891__, new_new_n34892__, new_new_n34893__,
    new_new_n34894__, new_new_n34895__, new_new_n34896__, new_new_n34897__,
    new_new_n34898__, new_new_n34899__, new_new_n34900__, new_new_n34901__,
    new_new_n34902__, new_new_n34903__, new_new_n34904__, new_new_n34905__,
    new_new_n34906__, new_new_n34907__, new_new_n34908__, new_new_n34909__,
    new_new_n34910__, new_new_n34911__, new_new_n34912__, new_new_n34913__,
    new_new_n34914__, new_new_n34915__, new_new_n34916__, new_new_n34917__,
    new_new_n34918__, new_new_n34919__, new_new_n34920__, new_new_n34921__,
    new_new_n34922__, new_new_n34923__, new_new_n34924__, new_new_n34925__,
    new_new_n34926__, new_new_n34927__, new_new_n34929__, new_new_n34930__,
    new_new_n34931__, new_new_n34932__, new_new_n34933__, new_new_n34934__,
    new_new_n34935__, new_new_n34936__, new_new_n34937__, new_new_n34938__,
    new_new_n34939__, new_new_n34940__, new_new_n34941__, new_new_n34942__,
    new_new_n34943__, new_new_n34944__, new_new_n34945__, new_new_n34946__,
    new_new_n34947__, new_new_n34948__, new_new_n34949__, new_new_n34950__,
    new_new_n34951__, new_new_n34952__, new_new_n34953__, new_new_n34954__,
    new_new_n34955__, new_new_n34956__, new_new_n34957__, new_new_n34958__,
    new_new_n34959__, new_new_n34960__, new_new_n34961__, new_new_n34962__,
    new_new_n34963__, new_new_n34964__, new_new_n34965__, new_new_n34966__,
    new_new_n34967__, new_new_n34968__, new_new_n34969__, new_new_n34970__,
    new_new_n34971__, new_new_n34972__, new_new_n34973__, new_new_n34974__,
    new_new_n34975__, new_new_n34976__, new_new_n34977__, new_new_n34978__,
    new_new_n34979__, new_new_n34980__, new_new_n34981__, new_new_n34982__,
    new_new_n34983__, new_new_n34984__, new_new_n34985__, new_new_n34986__,
    new_new_n34987__, new_new_n34988__, new_new_n34989__, new_new_n34990__,
    new_new_n34991__, new_new_n34992__, new_new_n34993__, new_new_n34994__,
    new_new_n34995__, new_new_n34996__, new_new_n34997__, new_new_n34998__,
    new_new_n34999__, new_new_n35000__, new_new_n35001__, new_new_n35002__,
    new_new_n35003__, new_new_n35004__, new_new_n35005__, new_new_n35006__,
    new_new_n35007__, new_new_n35008__, new_new_n35009__, new_new_n35010__,
    new_new_n35011__, new_new_n35012__, new_new_n35013__, new_new_n35014__,
    new_new_n35015__, new_new_n35016__, new_new_n35017__, new_new_n35018__,
    new_new_n35019__, new_new_n35020__, new_new_n35021__, new_new_n35022__,
    new_new_n35023__, new_new_n35024__, new_new_n35025__, new_new_n35026__,
    new_new_n35027__, new_new_n35028__, new_new_n35029__, new_new_n35030__,
    new_new_n35031__, new_new_n35032__, new_new_n35033__, new_new_n35034__,
    new_new_n35035__, new_new_n35036__, new_new_n35037__, new_new_n35038__,
    new_new_n35039__, new_new_n35040__, new_new_n35041__, new_new_n35042__,
    new_new_n35043__, new_new_n35044__, new_new_n35045__, new_new_n35046__,
    new_new_n35047__, new_new_n35048__, new_new_n35049__, new_new_n35050__,
    new_new_n35051__, new_new_n35052__, new_new_n35053__, new_new_n35054__,
    new_new_n35055__, new_new_n35056__, new_new_n35057__, new_new_n35058__,
    new_new_n35059__, new_new_n35060__, new_new_n35061__, new_new_n35062__,
    new_new_n35063__, new_new_n35064__, new_new_n35065__, new_new_n35066__,
    new_new_n35067__, new_new_n35068__, new_new_n35069__, new_new_n35070__,
    new_new_n35071__, new_new_n35072__, new_new_n35073__, new_new_n35074__,
    new_new_n35075__, new_new_n35076__, new_new_n35077__, new_new_n35078__,
    new_new_n35079__, new_new_n35080__, new_new_n35081__, new_new_n35082__,
    new_new_n35083__, new_new_n35084__, new_new_n35085__, new_new_n35086__,
    new_new_n35087__, new_new_n35088__, new_new_n35089__, new_new_n35090__,
    new_new_n35091__, new_new_n35092__, new_new_n35093__, new_new_n35094__,
    new_new_n35095__, new_new_n35096__, new_new_n35097__, new_new_n35098__,
    new_new_n35099__, new_new_n35100__, new_new_n35101__, new_new_n35102__,
    new_new_n35103__, new_new_n35104__, new_new_n35105__, new_new_n35106__,
    new_new_n35107__, new_new_n35108__, new_new_n35109__, new_new_n35110__,
    new_new_n35111__, new_new_n35112__, new_new_n35113__, new_new_n35114__,
    new_new_n35115__, new_new_n35116__, new_new_n35117__, new_new_n35118__,
    new_new_n35119__, new_new_n35120__, new_new_n35121__, new_new_n35122__,
    new_new_n35123__, new_new_n35124__, new_new_n35125__, new_new_n35126__,
    new_new_n35127__, new_new_n35128__, new_new_n35129__, new_new_n35130__,
    new_new_n35131__, new_new_n35132__, new_new_n35133__, new_new_n35134__,
    new_new_n35135__, new_new_n35136__, new_new_n35137__, new_new_n35138__,
    new_new_n35139__, new_new_n35140__, new_new_n35141__, new_new_n35142__,
    new_new_n35143__, new_new_n35144__, new_new_n35145__, new_new_n35146__,
    new_new_n35147__, new_new_n35148__, new_new_n35149__, new_new_n35150__,
    new_new_n35151__, new_new_n35152__, new_new_n35153__, new_new_n35154__,
    new_new_n35155__, new_new_n35156__, new_new_n35157__, new_new_n35158__,
    new_new_n35159__, new_new_n35160__, new_new_n35161__, new_new_n35162__,
    new_new_n35164__, new_new_n35165__, new_new_n35166__, new_new_n35167__,
    new_new_n35168__, new_new_n35169__, new_new_n35170__, new_new_n35171__,
    new_new_n35172__, new_new_n35173__, new_new_n35174__, new_new_n35175__,
    new_new_n35176__, new_new_n35177__, new_new_n35178__, new_new_n35179__,
    new_new_n35180__, new_new_n35181__, new_new_n35182__, new_new_n35183__,
    new_new_n35184__, new_new_n35185__, new_new_n35186__, new_new_n35187__,
    new_new_n35188__, new_new_n35189__, new_new_n35190__, new_new_n35191__,
    new_new_n35192__, new_new_n35193__, new_new_n35194__, new_new_n35195__,
    new_new_n35196__, new_new_n35197__, new_new_n35198__, new_new_n35199__,
    new_new_n35200__, new_new_n35201__, new_new_n35202__, new_new_n35203__,
    new_new_n35204__, new_new_n35205__, new_new_n35206__, new_new_n35207__,
    new_new_n35208__, new_new_n35209__, new_new_n35210__, new_new_n35211__,
    new_new_n35212__, new_new_n35213__, new_new_n35214__, new_new_n35215__,
    new_new_n35216__, new_new_n35217__, new_new_n35218__, new_new_n35219__,
    new_new_n35220__, new_new_n35221__, new_new_n35222__, new_new_n35223__,
    new_new_n35224__, new_new_n35225__, new_new_n35226__, new_new_n35227__,
    new_new_n35228__, new_new_n35229__, new_new_n35230__, new_new_n35231__,
    new_new_n35232__, new_new_n35233__, new_new_n35234__, new_new_n35235__,
    new_new_n35236__, new_new_n35237__, new_new_n35238__, new_new_n35239__,
    new_new_n35240__, new_new_n35241__, new_new_n35242__, new_new_n35243__,
    new_new_n35244__, new_new_n35245__, new_new_n35246__, new_new_n35247__,
    new_new_n35248__, new_new_n35249__, new_new_n35250__, new_new_n35251__,
    new_new_n35252__, new_new_n35253__, new_new_n35254__, new_new_n35255__,
    new_new_n35256__, new_new_n35257__, new_new_n35258__, new_new_n35259__,
    new_new_n35260__, new_new_n35261__, new_new_n35262__, new_new_n35263__,
    new_new_n35264__, new_new_n35265__, new_new_n35266__, new_new_n35267__,
    new_new_n35268__, new_new_n35269__, new_new_n35270__, new_new_n35271__,
    new_new_n35272__, new_new_n35273__, new_new_n35274__, new_new_n35275__,
    new_new_n35276__, new_new_n35277__, new_new_n35278__, new_new_n35279__,
    new_new_n35280__, new_new_n35281__, new_new_n35282__, new_new_n35283__,
    new_new_n35284__, new_new_n35285__, new_new_n35286__, new_new_n35287__,
    new_new_n35288__, new_new_n35289__, new_new_n35290__, new_new_n35291__,
    new_new_n35292__, new_new_n35293__, new_new_n35294__, new_new_n35295__,
    new_new_n35296__, new_new_n35297__, new_new_n35298__, new_new_n35299__,
    new_new_n35300__, new_new_n35301__, new_new_n35302__, new_new_n35303__,
    new_new_n35304__, new_new_n35305__, new_new_n35306__, new_new_n35307__,
    new_new_n35308__, new_new_n35309__, new_new_n35310__, new_new_n35311__,
    new_new_n35312__, new_new_n35313__, new_new_n35314__, new_new_n35315__,
    new_new_n35316__, new_new_n35317__, new_new_n35318__, new_new_n35319__,
    new_new_n35320__, new_new_n35321__, new_new_n35322__, new_new_n35323__,
    new_new_n35324__, new_new_n35325__, new_new_n35326__, new_new_n35327__,
    new_new_n35328__, new_new_n35329__, new_new_n35330__, new_new_n35331__,
    new_new_n35332__, new_new_n35333__, new_new_n35334__, new_new_n35335__,
    new_new_n35336__, new_new_n35337__, new_new_n35338__, new_new_n35339__,
    new_new_n35340__, new_new_n35341__, new_new_n35342__, new_new_n35343__,
    new_new_n35344__, new_new_n35345__, new_new_n35346__, new_new_n35347__,
    new_new_n35348__, new_new_n35349__, new_new_n35350__, new_new_n35351__,
    new_new_n35352__, new_new_n35353__, new_new_n35354__, new_new_n35355__,
    new_new_n35356__, new_new_n35357__, new_new_n35358__, new_new_n35359__,
    new_new_n35360__, new_new_n35361__, new_new_n35362__, new_new_n35363__,
    new_new_n35364__, new_new_n35365__, new_new_n35366__, new_new_n35367__,
    new_new_n35368__, new_new_n35369__, new_new_n35370__, new_new_n35371__,
    new_new_n35372__, new_new_n35373__, new_new_n35374__, new_new_n35375__,
    new_new_n35376__, new_new_n35377__, new_new_n35378__, new_new_n35379__,
    new_new_n35380__, new_new_n35381__, new_new_n35382__, new_new_n35383__,
    new_new_n35384__, new_new_n35385__, new_new_n35386__, new_new_n35387__,
    new_new_n35388__, new_new_n35389__, new_new_n35390__, new_new_n35391__,
    new_new_n35392__, new_new_n35393__, new_new_n35394__, new_new_n35395__,
    new_new_n35396__, new_new_n35397__, new_new_n35398__, new_new_n35399__,
    new_new_n35400__, new_new_n35401__, new_new_n35402__, new_new_n35403__,
    new_new_n35404__, new_new_n35405__, new_new_n35406__, new_new_n35407__,
    new_new_n35408__, new_new_n35409__, new_new_n35410__, new_new_n35411__,
    new_new_n35412__, new_new_n35413__, new_new_n35414__, new_new_n35415__,
    new_new_n35416__, new_new_n35417__, new_new_n35418__, new_new_n35419__,
    new_new_n35420__, new_new_n35421__, new_new_n35422__, new_new_n35423__,
    new_new_n35425__, new_new_n35426__, new_new_n35427__, new_new_n35428__,
    new_new_n35429__, new_new_n35430__, new_new_n35431__, new_new_n35432__,
    new_new_n35433__, new_new_n35434__, new_new_n35435__, new_new_n35436__,
    new_new_n35437__, new_new_n35438__, new_new_n35439__, new_new_n35440__,
    new_new_n35441__, new_new_n35442__, new_new_n35443__, new_new_n35444__,
    new_new_n35445__, new_new_n35446__, new_new_n35447__, new_new_n35448__,
    new_new_n35449__, new_new_n35450__, new_new_n35451__, new_new_n35452__,
    new_new_n35453__, new_new_n35454__, new_new_n35455__, new_new_n35456__,
    new_new_n35457__, new_new_n35458__, new_new_n35459__, new_new_n35460__,
    new_new_n35461__, new_new_n35462__, new_new_n35463__, new_new_n35464__,
    new_new_n35465__, new_new_n35466__, new_new_n35467__, new_new_n35468__,
    new_new_n35469__, new_new_n35470__, new_new_n35471__, new_new_n35472__,
    new_new_n35473__, new_new_n35474__, new_new_n35475__, new_new_n35476__,
    new_new_n35477__, new_new_n35478__, new_new_n35479__, new_new_n35480__,
    new_new_n35481__, new_new_n35482__, new_new_n35483__, new_new_n35484__,
    new_new_n35485__, new_new_n35486__, new_new_n35487__, new_new_n35488__,
    new_new_n35489__, new_new_n35490__, new_new_n35491__, new_new_n35492__,
    new_new_n35493__, new_new_n35494__, new_new_n35495__, new_new_n35496__,
    new_new_n35497__, new_new_n35498__, new_new_n35499__, new_new_n35500__,
    new_new_n35501__, new_new_n35502__, new_new_n35503__, new_new_n35504__,
    new_new_n35505__, new_new_n35506__, new_new_n35507__, new_new_n35508__,
    new_new_n35509__, new_new_n35510__, new_new_n35511__, new_new_n35512__,
    new_new_n35513__, new_new_n35514__, new_new_n35515__, new_new_n35516__,
    new_new_n35517__, new_new_n35518__, new_new_n35519__, new_new_n35520__,
    new_new_n35521__, new_new_n35522__, new_new_n35523__, new_new_n35524__,
    new_new_n35525__, new_new_n35526__, new_new_n35527__, new_new_n35528__,
    new_new_n35529__, new_new_n35530__, new_new_n35531__, new_new_n35532__,
    new_new_n35533__, new_new_n35534__, new_new_n35535__, new_new_n35536__,
    new_new_n35537__, new_new_n35538__, new_new_n35539__, new_new_n35540__,
    new_new_n35541__, new_new_n35542__, new_new_n35543__, new_new_n35544__,
    new_new_n35545__, new_new_n35546__, new_new_n35547__, new_new_n35548__,
    new_new_n35549__, new_new_n35550__, new_new_n35551__, new_new_n35552__,
    new_new_n35553__, new_new_n35554__, new_new_n35555__, new_new_n35556__,
    new_new_n35557__, new_new_n35558__, new_new_n35559__, new_new_n35560__,
    new_new_n35561__, new_new_n35562__, new_new_n35563__, new_new_n35564__,
    new_new_n35565__, new_new_n35566__, new_new_n35567__, new_new_n35568__,
    new_new_n35569__, new_new_n35570__, new_new_n35571__, new_new_n35572__,
    new_new_n35573__, new_new_n35574__, new_new_n35575__, new_new_n35576__,
    new_new_n35577__, new_new_n35578__, new_new_n35579__, new_new_n35580__,
    new_new_n35581__, new_new_n35582__, new_new_n35583__, new_new_n35584__,
    new_new_n35585__, new_new_n35586__, new_new_n35587__, new_new_n35588__,
    new_new_n35589__, new_new_n35590__, new_new_n35591__, new_new_n35592__,
    new_new_n35593__, new_new_n35594__, new_new_n35595__, new_new_n35596__,
    new_new_n35597__, new_new_n35598__, new_new_n35599__, new_new_n35600__,
    new_new_n35601__, new_new_n35602__, new_new_n35603__, new_new_n35604__,
    new_new_n35605__, new_new_n35606__, new_new_n35607__, new_new_n35608__,
    new_new_n35609__, new_new_n35610__, new_new_n35611__, new_new_n35612__,
    new_new_n35613__, new_new_n35614__, new_new_n35615__, new_new_n35616__,
    new_new_n35617__, new_new_n35618__, new_new_n35619__, new_new_n35620__,
    new_new_n35621__, new_new_n35622__, new_new_n35623__, new_new_n35624__,
    new_new_n35625__, new_new_n35626__, new_new_n35627__, new_new_n35628__,
    new_new_n35629__, new_new_n35630__, new_new_n35631__, new_new_n35632__,
    new_new_n35633__, new_new_n35634__, new_new_n35635__, new_new_n35636__,
    new_new_n35637__, new_new_n35638__, new_new_n35639__, new_new_n35640__,
    new_new_n35641__, new_new_n35642__, new_new_n35643__, new_new_n35644__,
    new_new_n35645__, new_new_n35646__, new_new_n35647__, new_new_n35648__,
    new_new_n35649__, new_new_n35650__, new_new_n35651__, new_new_n35652__,
    new_new_n35653__, new_new_n35654__, new_new_n35655__, new_new_n35656__,
    new_new_n35657__, new_new_n35658__, new_new_n35659__, new_new_n35660__,
    new_new_n35661__, new_new_n35663__, new_new_n35664__, new_new_n35665__,
    new_new_n35666__, new_new_n35667__, new_new_n35668__, new_new_n35669__,
    new_new_n35670__, new_new_n35671__, new_new_n35672__, new_new_n35673__,
    new_new_n35674__, new_new_n35675__, new_new_n35676__, new_new_n35677__,
    new_new_n35678__, new_new_n35679__, new_new_n35680__, new_new_n35681__,
    new_new_n35682__, new_new_n35683__, new_new_n35684__, new_new_n35685__,
    new_new_n35686__, new_new_n35687__, new_new_n35688__, new_new_n35689__,
    new_new_n35690__, new_new_n35691__, new_new_n35692__, new_new_n35693__,
    new_new_n35694__, new_new_n35695__, new_new_n35696__, new_new_n35697__,
    new_new_n35698__, new_new_n35699__, new_new_n35700__, new_new_n35701__,
    new_new_n35702__, new_new_n35703__, new_new_n35704__, new_new_n35705__,
    new_new_n35706__, new_new_n35707__, new_new_n35708__, new_new_n35709__,
    new_new_n35710__, new_new_n35711__, new_new_n35712__, new_new_n35713__,
    new_new_n35714__, new_new_n35715__, new_new_n35716__, new_new_n35717__,
    new_new_n35718__, new_new_n35719__, new_new_n35720__, new_new_n35721__,
    new_new_n35722__, new_new_n35723__, new_new_n35724__, new_new_n35725__,
    new_new_n35726__, new_new_n35727__, new_new_n35728__, new_new_n35729__,
    new_new_n35730__, new_new_n35731__, new_new_n35732__, new_new_n35733__,
    new_new_n35734__, new_new_n35735__, new_new_n35736__, new_new_n35737__,
    new_new_n35738__, new_new_n35739__, new_new_n35740__, new_new_n35741__,
    new_new_n35742__, new_new_n35743__, new_new_n35744__, new_new_n35745__,
    new_new_n35746__, new_new_n35747__, new_new_n35748__, new_new_n35749__,
    new_new_n35750__, new_new_n35751__, new_new_n35752__, new_new_n35753__,
    new_new_n35754__, new_new_n35755__, new_new_n35756__, new_new_n35757__,
    new_new_n35758__, new_new_n35759__, new_new_n35760__, new_new_n35761__,
    new_new_n35762__, new_new_n35763__, new_new_n35764__, new_new_n35765__,
    new_new_n35766__, new_new_n35767__, new_new_n35768__, new_new_n35769__,
    new_new_n35770__, new_new_n35771__, new_new_n35772__, new_new_n35773__,
    new_new_n35774__, new_new_n35775__, new_new_n35776__, new_new_n35777__,
    new_new_n35778__, new_new_n35779__, new_new_n35780__, new_new_n35781__,
    new_new_n35782__, new_new_n35783__, new_new_n35784__, new_new_n35785__,
    new_new_n35786__, new_new_n35787__, new_new_n35788__, new_new_n35789__,
    new_new_n35790__, new_new_n35791__, new_new_n35792__, new_new_n35793__,
    new_new_n35794__, new_new_n35795__, new_new_n35796__, new_new_n35797__,
    new_new_n35798__, new_new_n35799__, new_new_n35800__, new_new_n35801__,
    new_new_n35802__, new_new_n35803__, new_new_n35804__, new_new_n35805__,
    new_new_n35806__, new_new_n35807__, new_new_n35808__, new_new_n35809__,
    new_new_n35810__, new_new_n35811__, new_new_n35812__, new_new_n35813__,
    new_new_n35814__, new_new_n35815__, new_new_n35816__, new_new_n35817__,
    new_new_n35818__, new_new_n35819__, new_new_n35820__, new_new_n35821__,
    new_new_n35822__, new_new_n35823__, new_new_n35824__, new_new_n35825__,
    new_new_n35826__, new_new_n35827__, new_new_n35828__, new_new_n35829__,
    new_new_n35830__, new_new_n35831__, new_new_n35832__, new_new_n35833__,
    new_new_n35834__, new_new_n35835__, new_new_n35836__, new_new_n35837__,
    new_new_n35838__, new_new_n35839__, new_new_n35840__, new_new_n35841__,
    new_new_n35842__, new_new_n35843__, new_new_n35844__, new_new_n35845__,
    new_new_n35846__, new_new_n35847__, new_new_n35848__, new_new_n35849__,
    new_new_n35850__, new_new_n35851__, new_new_n35852__, new_new_n35853__,
    new_new_n35854__, new_new_n35855__, new_new_n35856__, new_new_n35857__,
    new_new_n35858__, new_new_n35859__, new_new_n35860__, new_new_n35861__,
    new_new_n35862__, new_new_n35863__, new_new_n35864__, new_new_n35865__,
    new_new_n35866__, new_new_n35867__, new_new_n35868__, new_new_n35869__,
    new_new_n35870__, new_new_n35871__, new_new_n35872__, new_new_n35873__,
    new_new_n35874__, new_new_n35875__, new_new_n35877__, new_new_n35878__,
    new_new_n35879__, new_new_n35880__, new_new_n35881__, new_new_n35882__,
    new_new_n35883__, new_new_n35884__, new_new_n35885__, new_new_n35886__,
    new_new_n35887__, new_new_n35888__, new_new_n35889__, new_new_n35890__,
    new_new_n35891__, new_new_n35892__, new_new_n35893__, new_new_n35894__,
    new_new_n35895__, new_new_n35896__, new_new_n35897__, new_new_n35898__,
    new_new_n35899__, new_new_n35900__, new_new_n35901__, new_new_n35902__,
    new_new_n35903__, new_new_n35904__, new_new_n35905__, new_new_n35906__,
    new_new_n35907__, new_new_n35908__, new_new_n35909__, new_new_n35910__,
    new_new_n35911__, new_new_n35912__, new_new_n35913__, new_new_n35914__,
    new_new_n35915__, new_new_n35916__, new_new_n35917__, new_new_n35918__,
    new_new_n35919__, new_new_n35920__, new_new_n35921__, new_new_n35922__,
    new_new_n35923__, new_new_n35924__, new_new_n35925__, new_new_n35926__,
    new_new_n35927__, new_new_n35928__, new_new_n35929__, new_new_n35930__,
    new_new_n35931__, new_new_n35932__, new_new_n35933__, new_new_n35934__,
    new_new_n35935__, new_new_n35936__, new_new_n35937__, new_new_n35938__,
    new_new_n35939__, new_new_n35940__, new_new_n35941__, new_new_n35942__,
    new_new_n35943__, new_new_n35944__, new_new_n35945__, new_new_n35946__,
    new_new_n35947__, new_new_n35948__, new_new_n35949__, new_new_n35950__,
    new_new_n35951__, new_new_n35952__, new_new_n35953__, new_new_n35954__,
    new_new_n35955__, new_new_n35956__, new_new_n35957__, new_new_n35958__,
    new_new_n35959__, new_new_n35960__, new_new_n35961__, new_new_n35962__,
    new_new_n35963__, new_new_n35964__, new_new_n35965__, new_new_n35966__,
    new_new_n35967__, new_new_n35968__, new_new_n35969__, new_new_n35970__,
    new_new_n35971__, new_new_n35972__, new_new_n35973__, new_new_n35974__,
    new_new_n35975__, new_new_n35976__, new_new_n35977__, new_new_n35978__,
    new_new_n35979__, new_new_n35980__, new_new_n35981__, new_new_n35982__,
    new_new_n35983__, new_new_n35984__, new_new_n35985__, new_new_n35986__,
    new_new_n35987__, new_new_n35988__, new_new_n35989__, new_new_n35990__,
    new_new_n35991__, new_new_n35992__, new_new_n35993__, new_new_n35994__,
    new_new_n35995__, new_new_n35996__, new_new_n35997__, new_new_n35998__,
    new_new_n35999__, new_new_n36000__, new_new_n36001__, new_new_n36002__,
    new_new_n36003__, new_new_n36004__, new_new_n36005__, new_new_n36006__,
    new_new_n36007__, new_new_n36008__, new_new_n36009__, new_new_n36010__,
    new_new_n36011__, new_new_n36012__, new_new_n36013__, new_new_n36014__,
    new_new_n36015__, new_new_n36016__, new_new_n36017__, new_new_n36018__,
    new_new_n36019__, new_new_n36020__, new_new_n36021__, new_new_n36022__,
    new_new_n36023__, new_new_n36024__, new_new_n36025__, new_new_n36026__,
    new_new_n36027__, new_new_n36028__, new_new_n36029__, new_new_n36030__,
    new_new_n36031__, new_new_n36032__, new_new_n36033__, new_new_n36034__,
    new_new_n36035__, new_new_n36036__, new_new_n36037__, new_new_n36038__,
    new_new_n36039__, new_new_n36040__, new_new_n36041__, new_new_n36042__,
    new_new_n36043__, new_new_n36044__, new_new_n36045__, new_new_n36046__,
    new_new_n36047__, new_new_n36048__, new_new_n36049__, new_new_n36050__,
    new_new_n36051__, new_new_n36052__, new_new_n36053__, new_new_n36054__,
    new_new_n36055__, new_new_n36056__, new_new_n36057__, new_new_n36058__,
    new_new_n36059__, new_new_n36060__, new_new_n36061__, new_new_n36062__,
    new_new_n36063__, new_new_n36064__, new_new_n36065__, new_new_n36066__,
    new_new_n36067__, new_new_n36068__, new_new_n36069__, new_new_n36070__,
    new_new_n36071__, new_new_n36072__, new_new_n36073__, new_new_n36074__,
    new_new_n36075__, new_new_n36076__, new_new_n36077__, new_new_n36078__,
    new_new_n36079__, new_new_n36080__, new_new_n36081__, new_new_n36082__,
    new_new_n36083__, new_new_n36084__, new_new_n36085__, new_new_n36086__,
    new_new_n36087__, new_new_n36088__, new_new_n36089__, new_new_n36090__,
    new_new_n36091__, new_new_n36092__, new_new_n36094__, new_new_n36095__,
    new_new_n36096__, new_new_n36097__, new_new_n36098__, new_new_n36099__,
    new_new_n36100__, new_new_n36101__, new_new_n36102__, new_new_n36103__,
    new_new_n36104__, new_new_n36105__, new_new_n36106__, new_new_n36107__,
    new_new_n36108__, new_new_n36109__, new_new_n36110__, new_new_n36111__,
    new_new_n36112__, new_new_n36113__, new_new_n36114__, new_new_n36115__,
    new_new_n36116__, new_new_n36117__, new_new_n36118__, new_new_n36119__,
    new_new_n36120__, new_new_n36121__, new_new_n36122__, new_new_n36123__,
    new_new_n36124__, new_new_n36125__, new_new_n36126__, new_new_n36127__,
    new_new_n36128__, new_new_n36129__, new_new_n36130__, new_new_n36131__,
    new_new_n36132__, new_new_n36133__, new_new_n36134__, new_new_n36135__,
    new_new_n36136__, new_new_n36137__, new_new_n36138__, new_new_n36139__,
    new_new_n36140__, new_new_n36141__, new_new_n36142__, new_new_n36143__,
    new_new_n36144__, new_new_n36145__, new_new_n36146__, new_new_n36147__,
    new_new_n36148__, new_new_n36149__, new_new_n36150__, new_new_n36151__,
    new_new_n36152__, new_new_n36153__, new_new_n36154__, new_new_n36155__,
    new_new_n36156__, new_new_n36157__, new_new_n36158__, new_new_n36159__,
    new_new_n36160__, new_new_n36161__, new_new_n36162__, new_new_n36163__,
    new_new_n36164__, new_new_n36165__, new_new_n36166__, new_new_n36167__,
    new_new_n36168__, new_new_n36169__, new_new_n36170__, new_new_n36171__,
    new_new_n36172__, new_new_n36173__, new_new_n36174__, new_new_n36175__,
    new_new_n36176__, new_new_n36177__, new_new_n36178__, new_new_n36179__,
    new_new_n36180__, new_new_n36181__, new_new_n36182__, new_new_n36183__,
    new_new_n36184__, new_new_n36185__, new_new_n36186__, new_new_n36187__,
    new_new_n36188__, new_new_n36189__, new_new_n36190__, new_new_n36191__,
    new_new_n36192__, new_new_n36193__, new_new_n36194__, new_new_n36195__,
    new_new_n36196__, new_new_n36197__, new_new_n36198__, new_new_n36199__,
    new_new_n36200__, new_new_n36201__, new_new_n36202__, new_new_n36203__,
    new_new_n36204__, new_new_n36205__, new_new_n36206__, new_new_n36207__,
    new_new_n36208__, new_new_n36209__, new_new_n36210__, new_new_n36211__,
    new_new_n36212__, new_new_n36213__, new_new_n36214__, new_new_n36215__,
    new_new_n36216__, new_new_n36217__, new_new_n36218__, new_new_n36219__,
    new_new_n36220__, new_new_n36221__, new_new_n36222__, new_new_n36223__,
    new_new_n36224__, new_new_n36225__, new_new_n36226__, new_new_n36227__,
    new_new_n36228__, new_new_n36229__, new_new_n36230__, new_new_n36231__,
    new_new_n36232__, new_new_n36233__, new_new_n36234__, new_new_n36235__,
    new_new_n36236__, new_new_n36237__, new_new_n36238__, new_new_n36239__,
    new_new_n36240__, new_new_n36241__, new_new_n36242__, new_new_n36243__,
    new_new_n36244__, new_new_n36245__, new_new_n36246__, new_new_n36247__,
    new_new_n36248__, new_new_n36249__, new_new_n36250__, new_new_n36251__,
    new_new_n36252__, new_new_n36253__, new_new_n36254__, new_new_n36255__,
    new_new_n36256__, new_new_n36257__, new_new_n36258__, new_new_n36259__,
    new_new_n36260__, new_new_n36261__, new_new_n36262__, new_new_n36263__,
    new_new_n36264__, new_new_n36265__, new_new_n36266__, new_new_n36267__,
    new_new_n36268__, new_new_n36269__, new_new_n36270__, new_new_n36271__,
    new_new_n36272__, new_new_n36273__, new_new_n36274__, new_new_n36275__,
    new_new_n36276__, new_new_n36277__, new_new_n36278__, new_new_n36279__,
    new_new_n36280__, new_new_n36281__, new_new_n36282__, new_new_n36283__,
    new_new_n36285__, new_new_n36286__, new_new_n36287__, new_new_n36288__,
    new_new_n36289__, new_new_n36290__, new_new_n36291__, new_new_n36292__,
    new_new_n36293__, new_new_n36294__, new_new_n36295__, new_new_n36296__,
    new_new_n36297__, new_new_n36298__, new_new_n36299__, new_new_n36300__,
    new_new_n36301__, new_new_n36302__, new_new_n36303__, new_new_n36304__,
    new_new_n36305__, new_new_n36306__, new_new_n36307__, new_new_n36308__,
    new_new_n36309__, new_new_n36310__, new_new_n36311__, new_new_n36312__,
    new_new_n36313__, new_new_n36314__, new_new_n36315__, new_new_n36316__,
    new_new_n36317__, new_new_n36318__, new_new_n36319__, new_new_n36320__,
    new_new_n36321__, new_new_n36322__, new_new_n36323__, new_new_n36324__,
    new_new_n36325__, new_new_n36326__, new_new_n36327__, new_new_n36328__,
    new_new_n36329__, new_new_n36330__, new_new_n36331__, new_new_n36332__,
    new_new_n36333__, new_new_n36334__, new_new_n36335__, new_new_n36336__,
    new_new_n36337__, new_new_n36338__, new_new_n36339__, new_new_n36340__,
    new_new_n36341__, new_new_n36342__, new_new_n36343__, new_new_n36344__,
    new_new_n36345__, new_new_n36346__, new_new_n36347__, new_new_n36348__,
    new_new_n36349__, new_new_n36350__, new_new_n36351__, new_new_n36352__,
    new_new_n36353__, new_new_n36354__, new_new_n36355__, new_new_n36356__,
    new_new_n36357__, new_new_n36358__, new_new_n36359__, new_new_n36360__,
    new_new_n36361__, new_new_n36362__, new_new_n36363__, new_new_n36364__,
    new_new_n36365__, new_new_n36366__, new_new_n36367__, new_new_n36368__,
    new_new_n36369__, new_new_n36370__, new_new_n36371__, new_new_n36372__,
    new_new_n36373__, new_new_n36374__, new_new_n36375__, new_new_n36376__,
    new_new_n36377__, new_new_n36378__, new_new_n36379__, new_new_n36380__,
    new_new_n36381__, new_new_n36382__, new_new_n36383__, new_new_n36384__,
    new_new_n36385__, new_new_n36386__, new_new_n36387__, new_new_n36388__,
    new_new_n36389__, new_new_n36390__, new_new_n36391__, new_new_n36392__,
    new_new_n36393__, new_new_n36394__, new_new_n36395__, new_new_n36396__,
    new_new_n36397__, new_new_n36398__, new_new_n36399__, new_new_n36400__,
    new_new_n36401__, new_new_n36402__, new_new_n36403__, new_new_n36404__,
    new_new_n36405__, new_new_n36406__, new_new_n36407__, new_new_n36408__,
    new_new_n36409__, new_new_n36410__, new_new_n36411__, new_new_n36412__,
    new_new_n36413__, new_new_n36414__, new_new_n36415__, new_new_n36416__,
    new_new_n36417__, new_new_n36418__, new_new_n36419__, new_new_n36420__,
    new_new_n36421__, new_new_n36422__, new_new_n36423__, new_new_n36424__,
    new_new_n36425__, new_new_n36426__, new_new_n36427__, new_new_n36428__,
    new_new_n36429__, new_new_n36430__, new_new_n36431__, new_new_n36432__,
    new_new_n36433__, new_new_n36434__, new_new_n36435__, new_new_n36436__,
    new_new_n36437__, new_new_n36438__, new_new_n36439__, new_new_n36440__,
    new_new_n36441__, new_new_n36442__, new_new_n36443__, new_new_n36444__,
    new_new_n36445__, new_new_n36446__, new_new_n36447__, new_new_n36448__,
    new_new_n36449__, new_new_n36450__, new_new_n36451__, new_new_n36452__,
    new_new_n36453__, new_new_n36454__, new_new_n36455__, new_new_n36456__,
    new_new_n36457__, new_new_n36458__, new_new_n36459__, new_new_n36460__,
    new_new_n36461__, new_new_n36462__, new_new_n36463__, new_new_n36464__,
    new_new_n36465__, new_new_n36466__, new_new_n36467__, new_new_n36468__,
    new_new_n36469__, new_new_n36470__, new_new_n36471__, new_new_n36472__,
    new_new_n36473__, new_new_n36474__, new_new_n36475__, new_new_n36476__,
    new_new_n36477__, new_new_n36478__, new_new_n36479__, new_new_n36480__,
    new_new_n36481__, new_new_n36482__, new_new_n36483__, new_new_n36484__,
    new_new_n36485__, new_new_n36486__, new_new_n36487__, new_new_n36488__,
    new_new_n36490__, new_new_n36491__, new_new_n36492__, new_new_n36493__,
    new_new_n36494__, new_new_n36495__, new_new_n36496__, new_new_n36497__,
    new_new_n36498__, new_new_n36499__, new_new_n36500__, new_new_n36501__,
    new_new_n36502__, new_new_n36503__, new_new_n36504__, new_new_n36505__,
    new_new_n36506__, new_new_n36507__, new_new_n36508__, new_new_n36509__,
    new_new_n36510__, new_new_n36511__, new_new_n36512__, new_new_n36513__,
    new_new_n36514__, new_new_n36515__, new_new_n36516__, new_new_n36517__,
    new_new_n36518__, new_new_n36519__, new_new_n36520__, new_new_n36521__,
    new_new_n36522__, new_new_n36523__, new_new_n36524__, new_new_n36525__,
    new_new_n36526__, new_new_n36527__, new_new_n36528__, new_new_n36529__,
    new_new_n36530__, new_new_n36531__, new_new_n36532__, new_new_n36533__,
    new_new_n36534__, new_new_n36535__, new_new_n36536__, new_new_n36537__,
    new_new_n36538__, new_new_n36539__, new_new_n36540__, new_new_n36541__,
    new_new_n36542__, new_new_n36543__, new_new_n36544__, new_new_n36545__,
    new_new_n36546__, new_new_n36547__, new_new_n36548__, new_new_n36549__,
    new_new_n36550__, new_new_n36551__, new_new_n36552__, new_new_n36553__,
    new_new_n36554__, new_new_n36555__, new_new_n36556__, new_new_n36557__,
    new_new_n36558__, new_new_n36559__, new_new_n36560__, new_new_n36561__,
    new_new_n36562__, new_new_n36563__, new_new_n36564__, new_new_n36565__,
    new_new_n36566__, new_new_n36567__, new_new_n36568__, new_new_n36569__,
    new_new_n36570__, new_new_n36571__, new_new_n36572__, new_new_n36573__,
    new_new_n36574__, new_new_n36575__, new_new_n36576__, new_new_n36577__,
    new_new_n36578__, new_new_n36579__, new_new_n36580__, new_new_n36581__,
    new_new_n36582__, new_new_n36583__, new_new_n36584__, new_new_n36585__,
    new_new_n36586__, new_new_n36587__, new_new_n36588__, new_new_n36589__,
    new_new_n36590__, new_new_n36591__, new_new_n36592__, new_new_n36593__,
    new_new_n36594__, new_new_n36595__, new_new_n36596__, new_new_n36597__,
    new_new_n36598__, new_new_n36599__, new_new_n36600__, new_new_n36601__,
    new_new_n36602__, new_new_n36603__, new_new_n36604__, new_new_n36605__,
    new_new_n36606__, new_new_n36607__, new_new_n36608__, new_new_n36609__,
    new_new_n36610__, new_new_n36611__, new_new_n36612__, new_new_n36613__,
    new_new_n36614__, new_new_n36615__, new_new_n36616__, new_new_n36617__,
    new_new_n36618__, new_new_n36619__, new_new_n36620__, new_new_n36621__,
    new_new_n36622__, new_new_n36623__, new_new_n36624__, new_new_n36625__,
    new_new_n36626__, new_new_n36627__, new_new_n36628__, new_new_n36629__,
    new_new_n36630__, new_new_n36631__, new_new_n36632__, new_new_n36633__,
    new_new_n36634__, new_new_n36635__, new_new_n36636__, new_new_n36637__,
    new_new_n36638__, new_new_n36639__, new_new_n36640__, new_new_n36641__,
    new_new_n36642__, new_new_n36643__, new_new_n36644__, new_new_n36645__,
    new_new_n36646__, new_new_n36647__, new_new_n36648__, new_new_n36649__,
    new_new_n36650__, new_new_n36651__, new_new_n36652__, new_new_n36653__,
    new_new_n36654__, new_new_n36655__, new_new_n36656__, new_new_n36657__,
    new_new_n36658__, new_new_n36659__, new_new_n36660__, new_new_n36661__,
    new_new_n36662__, new_new_n36663__, new_new_n36664__, new_new_n36665__,
    new_new_n36666__, new_new_n36667__, new_new_n36668__, new_new_n36669__,
    new_new_n36670__, new_new_n36671__, new_new_n36672__, new_new_n36673__,
    new_new_n36674__, new_new_n36675__, new_new_n36676__, new_new_n36677__,
    new_new_n36678__, new_new_n36679__, new_new_n36680__, new_new_n36682__,
    new_new_n36683__, new_new_n36684__, new_new_n36685__, new_new_n36686__,
    new_new_n36687__, new_new_n36688__, new_new_n36689__, new_new_n36690__,
    new_new_n36691__, new_new_n36692__, new_new_n36693__, new_new_n36694__,
    new_new_n36695__, new_new_n36696__, new_new_n36697__, new_new_n36698__,
    new_new_n36699__, new_new_n36700__, new_new_n36701__, new_new_n36702__,
    new_new_n36703__, new_new_n36704__, new_new_n36705__, new_new_n36706__,
    new_new_n36707__, new_new_n36708__, new_new_n36709__, new_new_n36710__,
    new_new_n36711__, new_new_n36712__, new_new_n36713__, new_new_n36714__,
    new_new_n36715__, new_new_n36716__, new_new_n36717__, new_new_n36718__,
    new_new_n36719__, new_new_n36720__, new_new_n36721__, new_new_n36722__,
    new_new_n36723__, new_new_n36724__, new_new_n36725__, new_new_n36726__,
    new_new_n36727__, new_new_n36728__, new_new_n36729__, new_new_n36730__,
    new_new_n36731__, new_new_n36732__, new_new_n36733__, new_new_n36734__,
    new_new_n36735__, new_new_n36736__, new_new_n36737__, new_new_n36738__,
    new_new_n36739__, new_new_n36740__, new_new_n36741__, new_new_n36742__,
    new_new_n36743__, new_new_n36744__, new_new_n36745__, new_new_n36746__,
    new_new_n36747__, new_new_n36748__, new_new_n36749__, new_new_n36750__,
    new_new_n36751__, new_new_n36752__, new_new_n36753__, new_new_n36754__,
    new_new_n36755__, new_new_n36756__, new_new_n36757__, new_new_n36758__,
    new_new_n36759__, new_new_n36760__, new_new_n36761__, new_new_n36762__,
    new_new_n36763__, new_new_n36764__, new_new_n36765__, new_new_n36766__,
    new_new_n36767__, new_new_n36768__, new_new_n36769__, new_new_n36770__,
    new_new_n36771__, new_new_n36772__, new_new_n36773__, new_new_n36774__,
    new_new_n36775__, new_new_n36776__, new_new_n36777__, new_new_n36778__,
    new_new_n36779__, new_new_n36780__, new_new_n36781__, new_new_n36782__,
    new_new_n36783__, new_new_n36784__, new_new_n36785__, new_new_n36786__,
    new_new_n36787__, new_new_n36788__, new_new_n36789__, new_new_n36790__,
    new_new_n36791__, new_new_n36792__, new_new_n36793__, new_new_n36794__,
    new_new_n36795__, new_new_n36796__, new_new_n36797__, new_new_n36798__,
    new_new_n36799__, new_new_n36800__, new_new_n36801__, new_new_n36802__,
    new_new_n36803__, new_new_n36804__, new_new_n36805__, new_new_n36806__,
    new_new_n36807__, new_new_n36808__, new_new_n36809__, new_new_n36810__,
    new_new_n36811__, new_new_n36812__, new_new_n36813__, new_new_n36814__,
    new_new_n36815__, new_new_n36816__, new_new_n36817__, new_new_n36818__,
    new_new_n36819__, new_new_n36820__, new_new_n36821__, new_new_n36822__,
    new_new_n36823__, new_new_n36824__, new_new_n36825__, new_new_n36826__,
    new_new_n36827__, new_new_n36828__, new_new_n36829__, new_new_n36830__,
    new_new_n36831__, new_new_n36832__, new_new_n36833__, new_new_n36834__,
    new_new_n36835__, new_new_n36836__, new_new_n36837__, new_new_n36838__,
    new_new_n36839__, new_new_n36840__, new_new_n36841__, new_new_n36842__,
    new_new_n36843__, new_new_n36844__, new_new_n36845__, new_new_n36846__,
    new_new_n36847__, new_new_n36848__, new_new_n36849__, new_new_n36850__,
    new_new_n36851__, new_new_n36852__, new_new_n36853__, new_new_n36854__,
    new_new_n36855__, new_new_n36856__, new_new_n36857__, new_new_n36858__,
    new_new_n36859__, new_new_n36860__, new_new_n36861__, new_new_n36862__,
    new_new_n36863__, new_new_n36864__, new_new_n36865__, new_new_n36866__,
    new_new_n36867__, new_new_n36868__, new_new_n36869__, new_new_n36870__,
    new_new_n36871__, new_new_n36872__, new_new_n36873__, new_new_n36874__,
    new_new_n36875__, new_new_n36876__, new_new_n36877__, new_new_n36878__,
    new_new_n36879__, new_new_n36881__, new_new_n36882__, new_new_n36883__,
    new_new_n36884__, new_new_n36885__, new_new_n36886__, new_new_n36887__,
    new_new_n36888__, new_new_n36889__, new_new_n36890__, new_new_n36891__,
    new_new_n36892__, new_new_n36893__, new_new_n36894__, new_new_n36895__,
    new_new_n36896__, new_new_n36897__, new_new_n36898__, new_new_n36899__,
    new_new_n36900__, new_new_n36901__, new_new_n36902__, new_new_n36903__,
    new_new_n36904__, new_new_n36905__, new_new_n36906__, new_new_n36907__,
    new_new_n36908__, new_new_n36909__, new_new_n36910__, new_new_n36911__,
    new_new_n36912__, new_new_n36913__, new_new_n36914__, new_new_n36915__,
    new_new_n36916__, new_new_n36917__, new_new_n36918__, new_new_n36919__,
    new_new_n36920__, new_new_n36921__, new_new_n36922__, new_new_n36923__,
    new_new_n36924__, new_new_n36925__, new_new_n36926__, new_new_n36927__,
    new_new_n36928__, new_new_n36929__, new_new_n36930__, new_new_n36931__,
    new_new_n36932__, new_new_n36933__, new_new_n36934__, new_new_n36935__,
    new_new_n36936__, new_new_n36937__, new_new_n36938__, new_new_n36939__,
    new_new_n36940__, new_new_n36941__, new_new_n36942__, new_new_n36943__,
    new_new_n36944__, new_new_n36945__, new_new_n36946__, new_new_n36947__,
    new_new_n36948__, new_new_n36949__, new_new_n36950__, new_new_n36951__,
    new_new_n36952__, new_new_n36953__, new_new_n36954__, new_new_n36955__,
    new_new_n36956__, new_new_n36957__, new_new_n36958__, new_new_n36959__,
    new_new_n36960__, new_new_n36961__, new_new_n36962__, new_new_n36963__,
    new_new_n36964__, new_new_n36965__, new_new_n36966__, new_new_n36967__,
    new_new_n36968__, new_new_n36969__, new_new_n36970__, new_new_n36971__,
    new_new_n36972__, new_new_n36973__, new_new_n36974__, new_new_n36975__,
    new_new_n36976__, new_new_n36977__, new_new_n36978__, new_new_n36979__,
    new_new_n36980__, new_new_n36981__, new_new_n36982__, new_new_n36983__,
    new_new_n36984__, new_new_n36985__, new_new_n36986__, new_new_n36987__,
    new_new_n36988__, new_new_n36989__, new_new_n36990__, new_new_n36991__,
    new_new_n36992__, new_new_n36993__, new_new_n36994__, new_new_n36995__,
    new_new_n36996__, new_new_n36997__, new_new_n36998__, new_new_n36999__,
    new_new_n37000__, new_new_n37001__, new_new_n37002__, new_new_n37003__,
    new_new_n37004__, new_new_n37005__, new_new_n37006__, new_new_n37007__,
    new_new_n37008__, new_new_n37009__, new_new_n37010__, new_new_n37011__,
    new_new_n37012__, new_new_n37013__, new_new_n37014__, new_new_n37015__,
    new_new_n37016__, new_new_n37017__, new_new_n37018__, new_new_n37019__,
    new_new_n37020__, new_new_n37021__, new_new_n37022__, new_new_n37023__,
    new_new_n37024__, new_new_n37025__, new_new_n37026__, new_new_n37027__,
    new_new_n37028__, new_new_n37029__, new_new_n37030__, new_new_n37031__,
    new_new_n37032__, new_new_n37033__, new_new_n37034__, new_new_n37035__,
    new_new_n37036__, new_new_n37037__, new_new_n37038__, new_new_n37039__,
    new_new_n37040__, new_new_n37041__, new_new_n37042__, new_new_n37043__,
    new_new_n37044__, new_new_n37045__, new_new_n37046__, new_new_n37047__,
    new_new_n37048__, new_new_n37049__, new_new_n37050__, new_new_n37051__,
    new_new_n37052__, new_new_n37053__, new_new_n37054__, new_new_n37055__,
    new_new_n37056__, new_new_n37058__, new_new_n37059__, new_new_n37060__,
    new_new_n37061__, new_new_n37062__, new_new_n37063__, new_new_n37064__,
    new_new_n37065__, new_new_n37066__, new_new_n37067__, new_new_n37068__,
    new_new_n37069__, new_new_n37070__, new_new_n37071__, new_new_n37072__,
    new_new_n37073__, new_new_n37074__, new_new_n37075__, new_new_n37076__,
    new_new_n37077__, new_new_n37078__, new_new_n37079__, new_new_n37080__,
    new_new_n37081__, new_new_n37082__, new_new_n37083__, new_new_n37084__,
    new_new_n37085__, new_new_n37086__, new_new_n37087__, new_new_n37088__,
    new_new_n37089__, new_new_n37090__, new_new_n37091__, new_new_n37092__,
    new_new_n37093__, new_new_n37094__, new_new_n37095__, new_new_n37096__,
    new_new_n37097__, new_new_n37098__, new_new_n37099__, new_new_n37100__,
    new_new_n37101__, new_new_n37102__, new_new_n37103__, new_new_n37104__,
    new_new_n37105__, new_new_n37106__, new_new_n37107__, new_new_n37108__,
    new_new_n37109__, new_new_n37110__, new_new_n37111__, new_new_n37112__,
    new_new_n37113__, new_new_n37114__, new_new_n37115__, new_new_n37116__,
    new_new_n37117__, new_new_n37118__, new_new_n37119__, new_new_n37120__,
    new_new_n37121__, new_new_n37122__, new_new_n37123__, new_new_n37124__,
    new_new_n37125__, new_new_n37126__, new_new_n37127__, new_new_n37128__,
    new_new_n37129__, new_new_n37130__, new_new_n37131__, new_new_n37132__,
    new_new_n37133__, new_new_n37134__, new_new_n37135__, new_new_n37136__,
    new_new_n37137__, new_new_n37138__, new_new_n37139__, new_new_n37140__,
    new_new_n37141__, new_new_n37142__, new_new_n37143__, new_new_n37144__,
    new_new_n37145__, new_new_n37146__, new_new_n37147__, new_new_n37148__,
    new_new_n37149__, new_new_n37150__, new_new_n37151__, new_new_n37152__,
    new_new_n37153__, new_new_n37154__, new_new_n37155__, new_new_n37156__,
    new_new_n37157__, new_new_n37158__, new_new_n37159__, new_new_n37160__,
    new_new_n37161__, new_new_n37162__, new_new_n37163__, new_new_n37164__,
    new_new_n37165__, new_new_n37166__, new_new_n37167__, new_new_n37168__,
    new_new_n37169__, new_new_n37170__, new_new_n37171__, new_new_n37172__,
    new_new_n37173__, new_new_n37174__, new_new_n37175__, new_new_n37176__,
    new_new_n37177__, new_new_n37178__, new_new_n37179__, new_new_n37180__,
    new_new_n37181__, new_new_n37182__, new_new_n37183__, new_new_n37184__,
    new_new_n37185__, new_new_n37186__, new_new_n37187__, new_new_n37188__,
    new_new_n37189__, new_new_n37190__, new_new_n37191__, new_new_n37192__,
    new_new_n37193__, new_new_n37194__, new_new_n37195__, new_new_n37196__,
    new_new_n37197__, new_new_n37198__, new_new_n37199__, new_new_n37200__,
    new_new_n37201__, new_new_n37202__, new_new_n37203__, new_new_n37204__,
    new_new_n37205__, new_new_n37206__, new_new_n37207__, new_new_n37208__,
    new_new_n37209__, new_new_n37210__, new_new_n37211__, new_new_n37212__,
    new_new_n37213__, new_new_n37214__, new_new_n37215__, new_new_n37216__,
    new_new_n37217__, new_new_n37218__, new_new_n37219__, new_new_n37220__,
    new_new_n37221__, new_new_n37222__, new_new_n37223__, new_new_n37224__,
    new_new_n37225__, new_new_n37226__, new_new_n37227__, new_new_n37228__,
    new_new_n37229__, new_new_n37230__, new_new_n37231__, new_new_n37232__,
    new_new_n37233__, new_new_n37234__, new_new_n37236__, new_new_n37237__,
    new_new_n37238__, new_new_n37239__, new_new_n37240__, new_new_n37241__,
    new_new_n37242__, new_new_n37243__, new_new_n37244__, new_new_n37245__,
    new_new_n37246__, new_new_n37247__, new_new_n37248__, new_new_n37249__,
    new_new_n37250__, new_new_n37251__, new_new_n37252__, new_new_n37253__,
    new_new_n37254__, new_new_n37255__, new_new_n37256__, new_new_n37257__,
    new_new_n37258__, new_new_n37259__, new_new_n37260__, new_new_n37261__,
    new_new_n37262__, new_new_n37263__, new_new_n37264__, new_new_n37265__,
    new_new_n37266__, new_new_n37267__, new_new_n37268__, new_new_n37269__,
    new_new_n37270__, new_new_n37271__, new_new_n37272__, new_new_n37273__,
    new_new_n37274__, new_new_n37275__, new_new_n37276__, new_new_n37277__,
    new_new_n37278__, new_new_n37279__, new_new_n37280__, new_new_n37281__,
    new_new_n37282__, new_new_n37283__, new_new_n37284__, new_new_n37285__,
    new_new_n37286__, new_new_n37287__, new_new_n37288__, new_new_n37289__,
    new_new_n37290__, new_new_n37291__, new_new_n37292__, new_new_n37293__,
    new_new_n37294__, new_new_n37295__, new_new_n37296__, new_new_n37297__,
    new_new_n37298__, new_new_n37299__, new_new_n37300__, new_new_n37301__,
    new_new_n37302__, new_new_n37303__, new_new_n37304__, new_new_n37305__,
    new_new_n37306__, new_new_n37307__, new_new_n37308__, new_new_n37309__,
    new_new_n37310__, new_new_n37311__, new_new_n37312__, new_new_n37313__,
    new_new_n37314__, new_new_n37315__, new_new_n37316__, new_new_n37317__,
    new_new_n37318__, new_new_n37319__, new_new_n37320__, new_new_n37321__,
    new_new_n37322__, new_new_n37323__, new_new_n37324__, new_new_n37325__,
    new_new_n37326__, new_new_n37327__, new_new_n37328__, new_new_n37329__,
    new_new_n37330__, new_new_n37331__, new_new_n37332__, new_new_n37333__,
    new_new_n37334__, new_new_n37335__, new_new_n37336__, new_new_n37337__,
    new_new_n37338__, new_new_n37339__, new_new_n37340__, new_new_n37341__,
    new_new_n37342__, new_new_n37343__, new_new_n37344__, new_new_n37345__,
    new_new_n37346__, new_new_n37347__, new_new_n37348__, new_new_n37349__,
    new_new_n37350__, new_new_n37351__, new_new_n37352__, new_new_n37353__,
    new_new_n37354__, new_new_n37355__, new_new_n37356__, new_new_n37357__,
    new_new_n37358__, new_new_n37359__, new_new_n37360__, new_new_n37361__,
    new_new_n37362__, new_new_n37363__, new_new_n37364__, new_new_n37365__,
    new_new_n37366__, new_new_n37367__, new_new_n37368__, new_new_n37369__,
    new_new_n37370__, new_new_n37371__, new_new_n37372__, new_new_n37373__,
    new_new_n37374__, new_new_n37375__, new_new_n37376__, new_new_n37378__,
    new_new_n37379__, new_new_n37380__, new_new_n37381__, new_new_n37382__,
    new_new_n37383__, new_new_n37384__, new_new_n37385__, new_new_n37386__,
    new_new_n37387__, new_new_n37388__, new_new_n37389__, new_new_n37390__,
    new_new_n37391__, new_new_n37392__, new_new_n37393__, new_new_n37394__,
    new_new_n37395__, new_new_n37396__, new_new_n37397__, new_new_n37398__,
    new_new_n37399__, new_new_n37400__, new_new_n37401__, new_new_n37402__,
    new_new_n37403__, new_new_n37404__, new_new_n37405__, new_new_n37406__,
    new_new_n37407__, new_new_n37408__, new_new_n37409__, new_new_n37410__,
    new_new_n37411__, new_new_n37412__, new_new_n37413__, new_new_n37414__,
    new_new_n37415__, new_new_n37416__, new_new_n37417__, new_new_n37418__,
    new_new_n37419__, new_new_n37420__, new_new_n37421__, new_new_n37422__,
    new_new_n37423__, new_new_n37424__, new_new_n37425__, new_new_n37426__,
    new_new_n37427__, new_new_n37428__, new_new_n37429__, new_new_n37430__,
    new_new_n37431__, new_new_n37432__, new_new_n37433__, new_new_n37434__,
    new_new_n37435__, new_new_n37436__, new_new_n37437__, new_new_n37438__,
    new_new_n37439__, new_new_n37440__, new_new_n37441__, new_new_n37442__,
    new_new_n37443__, new_new_n37444__, new_new_n37445__, new_new_n37446__,
    new_new_n37447__, new_new_n37448__, new_new_n37449__, new_new_n37450__,
    new_new_n37451__, new_new_n37452__, new_new_n37453__, new_new_n37454__,
    new_new_n37455__, new_new_n37456__, new_new_n37457__, new_new_n37458__,
    new_new_n37459__, new_new_n37460__, new_new_n37461__, new_new_n37462__,
    new_new_n37463__, new_new_n37464__, new_new_n37465__, new_new_n37466__,
    new_new_n37467__, new_new_n37468__, new_new_n37469__, new_new_n37470__,
    new_new_n37471__, new_new_n37472__, new_new_n37473__, new_new_n37474__,
    new_new_n37475__, new_new_n37476__, new_new_n37477__, new_new_n37478__,
    new_new_n37479__, new_new_n37480__, new_new_n37481__, new_new_n37482__,
    new_new_n37483__, new_new_n37484__, new_new_n37485__, new_new_n37486__,
    new_new_n37487__, new_new_n37488__, new_new_n37489__, new_new_n37490__,
    new_new_n37491__, new_new_n37492__, new_new_n37493__, new_new_n37494__,
    new_new_n37495__, new_new_n37496__, new_new_n37497__, new_new_n37498__,
    new_new_n37499__, new_new_n37500__, new_new_n37501__, new_new_n37502__,
    new_new_n37503__, new_new_n37504__, new_new_n37505__, new_new_n37506__,
    new_new_n37507__, new_new_n37508__, new_new_n37509__, new_new_n37510__,
    new_new_n37511__, new_new_n37512__, new_new_n37513__, new_new_n37514__,
    new_new_n37515__, new_new_n37516__, new_new_n37517__, new_new_n37518__,
    new_new_n37520__, new_new_n37521__, new_new_n37522__, new_new_n37523__,
    new_new_n37524__, new_new_n37525__, new_new_n37526__, new_new_n37527__,
    new_new_n37528__, new_new_n37529__, new_new_n37530__, new_new_n37531__,
    new_new_n37532__, new_new_n37533__, new_new_n37534__, new_new_n37535__,
    new_new_n37536__, new_new_n37537__, new_new_n37538__, new_new_n37539__,
    new_new_n37540__, new_new_n37541__, new_new_n37542__, new_new_n37543__,
    new_new_n37544__, new_new_n37545__, new_new_n37546__, new_new_n37547__,
    new_new_n37548__, new_new_n37549__, new_new_n37550__, new_new_n37551__,
    new_new_n37552__, new_new_n37553__, new_new_n37554__, new_new_n37555__,
    new_new_n37556__, new_new_n37557__, new_new_n37558__, new_new_n37559__,
    new_new_n37560__, new_new_n37561__, new_new_n37562__, new_new_n37563__,
    new_new_n37564__, new_new_n37565__, new_new_n37566__, new_new_n37567__,
    new_new_n37568__, new_new_n37569__, new_new_n37570__, new_new_n37571__,
    new_new_n37572__, new_new_n37573__, new_new_n37574__, new_new_n37575__,
    new_new_n37576__, new_new_n37577__, new_new_n37578__, new_new_n37579__,
    new_new_n37580__, new_new_n37581__, new_new_n37582__, new_new_n37583__,
    new_new_n37584__, new_new_n37585__, new_new_n37586__, new_new_n37587__,
    new_new_n37588__, new_new_n37589__, new_new_n37590__, new_new_n37591__,
    new_new_n37592__, new_new_n37593__, new_new_n37594__, new_new_n37595__,
    new_new_n37596__, new_new_n37597__, new_new_n37598__, new_new_n37599__,
    new_new_n37600__, new_new_n37601__, new_new_n37602__, new_new_n37603__,
    new_new_n37604__, new_new_n37605__, new_new_n37606__, new_new_n37607__,
    new_new_n37608__, new_new_n37609__, new_new_n37610__, new_new_n37611__,
    new_new_n37612__, new_new_n37613__, new_new_n37614__, new_new_n37615__,
    new_new_n37616__, new_new_n37617__, new_new_n37618__, new_new_n37619__,
    new_new_n37620__, new_new_n37621__, new_new_n37622__, new_new_n37623__,
    new_new_n37624__, new_new_n37625__, new_new_n37626__, new_new_n37627__,
    new_new_n37628__, new_new_n37629__, new_new_n37630__, new_new_n37631__,
    new_new_n37632__, new_new_n37633__, new_new_n37634__, new_new_n37635__,
    new_new_n37636__, new_new_n37637__, new_new_n37638__, new_new_n37639__,
    new_new_n37640__, new_new_n37641__, new_new_n37642__, new_new_n37643__,
    new_new_n37644__, new_new_n37645__, new_new_n37646__, new_new_n37647__,
    new_new_n37648__, new_new_n37649__, new_new_n37650__, new_new_n37651__,
    new_new_n37652__, new_new_n37653__, new_new_n37654__, new_new_n37655__,
    new_new_n37656__, new_new_n37657__, new_new_n37658__, new_new_n37659__,
    new_new_n37661__, new_new_n37662__, new_new_n37663__, new_new_n37664__,
    new_new_n37665__, new_new_n37666__, new_new_n37667__, new_new_n37668__,
    new_new_n37669__, new_new_n37670__, new_new_n37671__, new_new_n37672__,
    new_new_n37673__, new_new_n37674__, new_new_n37675__, new_new_n37676__,
    new_new_n37677__, new_new_n37678__, new_new_n37679__, new_new_n37680__,
    new_new_n37681__, new_new_n37682__, new_new_n37683__, new_new_n37684__,
    new_new_n37685__, new_new_n37686__, new_new_n37687__, new_new_n37688__,
    new_new_n37689__, new_new_n37690__, new_new_n37691__, new_new_n37692__,
    new_new_n37693__, new_new_n37694__, new_new_n37695__, new_new_n37696__,
    new_new_n37697__, new_new_n37698__, new_new_n37699__, new_new_n37700__,
    new_new_n37701__, new_new_n37702__, new_new_n37703__, new_new_n37704__,
    new_new_n37705__, new_new_n37706__, new_new_n37707__, new_new_n37708__,
    new_new_n37709__, new_new_n37710__, new_new_n37711__, new_new_n37712__,
    new_new_n37713__, new_new_n37714__, new_new_n37715__, new_new_n37716__,
    new_new_n37717__, new_new_n37718__, new_new_n37719__, new_new_n37720__,
    new_new_n37721__, new_new_n37722__, new_new_n37723__, new_new_n37724__,
    new_new_n37725__, new_new_n37726__, new_new_n37727__, new_new_n37728__,
    new_new_n37729__, new_new_n37730__, new_new_n37731__, new_new_n37732__,
    new_new_n37733__, new_new_n37734__, new_new_n37735__, new_new_n37736__,
    new_new_n37737__, new_new_n37738__, new_new_n37739__, new_new_n37740__,
    new_new_n37741__, new_new_n37742__, new_new_n37743__, new_new_n37744__,
    new_new_n37745__, new_new_n37746__, new_new_n37747__, new_new_n37748__,
    new_new_n37749__, new_new_n37750__, new_new_n37751__, new_new_n37752__,
    new_new_n37753__, new_new_n37754__, new_new_n37755__, new_new_n37756__,
    new_new_n37757__, new_new_n37758__, new_new_n37759__, new_new_n37760__,
    new_new_n37761__, new_new_n37762__, new_new_n37763__, new_new_n37764__,
    new_new_n37765__, new_new_n37766__, new_new_n37767__, new_new_n37768__,
    new_new_n37769__, new_new_n37770__, new_new_n37771__, new_new_n37772__,
    new_new_n37773__, new_new_n37774__, new_new_n37775__, new_new_n37776__,
    new_new_n37777__, new_new_n37778__, new_new_n37779__, new_new_n37780__,
    new_new_n37781__, new_new_n37782__, new_new_n37783__, new_new_n37784__,
    new_new_n37785__, new_new_n37786__, new_new_n37787__, new_new_n37788__,
    new_new_n37789__, new_new_n37790__, new_new_n37791__, new_new_n37792__,
    new_new_n37793__, new_new_n37794__, new_new_n37795__, new_new_n37796__,
    new_new_n37797__, new_new_n37798__, new_new_n37799__, new_new_n37800__,
    new_new_n37801__, new_new_n37802__, new_new_n37803__, new_new_n37804__,
    new_new_n37805__, new_new_n37806__, new_new_n37807__, new_new_n37808__,
    new_new_n37809__, new_new_n37810__, new_new_n37812__, new_new_n37813__,
    new_new_n37814__, new_new_n37815__, new_new_n37816__, new_new_n37817__,
    new_new_n37818__, new_new_n37819__, new_new_n37820__, new_new_n37821__,
    new_new_n37822__, new_new_n37823__, new_new_n37824__, new_new_n37825__,
    new_new_n37826__, new_new_n37827__, new_new_n37828__, new_new_n37829__,
    new_new_n37830__, new_new_n37831__, new_new_n37832__, new_new_n37833__,
    new_new_n37834__, new_new_n37835__, new_new_n37836__, new_new_n37837__,
    new_new_n37838__, new_new_n37839__, new_new_n37840__, new_new_n37841__,
    new_new_n37842__, new_new_n37843__, new_new_n37844__, new_new_n37845__,
    new_new_n37846__, new_new_n37847__, new_new_n37848__, new_new_n37849__,
    new_new_n37850__, new_new_n37851__, new_new_n37852__, new_new_n37853__,
    new_new_n37854__, new_new_n37855__, new_new_n37856__, new_new_n37857__,
    new_new_n37858__, new_new_n37859__, new_new_n37860__, new_new_n37861__,
    new_new_n37862__, new_new_n37863__, new_new_n37864__, new_new_n37865__,
    new_new_n37866__, new_new_n37867__, new_new_n37868__, new_new_n37869__,
    new_new_n37870__, new_new_n37871__, new_new_n37872__, new_new_n37873__,
    new_new_n37874__, new_new_n37875__, new_new_n37876__, new_new_n37877__,
    new_new_n37878__, new_new_n37879__, new_new_n37880__, new_new_n37881__,
    new_new_n37882__, new_new_n37883__, new_new_n37884__, new_new_n37885__,
    new_new_n37886__, new_new_n37887__, new_new_n37888__, new_new_n37889__,
    new_new_n37890__, new_new_n37891__, new_new_n37892__, new_new_n37893__,
    new_new_n37894__, new_new_n37895__, new_new_n37896__, new_new_n37897__,
    new_new_n37898__, new_new_n37899__, new_new_n37900__, new_new_n37901__,
    new_new_n37902__, new_new_n37903__, new_new_n37904__, new_new_n37905__,
    new_new_n37906__, new_new_n37907__, new_new_n37908__, new_new_n37909__,
    new_new_n37910__, new_new_n37911__, new_new_n37912__, new_new_n37913__,
    new_new_n37914__, new_new_n37915__, new_new_n37916__, new_new_n37917__,
    new_new_n37918__, new_new_n37919__, new_new_n37920__, new_new_n37921__,
    new_new_n37922__, new_new_n37923__, new_new_n37924__, new_new_n37925__,
    new_new_n37926__, new_new_n37927__, new_new_n37928__, new_new_n37929__,
    new_new_n37930__, new_new_n37931__, new_new_n37932__, new_new_n37933__,
    new_new_n37934__, new_new_n37935__, new_new_n37936__, new_new_n37937__,
    new_new_n37938__, new_new_n37939__, new_new_n37940__, new_new_n37941__,
    new_new_n37942__, new_new_n37943__, new_new_n37944__, new_new_n37945__,
    new_new_n37946__, new_new_n37947__, new_new_n37948__, new_new_n37949__,
    new_new_n37950__, new_new_n37951__, new_new_n37952__, new_new_n37953__,
    new_new_n37954__, new_new_n37955__, new_new_n37956__, new_new_n37957__,
    new_new_n37958__, new_new_n37959__, new_new_n37960__, new_new_n37961__,
    new_new_n37962__, new_new_n37963__, new_new_n37964__, new_new_n37965__,
    new_new_n37966__, new_new_n37967__, new_new_n37969__, new_new_n37970__,
    new_new_n37971__, new_new_n37972__, new_new_n37973__, new_new_n37974__,
    new_new_n37975__, new_new_n37976__, new_new_n37977__, new_new_n37978__,
    new_new_n37979__, new_new_n37980__, new_new_n37981__, new_new_n37982__,
    new_new_n37983__, new_new_n37984__, new_new_n37985__, new_new_n37986__,
    new_new_n37987__, new_new_n37988__, new_new_n37989__, new_new_n37990__,
    new_new_n37991__, new_new_n37992__, new_new_n37993__, new_new_n37994__,
    new_new_n37995__, new_new_n37996__, new_new_n37997__, new_new_n37998__,
    new_new_n37999__, new_new_n38000__, new_new_n38001__, new_new_n38002__,
    new_new_n38003__, new_new_n38004__, new_new_n38005__, new_new_n38006__,
    new_new_n38007__, new_new_n38008__, new_new_n38009__, new_new_n38010__,
    new_new_n38011__, new_new_n38012__, new_new_n38013__, new_new_n38014__,
    new_new_n38015__, new_new_n38016__, new_new_n38017__, new_new_n38018__,
    new_new_n38019__, new_new_n38020__, new_new_n38021__, new_new_n38022__,
    new_new_n38023__, new_new_n38024__, new_new_n38025__, new_new_n38026__,
    new_new_n38027__, new_new_n38028__, new_new_n38029__, new_new_n38030__,
    new_new_n38031__, new_new_n38032__, new_new_n38033__, new_new_n38034__,
    new_new_n38035__, new_new_n38036__, new_new_n38037__, new_new_n38038__,
    new_new_n38039__, new_new_n38040__, new_new_n38041__, new_new_n38042__,
    new_new_n38043__, new_new_n38044__, new_new_n38045__, new_new_n38046__,
    new_new_n38047__, new_new_n38048__, new_new_n38049__, new_new_n38050__,
    new_new_n38051__, new_new_n38052__, new_new_n38053__, new_new_n38054__,
    new_new_n38055__, new_new_n38056__, new_new_n38057__, new_new_n38058__,
    new_new_n38059__, new_new_n38060__, new_new_n38061__, new_new_n38062__,
    new_new_n38063__, new_new_n38064__, new_new_n38065__, new_new_n38066__,
    new_new_n38067__, new_new_n38068__, new_new_n38069__, new_new_n38070__,
    new_new_n38071__, new_new_n38072__, new_new_n38073__, new_new_n38074__,
    new_new_n38075__, new_new_n38076__, new_new_n38077__, new_new_n38078__,
    new_new_n38079__, new_new_n38080__, new_new_n38081__, new_new_n38082__,
    new_new_n38083__, new_new_n38084__, new_new_n38085__, new_new_n38086__,
    new_new_n38087__, new_new_n38088__, new_new_n38089__, new_new_n38090__,
    new_new_n38091__, new_new_n38093__, new_new_n38094__, new_new_n38095__,
    new_new_n38096__, new_new_n38097__, new_new_n38098__, new_new_n38099__,
    new_new_n38100__, new_new_n38101__, new_new_n38102__, new_new_n38103__,
    new_new_n38104__, new_new_n38105__, new_new_n38106__, new_new_n38107__,
    new_new_n38108__, new_new_n38109__, new_new_n38110__, new_new_n38111__,
    new_new_n38112__, new_new_n38113__, new_new_n38114__, new_new_n38115__,
    new_new_n38116__, new_new_n38117__, new_new_n38118__, new_new_n38119__,
    new_new_n38120__, new_new_n38121__, new_new_n38122__, new_new_n38123__,
    new_new_n38124__, new_new_n38125__, new_new_n38126__, new_new_n38127__,
    new_new_n38128__, new_new_n38129__, new_new_n38130__, new_new_n38131__,
    new_new_n38132__, new_new_n38133__, new_new_n38134__, new_new_n38135__,
    new_new_n38136__, new_new_n38137__, new_new_n38138__, new_new_n38139__,
    new_new_n38140__, new_new_n38141__, new_new_n38142__, new_new_n38143__,
    new_new_n38144__, new_new_n38145__, new_new_n38146__, new_new_n38147__,
    new_new_n38148__, new_new_n38149__, new_new_n38150__, new_new_n38151__,
    new_new_n38152__, new_new_n38153__, new_new_n38154__, new_new_n38155__,
    new_new_n38156__, new_new_n38157__, new_new_n38158__, new_new_n38159__,
    new_new_n38160__, new_new_n38161__, new_new_n38162__, new_new_n38163__,
    new_new_n38164__, new_new_n38165__, new_new_n38166__, new_new_n38167__,
    new_new_n38168__, new_new_n38169__, new_new_n38170__, new_new_n38171__,
    new_new_n38172__, new_new_n38173__, new_new_n38174__, new_new_n38175__,
    new_new_n38176__, new_new_n38177__, new_new_n38178__, new_new_n38179__,
    new_new_n38180__, new_new_n38181__, new_new_n38182__, new_new_n38183__,
    new_new_n38184__, new_new_n38185__, new_new_n38186__, new_new_n38187__,
    new_new_n38188__, new_new_n38189__, new_new_n38190__, new_new_n38191__,
    new_new_n38192__, new_new_n38193__, new_new_n38194__, new_new_n38195__,
    new_new_n38196__, new_new_n38197__, new_new_n38198__, new_new_n38199__,
    new_new_n38200__, new_new_n38201__, new_new_n38202__, new_new_n38203__,
    new_new_n38204__, new_new_n38205__, new_new_n38206__, new_new_n38207__,
    new_new_n38208__, new_new_n38209__, new_new_n38210__, new_new_n38211__,
    new_new_n38212__, new_new_n38213__, new_new_n38214__, new_new_n38215__,
    new_new_n38216__, new_new_n38217__, new_new_n38218__, new_new_n38219__,
    new_new_n38220__, new_new_n38222__, new_new_n38223__, new_new_n38224__,
    new_new_n38225__, new_new_n38226__, new_new_n38227__, new_new_n38228__,
    new_new_n38229__, new_new_n38230__, new_new_n38231__, new_new_n38232__,
    new_new_n38233__, new_new_n38234__, new_new_n38235__, new_new_n38236__,
    new_new_n38237__, new_new_n38238__, new_new_n38239__, new_new_n38240__,
    new_new_n38241__, new_new_n38242__, new_new_n38243__, new_new_n38244__,
    new_new_n38245__, new_new_n38246__, new_new_n38247__, new_new_n38248__,
    new_new_n38249__, new_new_n38250__, new_new_n38251__, new_new_n38252__,
    new_new_n38253__, new_new_n38254__, new_new_n38255__, new_new_n38256__,
    new_new_n38257__, new_new_n38258__, new_new_n38259__, new_new_n38260__,
    new_new_n38261__, new_new_n38262__, new_new_n38263__, new_new_n38264__,
    new_new_n38265__, new_new_n38266__, new_new_n38267__, new_new_n38268__,
    new_new_n38269__, new_new_n38270__, new_new_n38271__, new_new_n38272__,
    new_new_n38273__, new_new_n38274__, new_new_n38275__, new_new_n38276__,
    new_new_n38277__, new_new_n38278__, new_new_n38279__, new_new_n38280__,
    new_new_n38281__, new_new_n38282__, new_new_n38283__, new_new_n38284__,
    new_new_n38285__, new_new_n38286__, new_new_n38287__, new_new_n38288__,
    new_new_n38289__, new_new_n38290__, new_new_n38291__, new_new_n38292__,
    new_new_n38293__, new_new_n38294__, new_new_n38295__, new_new_n38296__,
    new_new_n38297__, new_new_n38298__, new_new_n38299__, new_new_n38300__,
    new_new_n38301__, new_new_n38302__, new_new_n38303__, new_new_n38304__,
    new_new_n38305__, new_new_n38306__, new_new_n38307__, new_new_n38308__,
    new_new_n38309__, new_new_n38310__, new_new_n38311__, new_new_n38312__,
    new_new_n38313__, new_new_n38314__, new_new_n38315__, new_new_n38316__,
    new_new_n38317__, new_new_n38318__, new_new_n38320__, new_new_n38321__,
    new_new_n38322__, new_new_n38323__, new_new_n38324__, new_new_n38325__,
    new_new_n38326__, new_new_n38327__, new_new_n38328__, new_new_n38329__,
    new_new_n38330__, new_new_n38331__, new_new_n38332__, new_new_n38333__,
    new_new_n38334__, new_new_n38335__, new_new_n38336__, new_new_n38337__,
    new_new_n38338__, new_new_n38339__, new_new_n38340__, new_new_n38341__,
    new_new_n38342__, new_new_n38343__, new_new_n38344__, new_new_n38345__,
    new_new_n38346__, new_new_n38347__, new_new_n38348__, new_new_n38349__,
    new_new_n38350__, new_new_n38351__, new_new_n38352__, new_new_n38353__,
    new_new_n38354__, new_new_n38355__, new_new_n38356__, new_new_n38357__,
    new_new_n38358__, new_new_n38359__, new_new_n38360__, new_new_n38361__,
    new_new_n38362__, new_new_n38363__, new_new_n38364__, new_new_n38365__,
    new_new_n38366__, new_new_n38367__, new_new_n38368__, new_new_n38369__,
    new_new_n38370__, new_new_n38371__, new_new_n38372__, new_new_n38373__,
    new_new_n38374__, new_new_n38375__, new_new_n38376__, new_new_n38377__,
    new_new_n38378__, new_new_n38379__, new_new_n38380__, new_new_n38381__,
    new_new_n38382__, new_new_n38383__, new_new_n38384__, new_new_n38385__,
    new_new_n38386__, new_new_n38387__, new_new_n38388__, new_new_n38389__,
    new_new_n38390__, new_new_n38391__, new_new_n38392__, new_new_n38393__,
    new_new_n38394__, new_new_n38395__, new_new_n38396__, new_new_n38397__,
    new_new_n38398__, new_new_n38399__, new_new_n38400__, new_new_n38401__,
    new_new_n38402__, new_new_n38403__, new_new_n38404__, new_new_n38405__,
    new_new_n38406__, new_new_n38407__, new_new_n38408__, new_new_n38409__,
    new_new_n38410__, new_new_n38411__, new_new_n38412__, new_new_n38413__,
    new_new_n38414__, new_new_n38415__, new_new_n38416__, new_new_n38417__,
    new_new_n38418__, new_new_n38419__, new_new_n38420__, new_new_n38421__,
    new_new_n38422__, new_new_n38423__, new_new_n38424__, new_new_n38425__,
    new_new_n38426__, new_new_n38427__, new_new_n38428__, new_new_n38429__,
    new_new_n38430__, new_new_n38431__, new_new_n38432__, new_new_n38433__,
    new_new_n38434__, new_new_n38435__, new_new_n38437__, new_new_n38438__,
    new_new_n38439__, new_new_n38440__, new_new_n38441__, new_new_n38442__,
    new_new_n38443__, new_new_n38444__, new_new_n38445__, new_new_n38446__,
    new_new_n38447__, new_new_n38448__, new_new_n38449__, new_new_n38450__,
    new_new_n38451__, new_new_n38452__, new_new_n38453__, new_new_n38454__,
    new_new_n38455__, new_new_n38456__, new_new_n38457__, new_new_n38458__,
    new_new_n38459__, new_new_n38460__, new_new_n38461__, new_new_n38462__,
    new_new_n38463__, new_new_n38464__, new_new_n38465__, new_new_n38466__,
    new_new_n38467__, new_new_n38468__, new_new_n38469__, new_new_n38470__,
    new_new_n38471__, new_new_n38472__, new_new_n38473__, new_new_n38474__,
    new_new_n38475__, new_new_n38476__, new_new_n38477__, new_new_n38478__,
    new_new_n38479__, new_new_n38480__, new_new_n38481__, new_new_n38482__,
    new_new_n38483__, new_new_n38484__, new_new_n38485__, new_new_n38486__,
    new_new_n38487__, new_new_n38488__, new_new_n38489__, new_new_n38490__,
    new_new_n38491__, new_new_n38492__, new_new_n38493__, new_new_n38494__,
    new_new_n38495__, new_new_n38496__, new_new_n38497__, new_new_n38498__,
    new_new_n38499__, new_new_n38500__, new_new_n38501__, new_new_n38502__,
    new_new_n38503__, new_new_n38504__, new_new_n38505__, new_new_n38506__,
    new_new_n38507__, new_new_n38508__, new_new_n38509__, new_new_n38510__,
    new_new_n38512__, new_new_n38513__, new_new_n38514__, new_new_n38515__,
    new_new_n38516__, new_new_n38517__, new_new_n38518__, new_new_n38519__,
    new_new_n38520__, new_new_n38521__, new_new_n38522__, new_new_n38523__,
    new_new_n38524__, new_new_n38525__, new_new_n38526__, new_new_n38527__,
    new_new_n38528__, new_new_n38529__, new_new_n38530__, new_new_n38531__,
    new_new_n38532__, new_new_n38533__, new_new_n38534__, new_new_n38535__,
    new_new_n38536__, new_new_n38537__, new_new_n38538__, new_new_n38539__,
    new_new_n38540__, new_new_n38541__, new_new_n38542__, new_new_n38543__,
    new_new_n38544__, new_new_n38545__, new_new_n38546__, new_new_n38547__,
    new_new_n38548__, new_new_n38549__, new_new_n38550__, new_new_n38551__,
    new_new_n38552__, new_new_n38553__, new_new_n38554__, new_new_n38555__,
    new_new_n38556__, new_new_n38557__, new_new_n38558__, new_new_n38559__,
    new_new_n38560__, new_new_n38561__, new_new_n38562__, new_new_n38563__,
    new_new_n38564__, new_new_n38565__, new_new_n38566__, new_new_n38567__,
    new_new_n38568__, new_new_n38569__, new_new_n38570__, new_new_n38571__,
    new_new_n38572__, new_new_n38573__, new_new_n38574__, new_new_n38575__,
    new_new_n38576__, new_new_n38577__, new_new_n38578__, new_new_n38579__,
    new_new_n38580__, new_new_n38581__, new_new_n38582__, new_new_n38583__,
    new_new_n38584__, new_new_n38585__, new_new_n38586__, new_new_n38587__,
    new_new_n38588__, new_new_n38589__, new_new_n38590__, new_new_n38591__,
    new_new_n38592__, new_new_n38593__, new_new_n38594__, new_new_n38595__,
    new_new_n38596__, new_new_n38597__, new_new_n38598__, new_new_n38599__,
    new_new_n38600__, new_new_n38601__, new_new_n38602__, new_new_n38603__;
  assign new_new_n65__ = pi27 & pi28;
  assign new_new_n66__ = pi26 & new_new_n65__;
  assign new_new_n67__ = ~pi27 & ~pi28;
  assign new_new_n68__ = ~pi26 & new_new_n67__;
  assign new_new_n69__ = ~pi29 & ~new_new_n68__;
  assign new_new_n70__ = ~new_new_n66__ & ~new_new_n69__;
  assign new_new_n71__ = ~pi29 & ~pi30;
  assign new_new_n72__ = new_new_n65__ & new_new_n71__;
  assign new_new_n73__ = pi23 & ~pi24;
  assign new_new_n74__ = pi25 & pi26;
  assign new_new_n75__ = new_new_n73__ & new_new_n74__;
  assign new_new_n76__ = new_new_n72__ & new_new_n75__;
  assign new_new_n77__ = ~pi27 & pi28;
  assign new_new_n78__ = new_new_n71__ & new_new_n77__;
  assign new_new_n79__ = pi24 & pi26;
  assign new_new_n80__ = pi23 & pi25;
  assign new_new_n81__ = new_new_n79__ & new_new_n80__;
  assign new_new_n82__ = new_new_n78__ & new_new_n81__;
  assign new_new_n83__ = ~new_new_n76__ & ~new_new_n82__;
  assign new_new_n84__ = pi27 & ~pi28;
  assign new_new_n85__ = new_new_n71__ & new_new_n84__;
  assign new_new_n86__ = pi25 & ~pi26;
  assign new_new_n87__ = new_new_n73__ & new_new_n86__;
  assign new_new_n88__ = new_new_n85__ & new_new_n87__;
  assign new_new_n89__ = ~pi24 & ~pi26;
  assign new_new_n90__ = ~pi23 & ~pi25;
  assign new_new_n91__ = new_new_n89__ & new_new_n90__;
  assign new_new_n92__ = new_new_n72__ & new_new_n91__;
  assign new_new_n93__ = ~new_new_n88__ & ~new_new_n92__;
  assign new_new_n94__ = ~pi29 & pi30;
  assign new_new_n95__ = new_new_n77__ & new_new_n94__;
  assign new_new_n96__ = new_new_n87__ & new_new_n95__;
  assign new_new_n97__ = new_new_n67__ & new_new_n71__;
  assign new_new_n98__ = ~pi25 & pi26;
  assign new_new_n99__ = pi23 & pi24;
  assign new_new_n100__ = new_new_n98__ & new_new_n99__;
  assign new_new_n101__ = new_new_n97__ & new_new_n100__;
  assign new_new_n102__ = ~new_new_n96__ & ~new_new_n101__;
  assign new_new_n103__ = new_new_n75__ & new_new_n78__;
  assign new_new_n104__ = ~pi23 & ~pi24;
  assign new_new_n105__ = new_new_n86__ & new_new_n104__;
  assign new_new_n106__ = new_new_n95__ & new_new_n105__;
  assign new_new_n107__ = ~new_new_n103__ & ~new_new_n106__;
  assign new_new_n108__ = new_new_n75__ & new_new_n85__;
  assign new_new_n109__ = ~pi23 & pi24;
  assign new_new_n110__ = ~new_new_n73__ & ~new_new_n109__;
  assign new_new_n111__ = ~pi24 & new_new_n110__;
  assign new_new_n112__ = ~pi23 & pi25;
  assign new_new_n113__ = pi26 & new_new_n112__;
  assign new_new_n114__ = ~new_new_n111__ & new_new_n113__;
  assign new_new_n115__ = new_new_n78__ & new_new_n114__;
  assign new_new_n116__ = ~new_new_n108__ & ~new_new_n115__;
  assign new_new_n117__ = ~pi24 & pi26;
  assign new_new_n118__ = new_new_n112__ & new_new_n117__;
  assign new_new_n119__ = new_new_n85__ & new_new_n118__;
  assign new_new_n120__ = new_new_n85__ & new_new_n100__;
  assign new_new_n121__ = ~new_new_n119__ & ~new_new_n120__;
  assign new_new_n122__ = new_new_n97__ & new_new_n104__;
  assign new_new_n123__ = pi26 & new_new_n122__;
  assign new_new_n124__ = pi25 & new_new_n123__;
  assign new_new_n125__ = pi29 & ~pi30;
  assign new_new_n126__ = new_new_n84__ & new_new_n125__;
  assign new_new_n127__ = new_new_n87__ & new_new_n126__;
  assign new_new_n128__ = pi24 & ~pi26;
  assign new_new_n129__ = new_new_n80__ & new_new_n128__;
  assign new_new_n130__ = new_new_n126__ & new_new_n129__;
  assign new_new_n131__ = ~new_new_n127__ & ~new_new_n130__;
  assign new_new_n132__ = new_new_n85__ & ~new_new_n91__;
  assign new_new_n133__ = pi24 & ~pi25;
  assign new_new_n134__ = ~pi23 & pi26;
  assign new_new_n135__ = new_new_n133__ & new_new_n134__;
  assign new_new_n136__ = new_new_n132__ & new_new_n135__;
  assign new_new_n137__ = new_new_n67__ & new_new_n125__;
  assign new_new_n138__ = new_new_n87__ & new_new_n137__;
  assign new_new_n139__ = pi23 & new_new_n128__;
  assign new_new_n140__ = ~pi24 & pi25;
  assign new_new_n141__ = ~new_new_n133__ & ~new_new_n140__;
  assign new_new_n142__ = new_new_n139__ & ~new_new_n141__;
  assign new_new_n143__ = new_new_n95__ & new_new_n142__;
  assign new_new_n144__ = ~new_new_n138__ & ~new_new_n143__;
  assign new_new_n145__ = pi24 & pi25;
  assign new_new_n146__ = pi23 & new_new_n145__;
  assign new_new_n147__ = new_new_n68__ & new_new_n125__;
  assign new_new_n148__ = new_new_n146__ & new_new_n147__;
  assign new_new_n149__ = new_new_n109__ & new_new_n137__;
  assign new_new_n150__ = new_new_n86__ & new_new_n149__;
  assign new_new_n151__ = ~pi29 & new_new_n65__;
  assign new_new_n152__ = pi23 & ~pi25;
  assign new_new_n153__ = new_new_n89__ & new_new_n152__;
  assign new_new_n154__ = new_new_n151__ & new_new_n153__;
  assign new_new_n155__ = ~pi30 & new_new_n154__;
  assign new_new_n156__ = ~new_new_n136__ & ~new_new_n148__;
  assign new_new_n157__ = ~new_new_n150__ & ~new_new_n155__;
  assign new_new_n158__ = new_new_n156__ & new_new_n157__;
  assign new_new_n159__ = new_new_n144__ & new_new_n158__;
  assign new_new_n160__ = new_new_n78__ & new_new_n129__;
  assign new_new_n161__ = pi29 & pi30;
  assign new_new_n162__ = new_new_n65__ & new_new_n161__;
  assign new_new_n163__ = new_new_n112__ & new_new_n128__;
  assign new_new_n164__ = new_new_n162__ & new_new_n163__;
  assign new_new_n165__ = new_new_n65__ & new_new_n125__;
  assign new_new_n166__ = new_new_n142__ & new_new_n165__;
  assign new_new_n167__ = ~new_new_n164__ & ~new_new_n166__;
  assign new_new_n168__ = new_new_n97__ & new_new_n129__;
  assign new_new_n169__ = new_new_n77__ & new_new_n161__;
  assign new_new_n170__ = pi23 & new_new_n169__;
  assign new_new_n171__ = new_new_n74__ & new_new_n170__;
  assign new_new_n172__ = pi26 & ~new_new_n90__;
  assign new_new_n173__ = ~pi26 & ~new_new_n112__;
  assign new_new_n174__ = pi24 & ~new_new_n173__;
  assign new_new_n175__ = new_new_n162__ & ~new_new_n172__;
  assign new_new_n176__ = ~new_new_n174__ & new_new_n175__;
  assign new_new_n177__ = ~new_new_n171__ & ~new_new_n176__;
  assign new_new_n178__ = ~new_new_n168__ & new_new_n177__;
  assign new_new_n179__ = new_new_n153__ & new_new_n165__;
  assign new_new_n180__ = new_new_n90__ & new_new_n128__;
  assign new_new_n181__ = pi27 & new_new_n125__;
  assign new_new_n182__ = new_new_n180__ & new_new_n181__;
  assign new_new_n183__ = pi28 & new_new_n182__;
  assign new_new_n184__ = ~new_new_n179__ & ~new_new_n183__;
  assign new_new_n185__ = ~new_new_n160__ & new_new_n167__;
  assign new_new_n186__ = new_new_n184__ & new_new_n185__;
  assign new_new_n187__ = new_new_n178__ & new_new_n186__;
  assign new_new_n188__ = new_new_n126__ & new_new_n152__;
  assign new_new_n189__ = new_new_n79__ & new_new_n188__;
  assign new_new_n190__ = pi24 & new_new_n86__;
  assign new_new_n191__ = ~pi23 & new_new_n97__;
  assign new_new_n192__ = new_new_n190__ & new_new_n191__;
  assign new_new_n193__ = ~new_new_n189__ & ~new_new_n192__;
  assign new_new_n194__ = pi26 & ~new_new_n145__;
  assign new_new_n195__ = new_new_n126__ & new_new_n194__;
  assign new_new_n196__ = new_new_n87__ & new_new_n97__;
  assign new_new_n197__ = new_new_n113__ & new_new_n169__;
  assign new_new_n198__ = ~new_new_n104__ & new_new_n197__;
  assign new_new_n199__ = ~new_new_n196__ & ~new_new_n198__;
  assign new_new_n200__ = new_new_n118__ & new_new_n169__;
  assign new_new_n201__ = ~pi23 & new_new_n126__;
  assign new_new_n202__ = new_new_n190__ & new_new_n201__;
  assign new_new_n203__ = ~new_new_n195__ & ~new_new_n200__;
  assign new_new_n204__ = ~new_new_n202__ & new_new_n203__;
  assign new_new_n205__ = new_new_n193__ & new_new_n204__;
  assign new_new_n206__ = new_new_n199__ & new_new_n205__;
  assign new_new_n207__ = new_new_n137__ & new_new_n180__;
  assign new_new_n208__ = new_new_n135__ & new_new_n162__;
  assign new_new_n209__ = new_new_n118__ & new_new_n162__;
  assign new_new_n210__ = ~new_new_n208__ & ~new_new_n209__;
  assign new_new_n211__ = new_new_n77__ & new_new_n125__;
  assign new_new_n212__ = new_new_n153__ & new_new_n211__;
  assign new_new_n213__ = new_new_n97__ & new_new_n135__;
  assign new_new_n214__ = ~new_new_n207__ & ~new_new_n212__;
  assign new_new_n215__ = ~new_new_n213__ & new_new_n214__;
  assign new_new_n216__ = new_new_n210__ & new_new_n215__;
  assign new_new_n217__ = new_new_n84__ & new_new_n94__;
  assign new_new_n218__ = new_new_n114__ & new_new_n217__;
  assign new_new_n219__ = pi27 & pi30;
  assign new_new_n220__ = pi28 & ~pi29;
  assign new_new_n221__ = new_new_n219__ & new_new_n220__;
  assign new_new_n222__ = new_new_n100__ & new_new_n221__;
  assign new_new_n223__ = ~pi25 & new_new_n73__;
  assign new_new_n224__ = new_new_n67__ & new_new_n161__;
  assign new_new_n225__ = ~pi26 & new_new_n224__;
  assign new_new_n226__ = new_new_n223__ & new_new_n225__;
  assign new_new_n227__ = ~new_new_n222__ & ~new_new_n226__;
  assign new_new_n228__ = ~new_new_n218__ & new_new_n227__;
  assign new_new_n229__ = new_new_n72__ & new_new_n81__;
  assign new_new_n230__ = ~pi30 & new_new_n84__;
  assign new_new_n231__ = new_new_n163__ & new_new_n230__;
  assign new_new_n232__ = ~pi29 & new_new_n231__;
  assign new_new_n233__ = ~new_new_n229__ & ~new_new_n232__;
  assign new_new_n234__ = new_new_n73__ & new_new_n98__;
  assign new_new_n235__ = new_new_n224__ & new_new_n234__;
  assign new_new_n236__ = ~pi28 & pi29;
  assign new_new_n237__ = new_new_n219__ & new_new_n236__;
  assign new_new_n238__ = new_new_n153__ & new_new_n237__;
  assign new_new_n239__ = ~new_new_n235__ & ~new_new_n238__;
  assign new_new_n240__ = new_new_n75__ & new_new_n221__;
  assign new_new_n241__ = new_new_n90__ & new_new_n117__;
  assign new_new_n242__ = new_new_n217__ & new_new_n241__;
  assign new_new_n243__ = ~new_new_n240__ & ~new_new_n242__;
  assign new_new_n244__ = new_new_n239__ & new_new_n243__;
  assign new_new_n245__ = new_new_n233__ & new_new_n244__;
  assign new_new_n246__ = new_new_n91__ & new_new_n137__;
  assign new_new_n247__ = new_new_n75__ & new_new_n224__;
  assign new_new_n248__ = new_new_n163__ & new_new_n165__;
  assign new_new_n249__ = new_new_n105__ & new_new_n137__;
  assign new_new_n250__ = new_new_n95__ & new_new_n153__;
  assign new_new_n251__ = new_new_n180__ & new_new_n211__;
  assign new_new_n252__ = new_new_n78__ & new_new_n118__;
  assign new_new_n253__ = new_new_n81__ & new_new_n217__;
  assign new_new_n254__ = new_new_n72__ & new_new_n114__;
  assign new_new_n255__ = new_new_n147__ & new_new_n223__;
  assign new_new_n256__ = ~new_new_n254__ & ~new_new_n255__;
  assign new_new_n257__ = ~pi26 & new_new_n217__;
  assign new_new_n258__ = new_new_n146__ & new_new_n257__;
  assign new_new_n259__ = new_new_n95__ & new_new_n180__;
  assign new_new_n260__ = new_new_n118__ & new_new_n217__;
  assign new_new_n261__ = ~new_new_n259__ & ~new_new_n260__;
  assign new_new_n262__ = new_new_n65__ & new_new_n100__;
  assign new_new_n263__ = new_new_n161__ & new_new_n262__;
  assign new_new_n264__ = ~pi26 & ~pi29;
  assign new_new_n265__ = new_new_n230__ & new_new_n264__;
  assign new_new_n266__ = new_new_n146__ & new_new_n265__;
  assign new_new_n267__ = new_new_n75__ & new_new_n165__;
  assign new_new_n268__ = pi26 & new_new_n224__;
  assign new_new_n269__ = pi23 & new_new_n133__;
  assign new_new_n270__ = new_new_n268__ & new_new_n269__;
  assign new_new_n271__ = new_new_n135__ & new_new_n217__;
  assign new_new_n272__ = pi24 & new_new_n74__;
  assign new_new_n273__ = pi23 & new_new_n165__;
  assign new_new_n274__ = new_new_n272__ & new_new_n273__;
  assign new_new_n275__ = ~new_new_n271__ & ~new_new_n274__;
  assign new_new_n276__ = new_new_n146__ & new_new_n225__;
  assign new_new_n277__ = new_new_n137__ & new_new_n142__;
  assign new_new_n278__ = ~pi23 & new_new_n89__;
  assign new_new_n279__ = ~new_new_n141__ & new_new_n278__;
  assign new_new_n280__ = new_new_n224__ & new_new_n279__;
  assign new_new_n281__ = ~new_new_n277__ & ~new_new_n280__;
  assign new_new_n282__ = new_new_n85__ & new_new_n241__;
  assign new_new_n283__ = new_new_n81__ & new_new_n162__;
  assign new_new_n284__ = new_new_n180__ & new_new_n224__;
  assign new_new_n285__ = new_new_n134__ & new_new_n165__;
  assign new_new_n286__ = new_new_n133__ & new_new_n285__;
  assign new_new_n287__ = ~new_new_n282__ & ~new_new_n283__;
  assign new_new_n288__ = ~new_new_n284__ & new_new_n287__;
  assign new_new_n289__ = ~new_new_n270__ & ~new_new_n276__;
  assign new_new_n290__ = ~new_new_n286__ & new_new_n289__;
  assign new_new_n291__ = new_new_n275__ & new_new_n288__;
  assign new_new_n292__ = new_new_n281__ & new_new_n291__;
  assign new_new_n293__ = new_new_n290__ & new_new_n292__;
  assign new_new_n294__ = new_new_n261__ & ~new_new_n267__;
  assign new_new_n295__ = ~new_new_n263__ & ~new_new_n266__;
  assign new_new_n296__ = new_new_n294__ & new_new_n295__;
  assign new_new_n297__ = new_new_n293__ & new_new_n296__;
  assign new_new_n298__ = new_new_n87__ & new_new_n217__;
  assign new_new_n299__ = ~new_new_n104__ & new_new_n113__;
  assign new_new_n300__ = new_new_n224__ & new_new_n299__;
  assign new_new_n301__ = ~new_new_n298__ & ~new_new_n300__;
  assign new_new_n302__ = new_new_n87__ & new_new_n165__;
  assign new_new_n303__ = ~pi24 & ~pi25;
  assign new_new_n304__ = ~pi23 & ~pi26;
  assign new_new_n305__ = new_new_n237__ & new_new_n304__;
  assign new_new_n306__ = new_new_n303__ & new_new_n305__;
  assign new_new_n307__ = ~new_new_n302__ & ~new_new_n306__;
  assign new_new_n308__ = new_new_n217__ & new_new_n234__;
  assign new_new_n309__ = new_new_n85__ & new_new_n234__;
  assign new_new_n310__ = ~new_new_n78__ & ~new_new_n162__;
  assign new_new_n311__ = new_new_n234__ & ~new_new_n310__;
  assign new_new_n312__ = new_new_n75__ & new_new_n162__;
  assign new_new_n313__ = new_new_n135__ & new_new_n224__;
  assign new_new_n314__ = ~new_new_n312__ & ~new_new_n313__;
  assign new_new_n315__ = new_new_n75__ & new_new_n217__;
  assign new_new_n316__ = new_new_n114__ & new_new_n221__;
  assign new_new_n317__ = new_new_n142__ & new_new_n217__;
  assign new_new_n318__ = ~new_new_n316__ & ~new_new_n317__;
  assign new_new_n319__ = pi23 & new_new_n303__;
  assign new_new_n320__ = new_new_n97__ & new_new_n319__;
  assign new_new_n321__ = pi26 & new_new_n320__;
  assign new_new_n322__ = new_new_n217__ & new_new_n279__;
  assign new_new_n323__ = ~new_new_n321__ & ~new_new_n322__;
  assign new_new_n324__ = new_new_n314__ & ~new_new_n315__;
  assign new_new_n325__ = new_new_n323__ & new_new_n324__;
  assign new_new_n326__ = new_new_n318__ & new_new_n325__;
  assign new_new_n327__ = new_new_n118__ & new_new_n221__;
  assign new_new_n328__ = pi23 & new_new_n221__;
  assign new_new_n329__ = new_new_n272__ & new_new_n328__;
  assign new_new_n330__ = ~new_new_n327__ & ~new_new_n329__;
  assign new_new_n331__ = new_new_n89__ & new_new_n224__;
  assign new_new_n332__ = new_new_n90__ & new_new_n331__;
  assign new_new_n333__ = ~new_new_n129__ & ~new_new_n241__;
  assign new_new_n334__ = new_new_n191__ & ~new_new_n333__;
  assign new_new_n335__ = new_new_n81__ & new_new_n126__;
  assign new_new_n336__ = new_new_n81__ & new_new_n224__;
  assign new_new_n337__ = ~new_new_n335__ & ~new_new_n336__;
  assign new_new_n338__ = new_new_n91__ & new_new_n94__;
  assign new_new_n339__ = ~pi27 & new_new_n338__;
  assign new_new_n340__ = ~new_new_n332__ & ~new_new_n334__;
  assign new_new_n341__ = new_new_n337__ & ~new_new_n339__;
  assign new_new_n342__ = new_new_n340__ & new_new_n341__;
  assign new_new_n343__ = new_new_n330__ & new_new_n342__;
  assign new_new_n344__ = new_new_n114__ & new_new_n126__;
  assign new_new_n345__ = ~pi24 & new_new_n98__;
  assign new_new_n346__ = new_new_n273__ & new_new_n345__;
  assign new_new_n347__ = ~new_new_n344__ & ~new_new_n346__;
  assign new_new_n348__ = new_new_n273__ & ~new_new_n333__;
  assign new_new_n349__ = ~pi23 & new_new_n303__;
  assign new_new_n350__ = new_new_n268__ & new_new_n349__;
  assign new_new_n351__ = new_new_n78__ & new_new_n135__;
  assign new_new_n352__ = new_new_n190__ & new_new_n224__;
  assign new_new_n353__ = ~pi23 & new_new_n352__;
  assign new_new_n354__ = ~new_new_n351__ & ~new_new_n353__;
  assign new_new_n355__ = ~new_new_n78__ & ~new_new_n165__;
  assign new_new_n356__ = new_new_n100__ & ~new_new_n355__;
  assign new_new_n357__ = ~new_new_n308__ & ~new_new_n309__;
  assign new_new_n358__ = ~new_new_n258__ & new_new_n357__;
  assign new_new_n359__ = ~new_new_n311__ & ~new_new_n348__;
  assign new_new_n360__ = ~new_new_n350__ & ~new_new_n356__;
  assign new_new_n361__ = new_new_n359__ & new_new_n360__;
  assign new_new_n362__ = new_new_n301__ & new_new_n358__;
  assign new_new_n363__ = new_new_n307__ & new_new_n354__;
  assign new_new_n364__ = new_new_n362__ & new_new_n363__;
  assign new_new_n365__ = new_new_n256__ & new_new_n361__;
  assign new_new_n366__ = new_new_n347__ & new_new_n365__;
  assign new_new_n367__ = new_new_n326__ & new_new_n364__;
  assign new_new_n368__ = new_new_n343__ & new_new_n367__;
  assign new_new_n369__ = new_new_n366__ & new_new_n368__;
  assign new_new_n370__ = new_new_n297__ & new_new_n369__;
  assign new_new_n371__ = ~pi23 & new_new_n140__;
  assign new_new_n372__ = new_new_n268__ & new_new_n371__;
  assign new_new_n373__ = new_new_n114__ & new_new_n162__;
  assign new_new_n374__ = new_new_n91__ & new_new_n211__;
  assign new_new_n375__ = new_new_n163__ & new_new_n217__;
  assign new_new_n376__ = ~new_new_n374__ & ~new_new_n375__;
  assign new_new_n377__ = ~new_new_n372__ & new_new_n376__;
  assign new_new_n378__ = ~new_new_n373__ & new_new_n377__;
  assign new_new_n379__ = new_new_n87__ & new_new_n224__;
  assign new_new_n380__ = new_new_n142__ & new_new_n224__;
  assign new_new_n381__ = ~new_new_n379__ & ~new_new_n380__;
  assign new_new_n382__ = new_new_n133__ & new_new_n305__;
  assign new_new_n383__ = new_new_n100__ & new_new_n217__;
  assign new_new_n384__ = new_new_n165__ & new_new_n241__;
  assign new_new_n385__ = new_new_n105__ & new_new_n165__;
  assign new_new_n386__ = ~new_new_n384__ & ~new_new_n385__;
  assign new_new_n387__ = ~new_new_n383__ & new_new_n386__;
  assign new_new_n388__ = new_new_n78__ & new_new_n241__;
  assign new_new_n389__ = ~pi25 & ~new_new_n99__;
  assign new_new_n390__ = new_new_n285__ & ~new_new_n389__;
  assign new_new_n391__ = ~new_new_n388__ & ~new_new_n390__;
  assign new_new_n392__ = new_new_n381__ & ~new_new_n382__;
  assign new_new_n393__ = new_new_n387__ & new_new_n391__;
  assign new_new_n394__ = new_new_n392__ & new_new_n393__;
  assign new_new_n395__ = ~new_new_n246__ & ~new_new_n247__;
  assign new_new_n396__ = ~new_new_n248__ & ~new_new_n249__;
  assign new_new_n397__ = ~new_new_n250__ & ~new_new_n251__;
  assign new_new_n398__ = ~new_new_n252__ & ~new_new_n253__;
  assign new_new_n399__ = new_new_n397__ & new_new_n398__;
  assign new_new_n400__ = new_new_n395__ & new_new_n396__;
  assign new_new_n401__ = new_new_n399__ & new_new_n400__;
  assign new_new_n402__ = new_new_n216__ & new_new_n401__;
  assign new_new_n403__ = new_new_n228__ & new_new_n245__;
  assign new_new_n404__ = new_new_n378__ & new_new_n403__;
  assign new_new_n405__ = new_new_n394__ & new_new_n402__;
  assign new_new_n406__ = new_new_n404__ & new_new_n405__;
  assign new_new_n407__ = new_new_n370__ & new_new_n406__;
  assign new_new_n408__ = new_new_n83__ & new_new_n93__;
  assign new_new_n409__ = new_new_n102__ & new_new_n107__;
  assign new_new_n410__ = new_new_n121__ & new_new_n131__;
  assign new_new_n411__ = new_new_n409__ & new_new_n410__;
  assign new_new_n412__ = ~new_new_n124__ & new_new_n408__;
  assign new_new_n413__ = new_new_n411__ & new_new_n412__;
  assign new_new_n414__ = new_new_n116__ & new_new_n413__;
  assign new_new_n415__ = new_new_n159__ & new_new_n206__;
  assign new_new_n416__ = new_new_n414__ & new_new_n415__;
  assign new_new_n417__ = new_new_n187__ & new_new_n416__;
  assign new_new_n418__ = new_new_n407__ & new_new_n417__;
  assign new_new_n419__ = pi25 & ~new_new_n104__;
  assign new_new_n420__ = new_new_n265__ & ~new_new_n419__;
  assign new_new_n421__ = ~new_new_n97__ & ~new_new_n420__;
  assign new_new_n422__ = new_new_n98__ & ~new_new_n99__;
  assign new_new_n423__ = ~new_new_n190__ & ~new_new_n422__;
  assign new_new_n424__ = new_new_n132__ & ~new_new_n423__;
  assign new_new_n425__ = new_new_n78__ & new_new_n153__;
  assign new_new_n426__ = new_new_n78__ & new_new_n139__;
  assign new_new_n427__ = ~new_new_n141__ & new_new_n426__;
  assign new_new_n428__ = ~new_new_n425__ & ~new_new_n427__;
  assign new_new_n429__ = pi26 & ~new_new_n104__;
  assign new_new_n430__ = ~pi25 & ~pi26;
  assign new_new_n431__ = ~new_new_n99__ & new_new_n430__;
  assign new_new_n432__ = ~new_new_n429__ & ~new_new_n431__;
  assign new_new_n433__ = ~pi26 & ~new_new_n110__;
  assign new_new_n434__ = pi24 & ~new_new_n74__;
  assign new_new_n435__ = ~new_new_n433__ & new_new_n434__;
  assign new_new_n436__ = ~new_new_n432__ & ~new_new_n435__;
  assign new_new_n437__ = new_new_n72__ & ~new_new_n436__;
  assign new_new_n438__ = new_new_n72__ & new_new_n234__;
  assign new_new_n439__ = new_new_n85__ & new_new_n114__;
  assign new_new_n440__ = ~new_new_n438__ & ~new_new_n439__;
  assign new_new_n441__ = new_new_n78__ & new_new_n100__;
  assign new_new_n442__ = ~new_new_n103__ & ~new_new_n441__;
  assign new_new_n443__ = ~pi23 & new_new_n430__;
  assign new_new_n444__ = new_new_n72__ & new_new_n443__;
  assign new_new_n445__ = new_new_n81__ & new_new_n85__;
  assign new_new_n446__ = ~pi23 & ~new_new_n79__;
  assign new_new_n447__ = ~new_new_n86__ & ~new_new_n98__;
  assign new_new_n448__ = ~pi24 & ~new_new_n447__;
  assign new_new_n449__ = ~new_new_n272__ & ~new_new_n446__;
  assign new_new_n450__ = ~new_new_n448__ & new_new_n449__;
  assign new_new_n451__ = new_new_n78__ & ~new_new_n450__;
  assign new_new_n452__ = ~new_new_n444__ & ~new_new_n445__;
  assign new_new_n453__ = ~new_new_n451__ & new_new_n452__;
  assign new_new_n454__ = new_new_n116__ & new_new_n453__;
  assign new_new_n455__ = ~new_new_n160__ & ~new_new_n351__;
  assign new_new_n456__ = new_new_n121__ & new_new_n455__;
  assign new_new_n457__ = ~new_new_n155__ & new_new_n442__;
  assign new_new_n458__ = new_new_n456__ & new_new_n457__;
  assign new_new_n459__ = new_new_n428__ & new_new_n458__;
  assign new_new_n460__ = ~new_new_n437__ & new_new_n440__;
  assign new_new_n461__ = new_new_n459__ & new_new_n460__;
  assign new_new_n462__ = new_new_n454__ & new_new_n461__;
  assign new_new_n463__ = ~new_new_n76__ & ~new_new_n88__;
  assign new_new_n464__ = ~new_new_n424__ & new_new_n463__;
  assign new_new_n465__ = new_new_n462__ & new_new_n464__;
  assign new_new_n466__ = new_new_n421__ & new_new_n465__;
  assign new_new_n467__ = new_new_n72__ & new_new_n79__;
  assign new_new_n468__ = ~new_new_n147__ & ~new_new_n467__;
  assign new_new_n469__ = pi25 & ~new_new_n468__;
  assign new_new_n470__ = ~new_new_n109__ & new_new_n137__;
  assign new_new_n471__ = ~new_new_n469__ & ~new_new_n470__;
  assign new_new_n472__ = new_new_n78__ & new_new_n163__;
  assign new_new_n473__ = new_new_n78__ & new_new_n105__;
  assign new_new_n474__ = ~new_new_n472__ & ~new_new_n473__;
  assign new_new_n475__ = ~new_new_n207__ & ~new_new_n427__;
  assign new_new_n476__ = new_new_n91__ & new_new_n126__;
  assign new_new_n477__ = ~pi28 & new_new_n182__;
  assign new_new_n478__ = ~new_new_n439__ & ~new_new_n477__;
  assign new_new_n479__ = new_new_n114__ & new_new_n137__;
  assign new_new_n480__ = new_new_n78__ & new_new_n91__;
  assign new_new_n481__ = ~new_new_n479__ & ~new_new_n480__;
  assign new_new_n482__ = new_new_n78__ & new_new_n180__;
  assign new_new_n483__ = new_new_n89__ & new_new_n188__;
  assign new_new_n484__ = ~new_new_n482__ & ~new_new_n483__;
  assign new_new_n485__ = ~new_new_n425__ & ~new_new_n445__;
  assign new_new_n486__ = new_new_n484__ & new_new_n485__;
  assign new_new_n487__ = new_new_n126__ & ~new_new_n141__;
  assign new_new_n488__ = new_new_n278__ & new_new_n487__;
  assign new_new_n489__ = new_new_n126__ & new_new_n142__;
  assign new_new_n490__ = ~new_new_n488__ & ~new_new_n489__;
  assign new_new_n491__ = ~new_new_n476__ & new_new_n490__;
  assign new_new_n492__ = new_new_n478__ & new_new_n491__;
  assign new_new_n493__ = new_new_n481__ & new_new_n486__;
  assign new_new_n494__ = new_new_n492__ & new_new_n493__;
  assign new_new_n495__ = new_new_n135__ & new_new_n137__;
  assign new_new_n496__ = new_new_n78__ & new_new_n87__;
  assign new_new_n497__ = ~new_new_n108__ & ~new_new_n496__;
  assign new_new_n498__ = new_new_n121__ & ~new_new_n495__;
  assign new_new_n499__ = new_new_n474__ & new_new_n497__;
  assign new_new_n500__ = new_new_n498__ & new_new_n499__;
  assign new_new_n501__ = new_new_n475__ & new_new_n500__;
  assign new_new_n502__ = new_new_n471__ & new_new_n501__;
  assign new_new_n503__ = new_new_n494__ & new_new_n502__;
  assign new_new_n504__ = new_new_n86__ & ~new_new_n110__;
  assign new_new_n505__ = ~new_new_n345__ & ~new_new_n504__;
  assign new_new_n506__ = new_new_n221__ & ~new_new_n505__;
  assign new_new_n507__ = pi28 & new_new_n338__;
  assign new_new_n508__ = pi27 & new_new_n507__;
  assign new_new_n509__ = new_new_n95__ & new_new_n129__;
  assign new_new_n510__ = new_new_n180__ & new_new_n217__;
  assign new_new_n511__ = new_new_n153__ & new_new_n221__;
  assign new_new_n512__ = pi25 & ~new_new_n110__;
  assign new_new_n513__ = pi26 & ~new_new_n73__;
  assign new_new_n514__ = ~new_new_n512__ & ~new_new_n513__;
  assign new_new_n515__ = new_new_n95__ & ~new_new_n514__;
  assign new_new_n516__ = ~new_new_n511__ & ~new_new_n515__;
  assign new_new_n517__ = pi26 & new_new_n95__;
  assign new_new_n518__ = ~new_new_n257__ & ~new_new_n517__;
  assign new_new_n519__ = new_new_n223__ & ~new_new_n518__;
  assign new_new_n520__ = pi26 & new_new_n110__;
  assign new_new_n521__ = new_new_n221__ & ~new_new_n303__;
  assign new_new_n522__ = ~new_new_n512__ & new_new_n521__;
  assign new_new_n523__ = ~new_new_n520__ & new_new_n522__;
  assign new_new_n524__ = new_new_n217__ & ~new_new_n431__;
  assign new_new_n525__ = ~pi26 & new_new_n303__;
  assign new_new_n526__ = new_new_n95__ & new_new_n525__;
  assign new_new_n527__ = ~new_new_n524__ & ~new_new_n526__;
  assign new_new_n528__ = ~new_new_n106__ & ~new_new_n259__;
  assign new_new_n529__ = ~new_new_n509__ & ~new_new_n510__;
  assign new_new_n530__ = new_new_n528__ & new_new_n529__;
  assign new_new_n531__ = ~new_new_n143__ & new_new_n527__;
  assign new_new_n532__ = new_new_n530__ & new_new_n531__;
  assign new_new_n533__ = ~new_new_n506__ & ~new_new_n508__;
  assign new_new_n534__ = ~new_new_n519__ & ~new_new_n523__;
  assign new_new_n535__ = new_new_n533__ & new_new_n534__;
  assign new_new_n536__ = new_new_n516__ & new_new_n532__;
  assign new_new_n537__ = new_new_n535__ & new_new_n536__;
  assign new_new_n538__ = ~new_new_n74__ & ~new_new_n77__;
  assign new_new_n539__ = new_new_n74__ & ~new_new_n84__;
  assign new_new_n540__ = new_new_n161__ & ~new_new_n538__;
  assign new_new_n541__ = ~new_new_n539__ & new_new_n540__;
  assign new_new_n542__ = ~new_new_n240__ & ~new_new_n276__;
  assign new_new_n543__ = ~new_new_n226__ & ~new_new_n284__;
  assign new_new_n544__ = new_new_n221__ & new_new_n513__;
  assign new_new_n545__ = ~new_new_n331__ & ~new_new_n544__;
  assign new_new_n546__ = pi25 & ~new_new_n545__;
  assign new_new_n547__ = new_new_n97__ & new_new_n430__;
  assign new_new_n548__ = ~new_new_n268__ & ~new_new_n305__;
  assign new_new_n549__ = pi24 & ~new_new_n548__;
  assign new_new_n550__ = ~new_new_n74__ & ~new_new_n430__;
  assign new_new_n551__ = ~new_new_n128__ & ~new_new_n134__;
  assign new_new_n552__ = new_new_n237__ & new_new_n551__;
  assign new_new_n553__ = new_new_n550__ & new_new_n552__;
  assign new_new_n554__ = ~new_new_n549__ & ~new_new_n553__;
  assign new_new_n555__ = ~pi25 & new_new_n134__;
  assign new_new_n556__ = ~new_new_n139__ & ~new_new_n555__;
  assign new_new_n557__ = new_new_n237__ & ~new_new_n556__;
  assign new_new_n558__ = ~pi25 & new_new_n237__;
  assign new_new_n559__ = ~new_new_n268__ & ~new_new_n558__;
  assign new_new_n560__ = ~pi24 & ~new_new_n152__;
  assign new_new_n561__ = ~new_new_n559__ & new_new_n560__;
  assign new_new_n562__ = ~new_new_n557__ & ~new_new_n561__;
  assign new_new_n563__ = new_new_n239__ & ~new_new_n547__;
  assign new_new_n564__ = new_new_n554__ & new_new_n563__;
  assign new_new_n565__ = new_new_n562__ & new_new_n564__;
  assign new_new_n566__ = new_new_n86__ & new_new_n122__;
  assign new_new_n567__ = ~new_new_n353__ & ~new_new_n380__;
  assign new_new_n568__ = ~new_new_n222__ & ~new_new_n332__;
  assign new_new_n569__ = ~new_new_n541__ & ~new_new_n566__;
  assign new_new_n570__ = new_new_n568__ & new_new_n569__;
  assign new_new_n571__ = new_new_n542__ & new_new_n543__;
  assign new_new_n572__ = ~new_new_n546__ & new_new_n567__;
  assign new_new_n573__ = new_new_n571__ & new_new_n572__;
  assign new_new_n574__ = new_new_n570__ & new_new_n573__;
  assign new_new_n575__ = new_new_n565__ & new_new_n574__;
  assign new_new_n576__ = ~new_new_n164__ & new_new_n178__;
  assign new_new_n577__ = new_new_n537__ & new_new_n576__;
  assign new_new_n578__ = new_new_n575__ & new_new_n577__;
  assign new_new_n579__ = new_new_n131__ & ~new_new_n160__;
  assign new_new_n580__ = ~new_new_n424__ & new_new_n579__;
  assign new_new_n581__ = new_new_n206__ & new_new_n580__;
  assign new_new_n582__ = new_new_n503__ & new_new_n581__;
  assign new_new_n583__ = new_new_n578__ & new_new_n582__;
  assign new_new_n584__ = new_new_n97__ & new_new_n241__;
  assign new_new_n585__ = new_new_n211__ & new_new_n234__;
  assign new_new_n586__ = new_new_n100__ & new_new_n137__;
  assign new_new_n587__ = pi25 & new_new_n211__;
  assign new_new_n588__ = new_new_n139__ & new_new_n587__;
  assign new_new_n589__ = ~new_new_n586__ & ~new_new_n588__;
  assign new_new_n590__ = new_new_n67__ & new_new_n118__;
  assign new_new_n591__ = new_new_n125__ & new_new_n590__;
  assign new_new_n592__ = ~new_new_n495__ & ~new_new_n591__;
  assign new_new_n593__ = ~new_new_n92__ & ~new_new_n106__;
  assign new_new_n594__ = ~pi23 & new_new_n211__;
  assign new_new_n595__ = new_new_n190__ & new_new_n594__;
  assign new_new_n596__ = ~new_new_n82__ & ~new_new_n351__;
  assign new_new_n597__ = new_new_n180__ & new_new_n221__;
  assign new_new_n598__ = ~new_new_n163__ & ~new_new_n241__;
  assign new_new_n599__ = new_new_n85__ & ~new_new_n598__;
  assign new_new_n600__ = new_new_n75__ & new_new_n211__;
  assign new_new_n601__ = ~new_new_n508__ & ~new_new_n600__;
  assign new_new_n602__ = new_new_n142__ & new_new_n211__;
  assign new_new_n603__ = new_new_n137__ & new_new_n234__;
  assign new_new_n604__ = new_new_n100__ & new_new_n211__;
  assign new_new_n605__ = ~new_new_n603__ & ~new_new_n604__;
  assign new_new_n606__ = new_new_n117__ & new_new_n594__;
  assign new_new_n607__ = ~pi25 & new_new_n606__;
  assign new_new_n608__ = ~new_new_n115__ & ~new_new_n607__;
  assign new_new_n609__ = ~new_new_n259__ & new_new_n608__;
  assign new_new_n610__ = ~new_new_n249__ & ~new_new_n597__;
  assign new_new_n611__ = new_new_n593__ & new_new_n610__;
  assign new_new_n612__ = ~new_new_n595__ & new_new_n596__;
  assign new_new_n613__ = ~new_new_n599__ & ~new_new_n602__;
  assign new_new_n614__ = new_new_n605__ & new_new_n613__;
  assign new_new_n615__ = new_new_n611__ & new_new_n612__;
  assign new_new_n616__ = ~new_new_n373__ & new_new_n589__;
  assign new_new_n617__ = new_new_n592__ & new_new_n616__;
  assign new_new_n618__ = new_new_n614__ & new_new_n615__;
  assign new_new_n619__ = new_new_n601__ & new_new_n618__;
  assign new_new_n620__ = new_new_n609__ & new_new_n617__;
  assign new_new_n621__ = new_new_n619__ & new_new_n620__;
  assign new_new_n622__ = new_new_n210__ & ~new_new_n309__;
  assign new_new_n623__ = ~new_new_n388__ & ~new_new_n509__;
  assign new_new_n624__ = new_new_n137__ & new_new_n241__;
  assign new_new_n625__ = ~new_new_n252__ & ~new_new_n624__;
  assign new_new_n626__ = ~new_new_n266__ & new_new_n625__;
  assign new_new_n627__ = new_new_n623__ & new_new_n626__;
  assign new_new_n628__ = ~new_new_n263__ & ~new_new_n283__;
  assign new_new_n629__ = ~new_new_n207__ & ~new_new_n312__;
  assign new_new_n630__ = pi25 & new_new_n606__;
  assign new_new_n631__ = new_new_n272__ & new_new_n594__;
  assign new_new_n632__ = new_new_n105__ & new_new_n211__;
  assign new_new_n633__ = ~new_new_n631__ & ~new_new_n632__;
  assign new_new_n634__ = new_new_n135__ & new_new_n211__;
  assign new_new_n635__ = new_new_n223__ & new_new_n517__;
  assign new_new_n636__ = ~new_new_n634__ & ~new_new_n635__;
  assign new_new_n637__ = new_new_n87__ & new_new_n211__;
  assign new_new_n638__ = ~new_new_n585__ & ~new_new_n637__;
  assign new_new_n639__ = ~new_new_n277__ & new_new_n638__;
  assign new_new_n640__ = ~new_new_n311__ & new_new_n442__;
  assign new_new_n641__ = new_new_n629__ & new_new_n640__;
  assign new_new_n642__ = new_new_n622__ & new_new_n639__;
  assign new_new_n643__ = new_new_n628__ & ~new_new_n630__;
  assign new_new_n644__ = new_new_n633__ & new_new_n636__;
  assign new_new_n645__ = new_new_n643__ & new_new_n644__;
  assign new_new_n646__ = new_new_n641__ & new_new_n642__;
  assign new_new_n647__ = new_new_n516__ & new_new_n627__;
  assign new_new_n648__ = new_new_n646__ & new_new_n647__;
  assign new_new_n649__ = new_new_n159__ & new_new_n645__;
  assign new_new_n650__ = new_new_n648__ & new_new_n649__;
  assign new_new_n651__ = new_new_n621__ & new_new_n650__;
  assign new_new_n652__ = new_new_n152__ & new_new_n523__;
  assign new_new_n653__ = ~new_new_n104__ & new_new_n165__;
  assign new_new_n654__ = ~new_new_n122__ & ~new_new_n653__;
  assign new_new_n655__ = new_new_n430__ & ~new_new_n654__;
  assign new_new_n656__ = new_new_n75__ & new_new_n97__;
  assign new_new_n657__ = new_new_n91__ & new_new_n165__;
  assign new_new_n658__ = new_new_n81__ & new_new_n211__;
  assign new_new_n659__ = ~new_new_n657__ & ~new_new_n658__;
  assign new_new_n660__ = ~new_new_n101__ & ~new_new_n213__;
  assign new_new_n661__ = ~new_new_n229__ & ~new_new_n246__;
  assign new_new_n662__ = ~new_new_n656__ & new_new_n661__;
  assign new_new_n663__ = ~new_new_n321__ & new_new_n660__;
  assign new_new_n664__ = new_new_n659__ & new_new_n663__;
  assign new_new_n665__ = ~new_new_n124__ & new_new_n662__;
  assign new_new_n666__ = ~new_new_n506__ & new_new_n665__;
  assign new_new_n667__ = new_new_n664__ & new_new_n666__;
  assign new_new_n668__ = ~pi24 & new_new_n523__;
  assign new_new_n669__ = ~new_new_n335__ & ~new_new_n668__;
  assign new_new_n670__ = new_new_n211__ & new_new_n525__;
  assign new_new_n671__ = new_new_n129__ & new_new_n221__;
  assign new_new_n672__ = ~new_new_n251__ & ~new_new_n671__;
  assign new_new_n673__ = new_new_n223__ & new_new_n257__;
  assign new_new_n674__ = ~new_new_n510__ & ~new_new_n673__;
  assign new_new_n675__ = ~pi26 & new_new_n320__;
  assign new_new_n676__ = new_new_n97__ & new_new_n114__;
  assign new_new_n677__ = ~new_new_n108__ & ~new_new_n584__;
  assign new_new_n678__ = ~new_new_n670__ & new_new_n677__;
  assign new_new_n679__ = new_new_n121__ & new_new_n527__;
  assign new_new_n680__ = new_new_n672__ & ~new_new_n675__;
  assign new_new_n681__ = new_new_n679__ & new_new_n680__;
  assign new_new_n682__ = ~new_new_n344__ & new_new_n678__;
  assign new_new_n683__ = ~new_new_n655__ & new_new_n674__;
  assign new_new_n684__ = ~new_new_n676__ & new_new_n683__;
  assign new_new_n685__ = new_new_n681__ & new_new_n682__;
  assign new_new_n686__ = new_new_n256__ & ~new_new_n652__;
  assign new_new_n687__ = new_new_n685__ & new_new_n686__;
  assign new_new_n688__ = new_new_n669__ & new_new_n684__;
  assign new_new_n689__ = new_new_n687__ & new_new_n688__;
  assign new_new_n690__ = new_new_n667__ & new_new_n689__;
  assign new_new_n691__ = new_new_n651__ & new_new_n690__;
  assign new_new_n692__ = new_new_n81__ & new_new_n95__;
  assign new_new_n693__ = new_new_n100__ & new_new_n165__;
  assign new_new_n694__ = new_new_n129__ & new_new_n237__;
  assign new_new_n695__ = ~new_new_n693__ & ~new_new_n694__;
  assign new_new_n696__ = new_new_n152__ & new_new_n467__;
  assign new_new_n697__ = ~new_new_n235__ & ~new_new_n696__;
  assign new_new_n698__ = new_new_n95__ & new_new_n163__;
  assign new_new_n699__ = ~new_new_n209__ & ~new_new_n698__;
  assign new_new_n700__ = new_new_n135__ & new_new_n237__;
  assign new_new_n701__ = new_new_n118__ & new_new_n237__;
  assign new_new_n702__ = ~new_new_n700__ & ~new_new_n701__;
  assign new_new_n703__ = ~new_new_n270__ & ~new_new_n692__;
  assign new_new_n704__ = ~new_new_n477__ & new_new_n695__;
  assign new_new_n705__ = new_new_n699__ & new_new_n702__;
  assign new_new_n706__ = new_new_n704__ & new_new_n705__;
  assign new_new_n707__ = new_new_n697__ & new_new_n703__;
  assign new_new_n708__ = new_new_n706__ & new_new_n707__;
  assign new_new_n709__ = ~new_new_n277__ & ~new_new_n508__;
  assign new_new_n710__ = ~new_new_n229__ & ~new_new_n267__;
  assign new_new_n711__ = ~new_new_n138__ & ~new_new_n511__;
  assign new_new_n712__ = ~new_new_n603__ & new_new_n711__;
  assign new_new_n713__ = new_new_n710__ & new_new_n712__;
  assign new_new_n714__ = new_new_n709__ & new_new_n713__;
  assign new_new_n715__ = new_new_n72__ & new_new_n241__;
  assign new_new_n716__ = ~new_new_n350__ & ~new_new_n715__;
  assign new_new_n717__ = new_new_n100__ & new_new_n169__;
  assign new_new_n718__ = new_new_n67__ & new_new_n94__;
  assign new_new_n719__ = new_new_n279__ & new_new_n718__;
  assign new_new_n720__ = ~new_new_n717__ & ~new_new_n719__;
  assign new_new_n721__ = new_new_n140__ & new_new_n285__;
  assign new_new_n722__ = ~new_new_n597__ & ~new_new_n721__;
  assign new_new_n723__ = new_new_n81__ & new_new_n97__;
  assign new_new_n724__ = new_new_n85__ & new_new_n105__;
  assign new_new_n725__ = ~new_new_n723__ & ~new_new_n724__;
  assign new_new_n726__ = ~new_new_n143__ & ~new_new_n315__;
  assign new_new_n727__ = new_new_n725__ & new_new_n726__;
  assign new_new_n728__ = new_new_n722__ & new_new_n727__;
  assign new_new_n729__ = new_new_n75__ & new_new_n169__;
  assign new_new_n730__ = ~new_new_n92__ & ~new_new_n729__;
  assign new_new_n731__ = new_new_n118__ & new_new_n151__;
  assign new_new_n732__ = ~pi30 & new_new_n731__;
  assign new_new_n733__ = ~new_new_n82__ & ~new_new_n732__;
  assign new_new_n734__ = ~new_new_n254__ & ~new_new_n353__;
  assign new_new_n735__ = ~new_new_n351__ & ~new_new_n673__;
  assign new_new_n736__ = ~new_new_n119__ & ~new_new_n383__;
  assign new_new_n737__ = ~new_new_n637__ & new_new_n736__;
  assign new_new_n738__ = new_new_n730__ & new_new_n737__;
  assign new_new_n739__ = ~new_new_n316__ & new_new_n733__;
  assign new_new_n740__ = new_new_n735__ & new_new_n739__;
  assign new_new_n741__ = new_new_n734__ & new_new_n738__;
  assign new_new_n742__ = new_new_n740__ & new_new_n741__;
  assign new_new_n743__ = ~new_new_n189__ & ~new_new_n202__;
  assign new_new_n744__ = ~new_new_n222__ & ~new_new_n372__;
  assign new_new_n745__ = ~new_new_n496__ & ~new_new_n510__;
  assign new_new_n746__ = new_new_n151__ & new_new_n180__;
  assign new_new_n747__ = ~pi30 & new_new_n746__;
  assign new_new_n748__ = ~new_new_n260__ & ~new_new_n747__;
  assign new_new_n749__ = new_new_n72__ & new_new_n87__;
  assign new_new_n750__ = ~new_new_n208__ & ~new_new_n495__;
  assign new_new_n751__ = ~new_new_n749__ & new_new_n750__;
  assign new_new_n752__ = ~new_new_n97__ & ~new_new_n237__;
  assign new_new_n753__ = new_new_n100__ & ~new_new_n752__;
  assign new_new_n754__ = ~new_new_n313__ & new_new_n745__;
  assign new_new_n755__ = ~new_new_n753__ & new_new_n754__;
  assign new_new_n756__ = new_new_n716__ & new_new_n720__;
  assign new_new_n757__ = new_new_n743__ & new_new_n744__;
  assign new_new_n758__ = new_new_n748__ & new_new_n751__;
  assign new_new_n759__ = new_new_n757__ & new_new_n758__;
  assign new_new_n760__ = new_new_n755__ & new_new_n756__;
  assign new_new_n761__ = new_new_n759__ & new_new_n760__;
  assign new_new_n762__ = new_new_n728__ & new_new_n761__;
  assign new_new_n763__ = new_new_n742__ & new_new_n762__;
  assign new_new_n764__ = ~new_new_n96__ & new_new_n542__;
  assign new_new_n765__ = ~new_new_n71__ & ~new_new_n161__;
  assign new_new_n766__ = new_new_n84__ & ~new_new_n765__;
  assign new_new_n767__ = new_new_n163__ & new_new_n766__;
  assign new_new_n768__ = new_new_n97__ & new_new_n180__;
  assign new_new_n769__ = ~new_new_n427__ & ~new_new_n768__;
  assign new_new_n770__ = ~new_new_n329__ & ~new_new_n767__;
  assign new_new_n771__ = new_new_n769__ & new_new_n770__;
  assign new_new_n772__ = new_new_n169__ & new_new_n241__;
  assign new_new_n773__ = ~new_new_n211__ & ~new_new_n718__;
  assign new_new_n774__ = new_new_n135__ & ~new_new_n773__;
  assign new_new_n775__ = ~new_new_n772__ & ~new_new_n774__;
  assign new_new_n776__ = new_new_n75__ & new_new_n137__;
  assign new_new_n777__ = ~new_new_n106__ & ~new_new_n776__;
  assign new_new_n778__ = new_new_n87__ & new_new_n237__;
  assign new_new_n779__ = ~new_new_n604__ & ~new_new_n778__;
  assign new_new_n780__ = new_new_n117__ & new_new_n718__;
  assign new_new_n781__ = new_new_n112__ & new_new_n780__;
  assign new_new_n782__ = ~new_new_n247__ & ~new_new_n781__;
  assign new_new_n783__ = new_new_n163__ & new_new_n169__;
  assign new_new_n784__ = ~new_new_n282__ & ~new_new_n335__;
  assign new_new_n785__ = new_new_n180__ & new_new_n718__;
  assign new_new_n786__ = ~new_new_n585__ & ~new_new_n785__;
  assign new_new_n787__ = ~new_new_n207__ & ~new_new_n388__;
  assign new_new_n788__ = ~new_new_n656__ & new_new_n787__;
  assign new_new_n789__ = new_new_n786__ & new_new_n788__;
  assign new_new_n790__ = ~new_new_n263__ & ~new_new_n783__;
  assign new_new_n791__ = new_new_n777__ & new_new_n779__;
  assign new_new_n792__ = new_new_n784__ & new_new_n791__;
  assign new_new_n793__ = new_new_n775__ & new_new_n790__;
  assign new_new_n794__ = new_new_n782__ & new_new_n793__;
  assign new_new_n795__ = new_new_n764__ & new_new_n792__;
  assign new_new_n796__ = new_new_n771__ & new_new_n789__;
  assign new_new_n797__ = new_new_n795__ & new_new_n796__;
  assign new_new_n798__ = new_new_n794__ & new_new_n797__;
  assign new_new_n799__ = ~new_new_n196__ & ~new_new_n584__;
  assign new_new_n800__ = new_new_n112__ & new_new_n169__;
  assign new_new_n801__ = ~new_new_n99__ & ~new_new_n104__;
  assign new_new_n802__ = ~new_new_n90__ & new_new_n162__;
  assign new_new_n803__ = new_new_n801__ & new_new_n802__;
  assign new_new_n804__ = ~new_new_n800__ & ~new_new_n803__;
  assign new_new_n805__ = pi26 & ~new_new_n804__;
  assign new_new_n806__ = new_new_n799__ & ~new_new_n805__;
  assign new_new_n807__ = new_new_n114__ & new_new_n230__;
  assign new_new_n808__ = new_new_n133__ & new_new_n328__;
  assign new_new_n809__ = ~new_new_n520__ & new_new_n808__;
  assign new_new_n810__ = ~new_new_n658__ & ~new_new_n809__;
  assign new_new_n811__ = new_new_n135__ & new_new_n221__;
  assign new_new_n812__ = new_new_n86__ & new_new_n165__;
  assign new_new_n813__ = ~new_new_n483__ & ~new_new_n602__;
  assign new_new_n814__ = pi29 & new_new_n84__;
  assign new_new_n815__ = new_new_n135__ & new_new_n814__;
  assign new_new_n816__ = ~pi30 & new_new_n815__;
  assign new_new_n817__ = ~new_new_n103__ & ~new_new_n425__;
  assign new_new_n818__ = ~new_new_n811__ & ~new_new_n812__;
  assign new_new_n819__ = new_new_n817__ & new_new_n818__;
  assign new_new_n820__ = ~new_new_n816__ & new_new_n819__;
  assign new_new_n821__ = new_new_n633__ & ~new_new_n807__;
  assign new_new_n822__ = new_new_n813__ & new_new_n821__;
  assign new_new_n823__ = new_new_n810__ & new_new_n820__;
  assign new_new_n824__ = new_new_n822__ & new_new_n823__;
  assign new_new_n825__ = new_new_n806__ & new_new_n824__;
  assign new_new_n826__ = new_new_n85__ & new_new_n180__;
  assign new_new_n827__ = ~new_new_n283__ & ~new_new_n826__;
  assign new_new_n828__ = new_new_n349__ & new_new_n517__;
  assign new_new_n829__ = new_new_n129__ & new_new_n169__;
  assign new_new_n830__ = ~new_new_n317__ & ~new_new_n509__;
  assign new_new_n831__ = ~new_new_n829__ & new_new_n830__;
  assign new_new_n832__ = ~new_new_n136__ & new_new_n827__;
  assign new_new_n833__ = ~new_new_n828__ & new_new_n832__;
  assign new_new_n834__ = new_new_n831__ & new_new_n833__;
  assign new_new_n835__ = new_new_n142__ & new_new_n718__;
  assign new_new_n836__ = ~new_new_n657__ & ~new_new_n835__;
  assign new_new_n837__ = new_new_n95__ & new_new_n114__;
  assign new_new_n838__ = new_new_n100__ & new_new_n718__;
  assign new_new_n839__ = ~new_new_n218__ & ~new_new_n838__;
  assign new_new_n840__ = ~new_new_n327__ & ~new_new_n438__;
  assign new_new_n841__ = new_new_n839__ & new_new_n840__;
  assign new_new_n842__ = new_new_n72__ & new_new_n142__;
  assign new_new_n843__ = new_new_n234__ & new_new_n237__;
  assign new_new_n844__ = ~new_new_n842__ & ~new_new_n843__;
  assign new_new_n845__ = new_new_n237__ & new_new_n241__;
  assign new_new_n846__ = new_new_n234__ & new_new_n718__;
  assign new_new_n847__ = ~new_new_n127__ & ~new_new_n846__;
  assign new_new_n848__ = ~new_new_n271__ & ~new_new_n845__;
  assign new_new_n849__ = new_new_n847__ & new_new_n848__;
  assign new_new_n850__ = ~new_new_n322__ & ~new_new_n479__;
  assign new_new_n851__ = new_new_n135__ & new_new_n169__;
  assign new_new_n852__ = ~new_new_n150__ & ~new_new_n851__;
  assign new_new_n853__ = new_new_n169__ & new_new_n234__;
  assign new_new_n854__ = ~new_new_n213__ & ~new_new_n374__;
  assign new_new_n855__ = ~new_new_n853__ & new_new_n854__;
  assign new_new_n856__ = new_new_n836__ & new_new_n855__;
  assign new_new_n857__ = ~new_new_n837__ & new_new_n844__;
  assign new_new_n858__ = new_new_n849__ & new_new_n852__;
  assign new_new_n859__ = new_new_n857__ & new_new_n858__;
  assign new_new_n860__ = new_new_n850__ & new_new_n856__;
  assign new_new_n861__ = new_new_n859__ & new_new_n860__;
  assign new_new_n862__ = new_new_n708__ & new_new_n714__;
  assign new_new_n863__ = new_new_n834__ & new_new_n841__;
  assign new_new_n864__ = new_new_n862__ & new_new_n863__;
  assign new_new_n865__ = new_new_n861__ & new_new_n864__;
  assign new_new_n866__ = new_new_n798__ & new_new_n825__;
  assign new_new_n867__ = new_new_n865__ & new_new_n866__;
  assign new_new_n868__ = new_new_n763__ & new_new_n867__;
  assign new_new_n869__ = new_new_n72__ & new_new_n279__;
  assign new_new_n870__ = ~new_new_n776__ & ~new_new_n869__;
  assign new_new_n871__ = new_new_n223__ & new_new_n265__;
  assign new_new_n872__ = ~new_new_n566__ & ~new_new_n871__;
  assign new_new_n873__ = ~new_new_n389__ & ~new_new_n419__;
  assign new_new_n874__ = new_new_n547__ & new_new_n873__;
  assign new_new_n875__ = new_new_n105__ & new_new_n237__;
  assign new_new_n876__ = ~new_new_n842__ & ~new_new_n875__;
  assign new_new_n877__ = new_new_n151__ & new_new_n163__;
  assign new_new_n878__ = ~pi30 & new_new_n877__;
  assign new_new_n879__ = new_new_n223__ & new_new_n718__;
  assign new_new_n880__ = ~new_new_n80__ & new_new_n211__;
  assign new_new_n881__ = ~new_new_n389__ & new_new_n880__;
  assign new_new_n882__ = ~new_new_n879__ & ~new_new_n881__;
  assign new_new_n883__ = ~pi26 & ~new_new_n882__;
  assign new_new_n884__ = new_new_n142__ & new_new_n237__;
  assign new_new_n885__ = ~new_new_n749__ & ~new_new_n884__;
  assign new_new_n886__ = ~new_new_n637__ & ~new_new_n878__;
  assign new_new_n887__ = ~new_new_n607__ & new_new_n886__;
  assign new_new_n888__ = new_new_n885__ & new_new_n887__;
  assign new_new_n889__ = ~new_new_n883__ & new_new_n888__;
  assign new_new_n890__ = new_new_n85__ & new_new_n91__;
  assign new_new_n891__ = new_new_n674__ & ~new_new_n890__;
  assign new_new_n892__ = pi23 & ~pi26;
  assign new_new_n893__ = new_new_n72__ & new_new_n145__;
  assign new_new_n894__ = new_new_n892__ & new_new_n893__;
  assign new_new_n895__ = pi26 & new_new_n523__;
  assign new_new_n896__ = new_new_n81__ & new_new_n137__;
  assign new_new_n897__ = ~new_new_n747__ & ~new_new_n768__;
  assign new_new_n898__ = ~new_new_n723__ & ~new_new_n896__;
  assign new_new_n899__ = ~new_new_n588__ & new_new_n898__;
  assign new_new_n900__ = ~new_new_n874__ & ~new_new_n894__;
  assign new_new_n901__ = new_new_n899__ & new_new_n900__;
  assign new_new_n902__ = new_new_n870__ & new_new_n872__;
  assign new_new_n903__ = new_new_n876__ & new_new_n897__;
  assign new_new_n904__ = new_new_n902__ & new_new_n903__;
  assign new_new_n905__ = new_new_n891__ & new_new_n901__;
  assign new_new_n906__ = ~new_new_n895__ & new_new_n905__;
  assign new_new_n907__ = new_new_n904__ & new_new_n906__;
  assign new_new_n908__ = new_new_n494__ & new_new_n889__;
  assign new_new_n909__ = new_new_n907__ & new_new_n908__;
  assign new_new_n910__ = new_new_n407__ & new_new_n909__;
  assign new_new_n911__ = ~new_new_n691__ & new_new_n910__;
  assign new_new_n912__ = ~new_new_n583__ & new_new_n911__;
  assign new_new_n913__ = ~new_new_n251__ & ~new_new_n673__;
  assign new_new_n914__ = ~new_new_n238__ & ~new_new_n248__;
  assign new_new_n915__ = ~new_new_n441__ & ~new_new_n624__;
  assign new_new_n916__ = new_new_n914__ & new_new_n915__;
  assign new_new_n917__ = ~new_new_n97__ & ~new_new_n211__;
  assign new_new_n918__ = new_new_n153__ & ~new_new_n917__;
  assign new_new_n919__ = new_new_n162__ & new_new_n279__;
  assign new_new_n920__ = ~pi25 & new_new_n97__;
  assign new_new_n921__ = new_new_n278__ & new_new_n920__;
  assign new_new_n922__ = ~new_new_n445__ & ~new_new_n843__;
  assign new_new_n923__ = ~new_new_n918__ & new_new_n922__;
  assign new_new_n924__ = ~new_new_n919__ & ~new_new_n921__;
  assign new_new_n925__ = new_new_n923__ & new_new_n924__;
  assign new_new_n926__ = new_new_n913__ & new_new_n916__;
  assign new_new_n927__ = new_new_n925__ & new_new_n926__;
  assign new_new_n928__ = ~new_new_n332__ & ~new_new_n344__;
  assign new_new_n929__ = ~new_new_n130__ & ~new_new_n168__;
  assign new_new_n930__ = ~new_new_n313__ & ~new_new_n826__;
  assign new_new_n931__ = new_new_n929__ & new_new_n930__;
  assign new_new_n932__ = ~new_new_n427__ & new_new_n931__;
  assign new_new_n933__ = new_new_n162__ & new_new_n234__;
  assign new_new_n934__ = ~new_new_n283__ & ~new_new_n933__;
  assign new_new_n935__ = new_new_n114__ & new_new_n237__;
  assign new_new_n936__ = ~new_new_n717__ & ~new_new_n935__;
  assign new_new_n937__ = new_new_n75__ & new_new_n237__;
  assign new_new_n938__ = ~new_new_n878__ & ~new_new_n937__;
  assign new_new_n939__ = new_new_n269__ & new_new_n517__;
  assign new_new_n940__ = new_new_n87__ & new_new_n162__;
  assign new_new_n941__ = ~new_new_n871__ & ~new_new_n940__;
  assign new_new_n942__ = new_new_n129__ & new_new_n718__;
  assign new_new_n943__ = ~new_new_n148__ & ~new_new_n942__;
  assign new_new_n944__ = ~new_new_n602__ & ~new_new_n634__;
  assign new_new_n945__ = new_new_n85__ & new_new_n142__;
  assign new_new_n946__ = ~new_new_n300__ & ~new_new_n945__;
  assign new_new_n947__ = new_new_n81__ & new_new_n718__;
  assign new_new_n948__ = ~new_new_n253__ & ~new_new_n700__;
  assign new_new_n949__ = ~new_new_n947__ & new_new_n948__;
  assign new_new_n950__ = new_new_n163__ & new_new_n237__;
  assign new_new_n951__ = ~new_new_n127__ & ~new_new_n671__;
  assign new_new_n952__ = new_new_n142__ & new_new_n169__;
  assign new_new_n953__ = ~new_new_n106__ & ~new_new_n595__;
  assign new_new_n954__ = ~new_new_n108__ & ~new_new_n811__;
  assign new_new_n955__ = ~new_new_n321__ & new_new_n954__;
  assign new_new_n956__ = ~new_new_n952__ & new_new_n955__;
  assign new_new_n957__ = new_new_n953__ & new_new_n956__;
  assign new_new_n958__ = pi26 & new_new_n140__;
  assign new_new_n959__ = new_new_n201__ & new_new_n958__;
  assign new_new_n960__ = ~new_new_n150__ & ~new_new_n959__;
  assign new_new_n961__ = new_new_n80__ & new_new_n780__;
  assign new_new_n962__ = ~new_new_n635__ & ~new_new_n961__;
  assign new_new_n963__ = new_new_n91__ & new_new_n162__;
  assign new_new_n964__ = ~new_new_n270__ & ~new_new_n963__;
  assign new_new_n965__ = ~new_new_n229__ & ~new_new_n382__;
  assign new_new_n966__ = ~new_new_n82__ & ~new_new_n179__;
  assign new_new_n967__ = ~new_new_n785__ & ~new_new_n838__;
  assign new_new_n968__ = ~new_new_n346__ & ~new_new_n950__;
  assign new_new_n969__ = new_new_n951__ & new_new_n966__;
  assign new_new_n970__ = new_new_n967__ & new_new_n969__;
  assign new_new_n971__ = ~new_new_n254__ & new_new_n968__;
  assign new_new_n972__ = ~new_new_n837__ & new_new_n941__;
  assign new_new_n973__ = new_new_n943__ & new_new_n944__;
  assign new_new_n974__ = new_new_n946__ & new_new_n949__;
  assign new_new_n975__ = new_new_n960__ & new_new_n962__;
  assign new_new_n976__ = new_new_n964__ & new_new_n965__;
  assign new_new_n977__ = new_new_n975__ & new_new_n976__;
  assign new_new_n978__ = new_new_n973__ & new_new_n974__;
  assign new_new_n979__ = new_new_n971__ & new_new_n972__;
  assign new_new_n980__ = new_new_n970__ & new_new_n979__;
  assign new_new_n981__ = new_new_n977__ & new_new_n978__;
  assign new_new_n982__ = new_new_n957__ & new_new_n981__;
  assign new_new_n983__ = new_new_n980__ & new_new_n982__;
  assign new_new_n984__ = ~new_new_n380__ & ~new_new_n783__;
  assign new_new_n985__ = ~new_new_n566__ & ~new_new_n676__;
  assign new_new_n986__ = ~new_new_n138__ & new_new_n984__;
  assign new_new_n987__ = new_new_n478__ & new_new_n986__;
  assign new_new_n988__ = new_new_n985__ & new_new_n987__;
  assign new_new_n989__ = ~new_new_n390__ & ~new_new_n631__;
  assign new_new_n990__ = new_new_n169__ & new_new_n180__;
  assign new_new_n991__ = ~pi26 & new_new_n110__;
  assign new_new_n992__ = new_new_n140__ & new_new_n221__;
  assign new_new_n993__ = new_new_n991__ & new_new_n992__;
  assign new_new_n994__ = ~new_new_n778__ & ~new_new_n993__;
  assign new_new_n995__ = new_new_n153__ & new_new_n162__;
  assign new_new_n996__ = new_new_n72__ & new_new_n135__;
  assign new_new_n997__ = ~new_new_n298__ & ~new_new_n489__;
  assign new_new_n998__ = ~new_new_n472__ & ~new_new_n588__;
  assign new_new_n999__ = ~new_new_n155__ & ~new_new_n250__;
  assign new_new_n1000__ = ~new_new_n143__ & ~new_new_n164__;
  assign new_new_n1001__ = ~new_new_n200__ & new_new_n1000__;
  assign new_new_n1002__ = new_new_n262__ & ~new_new_n765__;
  assign new_new_n1003__ = new_new_n170__ & new_new_n272__;
  assign new_new_n1004__ = ~new_new_n166__ & ~new_new_n600__;
  assign new_new_n1005__ = ~new_new_n242__ & ~new_new_n1003__;
  assign new_new_n1006__ = new_new_n1004__ & new_new_n1005__;
  assign new_new_n1007__ = new_new_n78__ & new_new_n234__;
  assign new_new_n1008__ = new_new_n67__ & new_new_n338__;
  assign new_new_n1009__ = new_new_n371__ & new_new_n517__;
  assign new_new_n1010__ = ~new_new_n208__ & ~new_new_n1009__;
  assign new_new_n1011__ = ~new_new_n101__ & ~new_new_n103__;
  assign new_new_n1012__ = ~new_new_n271__ & ~new_new_n385__;
  assign new_new_n1013__ = ~new_new_n657__ & ~new_new_n1007__;
  assign new_new_n1014__ = new_new_n1012__ & new_new_n1013__;
  assign new_new_n1015__ = ~new_new_n280__ & new_new_n1011__;
  assign new_new_n1016__ = ~new_new_n1008__ & new_new_n1015__;
  assign new_new_n1017__ = new_new_n1010__ & new_new_n1014__;
  assign new_new_n1018__ = new_new_n1016__ & new_new_n1017__;
  assign new_new_n1019__ = new_new_n1006__ & new_new_n1018__;
  assign new_new_n1020__ = ~new_new_n249__ & ~new_new_n698__;
  assign new_new_n1021__ = ~new_new_n846__ & ~new_new_n995__;
  assign new_new_n1022__ = ~new_new_n996__ & new_new_n1021__;
  assign new_new_n1023__ = ~new_new_n835__ & new_new_n1020__;
  assign new_new_n1024__ = ~new_new_n1002__ & new_new_n1023__;
  assign new_new_n1025__ = new_new_n997__ & new_new_n1022__;
  assign new_new_n1026__ = new_new_n998__ & new_new_n999__;
  assign new_new_n1027__ = new_new_n1025__ & new_new_n1026__;
  assign new_new_n1028__ = new_new_n1001__ & new_new_n1024__;
  assign new_new_n1029__ = new_new_n1027__ & new_new_n1028__;
  assign new_new_n1030__ = new_new_n1019__ & new_new_n1029__;
  assign new_new_n1031__ = new_new_n163__ & new_new_n221__;
  assign new_new_n1032__ = ~new_new_n202__ & ~new_new_n1031__;
  assign new_new_n1033__ = new_new_n87__ & new_new_n718__;
  assign new_new_n1034__ = new_new_n75__ & new_new_n814__;
  assign new_new_n1035__ = ~pi30 & new_new_n1034__;
  assign new_new_n1036__ = ~new_new_n1033__ & ~new_new_n1035__;
  assign new_new_n1037__ = ~new_new_n693__ & ~new_new_n869__;
  assign new_new_n1038__ = ~new_new_n260__ & ~new_new_n488__;
  assign new_new_n1039__ = new_new_n1036__ & new_new_n1038__;
  assign new_new_n1040__ = new_new_n1037__ & new_new_n1039__;
  assign new_new_n1041__ = ~new_new_n482__ & ~new_new_n511__;
  assign new_new_n1042__ = ~new_new_n829__ & ~new_new_n990__;
  assign new_new_n1043__ = new_new_n1041__ & new_new_n1042__;
  assign new_new_n1044__ = ~new_new_n317__ & ~new_new_n353__;
  assign new_new_n1045__ = ~new_new_n894__ & new_new_n934__;
  assign new_new_n1046__ = ~new_new_n939__ & new_new_n1045__;
  assign new_new_n1047__ = new_new_n1043__ & new_new_n1044__;
  assign new_new_n1048__ = new_new_n542__ & new_new_n938__;
  assign new_new_n1049__ = new_new_n989__ & new_new_n994__;
  assign new_new_n1050__ = new_new_n1032__ & new_new_n1049__;
  assign new_new_n1051__ = new_new_n1047__ & new_new_n1048__;
  assign new_new_n1052__ = new_new_n928__ & new_new_n1046__;
  assign new_new_n1053__ = new_new_n932__ & new_new_n936__;
  assign new_new_n1054__ = new_new_n1052__ & new_new_n1053__;
  assign new_new_n1055__ = new_new_n1050__ & new_new_n1051__;
  assign new_new_n1056__ = new_new_n927__ & new_new_n1040__;
  assign new_new_n1057__ = new_new_n1055__ & new_new_n1056__;
  assign new_new_n1058__ = new_new_n988__ & new_new_n1054__;
  assign new_new_n1059__ = new_new_n1057__ & new_new_n1058__;
  assign new_new_n1060__ = new_new_n1030__ & new_new_n1059__;
  assign new_new_n1061__ = new_new_n983__ & new_new_n1060__;
  assign new_new_n1062__ = ~new_new_n282__ & ~new_new_n584__;
  assign new_new_n1063__ = ~new_new_n246__ & new_new_n1062__;
  assign new_new_n1064__ = new_new_n201__ & new_new_n345__;
  assign new_new_n1065__ = ~new_new_n212__ & ~new_new_n1064__;
  assign new_new_n1066__ = ~new_new_n375__ & ~new_new_n776__;
  assign new_new_n1067__ = new_new_n1063__ & new_new_n1066__;
  assign new_new_n1068__ = new_new_n1065__ & new_new_n1067__;
  assign new_new_n1069__ = ~new_new_n585__ & ~new_new_n749__;
  assign new_new_n1070__ = new_new_n163__ & new_new_n718__;
  assign new_new_n1071__ = ~new_new_n845__ & ~new_new_n1070__;
  assign new_new_n1072__ = pi24 & ~new_new_n90__;
  assign new_new_n1073__ = new_new_n285__ & new_new_n1072__;
  assign new_new_n1074__ = ~new_new_n631__ & ~new_new_n1073__;
  assign new_new_n1075__ = ~new_new_n136__ & ~new_new_n258__;
  assign new_new_n1076__ = ~new_new_n747__ & new_new_n1075__;
  assign new_new_n1077__ = ~new_new_n336__ & ~new_new_n586__;
  assign new_new_n1078__ = ~new_new_n274__ & ~new_new_n961__;
  assign new_new_n1079__ = new_new_n1077__ & new_new_n1078__;
  assign new_new_n1080__ = new_new_n81__ & new_new_n237__;
  assign new_new_n1081__ = new_new_n153__ & new_new_n169__;
  assign new_new_n1082__ = ~new_new_n1080__ & ~new_new_n1081__;
  assign new_new_n1083__ = ~new_new_n271__ & ~new_new_n351__;
  assign new_new_n1084__ = ~new_new_n76__ & ~new_new_n115__;
  assign new_new_n1085__ = ~new_new_n127__ & ~new_new_n603__;
  assign new_new_n1086__ = ~new_new_n253__ & ~new_new_n472__;
  assign new_new_n1087__ = ~new_new_n473__ & ~new_new_n933__;
  assign new_new_n1088__ = new_new_n1086__ & new_new_n1087__;
  assign new_new_n1089__ = ~new_new_n226__ & new_new_n1085__;
  assign new_new_n1090__ = new_new_n1088__ & new_new_n1089__;
  assign new_new_n1091__ = new_new_n813__ & new_new_n938__;
  assign new_new_n1092__ = new_new_n1090__ & new_new_n1091__;
  assign new_new_n1093__ = new_new_n1084__ & new_new_n1092__;
  assign new_new_n1094__ = new_new_n135__ & new_new_n718__;
  assign new_new_n1095__ = ~new_new_n298__ & ~new_new_n1094__;
  assign new_new_n1096__ = ~new_new_n846__ & ~new_new_n993__;
  assign new_new_n1097__ = ~new_new_n148__ & ~new_new_n896__;
  assign new_new_n1098__ = ~new_new_n208__ & ~new_new_n778__;
  assign new_new_n1099__ = ~new_new_n306__ & new_new_n1098__;
  assign new_new_n1100__ = ~new_new_n816__ & new_new_n1095__;
  assign new_new_n1101__ = new_new_n1099__ & new_new_n1100__;
  assign new_new_n1102__ = ~new_new_n373__ & new_new_n1096__;
  assign new_new_n1103__ = new_new_n1097__ & new_new_n1102__;
  assign new_new_n1104__ = new_new_n1101__ & new_new_n1103__;
  assign new_new_n1105__ = new_new_n114__ & new_new_n718__;
  assign new_new_n1106__ = ~new_new_n694__ & ~new_new_n1033__;
  assign new_new_n1107__ = ~new_new_n97__ & ~new_new_n169__;
  assign new_new_n1108__ = new_new_n129__ & ~new_new_n1107__;
  assign new_new_n1109__ = new_new_n91__ & new_new_n169__;
  assign new_new_n1110__ = ~new_new_n945__ & ~new_new_n1109__;
  assign new_new_n1111__ = ~new_new_n276__ & ~new_new_n350__;
  assign new_new_n1112__ = ~new_new_n441__ & ~new_new_n630__;
  assign new_new_n1113__ = new_new_n95__ & new_new_n135__;
  assign new_new_n1114__ = ~new_new_n183__ & ~new_new_n1113__;
  assign new_new_n1115__ = ~new_new_n130__ & ~new_new_n496__;
  assign new_new_n1116__ = ~new_new_n768__ & new_new_n1115__;
  assign new_new_n1117__ = ~new_new_n232__ & ~new_new_n635__;
  assign new_new_n1118__ = new_new_n966__ & new_new_n1106__;
  assign new_new_n1119__ = ~new_new_n1108__ & new_new_n1118__;
  assign new_new_n1120__ = new_new_n1116__ & new_new_n1117__;
  assign new_new_n1121__ = ~new_new_n1105__ & new_new_n1110__;
  assign new_new_n1122__ = new_new_n1111__ & new_new_n1114__;
  assign new_new_n1123__ = new_new_n1121__ & new_new_n1122__;
  assign new_new_n1124__ = new_new_n1119__ & new_new_n1120__;
  assign new_new_n1125__ = new_new_n1112__ & new_new_n1124__;
  assign new_new_n1126__ = new_new_n1123__ & new_new_n1125__;
  assign new_new_n1127__ = new_new_n1093__ & new_new_n1104__;
  assign new_new_n1128__ = new_new_n1126__ & new_new_n1127__;
  assign new_new_n1129__ = ~new_new_n95__ & ~new_new_n165__;
  assign new_new_n1130__ = new_new_n105__ & ~new_new_n1129__;
  assign new_new_n1131__ = ~new_new_n508__ & ~new_new_n673__;
  assign new_new_n1132__ = ~new_new_n138__ & ~new_new_n196__;
  assign new_new_n1133__ = ~new_new_n309__ & ~new_new_n384__;
  assign new_new_n1134__ = ~new_new_n995__ & new_new_n1133__;
  assign new_new_n1135__ = new_new_n1082__ & new_new_n1132__;
  assign new_new_n1136__ = new_new_n1083__ & ~new_new_n1130__;
  assign new_new_n1137__ = new_new_n1135__ & new_new_n1136__;
  assign new_new_n1138__ = ~new_new_n124__ & new_new_n1134__;
  assign new_new_n1139__ = new_new_n1137__ & new_new_n1138__;
  assign new_new_n1140__ = new_new_n1131__ & new_new_n1139__;
  assign new_new_n1141__ = new_new_n1128__ & new_new_n1140__;
  assign new_new_n1142__ = ~new_new_n143__ & ~new_new_n312__;
  assign new_new_n1143__ = ~new_new_n263__ & ~new_new_n489__;
  assign new_new_n1144__ = ~new_new_n715__ & new_new_n928__;
  assign new_new_n1145__ = ~new_new_n266__ & ~new_new_n963__;
  assign new_new_n1146__ = ~new_new_n675__ & ~new_new_n950__;
  assign new_new_n1147__ = ~new_new_n935__ & new_new_n1146__;
  assign new_new_n1148__ = ~new_new_n895__ & new_new_n1147__;
  assign new_new_n1149__ = new_new_n121__ & ~new_new_n254__;
  assign new_new_n1150__ = ~new_new_n353__ & ~new_new_n959__;
  assign new_new_n1151__ = new_new_n142__ & new_new_n162__;
  assign new_new_n1152__ = ~new_new_n837__ & ~new_new_n1151__;
  assign new_new_n1153__ = ~new_new_n101__ & ~new_new_n696__;
  assign new_new_n1154__ = ~new_new_n284__ & ~new_new_n692__;
  assign new_new_n1155__ = ~new_new_n300__ & new_new_n1154__;
  assign new_new_n1156__ = ~new_new_n96__ & ~new_new_n632__;
  assign new_new_n1157__ = ~new_new_n209__ & ~new_new_n1003__;
  assign new_new_n1158__ = ~new_new_n445__ & ~new_new_n566__;
  assign new_new_n1159__ = ~new_new_n785__ & ~new_new_n853__;
  assign new_new_n1160__ = new_new_n1158__ & new_new_n1159__;
  assign new_new_n1161__ = ~new_new_n222__ & ~new_new_n439__;
  assign new_new_n1162__ = new_new_n87__ & new_new_n221__;
  assign new_new_n1163__ = ~new_new_n693__ & ~new_new_n1162__;
  assign new_new_n1164__ = ~new_new_n235__ & ~new_new_n595__;
  assign new_new_n1165__ = ~new_new_n85__ & ~new_new_n137__;
  assign new_new_n1166__ = new_new_n180__ & ~new_new_n1165__;
  assign new_new_n1167__ = new_new_n77__ & new_new_n338__;
  assign new_new_n1168__ = ~new_new_n658__ & ~new_new_n1167__;
  assign new_new_n1169__ = ~new_new_n302__ & ~new_new_n383__;
  assign new_new_n1170__ = ~new_new_n656__ & ~new_new_n851__;
  assign new_new_n1171__ = ~new_new_n88__ & ~new_new_n108__;
  assign new_new_n1172__ = ~new_new_n335__ & new_new_n1171__;
  assign new_new_n1173__ = new_new_n1169__ & new_new_n1170__;
  assign new_new_n1174__ = new_new_n1172__ & new_new_n1173__;
  assign new_new_n1175__ = new_new_n1168__ & new_new_n1174__;
  assign new_new_n1176__ = new_new_n162__ & new_new_n180__;
  assign new_new_n1177__ = ~new_new_n327__ & ~new_new_n1176__;
  assign new_new_n1178__ = ~new_new_n510__ & ~new_new_n772__;
  assign new_new_n1179__ = new_new_n1156__ & new_new_n1178__;
  assign new_new_n1180__ = new_new_n1163__ & ~new_new_n1166__;
  assign new_new_n1181__ = new_new_n1177__ & new_new_n1180__;
  assign new_new_n1182__ = new_new_n1150__ & new_new_n1179__;
  assign new_new_n1183__ = new_new_n1153__ & new_new_n1155__;
  assign new_new_n1184__ = new_new_n1157__ & new_new_n1164__;
  assign new_new_n1185__ = new_new_n1183__ & new_new_n1184__;
  assign new_new_n1186__ = new_new_n1181__ & new_new_n1182__;
  assign new_new_n1187__ = new_new_n1149__ & new_new_n1152__;
  assign new_new_n1188__ = new_new_n1160__ & new_new_n1161__;
  assign new_new_n1189__ = new_new_n1187__ & new_new_n1188__;
  assign new_new_n1190__ = new_new_n1185__ & new_new_n1186__;
  assign new_new_n1191__ = new_new_n1175__ & new_new_n1190__;
  assign new_new_n1192__ = new_new_n1189__ & new_new_n1191__;
  assign new_new_n1193__ = ~new_new_n724__ & ~new_new_n783__;
  assign new_new_n1194__ = ~new_new_n871__ & new_new_n1193__;
  assign new_new_n1195__ = new_new_n1069__ & new_new_n1071__;
  assign new_new_n1196__ = new_new_n1194__ & new_new_n1195__;
  assign new_new_n1197__ = new_new_n1074__ & new_new_n1142__;
  assign new_new_n1198__ = new_new_n1143__ & new_new_n1145__;
  assign new_new_n1199__ = new_new_n1197__ & new_new_n1198__;
  assign new_new_n1200__ = new_new_n1076__ & new_new_n1196__;
  assign new_new_n1201__ = new_new_n1079__ & new_new_n1200__;
  assign new_new_n1202__ = new_new_n1068__ & new_new_n1199__;
  assign new_new_n1203__ = new_new_n1144__ & new_new_n1148__;
  assign new_new_n1204__ = new_new_n1202__ & new_new_n1203__;
  assign new_new_n1205__ = new_new_n1201__ & new_new_n1204__;
  assign new_new_n1206__ = new_new_n1192__ & new_new_n1205__;
  assign new_new_n1207__ = new_new_n1141__ & new_new_n1206__;
  assign new_new_n1208__ = ~new_new_n868__ & ~new_new_n1207__;
  assign new_new_n1209__ = ~new_new_n385__ & new_new_n1154__;
  assign new_new_n1210__ = new_new_n162__ & new_new_n241__;
  assign new_new_n1211__ = ~new_new_n772__ & ~new_new_n1210__;
  assign new_new_n1212__ = new_new_n100__ & new_new_n237__;
  assign new_new_n1213__ = ~new_new_n213__ & ~new_new_n1212__;
  assign new_new_n1214__ = ~new_new_n495__ & ~new_new_n496__;
  assign new_new_n1215__ = ~new_new_n632__ & ~new_new_n721__;
  assign new_new_n1216__ = ~new_new_n183__ & ~new_new_n246__;
  assign new_new_n1217__ = new_new_n117__ & new_new_n188__;
  assign new_new_n1218__ = ~new_new_n238__ & ~new_new_n476__;
  assign new_new_n1219__ = ~new_new_n871__ & ~new_new_n1033__;
  assign new_new_n1220__ = ~new_new_n1217__ & new_new_n1218__;
  assign new_new_n1221__ = new_new_n1219__ & new_new_n1220__;
  assign new_new_n1222__ = new_new_n985__ & new_new_n1221__;
  assign new_new_n1223__ = ~new_new_n375__ & ~new_new_n894__;
  assign new_new_n1224__ = ~new_new_n271__ & ~new_new_n1113__;
  assign new_new_n1225__ = ~new_new_n322__ & ~new_new_n884__;
  assign new_new_n1226__ = ~new_new_n136__ & ~new_new_n189__;
  assign new_new_n1227__ = ~new_new_n248__ & ~new_new_n286__;
  assign new_new_n1228__ = ~new_new_n747__ & new_new_n1227__;
  assign new_new_n1229__ = new_new_n1226__ & new_new_n1228__;
  assign new_new_n1230__ = ~new_new_n631__ & ~new_new_n890__;
  assign new_new_n1231__ = ~new_new_n143__ & ~new_new_n309__;
  assign new_new_n1232__ = ~new_new_n869__ & new_new_n1224__;
  assign new_new_n1233__ = new_new_n1231__ & new_new_n1232__;
  assign new_new_n1234__ = new_new_n1164__ & new_new_n1225__;
  assign new_new_n1235__ = new_new_n1230__ & new_new_n1234__;
  assign new_new_n1236__ = new_new_n1233__ & new_new_n1235__;
  assign new_new_n1237__ = new_new_n1229__ & new_new_n1236__;
  assign new_new_n1238__ = ~new_new_n103__ & new_new_n131__;
  assign new_new_n1239__ = new_new_n1211__ & new_new_n1213__;
  assign new_new_n1240__ = new_new_n1214__ & new_new_n1239__;
  assign new_new_n1241__ = new_new_n1209__ & new_new_n1238__;
  assign new_new_n1242__ = new_new_n1215__ & new_new_n1216__;
  assign new_new_n1243__ = new_new_n1223__ & new_new_n1242__;
  assign new_new_n1244__ = new_new_n1240__ & new_new_n1241__;
  assign new_new_n1245__ = new_new_n764__ & new_new_n1244__;
  assign new_new_n1246__ = new_new_n1148__ & new_new_n1243__;
  assign new_new_n1247__ = new_new_n1222__ & new_new_n1246__;
  assign new_new_n1248__ = new_new_n1245__ & new_new_n1247__;
  assign new_new_n1249__ = new_new_n1237__ & new_new_n1248__;
  assign new_new_n1250__ = ~new_new_n344__ & ~new_new_n603__;
  assign new_new_n1251__ = ~new_new_n382__ & ~new_new_n843__;
  assign new_new_n1252__ = ~new_new_n266__ & ~new_new_n350__;
  assign new_new_n1253__ = ~new_new_n317__ & ~new_new_n919__;
  assign new_new_n1254__ = ~new_new_n124__ & ~new_new_n308__;
  assign new_new_n1255__ = ~new_new_n993__ & new_new_n1254__;
  assign new_new_n1256__ = ~new_new_n483__ & ~new_new_n658__;
  assign new_new_n1257__ = ~new_new_n229__ & ~new_new_n937__;
  assign new_new_n1258__ = ~new_new_n701__ & ~new_new_n853__;
  assign new_new_n1259__ = new_new_n638__ & new_new_n1258__;
  assign new_new_n1260__ = ~new_new_n155__ & ~new_new_n311__;
  assign new_new_n1261__ = new_new_n672__ & new_new_n1260__;
  assign new_new_n1262__ = new_new_n1259__ & new_new_n1261__;
  assign new_new_n1263__ = ~new_new_n384__ & ~new_new_n829__;
  assign new_new_n1264__ = ~new_new_n89__ & ~new_new_n429__;
  assign new_new_n1265__ = new_new_n920__ & new_new_n1264__;
  assign new_new_n1266__ = ~new_new_n192__ & ~new_new_n488__;
  assign new_new_n1267__ = ~new_new_n1265__ & new_new_n1266__;
  assign new_new_n1268__ = ~new_new_n835__ & ~new_new_n1080__;
  assign new_new_n1269__ = new_new_n1077__ & new_new_n1257__;
  assign new_new_n1270__ = new_new_n1263__ & new_new_n1269__;
  assign new_new_n1271__ = ~new_new_n316__ & new_new_n1268__;
  assign new_new_n1272__ = new_new_n944__ & new_new_n984__;
  assign new_new_n1273__ = new_new_n1251__ & new_new_n1252__;
  assign new_new_n1274__ = new_new_n1253__ & new_new_n1256__;
  assign new_new_n1275__ = new_new_n1273__ & new_new_n1274__;
  assign new_new_n1276__ = new_new_n1271__ & new_new_n1272__;
  assign new_new_n1277__ = new_new_n1250__ & new_new_n1270__;
  assign new_new_n1278__ = new_new_n1267__ & new_new_n1277__;
  assign new_new_n1279__ = new_new_n1275__ & new_new_n1276__;
  assign new_new_n1280__ = new_new_n1255__ & new_new_n1262__;
  assign new_new_n1281__ = new_new_n1279__ & new_new_n1280__;
  assign new_new_n1282__ = new_new_n1278__ & new_new_n1281__;
  assign new_new_n1283__ = ~new_new_n179__ & ~new_new_n274__;
  assign new_new_n1284__ = ~new_new_n119__ & ~new_new_n472__;
  assign new_new_n1285__ = ~new_new_n267__ & ~new_new_n315__;
  assign new_new_n1286__ = ~new_new_n694__ & ~new_new_n1031__;
  assign new_new_n1287__ = ~new_new_n198__ & new_new_n1286__;
  assign new_new_n1288__ = ~new_new_n599__ & new_new_n1284__;
  assign new_new_n1289__ = new_new_n1285__ & new_new_n1288__;
  assign new_new_n1290__ = new_new_n1287__ & new_new_n1289__;
  assign new_new_n1291__ = new_new_n75__ & new_new_n95__;
  assign new_new_n1292__ = ~new_new_n511__ & ~new_new_n1003__;
  assign new_new_n1293__ = ~new_new_n700__ & new_new_n1292__;
  assign new_new_n1294__ = ~new_new_n226__ & ~new_new_n509__;
  assign new_new_n1295__ = ~new_new_n298__ & ~new_new_n1151__;
  assign new_new_n1296__ = ~new_new_n306__ & ~new_new_n875__;
  assign new_new_n1297__ = ~new_new_n249__ & ~new_new_n388__;
  assign new_new_n1298__ = ~new_new_n845__ & ~new_new_n896__;
  assign new_new_n1299__ = ~new_new_n1291__ & new_new_n1298__;
  assign new_new_n1300__ = ~new_new_n353__ & new_new_n1297__;
  assign new_new_n1301__ = new_new_n1299__ & new_new_n1300__;
  assign new_new_n1302__ = new_new_n1294__ & new_new_n1295__;
  assign new_new_n1303__ = new_new_n1296__ & new_new_n1302__;
  assign new_new_n1304__ = new_new_n1293__ & new_new_n1301__;
  assign new_new_n1305__ = new_new_n1303__ & new_new_n1304__;
  assign new_new_n1306__ = ~new_new_n778__ & ~new_new_n1166__;
  assign new_new_n1307__ = ~new_new_n150__ & ~new_new_n878__;
  assign new_new_n1308__ = new_new_n118__ & ~new_new_n310__;
  assign new_new_n1309__ = ~new_new_n312__ & ~new_new_n1109__;
  assign new_new_n1310__ = ~new_new_n321__ & ~new_new_n1167__;
  assign new_new_n1311__ = ~new_new_n588__ & ~new_new_n719__;
  assign new_new_n1312__ = new_new_n725__ & ~new_new_n1008__;
  assign new_new_n1313__ = ~new_new_n1308__ & new_new_n1309__;
  assign new_new_n1314__ = new_new_n1312__ & new_new_n1313__;
  assign new_new_n1315__ = ~new_new_n439__ & new_new_n1311__;
  assign new_new_n1316__ = new_new_n1283__ & new_new_n1306__;
  assign new_new_n1317__ = new_new_n1307__ & new_new_n1310__;
  assign new_new_n1318__ = new_new_n1316__ & new_new_n1317__;
  assign new_new_n1319__ = new_new_n1314__ & new_new_n1315__;
  assign new_new_n1320__ = new_new_n608__ & new_new_n1319__;
  assign new_new_n1321__ = new_new_n1290__ & new_new_n1318__;
  assign new_new_n1322__ = new_new_n1320__ & new_new_n1321__;
  assign new_new_n1323__ = new_new_n1305__ & new_new_n1322__;
  assign new_new_n1324__ = new_new_n1282__ & new_new_n1323__;
  assign new_new_n1325__ = new_new_n1249__ & new_new_n1324__;
  assign new_new_n1326__ = ~new_new_n322__ & ~new_new_n346__;
  assign new_new_n1327__ = new_new_n265__ & new_new_n512__;
  assign new_new_n1328__ = ~new_new_n213__ & ~new_new_n388__;
  assign new_new_n1329__ = ~new_new_n1327__ & new_new_n1328__;
  assign new_new_n1330__ = ~new_new_n229__ & ~new_new_n894__;
  assign new_new_n1331__ = ~new_new_n198__ & ~new_new_n853__;
  assign new_new_n1332__ = ~new_new_n283__ & ~new_new_n308__;
  assign new_new_n1333__ = ~new_new_n120__ & ~new_new_n240__;
  assign new_new_n1334__ = ~new_new_n164__ & ~new_new_n332__;
  assign new_new_n1335__ = ~new_new_n606__ & new_new_n1333__;
  assign new_new_n1336__ = new_new_n1334__ & new_new_n1335__;
  assign new_new_n1337__ = ~new_new_n375__ & ~new_new_n772__;
  assign new_new_n1338__ = ~new_new_n316__ & ~new_new_n600__;
  assign new_new_n1339__ = ~new_new_n274__ & ~new_new_n284__;
  assign new_new_n1340__ = ~new_new_n148__ & ~new_new_n242__;
  assign new_new_n1341__ = ~new_new_n136__ & ~new_new_n952__;
  assign new_new_n1342__ = ~new_new_n260__ & ~new_new_n313__;
  assign new_new_n1343__ = new_new_n153__ & new_new_n718__;
  assign new_new_n1344__ = ~new_new_n130__ & ~new_new_n335__;
  assign new_new_n1345__ = ~new_new_n1094__ & ~new_new_n1176__;
  assign new_new_n1346__ = ~new_new_n1343__ & new_new_n1345__;
  assign new_new_n1347__ = ~new_new_n878__ & new_new_n1344__;
  assign new_new_n1348__ = new_new_n1342__ & new_new_n1347__;
  assign new_new_n1349__ = new_new_n1339__ & new_new_n1346__;
  assign new_new_n1350__ = new_new_n1340__ & new_new_n1341__;
  assign new_new_n1351__ = new_new_n1349__ & new_new_n1350__;
  assign new_new_n1352__ = new_new_n1338__ & new_new_n1348__;
  assign new_new_n1353__ = new_new_n1351__ & new_new_n1352__;
  assign new_new_n1354__ = ~new_new_n634__ & ~new_new_n671__;
  assign new_new_n1355__ = ~new_new_n258__ & new_new_n1354__;
  assign new_new_n1356__ = ~new_new_n993__ & ~new_new_n1008__;
  assign new_new_n1357__ = new_new_n1332__ & new_new_n1337__;
  assign new_new_n1358__ = new_new_n1356__ & new_new_n1357__;
  assign new_new_n1359__ = new_new_n1326__ & new_new_n1355__;
  assign new_new_n1360__ = new_new_n1329__ & new_new_n1330__;
  assign new_new_n1361__ = new_new_n1331__ & new_new_n1360__;
  assign new_new_n1362__ = new_new_n1358__ & new_new_n1359__;
  assign new_new_n1363__ = new_new_n1336__ & new_new_n1362__;
  assign new_new_n1364__ = new_new_n1361__ & new_new_n1363__;
  assign new_new_n1365__ = new_new_n1353__ & new_new_n1364__;
  assign new_new_n1366__ = ~new_new_n597__ & ~new_new_n996__;
  assign new_new_n1367__ = ~new_new_n246__ & ~new_new_n933__;
  assign new_new_n1368__ = ~new_new_n603__ & ~new_new_n875__;
  assign new_new_n1369__ = ~new_new_n373__ & ~new_new_n385__;
  assign new_new_n1370__ = ~new_new_n694__ & ~new_new_n1210__;
  assign new_new_n1371__ = ~new_new_n692__ & ~new_new_n1113__;
  assign new_new_n1372__ = new_new_n91__ & new_new_n217__;
  assign new_new_n1373__ = ~new_new_n947__ & ~new_new_n1372__;
  assign new_new_n1374__ = ~new_new_n921__ & new_new_n1366__;
  assign new_new_n1375__ = new_new_n1367__ & new_new_n1368__;
  assign new_new_n1376__ = new_new_n1370__ & new_new_n1371__;
  assign new_new_n1377__ = new_new_n1373__ & new_new_n1376__;
  assign new_new_n1378__ = new_new_n1374__ & new_new_n1375__;
  assign new_new_n1379__ = new_new_n1377__ & new_new_n1378__;
  assign new_new_n1380__ = new_new_n1369__ & new_new_n1379__;
  assign new_new_n1381__ = ~new_new_n124__ & ~new_new_n845__;
  assign new_new_n1382__ = ~new_new_n127__ & ~new_new_n729__;
  assign new_new_n1383__ = ~new_new_n637__ & ~new_new_n658__;
  assign new_new_n1384__ = ~new_new_n479__ & ~new_new_n656__;
  assign new_new_n1385__ = ~new_new_n183__ & ~new_new_n383__;
  assign new_new_n1386__ = ~new_new_n329__ & ~new_new_n353__;
  assign new_new_n1387__ = new_new_n702__ & new_new_n1382__;
  assign new_new_n1388__ = new_new_n1383__ & new_new_n1387__;
  assign new_new_n1389__ = new_new_n1385__ & new_new_n1386__;
  assign new_new_n1390__ = new_new_n998__ & new_new_n1389__;
  assign new_new_n1391__ = new_new_n1381__ & new_new_n1388__;
  assign new_new_n1392__ = new_new_n1384__ & new_new_n1391__;
  assign new_new_n1393__ = new_new_n1390__ & new_new_n1392__;
  assign new_new_n1394__ = ~new_new_n336__ & ~new_new_n507__;
  assign new_new_n1395__ = ~new_new_n635__ & ~new_new_n1070__;
  assign new_new_n1396__ = new_new_n1394__ & new_new_n1395__;
  assign new_new_n1397__ = ~new_new_n321__ & ~new_new_n344__;
  assign new_new_n1398__ = new_new_n129__ & new_new_n162__;
  assign new_new_n1399__ = ~new_new_n350__ & ~new_new_n1398__;
  assign new_new_n1400__ = ~new_new_n115__ & ~new_new_n846__;
  assign new_new_n1401__ = ~new_new_n372__ & ~new_new_n871__;
  assign new_new_n1402__ = ~new_new_n96__ & ~new_new_n950__;
  assign new_new_n1403__ = ~new_new_n1212__ & new_new_n1402__;
  assign new_new_n1404__ = new_new_n1399__ & new_new_n1403__;
  assign new_new_n1405__ = new_new_n1401__ & new_new_n1404__;
  assign new_new_n1406__ = new_new_n1397__ & new_new_n1400__;
  assign new_new_n1407__ = new_new_n1405__ & new_new_n1406__;
  assign new_new_n1408__ = ~new_new_n169__ & ~new_new_n718__;
  assign new_new_n1409__ = new_new_n87__ & ~new_new_n1408__;
  assign new_new_n1410__ = ~new_new_n302__ & ~new_new_n843__;
  assign new_new_n1411__ = ~new_new_n92__ & ~new_new_n138__;
  assign new_new_n1412__ = ~new_new_n251__ & ~new_new_n252__;
  assign new_new_n1413__ = ~new_new_n495__ & ~new_new_n584__;
  assign new_new_n1414__ = ~new_new_n1031__ & ~new_new_n1080__;
  assign new_new_n1415__ = new_new_n1413__ & new_new_n1414__;
  assign new_new_n1416__ = new_new_n1411__ & new_new_n1412__;
  assign new_new_n1417__ = ~new_new_n566__ & ~new_new_n1409__;
  assign new_new_n1418__ = new_new_n1410__ & new_new_n1417__;
  assign new_new_n1419__ = new_new_n1415__ & new_new_n1416__;
  assign new_new_n1420__ = new_new_n633__ & new_new_n1419__;
  assign new_new_n1421__ = new_new_n1418__ & new_new_n1420__;
  assign new_new_n1422__ = ~new_new_n696__ & ~new_new_n717__;
  assign new_new_n1423__ = ~new_new_n476__ & ~new_new_n778__;
  assign new_new_n1424__ = ~new_new_n715__ & ~new_new_n1109__;
  assign new_new_n1425__ = ~new_new_n106__ & ~new_new_n168__;
  assign new_new_n1426__ = ~new_new_n959__ & new_new_n1425__;
  assign new_new_n1427__ = new_new_n622__ & new_new_n1426__;
  assign new_new_n1428__ = ~new_new_n835__ & ~new_new_n939__;
  assign new_new_n1429__ = ~new_new_n884__ & ~new_new_n945__;
  assign new_new_n1430__ = new_new_n1428__ & new_new_n1429__;
  assign new_new_n1431__ = ~new_new_n895__ & new_new_n1430__;
  assign new_new_n1432__ = ~new_new_n312__ & ~new_new_n374__;
  assign new_new_n1433__ = new_new_n725__ & new_new_n1432__;
  assign new_new_n1434__ = ~new_new_n816__ & new_new_n1433__;
  assign new_new_n1435__ = ~new_new_n731__ & ~new_new_n995__;
  assign new_new_n1436__ = ~new_new_n286__ & new_new_n1435__;
  assign new_new_n1437__ = new_new_n1423__ & new_new_n1424__;
  assign new_new_n1438__ = new_new_n1436__ & new_new_n1437__;
  assign new_new_n1439__ = new_new_n1422__ & new_new_n1438__;
  assign new_new_n1440__ = new_new_n256__ & new_new_n1161__;
  assign new_new_n1441__ = new_new_n1427__ & new_new_n1434__;
  assign new_new_n1442__ = new_new_n1440__ & new_new_n1441__;
  assign new_new_n1443__ = new_new_n1431__ & new_new_n1439__;
  assign new_new_n1444__ = new_new_n1442__ & new_new_n1443__;
  assign new_new_n1445__ = new_new_n1407__ & new_new_n1421__;
  assign new_new_n1446__ = new_new_n1444__ & new_new_n1445__;
  assign new_new_n1447__ = ~new_new_n510__ & ~new_new_n721__;
  assign new_new_n1448__ = ~new_new_n259__ & ~new_new_n591__;
  assign new_new_n1449__ = ~new_new_n379__ & ~new_new_n776__;
  assign new_new_n1450__ = ~new_new_n315__ & ~new_new_n1217__;
  assign new_new_n1451__ = ~new_new_n657__ & ~new_new_n1064__;
  assign new_new_n1452__ = ~new_new_n282__ & ~new_new_n785__;
  assign new_new_n1453__ = new_new_n1011__ & new_new_n1452__;
  assign new_new_n1454__ = ~new_new_n150__ & ~new_new_n226__;
  assign new_new_n1455__ = ~new_new_n263__ & new_new_n1449__;
  assign new_new_n1456__ = new_new_n1454__ & new_new_n1455__;
  assign new_new_n1457__ = new_new_n1447__ & new_new_n1453__;
  assign new_new_n1458__ = new_new_n1448__ & new_new_n1450__;
  assign new_new_n1459__ = new_new_n1451__ & new_new_n1458__;
  assign new_new_n1460__ = new_new_n1456__ & new_new_n1457__;
  assign new_new_n1461__ = new_new_n1396__ & new_new_n1460__;
  assign new_new_n1462__ = new_new_n1459__ & new_new_n1461__;
  assign new_new_n1463__ = new_new_n1380__ & new_new_n1462__;
  assign new_new_n1464__ = new_new_n1393__ & new_new_n1463__;
  assign new_new_n1465__ = new_new_n1365__ & new_new_n1446__;
  assign new_new_n1466__ = new_new_n1464__ & new_new_n1465__;
  assign new_new_n1467__ = new_new_n1325__ & new_new_n1466__;
  assign new_new_n1468__ = ~new_new_n263__ & ~new_new_n1109__;
  assign new_new_n1469__ = ~new_new_n336__ & ~new_new_n1031__;
  assign new_new_n1470__ = ~new_new_n313__ & ~new_new_n511__;
  assign new_new_n1471__ = ~new_new_n222__ & ~new_new_n635__;
  assign new_new_n1472__ = ~new_new_n232__ & ~new_new_n729__;
  assign new_new_n1473__ = ~new_new_n719__ & ~new_new_n835__;
  assign new_new_n1474__ = ~new_new_n260__ & ~new_new_n298__;
  assign new_new_n1475__ = ~new_new_n335__ & ~new_new_n634__;
  assign new_new_n1476__ = ~new_new_n1080__ & new_new_n1475__;
  assign new_new_n1477__ = new_new_n1474__ & new_new_n1476__;
  assign new_new_n1478__ = ~new_new_n254__ & ~new_new_n479__;
  assign new_new_n1479__ = new_new_n1473__ & new_new_n1478__;
  assign new_new_n1480__ = new_new_n1477__ & new_new_n1479__;
  assign new_new_n1481__ = ~new_new_n280__ & ~new_new_n658__;
  assign new_new_n1482__ = ~new_new_n242__ & ~new_new_n266__;
  assign new_new_n1483__ = pi23 & new_new_n430__;
  assign new_new_n1484__ = new_new_n718__ & new_new_n1483__;
  assign new_new_n1485__ = ~new_new_n197__ & ~new_new_n1484__;
  assign new_new_n1486__ = ~pi24 & ~new_new_n1485__;
  assign new_new_n1487__ = ~new_new_n306__ & ~new_new_n919__;
  assign new_new_n1488__ = ~new_new_n673__ & new_new_n1469__;
  assign new_new_n1489__ = new_new_n1470__ & new_new_n1488__;
  assign new_new_n1490__ = new_new_n1037__ & new_new_n1468__;
  assign new_new_n1491__ = new_new_n1471__ & new_new_n1472__;
  assign new_new_n1492__ = new_new_n1481__ & new_new_n1482__;
  assign new_new_n1493__ = ~new_new_n1486__ & new_new_n1487__;
  assign new_new_n1494__ = new_new_n1492__ & new_new_n1493__;
  assign new_new_n1495__ = new_new_n1490__ & new_new_n1491__;
  assign new_new_n1496__ = new_new_n1489__ & new_new_n1495__;
  assign new_new_n1497__ = new_new_n1494__ & new_new_n1496__;
  assign new_new_n1498__ = new_new_n1480__ & new_new_n1497__;
  assign new_new_n1499__ = ~new_new_n270__ & ~new_new_n939__;
  assign new_new_n1500__ = ~new_new_n252__ & ~new_new_n749__;
  assign new_new_n1501__ = ~new_new_n776__ & ~new_new_n1176__;
  assign new_new_n1502__ = new_new_n1500__ & new_new_n1501__;
  assign new_new_n1503__ = new_new_n1150__ & new_new_n1502__;
  assign new_new_n1504__ = new_new_n1499__ & new_new_n1503__;
  assign new_new_n1505__ = ~new_new_n240__ & ~new_new_n853__;
  assign new_new_n1506__ = new_new_n90__ & new_new_n780__;
  assign new_new_n1507__ = new_new_n169__ & new_new_n279__;
  assign new_new_n1508__ = ~new_new_n1506__ & ~new_new_n1507__;
  assign new_new_n1509__ = ~new_new_n445__ & ~new_new_n585__;
  assign new_new_n1510__ = ~new_new_n283__ & ~new_new_n510__;
  assign new_new_n1511__ = ~new_new_n584__ & ~new_new_n715__;
  assign new_new_n1512__ = new_new_n129__ & ~new_new_n310__;
  assign new_new_n1513__ = ~new_new_n375__ & ~new_new_n1003__;
  assign new_new_n1514__ = ~new_new_n438__ & ~new_new_n935__;
  assign new_new_n1515__ = new_new_n87__ & new_new_n169__;
  assign new_new_n1516__ = ~new_new_n489__ & ~new_new_n1515__;
  assign new_new_n1517__ = ~new_new_n166__ & ~new_new_n1070__;
  assign new_new_n1518__ = ~new_new_n238__ & new_new_n1224__;
  assign new_new_n1519__ = ~new_new_n676__ & new_new_n1518__;
  assign new_new_n1520__ = new_new_n1516__ & new_new_n1517__;
  assign new_new_n1521__ = new_new_n1519__ & new_new_n1520__;
  assign new_new_n1522__ = ~new_new_n213__ & ~new_new_n1162__;
  assign new_new_n1523__ = ~new_new_n747__ & ~new_new_n826__;
  assign new_new_n1524__ = ~new_new_n136__ & ~new_new_n251__;
  assign new_new_n1525__ = ~new_new_n329__ & new_new_n1524__;
  assign new_new_n1526__ = new_new_n943__ & new_new_n1525__;
  assign new_new_n1527__ = ~new_new_n320__ & ~new_new_n351__;
  assign new_new_n1528__ = ~new_new_n600__ & new_new_n1527__;
  assign new_new_n1529__ = ~new_new_n274__ & ~new_new_n276__;
  assign new_new_n1530__ = ~new_new_n382__ & new_new_n1522__;
  assign new_new_n1531__ = new_new_n1529__ & new_new_n1530__;
  assign new_new_n1532__ = new_new_n1216__ & new_new_n1528__;
  assign new_new_n1533__ = new_new_n1448__ & new_new_n1523__;
  assign new_new_n1534__ = new_new_n1532__ & new_new_n1533__;
  assign new_new_n1535__ = new_new_n1514__ & new_new_n1531__;
  assign new_new_n1536__ = new_new_n1534__ & new_new_n1535__;
  assign new_new_n1537__ = new_new_n1521__ & new_new_n1526__;
  assign new_new_n1538__ = new_new_n1536__ & new_new_n1537__;
  assign new_new_n1539__ = new_new_n506__ & ~new_new_n801__;
  assign new_new_n1540__ = ~new_new_n103__ & ~new_new_n597__;
  assign new_new_n1541__ = ~new_new_n842__ & new_new_n1540__;
  assign new_new_n1542__ = new_new_n1505__ & new_new_n1509__;
  assign new_new_n1543__ = new_new_n1510__ & new_new_n1511__;
  assign new_new_n1544__ = ~new_new_n1512__ & new_new_n1543__;
  assign new_new_n1545__ = new_new_n1541__ & new_new_n1542__;
  assign new_new_n1546__ = new_new_n391__ & new_new_n743__;
  assign new_new_n1547__ = new_new_n1142__ & new_new_n1508__;
  assign new_new_n1548__ = new_new_n1513__ & new_new_n1547__;
  assign new_new_n1549__ = new_new_n1545__ & new_new_n1546__;
  assign new_new_n1550__ = ~new_new_n1539__ & new_new_n1544__;
  assign new_new_n1551__ = new_new_n1549__ & new_new_n1550__;
  assign new_new_n1552__ = new_new_n1504__ & new_new_n1548__;
  assign new_new_n1553__ = new_new_n1551__ & new_new_n1552__;
  assign new_new_n1554__ = new_new_n1093__ & new_new_n1553__;
  assign new_new_n1555__ = new_new_n1538__ & new_new_n1554__;
  assign new_new_n1556__ = new_new_n1498__ & new_new_n1555__;
  assign new_new_n1557__ = ~new_new_n1467__ & ~new_new_n1556__;
  assign new_new_n1558__ = ~new_new_n375__ & ~new_new_n990__;
  assign new_new_n1559__ = ~new_new_n196__ & ~new_new_n1291__;
  assign new_new_n1560__ = ~new_new_n509__ & ~new_new_n996__;
  assign new_new_n1561__ = new_new_n1558__ & new_new_n1560__;
  assign new_new_n1562__ = new_new_n1559__ & new_new_n1561__;
  assign new_new_n1563__ = ~new_new_n238__ & ~new_new_n896__;
  assign new_new_n1564__ = ~new_new_n160__ & ~new_new_n595__;
  assign new_new_n1565__ = ~new_new_n106__ & ~new_new_n164__;
  assign new_new_n1566__ = ~new_new_n816__ & ~new_new_n837__;
  assign new_new_n1567__ = new_new_n141__ & new_new_n718__;
  assign new_new_n1568__ = new_new_n433__ & new_new_n1567__;
  assign new_new_n1569__ = ~new_new_n668__ & ~new_new_n835__;
  assign new_new_n1570__ = ~new_new_n108__ & ~new_new_n379__;
  assign new_new_n1571__ = ~new_new_n92__ & ~new_new_n724__;
  assign new_new_n1572__ = ~new_new_n130__ & ~new_new_n871__;
  assign new_new_n1573__ = ~new_new_n134__ & ~new_new_n892__;
  assign new_new_n1574__ = new_new_n169__ & new_new_n1573__;
  assign new_new_n1575__ = new_new_n873__ & new_new_n1574__;
  assign new_new_n1576__ = ~new_new_n311__ & new_new_n1570__;
  assign new_new_n1577__ = new_new_n1571__ & ~new_new_n1575__;
  assign new_new_n1578__ = new_new_n1576__ & new_new_n1577__;
  assign new_new_n1579__ = new_new_n1572__ & new_new_n1578__;
  assign new_new_n1580__ = ~new_new_n313__ & ~new_new_n472__;
  assign new_new_n1581__ = ~new_new_n591__ & new_new_n1580__;
  assign new_new_n1582__ = ~new_new_n635__ & ~new_new_n842__;
  assign new_new_n1583__ = ~new_new_n894__ & new_new_n1154__;
  assign new_new_n1584__ = new_new_n1423__ & new_new_n1563__;
  assign new_new_n1585__ = new_new_n1565__ & ~new_new_n1568__;
  assign new_new_n1586__ = new_new_n1584__ & new_new_n1585__;
  assign new_new_n1587__ = new_new_n1582__ & new_new_n1583__;
  assign new_new_n1588__ = ~new_new_n344__ & new_new_n1581__;
  assign new_new_n1589__ = new_new_n628__ & new_new_n1564__;
  assign new_new_n1590__ = new_new_n1588__ & new_new_n1589__;
  assign new_new_n1591__ = new_new_n1586__ & new_new_n1587__;
  assign new_new_n1592__ = new_new_n734__ & new_new_n1566__;
  assign new_new_n1593__ = new_new_n1591__ & new_new_n1592__;
  assign new_new_n1594__ = new_new_n1569__ & new_new_n1590__;
  assign new_new_n1595__ = new_new_n1579__ & new_new_n1594__;
  assign new_new_n1596__ = new_new_n1593__ & new_new_n1595__;
  assign new_new_n1597__ = ~new_new_n212__ & ~new_new_n480__;
  assign new_new_n1598__ = ~new_new_n235__ & ~new_new_n809__;
  assign new_new_n1599__ = ~new_new_n306__ & ~new_new_n600__;
  assign new_new_n1600__ = ~new_new_n335__ & ~new_new_n1113__;
  assign new_new_n1601__ = ~new_new_n427__ & new_new_n1600__;
  assign new_new_n1602__ = new_new_n1597__ & new_new_n1601__;
  assign new_new_n1603__ = ~new_new_n607__ & new_new_n1599__;
  assign new_new_n1604__ = new_new_n1602__ & new_new_n1603__;
  assign new_new_n1605__ = new_new_n1598__ & new_new_n1604__;
  assign new_new_n1606__ = ~new_new_n441__ & ~new_new_n875__;
  assign new_new_n1607__ = ~new_new_n179__ & ~new_new_n597__;
  assign new_new_n1608__ = ~new_new_n1105__ & new_new_n1607__;
  assign new_new_n1609__ = ~new_new_n312__ & ~new_new_n772__;
  assign new_new_n1610__ = new_new_n1608__ & new_new_n1609__;
  assign new_new_n1611__ = ~new_new_n255__ & ~new_new_n878__;
  assign new_new_n1612__ = ~new_new_n213__ & ~new_new_n1035__;
  assign new_new_n1613__ = ~new_new_n101__ & ~new_new_n222__;
  assign new_new_n1614__ = ~new_new_n271__ & ~new_new_n388__;
  assign new_new_n1615__ = ~new_new_n700__ & ~new_new_n1031__;
  assign new_new_n1616__ = ~new_new_n1210__ & new_new_n1615__;
  assign new_new_n1617__ = new_new_n1613__ & new_new_n1614__;
  assign new_new_n1618__ = new_new_n210__ & new_new_n261__;
  assign new_new_n1619__ = new_new_n1606__ & new_new_n1618__;
  assign new_new_n1620__ = new_new_n1616__ & new_new_n1617__;
  assign new_new_n1621__ = new_new_n1611__ & new_new_n1612__;
  assign new_new_n1622__ = new_new_n1620__ & new_new_n1621__;
  assign new_new_n1623__ = new_new_n1076__ & new_new_n1619__;
  assign new_new_n1624__ = new_new_n1622__ & new_new_n1623__;
  assign new_new_n1625__ = new_new_n1610__ & new_new_n1624__;
  assign new_new_n1626__ = new_new_n1605__ & new_new_n1625__;
  assign new_new_n1627__ = ~new_new_n88__ & ~new_new_n479__;
  assign new_new_n1628__ = ~new_new_n658__ & ~new_new_n729__;
  assign new_new_n1629__ = ~new_new_n247__ & ~new_new_n496__;
  assign new_new_n1630__ = ~new_new_n253__ & ~new_new_n286__;
  assign new_new_n1631__ = ~new_new_n82__ & ~new_new_n252__;
  assign new_new_n1632__ = new_new_n91__ & ~new_new_n773__;
  assign new_new_n1633__ = ~new_new_n719__ & ~new_new_n1632__;
  assign new_new_n1634__ = ~new_new_n1166__ & new_new_n1633__;
  assign new_new_n1635__ = new_new_n1131__ & new_new_n1634__;
  assign new_new_n1636__ = ~new_new_n385__ & ~new_new_n488__;
  assign new_new_n1637__ = ~new_new_n226__ & ~new_new_n732__;
  assign new_new_n1638__ = new_new_n137__ & ~new_new_n598__;
  assign new_new_n1639__ = ~new_new_n250__ & ~new_new_n384__;
  assign new_new_n1640__ = ~new_new_n656__ & ~new_new_n701__;
  assign new_new_n1641__ = ~new_new_n1638__ & new_new_n1640__;
  assign new_new_n1642__ = new_new_n1639__ & new_new_n1641__;
  assign new_new_n1643__ = new_new_n1636__ & new_new_n1637__;
  assign new_new_n1644__ = new_new_n1642__ & new_new_n1643__;
  assign new_new_n1645__ = ~new_new_n322__ & ~new_new_n942__;
  assign new_new_n1646__ = ~new_new_n309__ & ~new_new_n829__;
  assign new_new_n1647__ = new_new_n121__ & new_new_n1646__;
  assign new_new_n1648__ = ~new_new_n919__ & ~new_new_n939__;
  assign new_new_n1649__ = new_new_n1628__ & new_new_n1629__;
  assign new_new_n1650__ = new_new_n1631__ & new_new_n1649__;
  assign new_new_n1651__ = new_new_n1647__ & new_new_n1648__;
  assign new_new_n1652__ = new_new_n1630__ & new_new_n1645__;
  assign new_new_n1653__ = new_new_n1651__ & new_new_n1652__;
  assign new_new_n1654__ = new_new_n1562__ & new_new_n1650__;
  assign new_new_n1655__ = new_new_n1627__ & new_new_n1654__;
  assign new_new_n1656__ = new_new_n1635__ & new_new_n1653__;
  assign new_new_n1657__ = new_new_n1644__ & new_new_n1656__;
  assign new_new_n1658__ = new_new_n1655__ & new_new_n1657__;
  assign new_new_n1659__ = new_new_n1596__ & new_new_n1658__;
  assign new_new_n1660__ = new_new_n1626__ & new_new_n1659__;
  assign new_new_n1661__ = ~new_new_n160__ & ~new_new_n961__;
  assign new_new_n1662__ = ~new_new_n935__ & ~new_new_n1151__;
  assign new_new_n1663__ = ~new_new_n298__ & ~new_new_n657__;
  assign new_new_n1664__ = ~new_new_n1031__ & new_new_n1663__;
  assign new_new_n1665__ = ~new_new_n427__ & ~new_new_n693__;
  assign new_new_n1666__ = ~new_new_n315__ & ~new_new_n715__;
  assign new_new_n1667__ = ~new_new_n1372__ & new_new_n1666__;
  assign new_new_n1668__ = ~new_new_n143__ & ~new_new_n255__;
  assign new_new_n1669__ = ~new_new_n353__ & new_new_n730__;
  assign new_new_n1670__ = ~new_new_n952__ & new_new_n1669__;
  assign new_new_n1671__ = new_new_n1667__ & new_new_n1668__;
  assign new_new_n1672__ = new_new_n1661__ & new_new_n1664__;
  assign new_new_n1673__ = new_new_n1665__ & new_new_n1672__;
  assign new_new_n1674__ = new_new_n1670__ & new_new_n1671__;
  assign new_new_n1675__ = new_new_n1662__ & new_new_n1674__;
  assign new_new_n1676__ = new_new_n1673__ & new_new_n1675__;
  assign new_new_n1677__ = ~new_new_n445__ & ~new_new_n1003__;
  assign new_new_n1678__ = ~new_new_n200__ & ~new_new_n511__;
  assign new_new_n1679__ = ~new_new_n586__ & ~new_new_n591__;
  assign new_new_n1680__ = ~new_new_n150__ & ~new_new_n309__;
  assign new_new_n1681__ = new_new_n1627__ & new_new_n1680__;
  assign new_new_n1682__ = ~new_new_n164__ & ~new_new_n248__;
  assign new_new_n1683__ = ~new_new_n624__ & ~new_new_n1109__;
  assign new_new_n1684__ = ~new_new_n1113__ & new_new_n1683__;
  assign new_new_n1685__ = ~new_new_n1166__ & new_new_n1682__;
  assign new_new_n1686__ = new_new_n1263__ & ~new_new_n1265__;
  assign new_new_n1687__ = new_new_n1678__ & new_new_n1686__;
  assign new_new_n1688__ = new_new_n1684__ & new_new_n1685__;
  assign new_new_n1689__ = ~new_new_n115__ & ~new_new_n344__;
  assign new_new_n1690__ = new_new_n782__ & new_new_n1677__;
  assign new_new_n1691__ = new_new_n1679__ & new_new_n1690__;
  assign new_new_n1692__ = new_new_n1688__ & new_new_n1689__;
  assign new_new_n1693__ = new_new_n1396__ & new_new_n1687__;
  assign new_new_n1694__ = ~new_new_n1539__ & new_new_n1693__;
  assign new_new_n1695__ = new_new_n1691__ & new_new_n1692__;
  assign new_new_n1696__ = new_new_n1431__ & new_new_n1681__;
  assign new_new_n1697__ = new_new_n1695__ & new_new_n1696__;
  assign new_new_n1698__ = new_new_n293__ & new_new_n1694__;
  assign new_new_n1699__ = new_new_n1697__ & new_new_n1698__;
  assign new_new_n1700__ = ~new_new_n72__ & ~new_new_n718__;
  assign new_new_n1701__ = new_new_n180__ & ~new_new_n1700__;
  assign new_new_n1702__ = ~new_new_n101__ & ~new_new_n846__;
  assign new_new_n1703__ = ~new_new_n106__ & ~new_new_n306__;
  assign new_new_n1704__ = ~new_new_n483__ & ~new_new_n837__;
  assign new_new_n1705__ = ~new_new_n480__ & ~new_new_n595__;
  assign new_new_n1706__ = ~new_new_n267__ & ~new_new_n772__;
  assign new_new_n1707__ = ~new_new_n838__ & new_new_n1706__;
  assign new_new_n1708__ = new_new_n1705__ & new_new_n1707__;
  assign new_new_n1709__ = ~new_new_n776__ & ~new_new_n890__;
  assign new_new_n1710__ = ~new_new_n942__ & new_new_n1709__;
  assign new_new_n1711__ = ~new_new_n995__ & ~new_new_n1162__;
  assign new_new_n1712__ = ~new_new_n249__ & ~new_new_n348__;
  assign new_new_n1713__ = ~new_new_n253__ & ~new_new_n698__;
  assign new_new_n1714__ = ~new_new_n701__ & ~new_new_n749__;
  assign new_new_n1715__ = new_new_n1711__ & new_new_n1714__;
  assign new_new_n1716__ = new_new_n1713__ & new_new_n1715__;
  assign new_new_n1717__ = new_new_n1712__ & new_new_n1716__;
  assign new_new_n1718__ = ~new_new_n335__ & ~new_new_n495__;
  assign new_new_n1719__ = ~new_new_n990__ & new_new_n1718__;
  assign new_new_n1720__ = ~new_new_n232__ & ~new_new_n878__;
  assign new_new_n1721__ = new_new_n1213__ & ~new_new_n1701__;
  assign new_new_n1722__ = new_new_n1702__ & new_new_n1721__;
  assign new_new_n1723__ = new_new_n1719__ & new_new_n1720__;
  assign new_new_n1724__ = ~new_new_n630__ & ~new_new_n1105__;
  assign new_new_n1725__ = new_new_n1215__ & new_new_n1399__;
  assign new_new_n1726__ = new_new_n1703__ & new_new_n1710__;
  assign new_new_n1727__ = new_new_n1725__ & new_new_n1726__;
  assign new_new_n1728__ = new_new_n1723__ & new_new_n1724__;
  assign new_new_n1729__ = new_new_n378__ & new_new_n1722__;
  assign new_new_n1730__ = new_new_n985__ & new_new_n1704__;
  assign new_new_n1731__ = new_new_n1708__ & new_new_n1730__;
  assign new_new_n1732__ = new_new_n1728__ & new_new_n1729__;
  assign new_new_n1733__ = new_new_n1717__ & new_new_n1727__;
  assign new_new_n1734__ = new_new_n1732__ & new_new_n1733__;
  assign new_new_n1735__ = new_new_n1731__ & new_new_n1734__;
  assign new_new_n1736__ = new_new_n1676__ & new_new_n1735__;
  assign new_new_n1737__ = new_new_n1699__ & new_new_n1736__;
  assign new_new_n1738__ = ~new_new_n1556__ & ~new_new_n1737__;
  assign new_new_n1739__ = ~new_new_n1325__ & ~new_new_n1466__;
  assign new_new_n1740__ = ~new_new_n238__ & ~new_new_n749__;
  assign new_new_n1741__ = ~new_new_n96__ & ~new_new_n248__;
  assign new_new_n1742__ = ~new_new_n604__ & ~new_new_n624__;
  assign new_new_n1743__ = ~new_new_n226__ & ~new_new_n252__;
  assign new_new_n1744__ = ~new_new_n271__ & ~new_new_n438__;
  assign new_new_n1745__ = new_new_n1743__ & new_new_n1744__;
  assign new_new_n1746__ = ~new_new_n510__ & ~new_new_n829__;
  assign new_new_n1747__ = ~new_new_n1008__ & new_new_n1746__;
  assign new_new_n1748__ = ~new_new_n258__ & ~new_new_n869__;
  assign new_new_n1749__ = ~new_new_n380__ & new_new_n1448__;
  assign new_new_n1750__ = ~new_new_n148__ & ~new_new_n312__;
  assign new_new_n1751__ = ~new_new_n250__ & ~new_new_n332__;
  assign new_new_n1752__ = new_new_n1750__ & new_new_n1751__;
  assign new_new_n1753__ = ~new_new_n82__ & ~new_new_n101__;
  assign new_new_n1754__ = ~new_new_n280__ & new_new_n1753__;
  assign new_new_n1755__ = ~new_new_n884__ & new_new_n1740__;
  assign new_new_n1756__ = new_new_n1741__ & new_new_n1742__;
  assign new_new_n1757__ = new_new_n1755__ & new_new_n1756__;
  assign new_new_n1758__ = ~new_new_n607__ & new_new_n1754__;
  assign new_new_n1759__ = new_new_n1747__ & new_new_n1748__;
  assign new_new_n1760__ = new_new_n1758__ & new_new_n1759__;
  assign new_new_n1761__ = new_new_n347__ & new_new_n1757__;
  assign new_new_n1762__ = new_new_n985__ & new_new_n1708__;
  assign new_new_n1763__ = new_new_n1745__ & new_new_n1749__;
  assign new_new_n1764__ = new_new_n1752__ & new_new_n1763__;
  assign new_new_n1765__ = new_new_n1761__ & new_new_n1762__;
  assign new_new_n1766__ = new_new_n1760__ & new_new_n1765__;
  assign new_new_n1767__ = new_new_n1764__ & new_new_n1766__;
  assign new_new_n1768__ = ~new_new_n160__ & ~new_new_n222__;
  assign new_new_n1769__ = ~new_new_n375__ & ~new_new_n445__;
  assign new_new_n1770__ = new_new_n1768__ & new_new_n1769__;
  assign new_new_n1771__ = new_new_n1487__ & new_new_n1770__;
  assign new_new_n1772__ = ~new_new_n509__ & ~new_new_n1105__;
  assign new_new_n1773__ = ~new_new_n384__ & ~new_new_n584__;
  assign new_new_n1774__ = ~new_new_n776__ & ~new_new_n837__;
  assign new_new_n1775__ = ~new_new_n816__ & ~new_new_n890__;
  assign new_new_n1776__ = new_new_n1774__ & new_new_n1775__;
  assign new_new_n1777__ = ~new_new_n166__ & ~new_new_n235__;
  assign new_new_n1778__ = ~new_new_n247__ & ~new_new_n276__;
  assign new_new_n1779__ = ~new_new_n92__ & ~new_new_n212__;
  assign new_new_n1780__ = ~new_new_n374__ & ~new_new_n473__;
  assign new_new_n1781__ = ~new_new_n698__ & new_new_n1780__;
  assign new_new_n1782__ = ~new_new_n143__ & new_new_n1779__;
  assign new_new_n1783__ = ~new_new_n781__ & ~new_new_n939__;
  assign new_new_n1784__ = ~new_new_n1506__ & new_new_n1773__;
  assign new_new_n1785__ = new_new_n1783__ & new_new_n1784__;
  assign new_new_n1786__ = new_new_n1781__ & new_new_n1782__;
  assign new_new_n1787__ = ~new_new_n254__ & new_new_n1523__;
  assign new_new_n1788__ = new_new_n1777__ & new_new_n1778__;
  assign new_new_n1789__ = new_new_n1787__ & new_new_n1788__;
  assign new_new_n1790__ = new_new_n1785__ & new_new_n1786__;
  assign new_new_n1791__ = new_new_n1427__ & new_new_n1772__;
  assign new_new_n1792__ = new_new_n1790__ & new_new_n1791__;
  assign new_new_n1793__ = new_new_n1776__ & new_new_n1789__;
  assign new_new_n1794__ = new_new_n1792__ & new_new_n1793__;
  assign new_new_n1795__ = new_new_n1380__ & new_new_n1794__;
  assign new_new_n1796__ = ~new_new_n137__ & new_new_n310__;
  assign new_new_n1797__ = new_new_n180__ & ~new_new_n1796__;
  assign new_new_n1798__ = ~new_new_n108__ & ~new_new_n382__;
  assign new_new_n1799__ = ~new_new_n602__ & ~new_new_n1003__;
  assign new_new_n1800__ = new_new_n1798__ & new_new_n1799__;
  assign new_new_n1801__ = new_new_n1712__ & ~new_new_n1797__;
  assign new_new_n1802__ = new_new_n1800__ & new_new_n1801__;
  assign new_new_n1803__ = ~new_new_n439__ & ~new_new_n489__;
  assign new_new_n1804__ = ~new_new_n119__ & ~new_new_n255__;
  assign new_new_n1805__ = ~new_new_n76__ & ~new_new_n630__;
  assign new_new_n1806__ = ~new_new_n266__ & ~new_new_n1398__;
  assign new_new_n1807__ = ~new_new_n213__ & ~new_new_n1007__;
  assign new_new_n1808__ = ~new_new_n671__ & ~new_new_n717__;
  assign new_new_n1809__ = ~new_new_n1515__ & new_new_n1808__;
  assign new_new_n1810__ = ~new_new_n202__ & ~new_new_n1073__;
  assign new_new_n1811__ = new_new_n1807__ & new_new_n1810__;
  assign new_new_n1812__ = new_new_n1473__ & new_new_n1809__;
  assign new_new_n1813__ = new_new_n1572__ & new_new_n1804__;
  assign new_new_n1814__ = new_new_n1806__ & new_new_n1813__;
  assign new_new_n1815__ = new_new_n1811__ & new_new_n1812__;
  assign new_new_n1816__ = new_new_n1771__ & new_new_n1803__;
  assign new_new_n1817__ = new_new_n1805__ & new_new_n1816__;
  assign new_new_n1818__ = new_new_n1814__ & new_new_n1815__;
  assign new_new_n1819__ = new_new_n1802__ & new_new_n1818__;
  assign new_new_n1820__ = new_new_n1817__ & new_new_n1819__;
  assign new_new_n1821__ = new_new_n1393__ & new_new_n1820__;
  assign new_new_n1822__ = new_new_n1767__ & new_new_n1795__;
  assign new_new_n1823__ = new_new_n1821__ & new_new_n1822__;
  assign new_new_n1824__ = new_new_n1660__ & new_new_n1823__;
  assign new_new_n1825__ = ~new_new_n327__ & ~new_new_n673__;
  assign new_new_n1826__ = ~new_new_n218__ & ~new_new_n894__;
  assign new_new_n1827__ = ~new_new_n586__ & ~new_new_n939__;
  assign new_new_n1828__ = ~new_new_n477__ & ~new_new_n851__;
  assign new_new_n1829__ = ~new_new_n251__ & ~new_new_n811__;
  assign new_new_n1830__ = ~new_new_n235__ & ~new_new_n1291__;
  assign new_new_n1831__ = ~new_new_n473__ & ~new_new_n1151__;
  assign new_new_n1832__ = new_new_n1829__ & new_new_n1830__;
  assign new_new_n1833__ = new_new_n1831__ & new_new_n1832__;
  assign new_new_n1834__ = ~new_new_n508__ & new_new_n1451__;
  assign new_new_n1835__ = new_new_n1825__ & new_new_n1827__;
  assign new_new_n1836__ = new_new_n1828__ & new_new_n1835__;
  assign new_new_n1837__ = new_new_n1833__ & new_new_n1834__;
  assign new_new_n1838__ = new_new_n1826__ & new_new_n1837__;
  assign new_new_n1839__ = new_new_n1836__ & new_new_n1838__;
  assign new_new_n1840__ = ~new_new_n353__ & ~new_new_n1210__;
  assign new_new_n1841__ = ~new_new_n1166__ & new_new_n1214__;
  assign new_new_n1842__ = ~new_new_n119__ & ~new_new_n511__;
  assign new_new_n1843__ = ~new_new_n276__ & new_new_n1842__;
  assign new_new_n1844__ = ~new_new_n306__ & new_new_n1843__;
  assign new_new_n1845__ = ~new_new_n809__ & new_new_n1844__;
  assign new_new_n1846__ = ~new_new_n130__ & ~new_new_n631__;
  assign new_new_n1847__ = ~new_new_n155__ & ~new_new_n488__;
  assign new_new_n1848__ = ~new_new_n348__ & ~new_new_n385__;
  assign new_new_n1849__ = ~new_new_n372__ & ~new_new_n1009__;
  assign new_new_n1850__ = ~new_new_n732__ & new_new_n1849__;
  assign new_new_n1851__ = ~new_new_n92__ & ~new_new_n242__;
  assign new_new_n1852__ = ~new_new_n313__ & ~new_new_n698__;
  assign new_new_n1853__ = ~new_new_n1034__ & new_new_n1852__;
  assign new_new_n1854__ = ~new_new_n816__ & new_new_n1851__;
  assign new_new_n1855__ = ~new_new_n993__ & new_new_n1854__;
  assign new_new_n1856__ = new_new_n1853__ & new_new_n1855__;
  assign new_new_n1857__ = new_new_n1850__ & new_new_n1856__;
  assign new_new_n1858__ = ~new_new_n375__ & ~new_new_n1081__;
  assign new_new_n1859__ = ~new_new_n213__ & ~new_new_n768__;
  assign new_new_n1860__ = ~new_new_n88__ & new_new_n1859__;
  assign new_new_n1861__ = new_new_n1450__ & new_new_n1860__;
  assign new_new_n1862__ = ~new_new_n192__ & ~new_new_n246__;
  assign new_new_n1863__ = ~new_new_n317__ & ~new_new_n602__;
  assign new_new_n1864__ = new_new_n1858__ & new_new_n1863__;
  assign new_new_n1865__ = new_new_n1661__ & new_new_n1862__;
  assign new_new_n1866__ = new_new_n1840__ & new_new_n1841__;
  assign new_new_n1867__ = new_new_n1846__ & new_new_n1847__;
  assign new_new_n1868__ = new_new_n1848__ & new_new_n1867__;
  assign new_new_n1869__ = new_new_n1865__ & new_new_n1866__;
  assign new_new_n1870__ = new_new_n1861__ & new_new_n1864__;
  assign new_new_n1871__ = new_new_n1869__ & new_new_n1870__;
  assign new_new_n1872__ = new_new_n1845__ & new_new_n1868__;
  assign new_new_n1873__ = new_new_n1871__ & new_new_n1872__;
  assign new_new_n1874__ = new_new_n1857__ & new_new_n1873__;
  assign new_new_n1875__ = ~new_new_n189__ & ~new_new_n585__;
  assign new_new_n1876__ = ~new_new_n120__ & ~new_new_n747__;
  assign new_new_n1877__ = new_new_n1606__ & new_new_n1876__;
  assign new_new_n1878__ = new_new_n946__ & new_new_n1875__;
  assign new_new_n1879__ = new_new_n1877__ & new_new_n1878__;
  assign new_new_n1880__ = ~new_new_n78__ & ~new_new_n718__;
  assign new_new_n1881__ = new_new_n153__ & ~new_new_n1880__;
  assign new_new_n1882__ = new_new_n1366__ & ~new_new_n1881__;
  assign new_new_n1883__ = new_new_n1517__ & new_new_n1882__;
  assign new_new_n1884__ = ~new_new_n696__ & ~new_new_n843__;
  assign new_new_n1885__ = ~new_new_n103__ & ~new_new_n198__;
  assign new_new_n1886__ = ~new_new_n168__ & ~new_new_n309__;
  assign new_new_n1887__ = ~new_new_n320__ & ~new_new_n670__;
  assign new_new_n1888__ = new_new_n898__ & ~new_new_n950__;
  assign new_new_n1889__ = new_new_n1886__ & new_new_n1887__;
  assign new_new_n1890__ = ~new_new_n150__ & ~new_new_n274__;
  assign new_new_n1891__ = ~new_new_n635__ & new_new_n1373__;
  assign new_new_n1892__ = new_new_n1890__ & new_new_n1891__;
  assign new_new_n1893__ = new_new_n1888__ & new_new_n1889__;
  assign new_new_n1894__ = new_new_n1710__ & new_new_n1884__;
  assign new_new_n1895__ = new_new_n1885__ & new_new_n1894__;
  assign new_new_n1896__ = new_new_n1892__ & new_new_n1893__;
  assign new_new_n1897__ = new_new_n1883__ & new_new_n1896__;
  assign new_new_n1898__ = new_new_n1879__ & new_new_n1895__;
  assign new_new_n1899__ = new_new_n1897__ & new_new_n1898__;
  assign new_new_n1900__ = new_new_n1839__ & new_new_n1899__;
  assign new_new_n1901__ = new_new_n1767__ & new_new_n1900__;
  assign new_new_n1902__ = new_new_n1874__ & new_new_n1901__;
  assign new_new_n1903__ = ~new_new_n127__ & ~new_new_n1094__;
  assign new_new_n1904__ = ~new_new_n88__ & ~new_new_n160__;
  assign new_new_n1905__ = ~new_new_n632__ & ~new_new_n1506__;
  assign new_new_n1906__ = ~new_new_n781__ & new_new_n1904__;
  assign new_new_n1907__ = new_new_n1905__ & new_new_n1906__;
  assign new_new_n1908__ = ~new_new_n1539__ & new_new_n1907__;
  assign new_new_n1909__ = ~new_new_n252__ & ~new_new_n425__;
  assign new_new_n1910__ = ~new_new_n212__ & ~new_new_n495__;
  assign new_new_n1911__ = ~new_new_n995__ & new_new_n1910__;
  assign new_new_n1912__ = ~new_new_n255__ & ~new_new_n1035__;
  assign new_new_n1913__ = new_new_n1903__ & new_new_n1909__;
  assign new_new_n1914__ = new_new_n1912__ & new_new_n1913__;
  assign new_new_n1915__ = new_new_n1911__ & new_new_n1914__;
  assign new_new_n1916__ = new_new_n1908__ & new_new_n1915__;
  assign new_new_n1917__ = ~new_new_n372__ & ~new_new_n783__;
  assign new_new_n1918__ = ~new_new_n179__ & ~new_new_n207__;
  assign new_new_n1919__ = ~new_new_n489__ & ~new_new_n1151__;
  assign new_new_n1920__ = ~new_new_n166__ & ~new_new_n309__;
  assign new_new_n1921__ = new_new_n162__ & ~new_new_n333__;
  assign new_new_n1922__ = ~new_new_n496__ & ~new_new_n586__;
  assign new_new_n1923__ = ~new_new_n247__ & ~new_new_n351__;
  assign new_new_n1924__ = ~new_new_n445__ & ~new_new_n937__;
  assign new_new_n1925__ = new_new_n1923__ & new_new_n1924__;
  assign new_new_n1926__ = new_new_n1922__ & new_new_n1925__;
  assign new_new_n1927__ = ~new_new_n630__ & new_new_n1926__;
  assign new_new_n1928__ = new_new_n1598__ & new_new_n1927__;
  assign new_new_n1929__ = ~new_new_n253__ & ~new_new_n327__;
  assign new_new_n1930__ = ~new_new_n282__ & ~new_new_n701__;
  assign new_new_n1931__ = ~new_new_n346__ & new_new_n1930__;
  assign new_new_n1932__ = new_new_n593__ & ~new_new_n952__;
  assign new_new_n1933__ = new_new_n1918__ & ~new_new_n1921__;
  assign new_new_n1934__ = new_new_n1929__ & new_new_n1933__;
  assign new_new_n1935__ = new_new_n1931__ & new_new_n1932__;
  assign new_new_n1936__ = new_new_n1917__ & new_new_n1919__;
  assign new_new_n1937__ = new_new_n1920__ & new_new_n1936__;
  assign new_new_n1938__ = new_new_n1934__ & new_new_n1935__;
  assign new_new_n1939__ = new_new_n1937__ & new_new_n1938__;
  assign new_new_n1940__ = new_new_n1916__ & new_new_n1939__;
  assign new_new_n1941__ = new_new_n1928__ & new_new_n1940__;
  assign new_new_n1942__ = ~new_new_n130__ & ~new_new_n692__;
  assign new_new_n1943__ = ~new_new_n286__ & ~new_new_n483__;
  assign new_new_n1944__ = ~new_new_n164__ & ~new_new_n996__;
  assign new_new_n1945__ = ~new_new_n263__ & ~new_new_n603__;
  assign new_new_n1946__ = ~new_new_n693__ & ~new_new_n1515__;
  assign new_new_n1947__ = ~new_new_n384__ & ~new_new_n595__;
  assign new_new_n1948__ = ~new_new_n76__ & ~new_new_n388__;
  assign new_new_n1949__ = ~new_new_n441__ & ~new_new_n584__;
  assign new_new_n1950__ = ~new_new_n597__ & ~new_new_n723__;
  assign new_new_n1951__ = ~new_new_n933__ & new_new_n1950__;
  assign new_new_n1952__ = new_new_n1948__ & new_new_n1949__;
  assign new_new_n1953__ = ~new_new_n591__ & new_new_n1946__;
  assign new_new_n1954__ = new_new_n1952__ & new_new_n1953__;
  assign new_new_n1955__ = ~new_new_n935__ & new_new_n1951__;
  assign new_new_n1956__ = new_new_n1945__ & new_new_n1947__;
  assign new_new_n1957__ = new_new_n1955__ & new_new_n1956__;
  assign new_new_n1958__ = ~new_new_n668__ & new_new_n1954__;
  assign new_new_n1959__ = new_new_n1957__ & new_new_n1958__;
  assign new_new_n1960__ = ~new_new_n251__ & ~new_new_n1007__;
  assign new_new_n1961__ = ~new_new_n192__ & ~new_new_n313__;
  assign new_new_n1962__ = new_new_n709__ & new_new_n1961__;
  assign new_new_n1963__ = new_new_n95__ & new_new_n1483__;
  assign new_new_n1964__ = new_new_n113__ & new_new_n126__;
  assign new_new_n1965__ = ~new_new_n1963__ & ~new_new_n1964__;
  assign new_new_n1966__ = ~pi24 & ~new_new_n1965__;
  assign new_new_n1967__ = ~new_new_n658__ & ~new_new_n1507__;
  assign new_new_n1968__ = ~new_new_n183__ & ~new_new_n283__;
  assign new_new_n1969__ = new_new_n1071__ & new_new_n1968__;
  assign new_new_n1970__ = ~new_new_n374__ & ~new_new_n945__;
  assign new_new_n1971__ = ~new_new_n198__ & ~new_new_n1212__;
  assign new_new_n1972__ = ~new_new_n119__ & ~new_new_n473__;
  assign new_new_n1973__ = ~new_new_n150__ & new_new_n1972__;
  assign new_new_n1974__ = new_new_n1971__ & new_new_n1973__;
  assign new_new_n1975__ = ~new_new_n274__ & ~new_new_n477__;
  assign new_new_n1976__ = ~new_new_n336__ & ~new_new_n950__;
  assign new_new_n1977__ = ~new_new_n721__ & new_new_n1976__;
  assign new_new_n1978__ = ~new_new_n816__ & ~new_new_n1073__;
  assign new_new_n1979__ = new_new_n1741__ & new_new_n1960__;
  assign new_new_n1980__ = new_new_n1978__ & new_new_n1979__;
  assign new_new_n1981__ = new_new_n1097__ & new_new_n1977__;
  assign new_new_n1982__ = new_new_n1230__ & new_new_n1252__;
  assign new_new_n1983__ = ~new_new_n1966__ & new_new_n1967__;
  assign new_new_n1984__ = new_new_n1970__ & new_new_n1975__;
  assign new_new_n1985__ = new_new_n1983__ & new_new_n1984__;
  assign new_new_n1986__ = new_new_n1981__ & new_new_n1982__;
  assign new_new_n1987__ = new_new_n1969__ & new_new_n1980__;
  assign new_new_n1988__ = new_new_n1974__ & new_new_n1987__;
  assign new_new_n1989__ = new_new_n1985__ & new_new_n1986__;
  assign new_new_n1990__ = new_new_n1962__ & new_new_n1989__;
  assign new_new_n1991__ = new_new_n1959__ & new_new_n1988__;
  assign new_new_n1992__ = new_new_n1990__ & new_new_n1991__;
  assign new_new_n1993__ = ~new_new_n566__ & ~new_new_n588__;
  assign new_new_n1994__ = ~new_new_n155__ & ~new_new_n1167__;
  assign new_new_n1995__ = ~new_new_n108__ & ~new_new_n189__;
  assign new_new_n1996__ = ~new_new_n202__ & new_new_n1645__;
  assign new_new_n1997__ = new_new_n1993__ & new_new_n1994__;
  assign new_new_n1998__ = new_new_n1995__ & new_new_n1997__;
  assign new_new_n1999__ = new_new_n1996__ & new_new_n1998__;
  assign new_new_n2000__ = ~new_new_n488__ & ~new_new_n657__;
  assign new_new_n2001__ = ~new_new_n246__ & ~new_new_n811__;
  assign new_new_n2002__ = ~new_new_n826__ & ~new_new_n1113__;
  assign new_new_n2003__ = ~new_new_n675__ & new_new_n2002__;
  assign new_new_n2004__ = ~new_new_n509__ & ~new_new_n828__;
  assign new_new_n2005__ = ~new_new_n768__ & ~new_new_n869__;
  assign new_new_n2006__ = ~new_new_n259__ & ~new_new_n637__;
  assign new_new_n2007__ = ~new_new_n427__ & new_new_n2006__;
  assign new_new_n2008__ = new_new_n967__ & new_new_n1069__;
  assign new_new_n2009__ = new_new_n1942__ & new_new_n1944__;
  assign new_new_n2010__ = new_new_n2001__ & new_new_n2009__;
  assign new_new_n2011__ = new_new_n2007__ & new_new_n2008__;
  assign new_new_n2012__ = new_new_n567__ & new_new_n941__;
  assign new_new_n2013__ = new_new_n1513__ & new_new_n1943__;
  assign new_new_n2014__ = new_new_n2000__ & new_new_n2003__;
  assign new_new_n2015__ = new_new_n2004__ & new_new_n2005__;
  assign new_new_n2016__ = new_new_n2014__ & new_new_n2015__;
  assign new_new_n2017__ = new_new_n2012__ & new_new_n2013__;
  assign new_new_n2018__ = new_new_n2010__ & new_new_n2011__;
  assign new_new_n2019__ = new_new_n2017__ & new_new_n2018__;
  assign new_new_n2020__ = new_new_n2016__ & new_new_n2019__;
  assign new_new_n2021__ = new_new_n1480__ & new_new_n1999__;
  assign new_new_n2022__ = new_new_n2020__ & new_new_n2021__;
  assign new_new_n2023__ = new_new_n1941__ & new_new_n2022__;
  assign new_new_n2024__ = new_new_n1992__ & new_new_n2023__;
  assign new_new_n2025__ = ~new_new_n276__ & ~new_new_n607__;
  assign new_new_n2026__ = ~new_new_n92__ & ~new_new_n1151__;
  assign new_new_n2027__ = ~new_new_n138__ & ~new_new_n242__;
  assign new_new_n2028__ = ~new_new_n1105__ & ~new_new_n1291__;
  assign new_new_n2029__ = ~new_new_n809__ & new_new_n2028__;
  assign new_new_n2030__ = ~new_new_n253__ & ~new_new_n260__;
  assign new_new_n2031__ = ~new_new_n630__ & new_new_n2030__;
  assign new_new_n2032__ = ~new_new_n284__ & ~new_new_n508__;
  assign new_new_n2033__ = ~new_new_n1081__ & ~new_new_n1176__;
  assign new_new_n2034__ = ~new_new_n198__ & ~new_new_n1007__;
  assign new_new_n2035__ = ~new_new_n200__ & ~new_new_n267__;
  assign new_new_n2036__ = ~new_new_n657__ & ~new_new_n1210__;
  assign new_new_n2037__ = new_new_n2035__ & new_new_n2036__;
  assign new_new_n2038__ = ~new_new_n286__ & ~new_new_n353__;
  assign new_new_n2039__ = ~new_new_n382__ & ~new_new_n732__;
  assign new_new_n2040__ = ~new_new_n842__ & ~new_new_n919__;
  assign new_new_n2041__ = new_new_n2039__ & new_new_n2040__;
  assign new_new_n2042__ = new_new_n2037__ & new_new_n2038__;
  assign new_new_n2043__ = ~new_new_n439__ & new_new_n1804__;
  assign new_new_n2044__ = ~new_new_n1966__ & new_new_n2034__;
  assign new_new_n2045__ = new_new_n2043__ & new_new_n2044__;
  assign new_new_n2046__ = new_new_n2041__ & new_new_n2042__;
  assign new_new_n2047__ = new_new_n2045__ & new_new_n2046__;
  assign new_new_n2048__ = ~new_new_n164__ & ~new_new_n385__;
  assign new_new_n2049__ = ~new_new_n1033__ & ~new_new_n1109__;
  assign new_new_n2050__ = new_new_n2048__ & new_new_n2049__;
  assign new_new_n2051__ = new_new_n474__ & new_new_n1740__;
  assign new_new_n2052__ = new_new_n2027__ & new_new_n2033__;
  assign new_new_n2053__ = new_new_n2051__ & new_new_n2052__;
  assign new_new_n2054__ = new_new_n1680__ & new_new_n2050__;
  assign new_new_n2055__ = new_new_n2026__ & new_new_n2054__;
  assign new_new_n2056__ = new_new_n2025__ & new_new_n2053__;
  assign new_new_n2057__ = new_new_n2031__ & new_new_n2032__;
  assign new_new_n2058__ = new_new_n2056__ & new_new_n2057__;
  assign new_new_n2059__ = new_new_n2029__ & new_new_n2055__;
  assign new_new_n2060__ = new_new_n2058__ & new_new_n2059__;
  assign new_new_n2061__ = new_new_n2047__ & new_new_n2060__;
  assign new_new_n2062__ = ~new_new_n263__ & new_new_n985__;
  assign new_new_n2063__ = new_new_n2061__ & new_new_n2062__;
  assign new_new_n2064__ = ~new_new_n350__ & ~new_new_n509__;
  assign new_new_n2065__ = ~new_new_n829__ & ~new_new_n1064__;
  assign new_new_n2066__ = ~new_new_n351__ & ~new_new_n483__;
  assign new_new_n2067__ = ~new_new_n209__ & ~new_new_n990__;
  assign new_new_n2068__ = ~new_new_n120__ & ~new_new_n441__;
  assign new_new_n2069__ = ~new_new_n247__ & ~new_new_n723__;
  assign new_new_n2070__ = ~new_new_n843__ & new_new_n2069__;
  assign new_new_n2071__ = new_new_n2067__ & new_new_n2068__;
  assign new_new_n2072__ = new_new_n2070__ & new_new_n2071__;
  assign new_new_n2073__ = new_new_n2064__ & new_new_n2065__;
  assign new_new_n2074__ = new_new_n2066__ & new_new_n2073__;
  assign new_new_n2075__ = new_new_n2072__ & new_new_n2074__;
  assign new_new_n2076__ = ~new_new_n329__ & ~new_new_n995__;
  assign new_new_n2077__ = ~new_new_n246__ & ~new_new_n947__;
  assign new_new_n2078__ = ~new_new_n312__ & ~new_new_n600__;
  assign new_new_n2079__ = ~new_new_n196__ & ~new_new_n693__;
  assign new_new_n2080__ = ~new_new_n127__ & ~new_new_n168__;
  assign new_new_n2081__ = ~new_new_n283__ & ~new_new_n327__;
  assign new_new_n2082__ = ~new_new_n715__ & ~new_new_n937__;
  assign new_new_n2083__ = new_new_n2081__ & new_new_n2082__;
  assign new_new_n2084__ = new_new_n2077__ & new_new_n2080__;
  assign new_new_n2085__ = new_new_n2078__ & new_new_n2079__;
  assign new_new_n2086__ = new_new_n2084__ & new_new_n2085__;
  assign new_new_n2087__ = new_new_n2076__ & new_new_n2083__;
  assign new_new_n2088__ = new_new_n2086__ & new_new_n2087__;
  assign new_new_n2089__ = ~new_new_n479__ & ~new_new_n884__;
  assign new_new_n2090__ = ~new_new_n282__ & ~new_new_n438__;
  assign new_new_n2091__ = new_new_n2089__ & new_new_n2090__;
  assign new_new_n2092__ = ~new_new_n373__ & ~new_new_n963__;
  assign new_new_n2093__ = ~new_new_n425__ & ~new_new_n875__;
  assign new_new_n2094__ = new_new_n80__ & new_new_n506__;
  assign new_new_n2095__ = ~new_new_n258__ & ~new_new_n656__;
  assign new_new_n2096__ = ~new_new_n921__ & new_new_n2095__;
  assign new_new_n2097__ = ~new_new_n2094__ & new_new_n2096__;
  assign new_new_n2098__ = ~new_new_n828__ & ~new_new_n835__;
  assign new_new_n2099__ = ~new_new_n315__ & ~new_new_n480__;
  assign new_new_n2100__ = ~new_new_n388__ & ~new_new_n445__;
  assign new_new_n2101__ = ~new_new_n700__ & ~new_new_n1343__;
  assign new_new_n2102__ = ~new_new_n202__ & new_new_n2101__;
  assign new_new_n2103__ = new_new_n337__ & new_new_n1449__;
  assign new_new_n2104__ = new_new_n1742__ & new_new_n1829__;
  assign new_new_n2105__ = new_new_n2099__ & new_new_n2100__;
  assign new_new_n2106__ = new_new_n2104__ & new_new_n2105__;
  assign new_new_n2107__ = new_new_n2102__ & new_new_n2103__;
  assign new_new_n2108__ = new_new_n490__ & new_new_n2098__;
  assign new_new_n2109__ = new_new_n2107__ & new_new_n2108__;
  assign new_new_n2110__ = new_new_n839__ & new_new_n2106__;
  assign new_new_n2111__ = new_new_n936__ & new_new_n1749__;
  assign new_new_n2112__ = new_new_n2110__ & new_new_n2111__;
  assign new_new_n2113__ = new_new_n1908__ & new_new_n2109__;
  assign new_new_n2114__ = new_new_n2097__ & new_new_n2113__;
  assign new_new_n2115__ = new_new_n2112__ & new_new_n2114__;
  assign new_new_n2116__ = ~new_new_n76__ & ~new_new_n476__;
  assign new_new_n2117__ = ~new_new_n313__ & ~new_new_n637__;
  assign new_new_n2118__ = ~new_new_n719__ & new_new_n2117__;
  assign new_new_n2119__ = ~new_new_n993__ & new_new_n2093__;
  assign new_new_n2120__ = new_new_n2116__ & new_new_n2119__;
  assign new_new_n2121__ = ~new_new_n254__ & new_new_n2118__;
  assign new_new_n2122__ = new_new_n1114__ & new_new_n1310__;
  assign new_new_n2123__ = new_new_n2121__ & new_new_n2122__;
  assign new_new_n2124__ = new_new_n2092__ & new_new_n2120__;
  assign new_new_n2125__ = new_new_n2123__ & new_new_n2124__;
  assign new_new_n2126__ = new_new_n2088__ & new_new_n2091__;
  assign new_new_n2127__ = new_new_n2125__ & new_new_n2126__;
  assign new_new_n2128__ = new_new_n2075__ & new_new_n2127__;
  assign new_new_n2129__ = new_new_n2115__ & new_new_n2128__;
  assign new_new_n2130__ = new_new_n2063__ & new_new_n2129__;
  assign new_new_n2131__ = ~new_new_n266__ & ~new_new_n719__;
  assign new_new_n2132__ = ~new_new_n657__ & ~new_new_n1217__;
  assign new_new_n2133__ = ~new_new_n676__ & new_new_n2132__;
  assign new_new_n2134__ = ~new_new_n380__ & ~new_new_n635__;
  assign new_new_n2135__ = ~new_new_n1701__ & new_new_n2134__;
  assign new_new_n2136__ = ~new_new_n479__ & new_new_n484__;
  assign new_new_n2137__ = new_new_n1707__ & new_new_n2131__;
  assign new_new_n2138__ = new_new_n2136__ & new_new_n2137__;
  assign new_new_n2139__ = new_new_n2133__ & new_new_n2135__;
  assign new_new_n2140__ = new_new_n2138__ & new_new_n2139__;
  assign new_new_n2141__ = new_new_n217__ & ~new_new_n598__;
  assign new_new_n2142__ = ~new_new_n166__ & new_new_n1424__;
  assign new_new_n2143__ = ~new_new_n155__ & ~new_new_n229__;
  assign new_new_n2144__ = ~new_new_n189__ & new_new_n2143__;
  assign new_new_n2145__ = ~new_new_n179__ & ~new_new_n286__;
  assign new_new_n2146__ = ~new_new_n673__ & ~new_new_n940__;
  assign new_new_n2147__ = ~new_new_n842__ & new_new_n1449__;
  assign new_new_n2148__ = ~new_new_n2141__ & new_new_n2147__;
  assign new_new_n2149__ = new_new_n744__ & new_new_n2146__;
  assign new_new_n2150__ = new_new_n1143__ & new_new_n1153__;
  assign new_new_n2151__ = ~new_new_n1966__ & new_new_n2142__;
  assign new_new_n2152__ = new_new_n2145__ & new_new_n2151__;
  assign new_new_n2153__ = new_new_n2149__ & new_new_n2150__;
  assign new_new_n2154__ = new_new_n2144__ & new_new_n2148__;
  assign new_new_n2155__ = new_new_n2153__ & new_new_n2154__;
  assign new_new_n2156__ = new_new_n2152__ & new_new_n2155__;
  assign new_new_n2157__ = new_new_n2140__ & new_new_n2156__;
  assign new_new_n2158__ = ~new_new_n351__ & ~new_new_n1372__;
  assign new_new_n2159__ = ~new_new_n477__ & ~new_new_n510__;
  assign new_new_n2160__ = ~new_new_n851__ & ~new_new_n990__;
  assign new_new_n2161__ = ~new_new_n637__ & ~new_new_n781__;
  assign new_new_n2162__ = ~new_new_n108__ & ~new_new_n385__;
  assign new_new_n2163__ = ~new_new_n1343__ & new_new_n2162__;
  assign new_new_n2164__ = ~new_new_n183__ & ~new_new_n1506__;
  assign new_new_n2165__ = new_new_n2163__ & new_new_n2164__;
  assign new_new_n2166__ = ~new_new_n335__ & ~new_new_n698__;
  assign new_new_n2167__ = ~new_new_n103__ & ~new_new_n874__;
  assign new_new_n2168__ = ~new_new_n212__ & ~new_new_n280__;
  assign new_new_n2169__ = ~new_new_n232__ & ~new_new_n1003__;
  assign new_new_n2170__ = new_new_n221__ & new_new_n234__;
  assign new_new_n2171__ = ~new_new_n890__ & ~new_new_n2170__;
  assign new_new_n2172__ = new_new_n2168__ & new_new_n2171__;
  assign new_new_n2173__ = new_new_n2169__ & new_new_n2172__;
  assign new_new_n2174__ = ~new_new_n597__ & ~new_new_n896__;
  assign new_new_n2175__ = ~new_new_n322__ & ~new_new_n473__;
  assign new_new_n2176__ = ~new_new_n120__ & ~new_new_n282__;
  assign new_new_n2177__ = ~new_new_n238__ & new_new_n2174__;
  assign new_new_n2178__ = new_new_n2176__ & new_new_n2177__;
  assign new_new_n2179__ = ~new_new_n809__ & new_new_n1487__;
  assign new_new_n2180__ = new_new_n2175__ & new_new_n2179__;
  assign new_new_n2181__ = new_new_n2178__ & new_new_n2180__;
  assign new_new_n2182__ = ~new_new_n76__ & ~new_new_n509__;
  assign new_new_n2183__ = ~new_new_n600__ & new_new_n2182__;
  assign new_new_n2184__ = ~new_new_n963__ & ~new_new_n1210__;
  assign new_new_n2185__ = ~new_new_n150__ & new_new_n2184__;
  assign new_new_n2186__ = ~new_new_n588__ & ~new_new_n1167__;
  assign new_new_n2187__ = new_new_n2166__ & new_new_n2186__;
  assign new_new_n2188__ = ~new_new_n935__ & new_new_n2185__;
  assign new_new_n2189__ = new_new_n2161__ & new_new_n2167__;
  assign new_new_n2190__ = new_new_n2183__ & new_new_n2189__;
  assign new_new_n2191__ = new_new_n2187__ & new_new_n2188__;
  assign new_new_n2192__ = new_new_n2165__ & new_new_n2191__;
  assign new_new_n2193__ = new_new_n2173__ & new_new_n2190__;
  assign new_new_n2194__ = new_new_n2192__ & new_new_n2193__;
  assign new_new_n2195__ = new_new_n2181__ & new_new_n2194__;
  assign new_new_n2196__ = ~new_new_n336__ & ~new_new_n871__;
  assign new_new_n2197__ = ~new_new_n828__ & ~new_new_n1398__;
  assign new_new_n2198__ = ~new_new_n200__ & ~new_new_n947__;
  assign new_new_n2199__ = ~new_new_n255__ & new_new_n2198__;
  assign new_new_n2200__ = ~new_new_n869__ & new_new_n2199__;
  assign new_new_n2201__ = new_new_n2197__ & new_new_n2200__;
  assign new_new_n2202__ = ~new_new_n441__ & ~new_new_n1507__;
  assign new_new_n2203__ = ~new_new_n1064__ & ~new_new_n1113__;
  assign new_new_n2204__ = new_new_n2202__ & new_new_n2203__;
  assign new_new_n2205__ = ~new_new_n445__ & ~new_new_n603__;
  assign new_new_n2206__ = ~new_new_n1176__ & new_new_n2205__;
  assign new_new_n2207__ = ~new_new_n321__ & ~new_new_n353__;
  assign new_new_n2208__ = ~new_new_n774__ & new_new_n827__;
  assign new_new_n2209__ = new_new_n1213__ & new_new_n1367__;
  assign new_new_n2210__ = new_new_n2158__ & new_new_n2160__;
  assign new_new_n2211__ = new_new_n2209__ & new_new_n2210__;
  assign new_new_n2212__ = new_new_n2207__ & new_new_n2208__;
  assign new_new_n2213__ = ~new_new_n373__ & new_new_n2206__;
  assign new_new_n2214__ = ~new_new_n837__ & new_new_n1078__;
  assign new_new_n2215__ = new_new_n2159__ & new_new_n2196__;
  assign new_new_n2216__ = new_new_n2214__ & new_new_n2215__;
  assign new_new_n2217__ = new_new_n2212__ & new_new_n2213__;
  assign new_new_n2218__ = new_new_n2204__ & new_new_n2211__;
  assign new_new_n2219__ = new_new_n2217__ & new_new_n2218__;
  assign new_new_n2220__ = new_new_n2201__ & new_new_n2216__;
  assign new_new_n2221__ = new_new_n2219__ & new_new_n2220__;
  assign new_new_n2222__ = new_new_n1421__ & new_new_n2221__;
  assign new_new_n2223__ = new_new_n2157__ & new_new_n2222__;
  assign new_new_n2224__ = new_new_n2195__ & new_new_n2223__;
  assign new_new_n2225__ = ~new_new_n2130__ & ~new_new_n2224__;
  assign new_new_n2226__ = ~new_new_n258__ & ~new_new_n1506__;
  assign new_new_n2227__ = ~new_new_n260__ & ~new_new_n473__;
  assign new_new_n2228__ = ~new_new_n846__ & ~new_new_n1291__;
  assign new_new_n2229__ = new_new_n2227__ & new_new_n2228__;
  assign new_new_n2230__ = ~new_new_n276__ & ~new_new_n332__;
  assign new_new_n2231__ = new_new_n799__ & new_new_n2230__;
  assign new_new_n2232__ = new_new_n2229__ & new_new_n2231__;
  assign new_new_n2233__ = ~new_new_n425__ & ~new_new_n851__;
  assign new_new_n2234__ = ~new_new_n778__ & ~new_new_n1081__;
  assign new_new_n2235__ = ~new_new_n694__ & ~new_new_n894__;
  assign new_new_n2236__ = ~new_new_n266__ & ~new_new_n631__;
  assign new_new_n2237__ = new_new_n1918__ & new_new_n2233__;
  assign new_new_n2238__ = new_new_n2234__ & new_new_n2237__;
  assign new_new_n2239__ = ~new_new_n373__ & new_new_n1142__;
  assign new_new_n2240__ = new_new_n1636__ & new_new_n2235__;
  assign new_new_n2241__ = new_new_n2236__ & new_new_n2240__;
  assign new_new_n2242__ = new_new_n2238__ & new_new_n2239__;
  assign new_new_n2243__ = new_new_n2241__ & new_new_n2242__;
  assign new_new_n2244__ = ~new_new_n198__ & ~new_new_n1109__;
  assign new_new_n2245__ = ~new_new_n202__ & new_new_n672__;
  assign new_new_n2246__ = new_new_n710__ & new_new_n948__;
  assign new_new_n2247__ = new_new_n1333__ & new_new_n2246__;
  assign new_new_n2248__ = new_new_n2244__ & new_new_n2245__;
  assign new_new_n2249__ = ~new_new_n508__ & new_new_n592__;
  assign new_new_n2250__ = new_new_n1153__ & new_new_n2226__;
  assign new_new_n2251__ = new_new_n2249__ & new_new_n2250__;
  assign new_new_n2252__ = new_new_n2247__ & new_new_n2248__;
  assign new_new_n2253__ = new_new_n2251__ & new_new_n2252__;
  assign new_new_n2254__ = new_new_n2232__ & new_new_n2253__;
  assign new_new_n2255__ = new_new_n2243__ & new_new_n2254__;
  assign new_new_n2256__ = ~new_new_n232__ & ~new_new_n263__;
  assign new_new_n2257__ = new_new_n2255__ & new_new_n2256__;
  assign new_new_n2258__ = ~new_new_n300__ & ~new_new_n940__;
  assign new_new_n2259__ = ~new_new_n632__ & ~new_new_n884__;
  assign new_new_n2260__ = ~new_new_n96__ & ~new_new_n242__;
  assign new_new_n2261__ = ~new_new_n246__ & ~new_new_n717__;
  assign new_new_n2262__ = ~new_new_n843__ & new_new_n2261__;
  assign new_new_n2263__ = ~new_new_n348__ & new_new_n2260__;
  assign new_new_n2264__ = new_new_n2262__ & new_new_n2263__;
  assign new_new_n2265__ = ~new_new_n88__ & ~new_new_n939__;
  assign new_new_n2266__ = ~new_new_n890__ & ~new_new_n921__;
  assign new_new_n2267__ = ~new_new_n298__ & ~new_new_n723__;
  assign new_new_n2268__ = ~new_new_n302__ & ~new_new_n853__;
  assign new_new_n2269__ = ~new_new_n336__ & ~new_new_n701__;
  assign new_new_n2270__ = ~new_new_n990__ & new_new_n2269__;
  assign new_new_n2271__ = new_new_n2268__ & new_new_n2270__;
  assign new_new_n2272__ = ~new_new_n200__ & ~new_new_n284__;
  assign new_new_n2273__ = ~new_new_n724__ & ~new_new_n937__;
  assign new_new_n2274__ = ~new_new_n995__ & new_new_n2273__;
  assign new_new_n2275__ = ~new_new_n155__ & new_new_n2272__;
  assign new_new_n2276__ = ~new_new_n277__ & ~new_new_n311__;
  assign new_new_n2277__ = ~new_new_n673__ & ~new_new_n721__;
  assign new_new_n2278__ = new_new_n1284__ & new_new_n2267__;
  assign new_new_n2279__ = new_new_n2277__ & new_new_n2278__;
  assign new_new_n2280__ = new_new_n2275__ & new_new_n2276__;
  assign new_new_n2281__ = new_new_n2265__ & new_new_n2274__;
  assign new_new_n2282__ = new_new_n2266__ & new_new_n2281__;
  assign new_new_n2283__ = new_new_n2279__ & new_new_n2280__;
  assign new_new_n2284__ = new_new_n2271__ & new_new_n2283__;
  assign new_new_n2285__ = new_new_n2282__ & new_new_n2284__;
  assign new_new_n2286__ = new_new_n1605__ & new_new_n2285__;
  assign new_new_n2287__ = ~new_new_n82__ & ~new_new_n445__;
  assign new_new_n2288__ = ~new_new_n327__ & ~new_new_n950__;
  assign new_new_n2289__ = ~new_new_n382__ & ~new_new_n829__;
  assign new_new_n2290__ = ~new_new_n315__ & ~new_new_n959__;
  assign new_new_n2291__ = ~new_new_n482__ & ~new_new_n772__;
  assign new_new_n2292__ = ~new_new_n842__ & new_new_n2291__;
  assign new_new_n2293__ = new_new_n2287__ & new_new_n2288__;
  assign new_new_n2294__ = new_new_n2292__ & new_new_n2293__;
  assign new_new_n2295__ = new_new_n1680__ & new_new_n2289__;
  assign new_new_n2296__ = new_new_n2290__ & new_new_n2295__;
  assign new_new_n2297__ = new_new_n228__ & new_new_n2294__;
  assign new_new_n2298__ = new_new_n2296__ & new_new_n2297__;
  assign new_new_n2299__ = ~new_new_n255__ & new_new_n1373__;
  assign new_new_n2300__ = new_new_n167__ & new_new_n2299__;
  assign new_new_n2301__ = new_new_n944__ & new_new_n1097__;
  assign new_new_n2302__ = new_new_n1292__ & new_new_n1633__;
  assign new_new_n2303__ = new_new_n1645__ & new_new_n2258__;
  assign new_new_n2304__ = new_new_n2259__ & new_new_n2303__;
  assign new_new_n2305__ = new_new_n2301__ & new_new_n2302__;
  assign new_new_n2306__ = ~new_new_n1539__ & new_new_n2300__;
  assign new_new_n2307__ = new_new_n2264__ & new_new_n2306__;
  assign new_new_n2308__ = new_new_n2304__ & new_new_n2305__;
  assign new_new_n2309__ = new_new_n2307__ & new_new_n2308__;
  assign new_new_n2310__ = new_new_n988__ & new_new_n2298__;
  assign new_new_n2311__ = new_new_n2309__ & new_new_n2310__;
  assign new_new_n2312__ = new_new_n2286__ & new_new_n2311__;
  assign new_new_n2313__ = new_new_n2257__ & new_new_n2312__;
  assign new_new_n2314__ = ~new_new_n441__ & ~new_new_n2170__;
  assign new_new_n2315__ = ~new_new_n251__ & ~new_new_n676__;
  assign new_new_n2316__ = ~new_new_n202__ & ~new_new_n259__;
  assign new_new_n2317__ = ~new_new_n388__ & ~new_new_n846__;
  assign new_new_n2318__ = ~new_new_n263__ & new_new_n2317__;
  assign new_new_n2319__ = new_new_n2314__ & new_new_n2318__;
  assign new_new_n2320__ = new_new_n2316__ & new_new_n2319__;
  assign new_new_n2321__ = new_new_n2315__ & new_new_n2320__;
  assign new_new_n2322__ = ~new_new_n842__ & ~new_new_n869__;
  assign new_new_n2323__ = ~new_new_n96__ & new_new_n2322__;
  assign new_new_n2324__ = ~new_new_n747__ & ~new_new_n772__;
  assign new_new_n2325__ = ~new_new_n327__ & ~new_new_n656__;
  assign new_new_n2326__ = new_new_n1004__ & new_new_n2325__;
  assign new_new_n2327__ = new_new_n2324__ & new_new_n2326__;
  assign new_new_n2328__ = ~new_new_n165__ & ~new_new_n718__;
  assign new_new_n2329__ = new_new_n241__ & ~new_new_n2328__;
  assign new_new_n2330__ = ~new_new_n229__ & ~new_new_n375__;
  assign new_new_n2331__ = ~new_new_n584__ & ~new_new_n894__;
  assign new_new_n2332__ = ~new_new_n723__ & ~new_new_n1212__;
  assign new_new_n2333__ = ~new_new_n253__ & ~new_new_n313__;
  assign new_new_n2334__ = ~new_new_n939__ & ~new_new_n940__;
  assign new_new_n2335__ = ~new_new_n602__ & ~new_new_n632__;
  assign new_new_n2336__ = ~new_new_n286__ & ~new_new_n372__;
  assign new_new_n2337__ = ~new_new_n315__ & ~new_new_n1151__;
  assign new_new_n2338__ = ~new_new_n316__ & new_new_n2337__;
  assign new_new_n2339__ = new_new_n1084__ & new_new_n2338__;
  assign new_new_n2340__ = ~new_new_n179__ & ~new_new_n1080__;
  assign new_new_n2341__ = ~new_new_n874__ & ~new_new_n921__;
  assign new_new_n2342__ = ~new_new_n160__ & ~new_new_n509__;
  assign new_new_n2343__ = ~new_new_n895__ & ~new_new_n963__;
  assign new_new_n2344__ = new_new_n163__ & ~new_new_n355__;
  assign new_new_n2345__ = ~new_new_n267__ & ~new_new_n309__;
  assign new_new_n2346__ = ~new_new_n488__ & new_new_n2345__;
  assign new_new_n2347__ = ~new_new_n945__ & new_new_n2342__;
  assign new_new_n2348__ = ~new_new_n2344__ & new_new_n2347__;
  assign new_new_n2349__ = ~new_new_n479__ & new_new_n2346__;
  assign new_new_n2350__ = new_new_n1394__ & new_new_n1705__;
  assign new_new_n2351__ = new_new_n2003__ & new_new_n2350__;
  assign new_new_n2352__ = new_new_n2348__ & new_new_n2349__;
  assign new_new_n2353__ = new_new_n2351__ & new_new_n2352__;
  assign new_new_n2354__ = new_new_n2343__ & new_new_n2353__;
  assign new_new_n2355__ = ~new_new_n425__ & ~new_new_n671__;
  assign new_new_n2356__ = ~new_new_n226__ & new_new_n2355__;
  assign new_new_n2357__ = new_new_n1169__ & new_new_n2340__;
  assign new_new_n2358__ = new_new_n2356__ & new_new_n2357__;
  assign new_new_n2359__ = new_new_n2334__ & new_new_n2335__;
  assign new_new_n2360__ = new_new_n2336__ & new_new_n2341__;
  assign new_new_n2361__ = new_new_n2359__ & new_new_n2360__;
  assign new_new_n2362__ = new_new_n1369__ & new_new_n2358__;
  assign new_new_n2363__ = new_new_n2361__ & new_new_n2362__;
  assign new_new_n2364__ = new_new_n708__ & new_new_n2339__;
  assign new_new_n2365__ = new_new_n2363__ & new_new_n2364__;
  assign new_new_n2366__ = new_new_n2354__ & new_new_n2365__;
  assign new_new_n2367__ = ~new_new_n103__ & ~new_new_n995__;
  assign new_new_n2368__ = ~new_new_n1033__ & new_new_n2367__;
  assign new_new_n2369__ = ~new_new_n719__ & new_new_n750__;
  assign new_new_n2370__ = new_new_n2332__ & new_new_n2333__;
  assign new_new_n2371__ = new_new_n2369__ & new_new_n2370__;
  assign new_new_n2372__ = ~new_new_n124__ & new_new_n2368__;
  assign new_new_n2373__ = new_new_n2331__ & new_new_n2372__;
  assign new_new_n2374__ = new_new_n2371__ & new_new_n2373__;
  assign new_new_n2375__ = new_new_n2366__ & new_new_n2374__;
  assign new_new_n2376__ = ~new_new_n280__ & ~new_new_n843__;
  assign new_new_n2377__ = ~new_new_n120__ & ~new_new_n198__;
  assign new_new_n2378__ = ~new_new_n183__ & ~new_new_n1291__;
  assign new_new_n2379__ = ~new_new_n1009__ & ~new_new_n1070__;
  assign new_new_n2380__ = ~new_new_n82__ & new_new_n2378__;
  assign new_new_n2381__ = new_new_n2379__ & new_new_n2380__;
  assign new_new_n2382__ = ~new_new_n321__ & ~new_new_n1162__;
  assign new_new_n2383__ = ~new_new_n271__ & ~new_new_n729__;
  assign new_new_n2384__ = ~new_new_n1176__ & new_new_n1423__;
  assign new_new_n2385__ = ~new_new_n255__ & ~new_new_n597__;
  assign new_new_n2386__ = ~new_new_n312__ & ~new_new_n322__;
  assign new_new_n2387__ = new_new_n2385__ & new_new_n2386__;
  assign new_new_n2388__ = ~new_new_n624__ & ~new_new_n776__;
  assign new_new_n2389__ = ~new_new_n851__ & ~new_new_n937__;
  assign new_new_n2390__ = new_new_n2388__ & new_new_n2389__;
  assign new_new_n2391__ = ~new_new_n353__ & ~new_new_n673__;
  assign new_new_n2392__ = ~new_new_n878__ & new_new_n2383__;
  assign new_new_n2393__ = new_new_n2391__ & new_new_n2392__;
  assign new_new_n2394__ = new_new_n2065__ & new_new_n2390__;
  assign new_new_n2395__ = new_new_n2376__ & new_new_n2377__;
  assign new_new_n2396__ = new_new_n2382__ & new_new_n2384__;
  assign new_new_n2397__ = new_new_n2395__ & new_new_n2396__;
  assign new_new_n2398__ = new_new_n2393__ & new_new_n2394__;
  assign new_new_n2399__ = new_new_n2387__ & new_new_n2398__;
  assign new_new_n2400__ = new_new_n159__ & new_new_n2397__;
  assign new_new_n2401__ = new_new_n2381__ & new_new_n2400__;
  assign new_new_n2402__ = new_new_n2399__ & new_new_n2401__;
  assign new_new_n2403__ = new_new_n114__ & ~new_new_n1700__;
  assign new_new_n2404__ = ~new_new_n838__ & ~new_new_n947__;
  assign new_new_n2405__ = ~new_new_n306__ & ~new_new_n715__;
  assign new_new_n2406__ = ~new_new_n721__ & ~new_new_n835__;
  assign new_new_n2407__ = ~new_new_n1073__ & new_new_n1368__;
  assign new_new_n2408__ = ~new_new_n2329__ & new_new_n2330__;
  assign new_new_n2409__ = new_new_n2404__ & new_new_n2408__;
  assign new_new_n2410__ = new_new_n2406__ & new_new_n2407__;
  assign new_new_n2411__ = ~new_new_n439__ & new_new_n2405__;
  assign new_new_n2412__ = new_new_n1712__ & ~new_new_n2403__;
  assign new_new_n2413__ = new_new_n2411__ & new_new_n2412__;
  assign new_new_n2414__ = new_new_n2409__ & new_new_n2410__;
  assign new_new_n2415__ = new_new_n2323__ & new_new_n2414__;
  assign new_new_n2416__ = new_new_n2327__ & new_new_n2413__;
  assign new_new_n2417__ = new_new_n2415__ & new_new_n2416__;
  assign new_new_n2418__ = new_new_n2321__ & new_new_n2417__;
  assign new_new_n2419__ = new_new_n2402__ & new_new_n2418__;
  assign new_new_n2420__ = new_new_n2375__ & new_new_n2419__;
  assign new_new_n2421__ = new_new_n2313__ & new_new_n2420__;
  assign new_new_n2422__ = new_new_n2225__ & ~new_new_n2421__;
  assign new_new_n2423__ = new_new_n2024__ & ~new_new_n2422__;
  assign new_new_n2424__ = ~new_new_n286__ & ~new_new_n477__;
  assign new_new_n2425__ = ~new_new_n482__ & ~new_new_n996__;
  assign new_new_n2426__ = ~new_new_n441__ & ~new_new_n853__;
  assign new_new_n2427__ = ~new_new_n249__ & ~new_new_n1507__;
  assign new_new_n2428__ = ~new_new_n271__ & ~new_new_n935__;
  assign new_new_n2429__ = ~new_new_n877__ & ~new_new_n921__;
  assign new_new_n2430__ = new_new_n2428__ & new_new_n2429__;
  assign new_new_n2431__ = ~new_new_n242__ & ~new_new_n588__;
  assign new_new_n2432__ = new_new_n2001__ & new_new_n2426__;
  assign new_new_n2433__ = new_new_n2431__ & new_new_n2432__;
  assign new_new_n2434__ = ~new_new_n1966__ & new_new_n2427__;
  assign new_new_n2435__ = new_new_n2433__ & new_new_n2434__;
  assign new_new_n2436__ = new_new_n1704__ & new_new_n2435__;
  assign new_new_n2437__ = new_new_n2430__ & new_new_n2436__;
  assign new_new_n2438__ = ~new_new_n247__ & ~new_new_n698__;
  assign new_new_n2439__ = ~new_new_n1398__ & new_new_n2438__;
  assign new_new_n2440__ = ~new_new_n160__ & ~new_new_n379__;
  assign new_new_n2441__ = ~new_new_n656__ & new_new_n2440__;
  assign new_new_n2442__ = ~new_new_n874__ & ~new_new_n918__;
  assign new_new_n2443__ = ~new_new_n1073__ & new_new_n2425__;
  assign new_new_n2444__ = new_new_n2442__ & new_new_n2443__;
  assign new_new_n2445__ = new_new_n769__ & new_new_n2441__;
  assign new_new_n2446__ = new_new_n1743__ & new_new_n1947__;
  assign new_new_n2447__ = new_new_n2424__ & new_new_n2439__;
  assign new_new_n2448__ = new_new_n2446__ & new_new_n2447__;
  assign new_new_n2449__ = new_new_n2444__ & new_new_n2445__;
  assign new_new_n2450__ = new_new_n2448__ & new_new_n2449__;
  assign new_new_n2451__ = new_new_n841__ & new_new_n2450__;
  assign new_new_n2452__ = new_new_n2437__ & new_new_n2451__;
  assign new_new_n2453__ = ~new_new_n235__ & ~new_new_n276__;
  assign new_new_n2454__ = ~new_new_n1151__ & ~new_new_n1217__;
  assign new_new_n2455__ = ~new_new_n635__ & ~new_new_n1080__;
  assign new_new_n2456__ = ~new_new_n96__ & ~new_new_n308__;
  assign new_new_n2457__ = ~new_new_n776__ & new_new_n2456__;
  assign new_new_n2458__ = new_new_n659__ & ~new_new_n884__;
  assign new_new_n2459__ = new_new_n2457__ & new_new_n2458__;
  assign new_new_n2460__ = new_new_n1680__ & new_new_n1945__;
  assign new_new_n2461__ = new_new_n2453__ & new_new_n2454__;
  assign new_new_n2462__ = new_new_n2455__ & new_new_n2461__;
  assign new_new_n2463__ = new_new_n2459__ & new_new_n2460__;
  assign new_new_n2464__ = new_new_n2462__ & new_new_n2463__;
  assign new_new_n2465__ = ~new_new_n332__ & ~new_new_n472__;
  assign new_new_n2466__ = new_new_n763__ & new_new_n2465__;
  assign new_new_n2467__ = ~new_new_n382__ & ~new_new_n896__;
  assign new_new_n2468__ = ~new_new_n209__ & ~new_new_n425__;
  assign new_new_n2469__ = ~new_new_n374__ & ~new_new_n1009__;
  assign new_new_n2470__ = ~new_new_n952__ & ~new_new_n1035__;
  assign new_new_n2471__ = ~new_new_n785__ & ~new_new_n945__;
  assign new_new_n2472__ = ~new_new_n1506__ & new_new_n2468__;
  assign new_new_n2473__ = new_new_n2471__ & new_new_n2472__;
  assign new_new_n2474__ = new_new_n2469__ & new_new_n2470__;
  assign new_new_n2475__ = new_new_n2473__ & new_new_n2474__;
  assign new_new_n2476__ = ~new_new_n138__ & ~new_new_n489__;
  assign new_new_n2477__ = ~new_new_n335__ & ~new_new_n1109__;
  assign new_new_n2478__ = ~new_new_n488__ & ~new_new_n1105__;
  assign new_new_n2479__ = ~new_new_n88__ & ~new_new_n1210__;
  assign new_new_n2480__ = ~new_new_n676__ & ~new_new_n774__;
  assign new_new_n2481__ = ~new_new_n266__ & ~new_new_n311__;
  assign new_new_n2482__ = ~new_new_n869__ & ~new_new_n1167__;
  assign new_new_n2483__ = new_new_n1711__ & new_new_n2160__;
  assign new_new_n2484__ = new_new_n2477__ & new_new_n2479__;
  assign new_new_n2485__ = new_new_n2483__ & new_new_n2484__;
  assign new_new_n2486__ = new_new_n2481__ & new_new_n2482__;
  assign new_new_n2487__ = new_new_n1155__ & new_new_n1326__;
  assign new_new_n2488__ = new_new_n2467__ & new_new_n2476__;
  assign new_new_n2489__ = new_new_n2487__ & new_new_n2488__;
  assign new_new_n2490__ = new_new_n2485__ & new_new_n2486__;
  assign new_new_n2491__ = new_new_n2478__ & new_new_n2480__;
  assign new_new_n2492__ = new_new_n2490__ & new_new_n2491__;
  assign new_new_n2493__ = new_new_n2475__ & new_new_n2489__;
  assign new_new_n2494__ = new_new_n2492__ & new_new_n2493__;
  assign new_new_n2495__ = new_new_n2464__ & new_new_n2494__;
  assign new_new_n2496__ = new_new_n2452__ & new_new_n2495__;
  assign new_new_n2497__ = new_new_n2466__ & new_new_n2496__;
  assign new_new_n2498__ = ~new_new_n2313__ & ~new_new_n2497__;
  assign new_new_n2499__ = ~new_new_n302__ & ~new_new_n939__;
  assign new_new_n2500__ = ~new_new_n308__ & ~new_new_n940__;
  assign new_new_n2501__ = ~new_new_n635__ & ~new_new_n838__;
  assign new_new_n2502__ = pi24 & ~new_new_n152__;
  assign new_new_n2503__ = ~new_new_n73__ & ~new_new_n2502__;
  assign new_new_n2504__ = new_new_n268__ & new_new_n2503__;
  assign new_new_n2505__ = ~new_new_n374__ & ~new_new_n696__;
  assign new_new_n2506__ = ~new_new_n252__ & ~new_new_n845__;
  assign new_new_n2507__ = ~new_new_n385__ & ~new_new_n1507__;
  assign new_new_n2508__ = ~new_new_n1212__ & ~new_new_n1217__;
  assign new_new_n2509__ = ~new_new_n232__ & ~new_new_n1162__;
  assign new_new_n2510__ = new_new_n1740__ & new_new_n2506__;
  assign new_new_n2511__ = new_new_n2509__ & new_new_n2510__;
  assign new_new_n2512__ = new_new_n2505__ & new_new_n2507__;
  assign new_new_n2513__ = new_new_n2508__ & new_new_n2512__;
  assign new_new_n2514__ = new_new_n2511__ & new_new_n2513__;
  assign new_new_n2515__ = ~new_new_n489__ & ~new_new_n496__;
  assign new_new_n2516__ = ~new_new_n248__ & ~new_new_n826__;
  assign new_new_n2517__ = new_new_n951__ & new_new_n2516__;
  assign new_new_n2518__ = new_new_n2515__ & new_new_n2517__;
  assign new_new_n2519__ = ~new_new_n200__ & ~new_new_n694__;
  assign new_new_n2520__ = ~new_new_n346__ & new_new_n2519__;
  assign new_new_n2521__ = ~new_new_n828__ & ~new_new_n842__;
  assign new_new_n2522__ = ~new_new_n1151__ & new_new_n2521__;
  assign new_new_n2523__ = new_new_n1158__ & new_new_n2520__;
  assign new_new_n2524__ = new_new_n2522__ & new_new_n2523__;
  assign new_new_n2525__ = ~new_new_n106__ & ~new_new_n637__;
  assign new_new_n2526__ = ~new_new_n778__ & ~new_new_n942__;
  assign new_new_n2527__ = new_new_n2525__ & new_new_n2526__;
  assign new_new_n2528__ = ~new_new_n202__ & ~new_new_n226__;
  assign new_new_n2529__ = ~new_new_n317__ & ~new_new_n816__;
  assign new_new_n2530__ = new_new_n1424__ & new_new_n2333__;
  assign new_new_n2531__ = new_new_n2529__ & new_new_n2530__;
  assign new_new_n2532__ = new_new_n2527__ & new_new_n2528__;
  assign new_new_n2533__ = new_new_n301__ & new_new_n2532__;
  assign new_new_n2534__ = new_new_n709__ & new_new_n2531__;
  assign new_new_n2535__ = new_new_n2518__ & new_new_n2534__;
  assign new_new_n2536__ = new_new_n2524__ & new_new_n2533__;
  assign new_new_n2537__ = new_new_n2535__ & new_new_n2536__;
  assign new_new_n2538__ = new_new_n2514__ & new_new_n2537__;
  assign new_new_n2539__ = ~new_new_n495__ & ~new_new_n673__;
  assign new_new_n2540__ = ~new_new_n896__ & ~new_new_n959__;
  assign new_new_n2541__ = ~new_new_n247__ & ~new_new_n947__;
  assign new_new_n2542__ = ~new_new_n952__ & new_new_n2541__;
  assign new_new_n2543__ = ~new_new_n124__ & new_new_n2542__;
  assign new_new_n2544__ = ~new_new_n586__ & ~new_new_n675__;
  assign new_new_n2545__ = ~new_new_n373__ & new_new_n2544__;
  assign new_new_n2546__ = new_new_n2543__ & new_new_n2545__;
  assign new_new_n2547__ = ~new_new_n168__ & ~new_new_n676__;
  assign new_new_n2548__ = ~new_new_n1064__ & ~new_new_n1081__;
  assign new_new_n2549__ = ~new_new_n96__ & ~new_new_n155__;
  assign new_new_n2550__ = ~new_new_n511__ & ~new_new_n732__;
  assign new_new_n2551__ = ~new_new_n1033__ & new_new_n2548__;
  assign new_new_n2552__ = new_new_n2549__ & new_new_n2550__;
  assign new_new_n2553__ = new_new_n2551__ & new_new_n2552__;
  assign new_new_n2554__ = new_new_n2547__ & new_new_n2553__;
  assign new_new_n2555__ = ~new_new_n192__ & ~new_new_n352__;
  assign new_new_n2556__ = ~new_new_n322__ & ~new_new_n874__;
  assign new_new_n2557__ = new_new_n2500__ & ~new_new_n2504__;
  assign new_new_n2558__ = new_new_n2556__ & new_new_n2557__;
  assign new_new_n2559__ = ~new_new_n218__ & new_new_n2555__;
  assign new_new_n2560__ = ~new_new_n837__ & new_new_n1875__;
  assign new_new_n2561__ = new_new_n2076__ & new_new_n2499__;
  assign new_new_n2562__ = new_new_n2501__ & new_new_n2539__;
  assign new_new_n2563__ = new_new_n2540__ & new_new_n2562__;
  assign new_new_n2564__ = new_new_n2560__ & new_new_n2561__;
  assign new_new_n2565__ = new_new_n2558__ & new_new_n2559__;
  assign new_new_n2566__ = new_new_n2564__ & new_new_n2565__;
  assign new_new_n2567__ = new_new_n1802__ & new_new_n2563__;
  assign new_new_n2568__ = new_new_n2546__ & new_new_n2567__;
  assign new_new_n2569__ = new_new_n2554__ & new_new_n2566__;
  assign new_new_n2570__ = new_new_n2568__ & new_new_n2569__;
  assign new_new_n2571__ = new_new_n1626__ & new_new_n2570__;
  assign new_new_n2572__ = new_new_n2538__ & new_new_n2571__;
  assign new_new_n2573__ = ~new_new_n2498__ & new_new_n2572__;
  assign new_new_n2574__ = ~new_new_n853__ & ~new_new_n1167__;
  assign new_new_n2575__ = ~new_new_n251__ & ~new_new_n717__;
  assign new_new_n2576__ = ~new_new_n235__ & ~new_new_n1094__;
  assign new_new_n2577__ = new_new_n163__ & ~new_new_n1408__;
  assign new_new_n2578__ = ~new_new_n298__ & ~new_new_n1343__;
  assign new_new_n2579__ = ~new_new_n921__ & new_new_n2578__;
  assign new_new_n2580__ = ~new_new_n2577__ & new_new_n2579__;
  assign new_new_n2581__ = ~new_new_n732__ & ~new_new_n996__;
  assign new_new_n2582__ = ~new_new_n566__ & ~new_new_n602__;
  assign new_new_n2583__ = ~new_new_n809__ & new_new_n2582__;
  assign new_new_n2584__ = new_new_n2581__ & new_new_n2583__;
  assign new_new_n2585__ = ~new_new_n82__ & ~new_new_n130__;
  assign new_new_n2586__ = ~new_new_n890__ & ~new_new_n1073__;
  assign new_new_n2587__ = ~new_new_n317__ & ~new_new_n724__;
  assign new_new_n2588__ = new_new_n1251__ & new_new_n2587__;
  assign new_new_n2589__ = ~new_new_n200__ & ~new_new_n253__;
  assign new_new_n2590__ = ~new_new_n208__ & ~new_new_n692__;
  assign new_new_n2591__ = ~new_new_n138__ & ~new_new_n207__;
  assign new_new_n2592__ = new_new_n107__ & new_new_n2591__;
  assign new_new_n2593__ = ~new_new_n595__ & ~new_new_n945__;
  assign new_new_n2594__ = new_new_n1342__ & new_new_n2585__;
  assign new_new_n2595__ = new_new_n2589__ & new_new_n2590__;
  assign new_new_n2596__ = new_new_n2594__ & new_new_n2595__;
  assign new_new_n2597__ = new_new_n2592__ & new_new_n2593__;
  assign new_new_n2598__ = new_new_n1612__ & new_new_n2586__;
  assign new_new_n2599__ = new_new_n2597__ & new_new_n2598__;
  assign new_new_n2600__ = new_new_n709__ & new_new_n2596__;
  assign new_new_n2601__ = new_new_n2588__ & new_new_n2600__;
  assign new_new_n2602__ = new_new_n2339__ & new_new_n2599__;
  assign new_new_n2603__ = new_new_n2343__ & new_new_n2602__;
  assign new_new_n2604__ = new_new_n2601__ & new_new_n2603__;
  assign new_new_n2605__ = ~new_new_n218__ & ~new_new_n630__;
  assign new_new_n2606__ = ~new_new_n209__ & ~new_new_n723__;
  assign new_new_n2607__ = ~new_new_n383__ & ~new_new_n1291__;
  assign new_new_n2608__ = ~new_new_n495__ & ~new_new_n604__;
  assign new_new_n2609__ = ~new_new_n637__ & ~new_new_n749__;
  assign new_new_n2610__ = ~new_new_n896__ & new_new_n2609__;
  assign new_new_n2611__ = ~new_new_n348__ & new_new_n2608__;
  assign new_new_n2612__ = new_new_n1904__ & new_new_n2606__;
  assign new_new_n2613__ = new_new_n2607__ & new_new_n2612__;
  assign new_new_n2614__ = new_new_n2610__ & new_new_n2611__;
  assign new_new_n2615__ = new_new_n852__ & new_new_n2614__;
  assign new_new_n2616__ = new_new_n1254__ & new_new_n2613__;
  assign new_new_n2617__ = new_new_n2605__ & new_new_n2616__;
  assign new_new_n2618__ = new_new_n2615__ & new_new_n2617__;
  assign new_new_n2619__ = ~new_new_n869__ & ~new_new_n919__;
  assign new_new_n2620__ = new_new_n256__ & ~new_new_n631__;
  assign new_new_n2621__ = ~new_new_n694__ & ~new_new_n990__;
  assign new_new_n2622__ = new_new_n847__ & new_new_n2621__;
  assign new_new_n2623__ = ~new_new_n993__ & new_new_n2575__;
  assign new_new_n2624__ = new_new_n2576__ & new_new_n2623__;
  assign new_new_n2625__ = new_new_n1111__ & new_new_n2622__;
  assign new_new_n2626__ = new_new_n1975__ & new_new_n2574__;
  assign new_new_n2627__ = new_new_n2619__ & new_new_n2626__;
  assign new_new_n2628__ = new_new_n2624__ & new_new_n2625__;
  assign new_new_n2629__ = new_new_n771__ & new_new_n2580__;
  assign new_new_n2630__ = new_new_n2628__ & new_new_n2629__;
  assign new_new_n2631__ = new_new_n2584__ & new_new_n2627__;
  assign new_new_n2632__ = new_new_n2620__ & new_new_n2631__;
  assign new_new_n2633__ = new_new_n2630__ & new_new_n2632__;
  assign new_new_n2634__ = new_new_n2618__ & new_new_n2633__;
  assign new_new_n2635__ = new_new_n2157__ & new_new_n2604__;
  assign new_new_n2636__ = new_new_n2634__ & new_new_n2635__;
  assign new_new_n2637__ = new_new_n2572__ & new_new_n2636__;
  assign new_new_n2638__ = new_new_n2313__ & new_new_n2497__;
  assign new_new_n2639__ = ~new_new_n284__ & ~new_new_n477__;
  assign new_new_n2640__ = ~new_new_n76__ & ~new_new_n749__;
  assign new_new_n2641__ = ~new_new_n280__ & ~new_new_n316__;
  assign new_new_n2642__ = ~new_new_n208__ & ~new_new_n845__;
  assign new_new_n2643__ = ~new_new_n597__ & ~new_new_n719__;
  assign new_new_n2644__ = ~new_new_n952__ & ~new_new_n1515__;
  assign new_new_n2645__ = new_new_n100__ & ~new_new_n2328__;
  assign new_new_n2646__ = ~new_new_n192__ & ~new_new_n385__;
  assign new_new_n2647__ = ~new_new_n747__ & new_new_n1062__;
  assign new_new_n2648__ = ~new_new_n2645__ & new_new_n2647__;
  assign new_new_n2649__ = new_new_n1142__ & new_new_n2646__;
  assign new_new_n2650__ = new_new_n2643__ & new_new_n2644__;
  assign new_new_n2651__ = new_new_n2649__ & new_new_n2650__;
  assign new_new_n2652__ = new_new_n2648__ & new_new_n2651__;
  assign new_new_n2653__ = ~new_new_n229__ & ~new_new_n631__;
  assign new_new_n2654__ = ~new_new_n990__ & ~new_new_n1033__;
  assign new_new_n2655__ = ~new_new_n961__ & new_new_n2654__;
  assign new_new_n2656__ = new_new_n852__ & new_new_n2655__;
  assign new_new_n2657__ = new_new_n2653__ & new_new_n2656__;
  assign new_new_n2658__ = ~new_new_n313__ & ~new_new_n1080__;
  assign new_new_n2659__ = ~new_new_n276__ & new_new_n2658__;
  assign new_new_n2660__ = ~new_new_n311__ & ~new_new_n1008__;
  assign new_new_n2661__ = new_new_n2640__ & new_new_n2642__;
  assign new_new_n2662__ = new_new_n2660__ & new_new_n2661__;
  assign new_new_n2663__ = new_new_n1664__ & new_new_n2659__;
  assign new_new_n2664__ = new_new_n1748__ & new_new_n1847__;
  assign new_new_n2665__ = new_new_n2639__ & new_new_n2664__;
  assign new_new_n2666__ = new_new_n2662__ & new_new_n2663__;
  assign new_new_n2667__ = new_new_n228__ & new_new_n2641__;
  assign new_new_n2668__ = new_new_n2666__ & new_new_n2667__;
  assign new_new_n2669__ = new_new_n2657__ & new_new_n2665__;
  assign new_new_n2670__ = new_new_n2668__ & new_new_n2669__;
  assign new_new_n2671__ = new_new_n2652__ & new_new_n2670__;
  assign new_new_n2672__ = ~pi29 & new_new_n219__;
  assign new_new_n2673__ = new_new_n81__ & new_new_n2672__;
  assign new_new_n2674__ = ~new_new_n120__ & ~new_new_n783__;
  assign new_new_n2675__ = ~new_new_n2673__ & new_new_n2674__;
  assign new_new_n2676__ = ~new_new_n317__ & new_new_n1083__;
  assign new_new_n2677__ = new_new_n2675__ & new_new_n2676__;
  assign new_new_n2678__ = ~new_new_n1539__ & new_new_n2677__;
  assign new_new_n2679__ = ~new_new_n940__ & ~new_new_n1212__;
  assign new_new_n2680__ = ~new_new_n717__ & ~new_new_n785__;
  assign new_new_n2681__ = ~new_new_n853__ & ~new_new_n937__;
  assign new_new_n2682__ = new_new_n2680__ & new_new_n2681__;
  assign new_new_n2683__ = ~new_new_n270__ & ~new_new_n919__;
  assign new_new_n2684__ = ~new_new_n945__ & ~new_new_n1009__;
  assign new_new_n2685__ = new_new_n1742__ & new_new_n2679__;
  assign new_new_n2686__ = new_new_n2684__ & new_new_n2685__;
  assign new_new_n2687__ = new_new_n2682__ & new_new_n2683__;
  assign new_new_n2688__ = ~new_new_n676__ & new_new_n733__;
  assign new_new_n2689__ = new_new_n994__ & new_new_n1599__;
  assign new_new_n2690__ = new_new_n1840__ & new_new_n2689__;
  assign new_new_n2691__ = new_new_n2687__ & new_new_n2688__;
  assign new_new_n2692__ = new_new_n2204__ & new_new_n2686__;
  assign new_new_n2693__ = new_new_n2691__ & new_new_n2692__;
  assign new_new_n2694__ = new_new_n2678__ & new_new_n2690__;
  assign new_new_n2695__ = new_new_n2693__ & new_new_n2694__;
  assign new_new_n2696__ = ~new_new_n112__ & ~new_new_n152__;
  assign new_new_n2697__ = new_new_n780__ & ~new_new_n2696__;
  assign new_new_n2698__ = ~new_new_n438__ & ~new_new_n724__;
  assign new_new_n2699__ = ~new_new_n255__ & new_new_n699__;
  assign new_new_n2700__ = new_new_n2698__ & new_new_n2699__;
  assign new_new_n2701__ = ~new_new_n124__ & ~new_new_n335__;
  assign new_new_n2702__ = ~new_new_n382__ & ~new_new_n1291__;
  assign new_new_n2703__ = new_new_n1397__ & new_new_n2702__;
  assign new_new_n2704__ = new_new_n2701__ & new_new_n2703__;
  assign new_new_n2705__ = ~new_new_n809__ & ~new_new_n874__;
  assign new_new_n2706__ = ~new_new_n671__ & new_new_n1449__;
  assign new_new_n2707__ = ~new_new_n701__ & ~new_new_n1081__;
  assign new_new_n2708__ = ~new_new_n101__ & ~new_new_n302__;
  assign new_new_n2709__ = new_new_n1168__ & new_new_n1741__;
  assign new_new_n2710__ = ~new_new_n247__ & ~new_new_n1506__;
  assign new_new_n2711__ = ~new_new_n260__ & ~new_new_n336__;
  assign new_new_n2712__ = ~new_new_n119__ & ~new_new_n829__;
  assign new_new_n2713__ = ~new_new_n168__ & ~new_new_n242__;
  assign new_new_n2714__ = ~new_new_n692__ & new_new_n2713__;
  assign new_new_n2715__ = ~new_new_n921__ & new_new_n2708__;
  assign new_new_n2716__ = new_new_n2711__ & new_new_n2712__;
  assign new_new_n2717__ = new_new_n2715__ & new_new_n2716__;
  assign new_new_n2718__ = ~new_new_n115__ & new_new_n2714__;
  assign new_new_n2719__ = ~new_new_n254__ & new_new_n2710__;
  assign new_new_n2720__ = new_new_n2718__ & new_new_n2719__;
  assign new_new_n2721__ = new_new_n2709__ & new_new_n2717__;
  assign new_new_n2722__ = new_new_n2720__ & new_new_n2721__;
  assign new_new_n2723__ = ~new_new_n372__ & ~new_new_n602__;
  assign new_new_n2724__ = new_new_n1510__ & ~new_new_n2697__;
  assign new_new_n2725__ = new_new_n2707__ & new_new_n2724__;
  assign new_new_n2726__ = new_new_n475__ & new_new_n2723__;
  assign new_new_n2727__ = ~new_new_n935__ & new_new_n1215__;
  assign new_new_n2728__ = new_new_n1777__ & new_new_n2706__;
  assign new_new_n2729__ = new_new_n2727__ & new_new_n2728__;
  assign new_new_n2730__ = new_new_n2725__ & new_new_n2726__;
  assign new_new_n2731__ = new_new_n2700__ & new_new_n2705__;
  assign new_new_n2732__ = new_new_n2730__ & new_new_n2731__;
  assign new_new_n2733__ = new_new_n2729__ & new_new_n2732__;
  assign new_new_n2734__ = new_new_n2704__ & new_new_n2722__;
  assign new_new_n2735__ = new_new_n2733__ & new_new_n2734__;
  assign new_new_n2736__ = new_new_n2695__ & new_new_n2735__;
  assign new_new_n2737__ = new_new_n2671__ & new_new_n2736__;
  assign new_new_n2738__ = new_new_n2638__ & new_new_n2737__;
  assign new_new_n2739__ = ~new_new_n2637__ & ~new_new_n2738__;
  assign new_new_n2740__ = ~new_new_n126__ & ~new_new_n594__;
  assign new_new_n2741__ = pi24 & ~new_new_n2740__;
  assign new_new_n2742__ = ~new_new_n201__ & ~new_new_n587__;
  assign new_new_n2743__ = ~new_new_n112__ & ~new_new_n2742__;
  assign new_new_n2744__ = ~new_new_n2741__ & ~new_new_n2743__;
  assign new_new_n2745__ = pi26 & ~new_new_n2744__;
  assign new_new_n2746__ = new_new_n112__ & new_new_n126__;
  assign new_new_n2747__ = ~new_new_n188__ & ~new_new_n211__;
  assign new_new_n2748__ = ~pi24 & ~new_new_n2747__;
  assign new_new_n2749__ = new_new_n211__ & ~new_new_n2696__;
  assign new_new_n2750__ = ~new_new_n2746__ & ~new_new_n2749__;
  assign new_new_n2751__ = ~new_new_n2748__ & new_new_n2750__;
  assign new_new_n2752__ = ~pi26 & ~new_new_n2751__;
  assign new_new_n2753__ = ~new_new_n2745__ & ~new_new_n2752__;
  assign new_new_n2754__ = ~new_new_n108__ & ~new_new_n351__;
  assign new_new_n2755__ = ~new_new_n479__ & ~new_new_n768__;
  assign new_new_n2756__ = ~new_new_n877__ & new_new_n2754__;
  assign new_new_n2757__ = new_new_n2755__ & new_new_n2756__;
  assign new_new_n2758__ = ~new_new_n719__ & ~new_new_n846__;
  assign new_new_n2759__ = pi23 & ~new_new_n194__;
  assign new_new_n2760__ = ~new_new_n303__ & ~new_new_n2759__;
  assign new_new_n2761__ = ~new_new_n134__ & new_new_n137__;
  assign new_new_n2762__ = ~new_new_n2760__ & new_new_n2761__;
  assign new_new_n2763__ = ~new_new_n286__ & ~new_new_n701__;
  assign new_new_n2764__ = ~new_new_n373__ & ~new_new_n894__;
  assign new_new_n2765__ = ~new_new_n300__ & ~new_new_n519__;
  assign new_new_n2766__ = new_new_n2763__ & new_new_n2765__;
  assign new_new_n2767__ = new_new_n2764__ & new_new_n2766__;
  assign new_new_n2768__ = ~new_new_n495__ & ~new_new_n692__;
  assign new_new_n2769__ = ~new_new_n350__ & ~new_new_n942__;
  assign new_new_n2770__ = ~new_new_n696__ & ~new_new_n724__;
  assign new_new_n2771__ = ~new_new_n274__ & ~new_new_n1176__;
  assign new_new_n2772__ = ~new_new_n196__ & ~new_new_n271__;
  assign new_new_n2773__ = ~new_new_n1008__ & new_new_n2772__;
  assign new_new_n2774__ = new_new_n1110__ & new_new_n2773__;
  assign new_new_n2775__ = new_new_n2769__ & new_new_n2770__;
  assign new_new_n2776__ = new_new_n2771__ & new_new_n2775__;
  assign new_new_n2777__ = new_new_n2774__ & new_new_n2776__;
  assign new_new_n2778__ = ~new_new_n270__ & ~new_new_n884__;
  assign new_new_n2779__ = ~new_new_n441__ & ~new_new_n749__;
  assign new_new_n2780__ = ~new_new_n1212__ & new_new_n2779__;
  assign new_new_n2781__ = ~new_new_n258__ & ~new_new_n781__;
  assign new_new_n2782__ = ~new_new_n1108__ & new_new_n2781__;
  assign new_new_n2783__ = ~new_new_n124__ & new_new_n2780__;
  assign new_new_n2784__ = new_new_n1848__ & new_new_n2196__;
  assign new_new_n2785__ = new_new_n2778__ & new_new_n2784__;
  assign new_new_n2786__ = new_new_n2782__ & new_new_n2783__;
  assign new_new_n2787__ = new_new_n2785__ & new_new_n2786__;
  assign new_new_n2788__ = new_new_n1845__ & new_new_n2787__;
  assign new_new_n2789__ = ~new_new_n835__ & ~new_new_n993__;
  assign new_new_n2790__ = new_new_n2788__ & new_new_n2789__;
  assign new_new_n2791__ = ~new_new_n439__ & ~new_new_n785__;
  assign new_new_n2792__ = ~pi25 & ~new_new_n95__;
  assign new_new_n2793__ = pi25 & ~new_new_n237__;
  assign new_new_n2794__ = new_new_n99__ & ~new_new_n2792__;
  assign new_new_n2795__ = ~new_new_n2793__ & new_new_n2794__;
  assign new_new_n2796__ = ~new_new_n566__ & ~new_new_n837__;
  assign new_new_n2797__ = ~new_new_n284__ & ~new_new_n315__;
  assign new_new_n2798__ = ~new_new_n427__ & new_new_n2797__;
  assign new_new_n2799__ = new_new_n1909__ & new_new_n2288__;
  assign new_new_n2800__ = new_new_n2798__ & new_new_n2799__;
  assign new_new_n2801__ = new_new_n2439__ & new_new_n2800__;
  assign new_new_n2802__ = new_new_n2796__ & new_new_n2801__;
  assign new_new_n2803__ = ~new_new_n82__ & ~new_new_n238__;
  assign new_new_n2804__ = ~new_new_n240__ & ~new_new_n845__;
  assign new_new_n2805__ = ~new_new_n937__ & new_new_n2804__;
  assign new_new_n2806__ = ~new_new_n317__ & new_new_n2803__;
  assign new_new_n2807__ = ~new_new_n321__ & new_new_n2067__;
  assign new_new_n2808__ = new_new_n2806__ & new_new_n2807__;
  assign new_new_n2809__ = ~new_new_n218__ & new_new_n2805__;
  assign new_new_n2810__ = new_new_n1329__ & new_new_n1482__;
  assign new_new_n2811__ = ~new_new_n2795__ & new_new_n2810__;
  assign new_new_n2812__ = new_new_n2808__ & new_new_n2809__;
  assign new_new_n2813__ = new_new_n936__ & new_new_n1001__;
  assign new_new_n2814__ = new_new_n1772__ & new_new_n2323__;
  assign new_new_n2815__ = new_new_n2791__ & new_new_n2814__;
  assign new_new_n2816__ = new_new_n2812__ & new_new_n2813__;
  assign new_new_n2817__ = new_new_n2811__ & new_new_n2816__;
  assign new_new_n2818__ = new_new_n2802__ & new_new_n2815__;
  assign new_new_n2819__ = new_new_n2817__ & new_new_n2818__;
  assign new_new_n2820__ = ~new_new_n332__ & ~new_new_n1009__;
  assign new_new_n2821__ = ~new_new_n155__ & ~new_new_n851__;
  assign new_new_n2822__ = ~new_new_n250__ & ~new_new_n496__;
  assign new_new_n2823__ = ~new_new_n92__ & ~new_new_n746__;
  assign new_new_n2824__ = ~new_new_n1167__ & new_new_n2823__;
  assign new_new_n2825__ = new_new_n2822__ & new_new_n2824__;
  assign new_new_n2826__ = new_new_n381__ & new_new_n949__;
  assign new_new_n2827__ = new_new_n2820__ & new_new_n2821__;
  assign new_new_n2828__ = new_new_n2826__ & new_new_n2827__;
  assign new_new_n2829__ = new_new_n2641__ & new_new_n2825__;
  assign new_new_n2830__ = new_new_n2828__ & new_new_n2829__;
  assign new_new_n2831__ = ~new_new_n106__ & ~new_new_n282__;
  assign new_new_n2832__ = ~new_new_n302__ & ~new_new_n893__;
  assign new_new_n2833__ = ~new_new_n933__ & ~new_new_n1343__;
  assign new_new_n2834__ = new_new_n2832__ & new_new_n2833__;
  assign new_new_n2835__ = ~new_new_n952__ & new_new_n2831__;
  assign new_new_n2836__ = ~new_new_n961__ & new_new_n2116__;
  assign new_new_n2837__ = new_new_n2768__ & new_new_n2836__;
  assign new_new_n2838__ = new_new_n2834__ & new_new_n2835__;
  assign new_new_n2839__ = new_new_n2758__ & ~new_new_n2762__;
  assign new_new_n2840__ = new_new_n2838__ & new_new_n2839__;
  assign new_new_n2841__ = new_new_n2837__ & new_new_n2840__;
  assign new_new_n2842__ = new_new_n2757__ & new_new_n2841__;
  assign new_new_n2843__ = new_new_n2753__ & new_new_n2767__;
  assign new_new_n2844__ = new_new_n2777__ & new_new_n2830__;
  assign new_new_n2845__ = new_new_n2843__ & new_new_n2844__;
  assign new_new_n2846__ = new_new_n2842__ & new_new_n2845__;
  assign new_new_n2847__ = new_new_n2790__ & new_new_n2819__;
  assign new_new_n2848__ = new_new_n2846__ & new_new_n2847__;
  assign new_new_n2849__ = ~new_new_n2737__ & ~new_new_n2848__;
  assign new_new_n2850__ = ~new_new_n602__ & ~new_new_n1507__;
  assign new_new_n2851__ = ~new_new_n143__ & ~new_new_n379__;
  assign new_new_n2852__ = ~new_new_n488__ & ~new_new_n2170__;
  assign new_new_n2853__ = ~new_new_n101__ & ~new_new_n235__;
  assign new_new_n2854__ = ~new_new_n258__ & new_new_n2853__;
  assign new_new_n2855__ = ~new_new_n828__ & ~new_new_n1009__;
  assign new_new_n2856__ = new_new_n1367__ & new_new_n1742__;
  assign new_new_n2857__ = new_new_n2855__ & new_new_n2856__;
  assign new_new_n2858__ = new_new_n2850__ & new_new_n2854__;
  assign new_new_n2859__ = new_new_n2851__ & new_new_n2852__;
  assign new_new_n2860__ = new_new_n2858__ & new_new_n2859__;
  assign new_new_n2861__ = new_new_n2518__ & new_new_n2857__;
  assign new_new_n2862__ = new_new_n2641__ & new_new_n2861__;
  assign new_new_n2863__ = new_new_n2546__ & new_new_n2860__;
  assign new_new_n2864__ = new_new_n2862__ & new_new_n2863__;
  assign new_new_n2865__ = new_new_n116__ & new_new_n2549__;
  assign new_new_n2866__ = ~new_new_n208__ & new_new_n1366__;
  assign new_new_n2867__ = ~new_new_n209__ & new_new_n2866__;
  assign new_new_n2868__ = ~new_new_n658__ & ~new_new_n785__;
  assign new_new_n2869__ = new_new_n193__ & ~new_new_n729__;
  assign new_new_n2870__ = new_new_n744__ & new_new_n2334__;
  assign new_new_n2871__ = new_new_n2869__ & new_new_n2870__;
  assign new_new_n2872__ = ~new_new_n767__ & ~new_new_n853__;
  assign new_new_n2873__ = ~new_new_n878__ & new_new_n1213__;
  assign new_new_n2874__ = ~new_new_n2697__ & new_new_n2868__;
  assign new_new_n2875__ = new_new_n2873__ & new_new_n2874__;
  assign new_new_n2876__ = new_new_n984__ & new_new_n2872__;
  assign new_new_n2877__ = new_new_n2875__ & new_new_n2876__;
  assign new_new_n2878__ = new_new_n347__ & new_new_n1434__;
  assign new_new_n2879__ = new_new_n2867__ & new_new_n2878__;
  assign new_new_n2880__ = new_new_n1526__ & new_new_n2877__;
  assign new_new_n2881__ = new_new_n2343__ & new_new_n2865__;
  assign new_new_n2882__ = new_new_n2871__ & new_new_n2881__;
  assign new_new_n2883__ = new_new_n2879__ & new_new_n2880__;
  assign new_new_n2884__ = new_new_n2882__ & new_new_n2883__;
  assign new_new_n2885__ = new_new_n2864__ & new_new_n2884__;
  assign new_new_n2886__ = new_new_n2063__ & new_new_n2885__;
  assign new_new_n2887__ = ~new_new_n2849__ & new_new_n2886__;
  assign new_new_n2888__ = ~new_new_n676__ & ~new_new_n694__;
  assign new_new_n2889__ = ~new_new_n781__ & ~new_new_n846__;
  assign new_new_n2890__ = ~new_new_n603__ & ~new_new_n933__;
  assign new_new_n2891__ = ~new_new_n990__ & ~new_new_n1070__;
  assign new_new_n2892__ = new_new_n2890__ & new_new_n2891__;
  assign new_new_n2893__ = new_new_n2889__ & new_new_n2892__;
  assign new_new_n2894__ = ~new_new_n284__ & ~new_new_n732__;
  assign new_new_n2895__ = ~new_new_n308__ & ~new_new_n379__;
  assign new_new_n2896__ = ~new_new_n92__ & ~new_new_n607__;
  assign new_new_n2897__ = ~new_new_n604__ & ~new_new_n768__;
  assign new_new_n2898__ = ~new_new_n483__ & new_new_n2897__;
  assign new_new_n2899__ = new_new_n2895__ & new_new_n2898__;
  assign new_new_n2900__ = ~new_new_n373__ & new_new_n1825__;
  assign new_new_n2901__ = new_new_n1905__ & new_new_n2316__;
  assign new_new_n2902__ = new_new_n2322__ & new_new_n2894__;
  assign new_new_n2903__ = new_new_n2901__ & new_new_n2902__;
  assign new_new_n2904__ = new_new_n2899__ & new_new_n2900__;
  assign new_new_n2905__ = new_new_n2888__ & new_new_n2893__;
  assign new_new_n2906__ = new_new_n2896__ & new_new_n2905__;
  assign new_new_n2907__ = new_new_n2903__ & new_new_n2904__;
  assign new_new_n2908__ = new_new_n2906__ & new_new_n2907__;
  assign new_new_n2909__ = ~new_new_n168__ & ~new_new_n1217__;
  assign new_new_n2910__ = ~new_new_n656__ & ~new_new_n698__;
  assign new_new_n2911__ = ~new_new_n1064__ & new_new_n2910__;
  assign new_new_n2912__ = new_new_n2909__ & new_new_n2911__;
  assign new_new_n2913__ = ~new_new_n148__ & ~new_new_n772__;
  assign new_new_n2914__ = ~new_new_n127__ & ~new_new_n482__;
  assign new_new_n2915__ = ~new_new_n749__ & new_new_n2914__;
  assign new_new_n2916__ = ~new_new_n280__ & ~new_new_n959__;
  assign new_new_n2917__ = new_new_n2915__ & new_new_n2916__;
  assign new_new_n2918__ = ~new_new_n218__ & new_new_n2917__;
  assign new_new_n2919__ = ~new_new_n427__ & ~new_new_n480__;
  assign new_new_n2920__ = ~new_new_n160__ & ~new_new_n246__;
  assign new_new_n2921__ = ~new_new_n671__ & ~new_new_n826__;
  assign new_new_n2922__ = new_new_n2920__ & new_new_n2921__;
  assign new_new_n2923__ = ~new_new_n263__ & ~new_new_n921__;
  assign new_new_n2924__ = new_new_n1944__ & new_new_n2923__;
  assign new_new_n2925__ = new_new_n716__ & new_new_n2922__;
  assign new_new_n2926__ = new_new_n2924__ & new_new_n2925__;
  assign new_new_n2927__ = new_new_n102__ & ~new_new_n1094__;
  assign new_new_n2928__ = ~new_new_n155__ & ~new_new_n183__;
  assign new_new_n2929__ = ~new_new_n276__ & ~new_new_n874__;
  assign new_new_n2930__ = new_new_n1082__ & new_new_n1469__;
  assign new_new_n2931__ = new_new_n2929__ & new_new_n2930__;
  assign new_new_n2932__ = new_new_n2927__ & new_new_n2928__;
  assign new_new_n2933__ = new_new_n744__ & new_new_n1747__;
  assign new_new_n2934__ = new_new_n2919__ & new_new_n2933__;
  assign new_new_n2935__ = new_new_n2931__ & new_new_n2932__;
  assign new_new_n2936__ = new_new_n1774__ & new_new_n2935__;
  assign new_new_n2937__ = new_new_n2918__ & new_new_n2934__;
  assign new_new_n2938__ = new_new_n2926__ & new_new_n2937__;
  assign new_new_n2939__ = new_new_n2936__ & new_new_n2938__;
  assign new_new_n2940__ = ~new_new_n286__ & new_new_n941__;
  assign new_new_n2941__ = new_new_n2939__ & new_new_n2940__;
  assign new_new_n2942__ = ~new_new_n320__ & ~new_new_n634__;
  assign new_new_n2943__ = ~new_new_n425__ & ~new_new_n785__;
  assign new_new_n2944__ = ~new_new_n335__ & ~new_new_n701__;
  assign new_new_n2945__ = ~new_new_n179__ & ~new_new_n309__;
  assign new_new_n2946__ = new_new_n474__ & new_new_n2945__;
  assign new_new_n2947__ = new_new_n2942__ & new_new_n2943__;
  assign new_new_n2948__ = new_new_n2944__ & new_new_n2947__;
  assign new_new_n2949__ = ~new_new_n344__ & new_new_n2946__;
  assign new_new_n2950__ = new_new_n916__ & ~new_new_n935__;
  assign new_new_n2951__ = new_new_n2515__ & new_new_n2913__;
  assign new_new_n2952__ = new_new_n2950__ & new_new_n2951__;
  assign new_new_n2953__ = new_new_n2948__ & new_new_n2949__;
  assign new_new_n2954__ = new_new_n1293__ & new_new_n2912__;
  assign new_new_n2955__ = new_new_n2953__ & new_new_n2954__;
  assign new_new_n2956__ = new_new_n2952__ & new_new_n2955__;
  assign new_new_n2957__ = new_new_n2652__ & new_new_n2956__;
  assign new_new_n2958__ = new_new_n2908__ & new_new_n2957__;
  assign new_new_n2959__ = new_new_n2604__ & new_new_n2958__;
  assign new_new_n2960__ = new_new_n2941__ & new_new_n2959__;
  assign new_new_n2961__ = new_new_n2737__ & new_new_n2848__;
  assign new_new_n2962__ = ~new_new_n488__ & ~new_new_n1073__;
  assign new_new_n2963__ = ~new_new_n238__ & ~new_new_n724__;
  assign new_new_n2964__ = ~new_new_n1210__ & new_new_n2963__;
  assign new_new_n2965__ = ~new_new_n380__ & ~new_new_n673__;
  assign new_new_n2966__ = ~new_new_n781__ & new_new_n2965__;
  assign new_new_n2967__ = ~new_new_n254__ & new_new_n2964__;
  assign new_new_n2968__ = new_new_n323__ & new_new_n2967__;
  assign new_new_n2969__ = new_new_n2966__ & new_new_n2968__;
  assign new_new_n2970__ = ~new_new_n624__ & ~new_new_n845__;
  assign new_new_n2971__ = ~new_new_n300__ & ~new_new_n473__;
  assign new_new_n2972__ = new_new_n2068__ & new_new_n2971__;
  assign new_new_n2973__ = new_new_n1679__ & new_new_n2972__;
  assign new_new_n2974__ = ~new_new_n138__ & ~new_new_n482__;
  assign new_new_n2975__ = ~new_new_n940__ & new_new_n2974__;
  assign new_new_n2976__ = ~new_new_n477__ & ~new_new_n1568__;
  assign new_new_n2977__ = ~new_new_n2329__ & new_new_n2707__;
  assign new_new_n2978__ = new_new_n2970__ & new_new_n2977__;
  assign new_new_n2979__ = new_new_n2975__ & new_new_n2976__;
  assign new_new_n2980__ = new_new_n2962__ & new_new_n2979__;
  assign new_new_n2981__ = new_new_n318__ & new_new_n2978__;
  assign new_new_n2982__ = new_new_n2896__ & new_new_n2981__;
  assign new_new_n2983__ = new_new_n669__ & new_new_n2980__;
  assign new_new_n2984__ = new_new_n2097__ & new_new_n2973__;
  assign new_new_n2985__ = new_new_n2983__ & new_new_n2984__;
  assign new_new_n2986__ = new_new_n2969__ & new_new_n2982__;
  assign new_new_n2987__ = new_new_n2985__ & new_new_n2986__;
  assign new_new_n2988__ = ~new_new_n189__ & ~new_new_n353__;
  assign new_new_n2989__ = ~new_new_n1035__ & new_new_n2988__;
  assign new_new_n2990__ = ~new_new_n115__ & ~new_new_n259__;
  assign new_new_n2991__ = ~new_new_n280__ & ~new_new_n919__;
  assign new_new_n2992__ = ~new_new_n119__ & ~new_new_n136__;
  assign new_new_n2993__ = ~new_new_n260__ & ~new_new_n816__;
  assign new_new_n2994__ = ~new_new_n208__ & ~new_new_n878__;
  assign new_new_n2995__ = new_new_n135__ & ~new_new_n1408__;
  assign new_new_n2996__ = ~new_new_n603__ & ~new_new_n778__;
  assign new_new_n2997__ = ~new_new_n1291__ & new_new_n2996__;
  assign new_new_n2998__ = ~new_new_n166__ & ~new_new_n274__;
  assign new_new_n2999__ = ~new_new_n2995__ & new_new_n2998__;
  assign new_new_n3000__ = new_new_n1705__ & new_new_n2997__;
  assign new_new_n3001__ = new_new_n2991__ & new_new_n2992__;
  assign new_new_n3002__ = new_new_n2993__ & new_new_n2994__;
  assign new_new_n3003__ = new_new_n3001__ & new_new_n3002__;
  assign new_new_n3004__ = new_new_n2999__ & new_new_n3000__;
  assign new_new_n3005__ = new_new_n2133__ & new_new_n2989__;
  assign new_new_n3006__ = new_new_n2990__ & new_new_n3005__;
  assign new_new_n3007__ = new_new_n3003__ & new_new_n3004__;
  assign new_new_n3008__ = new_new_n2088__ & new_new_n3007__;
  assign new_new_n3009__ = new_new_n3006__ & new_new_n3008__;
  assign new_new_n3010__ = ~new_new_n229__ & ~new_new_n996__;
  assign new_new_n3011__ = ~new_new_n374__ & ~new_new_n846__;
  assign new_new_n3012__ = new_new_n3010__ & new_new_n3011__;
  assign new_new_n3013__ = new_new_n163__ & new_new_n814__;
  assign new_new_n3014__ = ~pi25 & ~new_new_n304__;
  assign new_new_n3015__ = ~new_new_n79__ & ~new_new_n89__;
  assign new_new_n3016__ = new_new_n3014__ & new_new_n3015__;
  assign new_new_n3017__ = ~new_new_n278__ & ~new_new_n3016__;
  assign new_new_n3018__ = new_new_n169__ & ~new_new_n3017__;
  assign new_new_n3019__ = ~new_new_n1080__ & ~new_new_n3018__;
  assign new_new_n3020__ = ~new_new_n585__ & ~new_new_n838__;
  assign new_new_n3021__ = ~new_new_n106__ & new_new_n3020__;
  assign new_new_n3022__ = new_new_n1747__ & new_new_n3021__;
  assign new_new_n3023__ = ~new_new_n479__ & ~new_new_n961__;
  assign new_new_n3024__ = ~new_new_n198__ & ~new_new_n373__;
  assign new_new_n3025__ = ~new_new_n346__ & ~new_new_n809__;
  assign new_new_n3026__ = ~new_new_n348__ & ~new_new_n379__;
  assign new_new_n3027__ = ~new_new_n729__ & ~new_new_n869__;
  assign new_new_n3028__ = ~new_new_n277__ & ~new_new_n2170__;
  assign new_new_n3029__ = ~new_new_n306__ & ~new_new_n828__;
  assign new_new_n3030__ = new_new_n1631__ & new_new_n3029__;
  assign new_new_n3031__ = new_new_n3026__ & new_new_n3028__;
  assign new_new_n3032__ = new_new_n3027__ & new_new_n3031__;
  assign new_new_n3033__ = new_new_n1805__ & new_new_n3030__;
  assign new_new_n3034__ = new_new_n3024__ & new_new_n3025__;
  assign new_new_n3035__ = new_new_n3033__ & new_new_n3034__;
  assign new_new_n3036__ = new_new_n3032__ & new_new_n3035__;
  assign new_new_n3037__ = ~new_new_n179__ & ~new_new_n200__;
  assign new_new_n3038__ = ~new_new_n212__ & ~new_new_n658__;
  assign new_new_n3039__ = ~new_new_n890__ & ~new_new_n3013__;
  assign new_new_n3040__ = new_new_n3038__ & new_new_n3039__;
  assign new_new_n3041__ = ~new_new_n263__ & new_new_n3037__;
  assign new_new_n3042__ = ~new_new_n566__ & new_new_n1807__;
  assign new_new_n3043__ = new_new_n3041__ & new_new_n3042__;
  assign new_new_n3044__ = ~new_new_n439__ & new_new_n3040__;
  assign new_new_n3045__ = new_new_n2290__ & new_new_n2453__;
  assign new_new_n3046__ = new_new_n3012__ & new_new_n3045__;
  assign new_new_n3047__ = new_new_n3043__ & new_new_n3044__;
  assign new_new_n3048__ = new_new_n1774__ & new_new_n3019__;
  assign new_new_n3049__ = new_new_n3022__ & new_new_n3023__;
  assign new_new_n3050__ = new_new_n3048__ & new_new_n3049__;
  assign new_new_n3051__ = new_new_n3046__ & new_new_n3047__;
  assign new_new_n3052__ = new_new_n3050__ & new_new_n3051__;
  assign new_new_n3053__ = new_new_n3036__ & new_new_n3052__;
  assign new_new_n3054__ = new_new_n2987__ & new_new_n3053__;
  assign new_new_n3055__ = new_new_n3009__ & new_new_n3054__;
  assign new_new_n3056__ = ~new_new_n103__ & ~new_new_n196__;
  assign new_new_n3057__ = ~new_new_n166__ & ~new_new_n198__;
  assign new_new_n3058__ = ~new_new_n130__ & ~new_new_n845__;
  assign new_new_n3059__ = ~new_new_n842__ & ~new_new_n1035__;
  assign new_new_n3060__ = ~new_new_n472__ & ~new_new_n495__;
  assign new_new_n3061__ = ~new_new_n658__ & ~new_new_n843__;
  assign new_new_n3062__ = new_new_n3060__ & new_new_n3061__;
  assign new_new_n3063__ = ~new_new_n675__ & new_new_n725__;
  assign new_new_n3064__ = ~new_new_n781__ & ~new_new_n1217__;
  assign new_new_n3065__ = new_new_n3056__ & new_new_n3058__;
  assign new_new_n3066__ = new_new_n3064__ & new_new_n3065__;
  assign new_new_n3067__ = new_new_n3062__ & new_new_n3063__;
  assign new_new_n3068__ = ~new_new_n115__ & new_new_n743__;
  assign new_new_n3069__ = new_new_n962__ & new_new_n2235__;
  assign new_new_n3070__ = new_new_n3057__ & new_new_n3059__;
  assign new_new_n3071__ = new_new_n3069__ & new_new_n3070__;
  assign new_new_n3072__ = new_new_n3067__ & new_new_n3068__;
  assign new_new_n3073__ = new_new_n3066__ & new_new_n3072__;
  assign new_new_n3074__ = new_new_n1431__ & new_new_n3071__;
  assign new_new_n3075__ = new_new_n3073__ & new_new_n3074__;
  assign new_new_n3076__ = ~new_new_n192__ & ~new_new_n226__;
  assign new_new_n3077__ = ~new_new_n108__ & ~new_new_n212__;
  assign new_new_n3078__ = ~new_new_n473__ & ~new_new_n692__;
  assign new_new_n3079__ = ~new_new_n1398__ & new_new_n3078__;
  assign new_new_n3080__ = new_new_n629__ & ~new_new_n952__;
  assign new_new_n3081__ = new_new_n2268__ & new_new_n3077__;
  assign new_new_n3082__ = new_new_n3080__ & new_new_n3081__;
  assign new_new_n3083__ = ~new_new_n1486__ & new_new_n3079__;
  assign new_new_n3084__ = new_new_n2000__ & new_new_n2820__;
  assign new_new_n3085__ = new_new_n3076__ & new_new_n3084__;
  assign new_new_n3086__ = new_new_n3082__ & new_new_n3083__;
  assign new_new_n3087__ = new_new_n1772__ & new_new_n3086__;
  assign new_new_n3088__ = new_new_n1681__ & new_new_n3085__;
  assign new_new_n3089__ = new_new_n3087__ & new_new_n3088__;
  assign new_new_n3090__ = ~new_new_n630__ & new_new_n3089__;
  assign new_new_n3091__ = ~new_new_n270__ & ~new_new_n489__;
  assign new_new_n3092__ = new_new_n73__ & new_new_n587__;
  assign new_new_n3093__ = ~new_new_n950__ & ~new_new_n3092__;
  assign new_new_n3094__ = new_new_n2994__ & new_new_n3093__;
  assign new_new_n3095__ = new_new_n3091__ & new_new_n3094__;
  assign new_new_n3096__ = ~new_new_n251__ & ~new_new_n300__;
  assign new_new_n3097__ = ~new_new_n267__ & new_new_n967__;
  assign new_new_n3098__ = new_new_n1645__ & new_new_n3097__;
  assign new_new_n3099__ = ~new_new_n315__ & ~new_new_n439__;
  assign new_new_n3100__ = ~new_new_n298__ & ~new_new_n344__;
  assign new_new_n3101__ = ~new_new_n1162__ & ~new_new_n1506__;
  assign new_new_n3102__ = ~new_new_n283__ & ~new_new_n1372__;
  assign new_new_n3103__ = ~new_new_n249__ & ~new_new_n385__;
  assign new_new_n3104__ = ~new_new_n585__ & ~new_new_n783__;
  assign new_new_n3105__ = new_new_n3103__ & new_new_n3104__;
  assign new_new_n3106__ = new_new_n3102__ & new_new_n3105__;
  assign new_new_n3107__ = new_new_n1677__ & new_new_n2850__;
  assign new_new_n3108__ = new_new_n3101__ & new_new_n3107__;
  assign new_new_n3109__ = new_new_n3100__ & new_new_n3106__;
  assign new_new_n3110__ = new_new_n3108__ & new_new_n3109__;
  assign new_new_n3111__ = ~new_new_n82__ & ~new_new_n284__;
  assign new_new_n3112__ = ~new_new_n656__ & ~new_new_n778__;
  assign new_new_n3113__ = ~new_new_n896__ & new_new_n3112__;
  assign new_new_n3114__ = new_new_n2171__ & new_new_n3111__;
  assign new_new_n3115__ = new_new_n3113__ & new_new_n3114__;
  assign new_new_n3116__ = new_new_n2992__ & new_new_n3096__;
  assign new_new_n3117__ = new_new_n3115__ & new_new_n3116__;
  assign new_new_n3118__ = new_new_n245__ & new_new_n256__;
  assign new_new_n3119__ = new_new_n3098__ & new_new_n3099__;
  assign new_new_n3120__ = new_new_n3118__ & new_new_n3119__;
  assign new_new_n3121__ = new_new_n3095__ & new_new_n3117__;
  assign new_new_n3122__ = new_new_n3120__ & new_new_n3121__;
  assign new_new_n3123__ = new_new_n3110__ & new_new_n3122__;
  assign new_new_n3124__ = new_new_n3075__ & new_new_n3123__;
  assign new_new_n3125__ = new_new_n2939__ & new_new_n3090__;
  assign new_new_n3126__ = new_new_n3124__ & new_new_n3125__;
  assign new_new_n3127__ = ~new_new_n3055__ & ~new_new_n3126__;
  assign new_new_n3128__ = ~new_new_n693__ & ~new_new_n1109__;
  assign new_new_n3129__ = ~new_new_n196__ & ~new_new_n1035__;
  assign new_new_n3130__ = ~new_new_n441__ & ~new_new_n963__;
  assign new_new_n3131__ = ~new_new_n1080__ & new_new_n3130__;
  assign new_new_n3132__ = ~new_new_n1003__ & new_new_n3131__;
  assign new_new_n3133__ = ~new_new_n138__ & ~new_new_n476__;
  assign new_new_n3134__ = ~new_new_n427__ & new_new_n3133__;
  assign new_new_n3135__ = new_new_n1473__ & new_new_n3134__;
  assign new_new_n3136__ = new_new_n3129__ & new_new_n3135__;
  assign new_new_n3137__ = new_new_n3132__ & new_new_n3136__;
  assign new_new_n3138__ = ~new_new_n828__ & ~new_new_n1291__;
  assign new_new_n3139__ = ~new_new_n280__ & ~new_new_n937__;
  assign new_new_n3140__ = ~new_new_n115__ & ~new_new_n961__;
  assign new_new_n3141__ = ~new_new_n267__ & ~new_new_n480__;
  assign new_new_n3142__ = ~new_new_n940__ & ~new_new_n1007__;
  assign new_new_n3143__ = ~new_new_n1031__ & new_new_n3142__;
  assign new_new_n3144__ = ~new_new_n270__ & new_new_n497__;
  assign new_new_n3145__ = new_new_n1678__ & new_new_n3141__;
  assign new_new_n3146__ = new_new_n3144__ & new_new_n3145__;
  assign new_new_n3147__ = new_new_n744__ & new_new_n3143__;
  assign new_new_n3148__ = new_new_n2236__ & new_new_n3147__;
  assign new_new_n3149__ = new_new_n3140__ & new_new_n3146__;
  assign new_new_n3150__ = new_new_n3148__ & new_new_n3149__;
  assign new_new_n3151__ = ~new_new_n207__ & ~new_new_n731__;
  assign new_new_n3152__ = ~new_new_n783__ & new_new_n3151__;
  assign new_new_n3153__ = ~new_new_n488__ & new_new_n3128__;
  assign new_new_n3154__ = new_new_n3152__ & new_new_n3153__;
  assign new_new_n3155__ = ~new_new_n676__ & new_new_n946__;
  assign new_new_n3156__ = new_new_n1564__ & new_new_n3138__;
  assign new_new_n3157__ = new_new_n3139__ & new_new_n3156__;
  assign new_new_n3158__ = new_new_n3154__ & new_new_n3155__;
  assign new_new_n3159__ = new_new_n936__ & new_new_n3158__;
  assign new_new_n3160__ = new_new_n3157__ & new_new_n3159__;
  assign new_new_n3161__ = new_new_n3137__ & new_new_n3150__;
  assign new_new_n3162__ = new_new_n3160__ & new_new_n3161__;
  assign new_new_n3163__ = new_new_n1365__ & new_new_n3162__;
  assign new_new_n3164__ = new_new_n1795__ & new_new_n3163__;
  assign new_new_n3165__ = ~new_new_n2960__ & ~new_new_n3164__;
  assign new_new_n3166__ = ~new_new_n3127__ & ~new_new_n3165__;
  assign new_new_n3167__ = ~new_new_n1167__ & ~new_new_n1372__;
  assign new_new_n3168__ = ~new_new_n388__ & ~new_new_n1398__;
  assign new_new_n3169__ = ~new_new_n308__ & ~new_new_n427__;
  assign new_new_n3170__ = new_new_n3168__ & new_new_n3169__;
  assign new_new_n3171__ = ~new_new_n1539__ & new_new_n3170__;
  assign new_new_n3172__ = ~new_new_n143__ & ~new_new_n933__;
  assign new_new_n3173__ = ~new_new_n207__ & ~new_new_n1031__;
  assign new_new_n3174__ = ~new_new_n696__ & new_new_n3173__;
  assign new_new_n3175__ = ~new_new_n1064__ & new_new_n3174__;
  assign new_new_n3176__ = new_new_n3167__ & new_new_n3172__;
  assign new_new_n3177__ = new_new_n3175__ & new_new_n3176__;
  assign new_new_n3178__ = new_new_n3171__ & new_new_n3177__;
  assign new_new_n3179__ = ~new_new_n249__ & ~new_new_n624__;
  assign new_new_n3180__ = new_new_n1145__ & new_new_n1645__;
  assign new_new_n3181__ = ~new_new_n382__ & ~new_new_n1009__;
  assign new_new_n3182__ = ~new_new_n211__ & ~new_new_n328__;
  assign new_new_n3183__ = ~new_new_n333__ & ~new_new_n3182__;
  assign new_new_n3184__ = ~new_new_n1113__ & ~new_new_n1176__;
  assign new_new_n3185__ = ~new_new_n130__ & ~new_new_n258__;
  assign new_new_n3186__ = ~new_new_n137__ & ~new_new_n217__;
  assign new_new_n3187__ = new_new_n163__ & ~new_new_n3186__;
  assign new_new_n3188__ = ~new_new_n635__ & ~new_new_n723__;
  assign new_new_n3189__ = ~new_new_n675__ & new_new_n3184__;
  assign new_new_n3190__ = ~new_new_n3187__ & new_new_n3189__;
  assign new_new_n3191__ = new_new_n3185__ & new_new_n3188__;
  assign new_new_n3192__ = new_new_n3190__ & new_new_n3191__;
  assign new_new_n3193__ = ~new_new_n101__ & ~new_new_n242__;
  assign new_new_n3194__ = ~new_new_n103__ & ~new_new_n511__;
  assign new_new_n3195__ = ~new_new_n604__ & ~new_new_n729__;
  assign new_new_n3196__ = ~new_new_n336__ & ~new_new_n826__;
  assign new_new_n3197__ = ~new_new_n602__ & new_new_n3196__;
  assign new_new_n3198__ = new_new_n3193__ & new_new_n3194__;
  assign new_new_n3199__ = new_new_n3195__ & new_new_n3198__;
  assign new_new_n3200__ = ~new_new_n508__ & new_new_n3197__;
  assign new_new_n3201__ = new_new_n3199__ & new_new_n3200__;
  assign new_new_n3202__ = ~new_new_n348__ & ~new_new_n890__;
  assign new_new_n3203__ = ~new_new_n270__ & ~new_new_n379__;
  assign new_new_n3204__ = ~new_new_n298__ & ~new_new_n658__;
  assign new_new_n3205__ = ~new_new_n229__ & ~new_new_n700__;
  assign new_new_n3206__ = ~new_new_n252__ & ~new_new_n286__;
  assign new_new_n3207__ = ~new_new_n835__ & ~new_new_n1701__;
  assign new_new_n3208__ = new_new_n2476__ & new_new_n3207__;
  assign new_new_n3209__ = ~new_new_n476__ & ~new_new_n996__;
  assign new_new_n3210__ = ~new_new_n853__ & ~new_new_n2170__;
  assign new_new_n3211__ = ~new_new_n235__ & ~new_new_n317__;
  assign new_new_n3212__ = ~new_new_n160__ & ~new_new_n482__;
  assign new_new_n3213__ = ~new_new_n634__ & new_new_n3212__;
  assign new_new_n3214__ = ~new_new_n332__ & new_new_n1773__;
  assign new_new_n3215__ = new_new_n3209__ & new_new_n3210__;
  assign new_new_n3216__ = new_new_n3214__ & new_new_n3215__;
  assign new_new_n3217__ = ~new_new_n124__ & new_new_n3213__;
  assign new_new_n3218__ = new_new_n3206__ & new_new_n3211__;
  assign new_new_n3219__ = new_new_n3217__ & new_new_n3218__;
  assign new_new_n3220__ = new_new_n3208__ & new_new_n3216__;
  assign new_new_n3221__ = new_new_n3219__ & new_new_n3220__;
  assign new_new_n3222__ = ~new_new_n200__ & ~new_new_n692__;
  assign new_new_n3223__ = ~new_new_n749__ & ~new_new_n990__;
  assign new_new_n3224__ = new_new_n3222__ & new_new_n3223__;
  assign new_new_n3225__ = ~new_new_n993__ & new_new_n1169__;
  assign new_new_n3226__ = new_new_n2944__ & new_new_n3204__;
  assign new_new_n3227__ = new_new_n3205__ & new_new_n3226__;
  assign new_new_n3228__ = new_new_n3224__ & new_new_n3225__;
  assign new_new_n3229__ = ~new_new_n316__ & new_new_n2005__;
  assign new_new_n3230__ = new_new_n2161__ & new_new_n3202__;
  assign new_new_n3231__ = new_new_n3203__ & new_new_n3230__;
  assign new_new_n3232__ = new_new_n3228__ & new_new_n3229__;
  assign new_new_n3233__ = new_new_n1514__ & new_new_n3227__;
  assign new_new_n3234__ = new_new_n3232__ & new_new_n3233__;
  assign new_new_n3235__ = new_new_n3201__ & new_new_n3231__;
  assign new_new_n3236__ = new_new_n3234__ & new_new_n3235__;
  assign new_new_n3237__ = new_new_n3221__ & new_new_n3236__;
  assign new_new_n3238__ = ~new_new_n92__ & ~new_new_n96__;
  assign new_new_n3239__ = ~new_new_n108__ & ~new_new_n240__;
  assign new_new_n3240__ = ~new_new_n267__ & new_new_n1086__;
  assign new_new_n3241__ = new_new_n3238__ & new_new_n3239__;
  assign new_new_n3242__ = ~new_new_n721__ & new_new_n1214__;
  assign new_new_n3243__ = ~new_new_n1568__ & new_new_n3179__;
  assign new_new_n3244__ = new_new_n3242__ & new_new_n3243__;
  assign new_new_n3245__ = new_new_n3240__ & new_new_n3241__;
  assign new_new_n3246__ = new_new_n3181__ & ~new_new_n3183__;
  assign new_new_n3247__ = new_new_n3245__ & new_new_n3246__;
  assign new_new_n3248__ = new_new_n3180__ & new_new_n3244__;
  assign new_new_n3249__ = new_new_n3247__ & new_new_n3248__;
  assign new_new_n3250__ = new_new_n2620__ & new_new_n3192__;
  assign new_new_n3251__ = new_new_n3249__ & new_new_n3250__;
  assign new_new_n3252__ = new_new_n3178__ & new_new_n3251__;
  assign new_new_n3253__ = new_new_n3009__ & new_new_n3252__;
  assign new_new_n3254__ = new_new_n3237__ & new_new_n3253__;
  assign new_new_n3255__ = ~new_new_n3166__ & ~new_new_n3254__;
  assign new_new_n3256__ = ~new_new_n3126__ & ~new_new_n3164__;
  assign new_new_n3257__ = new_new_n2960__ & ~new_new_n3256__;
  assign new_new_n3258__ = ~new_new_n76__ & ~new_new_n282__;
  assign new_new_n3259__ = ~new_new_n254__ & ~new_new_n778__;
  assign new_new_n3260__ = ~new_new_n329__ & ~new_new_n896__;
  assign new_new_n3261__ = ~new_new_n249__ & new_new_n944__;
  assign new_new_n3262__ = ~new_new_n166__ & ~new_new_n658__;
  assign new_new_n3263__ = ~new_new_n250__ & ~new_new_n959__;
  assign new_new_n3264__ = ~new_new_n222__ & ~new_new_n259__;
  assign new_new_n3265__ = ~new_new_n441__ & new_new_n3264__;
  assign new_new_n3266__ = ~new_new_n350__ & ~new_new_n427__;
  assign new_new_n3267__ = ~new_new_n1009__ & new_new_n3266__;
  assign new_new_n3268__ = new_new_n1679__ & new_new_n3265__;
  assign new_new_n3269__ = new_new_n2161__ & new_new_n3262__;
  assign new_new_n3270__ = new_new_n3263__ & new_new_n3269__;
  assign new_new_n3271__ = new_new_n3267__ & new_new_n3268__;
  assign new_new_n3272__ = ~new_new_n668__ & new_new_n3271__;
  assign new_new_n3273__ = new_new_n3270__ & new_new_n3272__;
  assign new_new_n3274__ = ~new_new_n375__ & ~new_new_n878__;
  assign new_new_n3275__ = ~new_new_n1539__ & new_new_n3274__;
  assign new_new_n3276__ = ~new_new_n379__ & ~new_new_n635__;
  assign new_new_n3277__ = ~new_new_n719__ & ~new_new_n845__;
  assign new_new_n3278__ = ~new_new_n252__ & new_new_n3276__;
  assign new_new_n3279__ = new_new_n3277__ & new_new_n3278__;
  assign new_new_n3280__ = ~new_new_n657__ & ~new_new_n874__;
  assign new_new_n3281__ = new_new_n1145__ & new_new_n1263__;
  assign new_new_n3282__ = ~new_new_n673__ & ~new_new_n995__;
  assign new_new_n3283__ = ~new_new_n336__ & ~new_new_n783__;
  assign new_new_n3284__ = ~new_new_n1035__ & ~new_new_n1515__;
  assign new_new_n3285__ = ~new_new_n510__ & ~new_new_n846__;
  assign new_new_n3286__ = ~new_new_n835__ & new_new_n3285__;
  assign new_new_n3287__ = ~new_new_n952__ & new_new_n1332__;
  assign new_new_n3288__ = new_new_n1742__ & new_new_n3283__;
  assign new_new_n3289__ = new_new_n3287__ & new_new_n3288__;
  assign new_new_n3290__ = new_new_n3202__ & new_new_n3286__;
  assign new_new_n3291__ = new_new_n3282__ & new_new_n3284__;
  assign new_new_n3292__ = new_new_n3290__ & new_new_n3291__;
  assign new_new_n3293__ = new_new_n3289__ & new_new_n3292__;
  assign new_new_n3294__ = ~new_new_n595__ & ~new_new_n1372__;
  assign new_new_n3295__ = ~new_new_n309__ & ~new_new_n511__;
  assign new_new_n3296__ = ~new_new_n826__ & new_new_n3295__;
  assign new_new_n3297__ = ~new_new_n226__ & ~new_new_n306__;
  assign new_new_n3298__ = ~new_new_n321__ & new_new_n672__;
  assign new_new_n3299__ = new_new_n1284__ & new_new_n3298__;
  assign new_new_n3300__ = new_new_n3296__ & new_new_n3297__;
  assign new_new_n3301__ = new_new_n2852__ & new_new_n2911__;
  assign new_new_n3302__ = new_new_n3091__ & new_new_n3280__;
  assign new_new_n3303__ = new_new_n3294__ & new_new_n3302__;
  assign new_new_n3304__ = new_new_n3300__ & new_new_n3301__;
  assign new_new_n3305__ = new_new_n3281__ & new_new_n3299__;
  assign new_new_n3306__ = new_new_n3304__ & new_new_n3305__;
  assign new_new_n3307__ = new_new_n3275__ & new_new_n3303__;
  assign new_new_n3308__ = new_new_n3279__ & new_new_n3307__;
  assign new_new_n3309__ = new_new_n3293__ & new_new_n3306__;
  assign new_new_n3310__ = new_new_n3308__ & new_new_n3309__;
  assign new_new_n3311__ = ~new_new_n110__ & ~new_new_n550__;
  assign new_new_n3312__ = new_new_n587__ & new_new_n3311__;
  assign new_new_n3313__ = ~new_new_n843__ & ~new_new_n875__;
  assign new_new_n3314__ = new_new_n1565__ & new_new_n3313__;
  assign new_new_n3315__ = ~new_new_n3312__ & new_new_n3314__;
  assign new_new_n3316__ = ~new_new_n652__ & new_new_n3315__;
  assign new_new_n3317__ = ~new_new_n115__ & ~new_new_n218__;
  assign new_new_n3318__ = ~new_new_n150__ & ~new_new_n1031__;
  assign new_new_n3319__ = new_new_n1037__ & ~new_new_n1210__;
  assign new_new_n3320__ = ~new_new_n439__ & ~new_new_n884__;
  assign new_new_n3321__ = ~new_new_n138__ & ~new_new_n607__;
  assign new_new_n3322__ = ~new_new_n148__ & ~new_new_n715__;
  assign new_new_n3323__ = new_new_n275__ & new_new_n3322__;
  assign new_new_n3324__ = new_new_n3320__ & new_new_n3323__;
  assign new_new_n3325__ = new_new_n3321__ & new_new_n3324__;
  assign new_new_n3326__ = ~new_new_n209__ & ~new_new_n231__;
  assign new_new_n3327__ = ~new_new_n189__ & new_new_n3326__;
  assign new_new_n3328__ = ~new_new_n311__ & ~new_new_n919__;
  assign new_new_n3329__ = new_new_n1154__ & new_new_n3328__;
  assign new_new_n3330__ = ~new_new_n124__ & new_new_n3327__;
  assign new_new_n3331__ = new_new_n1422__ & new_new_n3318__;
  assign new_new_n3332__ = new_new_n3330__ & new_new_n3331__;
  assign new_new_n3333__ = new_new_n2028__ & new_new_n3329__;
  assign new_new_n3334__ = new_new_n3317__ & new_new_n3319__;
  assign new_new_n3335__ = new_new_n3333__ & new_new_n3334__;
  assign new_new_n3336__ = new_new_n3316__ & new_new_n3332__;
  assign new_new_n3337__ = new_new_n3335__ & new_new_n3336__;
  assign new_new_n3338__ = new_new_n3325__ & new_new_n3337__;
  assign new_new_n3339__ = ~new_new_n1212__ & new_new_n1903__;
  assign new_new_n3340__ = ~new_new_n143__ & ~new_new_n277__;
  assign new_new_n3341__ = ~new_new_n588__ & ~new_new_n921__;
  assign new_new_n3342__ = new_new_n2477__ & new_new_n3258__;
  assign new_new_n3343__ = new_new_n3341__ & new_new_n3342__;
  assign new_new_n3344__ = new_new_n3339__ & new_new_n3340__;
  assign new_new_n3345__ = new_new_n542__ & new_new_n2331__;
  assign new_new_n3346__ = new_new_n2821__ & new_new_n3260__;
  assign new_new_n3347__ = new_new_n3345__ & new_new_n3346__;
  assign new_new_n3348__ = new_new_n3343__ & new_new_n3344__;
  assign new_new_n3349__ = new_new_n486__ & new_new_n2641__;
  assign new_new_n3350__ = new_new_n3259__ & new_new_n3261__;
  assign new_new_n3351__ = new_new_n3349__ & new_new_n3350__;
  assign new_new_n3352__ = new_new_n3347__ & new_new_n3348__;
  assign new_new_n3353__ = new_new_n3351__ & new_new_n3352__;
  assign new_new_n3354__ = new_new_n3273__ & new_new_n3353__;
  assign new_new_n3355__ = new_new_n3310__ & new_new_n3354__;
  assign new_new_n3356__ = new_new_n3338__ & new_new_n3355__;
  assign new_new_n3357__ = ~new_new_n3055__ & ~new_new_n3164__;
  assign new_new_n3358__ = ~new_new_n3356__ & new_new_n3357__;
  assign new_new_n3359__ = new_new_n3126__ & ~new_new_n3358__;
  assign new_new_n3360__ = ~new_new_n3257__ & ~new_new_n3359__;
  assign new_new_n3361__ = ~new_new_n3255__ & ~new_new_n3360__;
  assign new_new_n3362__ = new_new_n2961__ & new_new_n3361__;
  assign new_new_n3363__ = ~new_new_n274__ & ~new_new_n1031__;
  assign new_new_n3364__ = ~new_new_n76__ & ~new_new_n385__;
  assign new_new_n3365__ = ~new_new_n329__ & new_new_n3364__;
  assign new_new_n3366__ = ~new_new_n119__ & ~new_new_n445__;
  assign new_new_n3367__ = ~new_new_n1035__ & new_new_n3366__;
  assign new_new_n3368__ = ~new_new_n240__ & ~new_new_n919__;
  assign new_new_n3369__ = ~new_new_n271__ & ~new_new_n372__;
  assign new_new_n3370__ = ~new_new_n698__ & ~new_new_n721__;
  assign new_new_n3371__ = ~new_new_n489__ & ~new_new_n933__;
  assign new_new_n3372__ = ~new_new_n1507__ & new_new_n3371__;
  assign new_new_n3373__ = new_new_n1164__ & new_new_n3370__;
  assign new_new_n3374__ = new_new_n3372__ & new_new_n3373__;
  assign new_new_n3375__ = ~new_new_n604__ & ~new_new_n1070__;
  assign new_new_n3376__ = new_new_n1680__ & new_new_n3375__;
  assign new_new_n3377__ = new_new_n3363__ & new_new_n3365__;
  assign new_new_n3378__ = new_new_n3367__ & new_new_n3368__;
  assign new_new_n3379__ = new_new_n3369__ & new_new_n3378__;
  assign new_new_n3380__ = new_new_n3376__ & new_new_n3377__;
  assign new_new_n3381__ = new_new_n1566__ & new_new_n3380__;
  assign new_new_n3382__ = new_new_n3374__ & new_new_n3379__;
  assign new_new_n3383__ = new_new_n3381__ & new_new_n3382__;
  assign new_new_n3384__ = new_new_n2969__ & new_new_n3383__;
  assign new_new_n3385__ = ~new_new_n853__ & new_new_n948__;
  assign new_new_n3386__ = ~new_new_n127__ & ~new_new_n878__;
  assign new_new_n3387__ = ~new_new_n768__ & ~new_new_n884__;
  assign new_new_n3388__ = ~new_new_n1176__ & new_new_n3386__;
  assign new_new_n3389__ = new_new_n3387__ & new_new_n3388__;
  assign new_new_n3390__ = ~new_new_n208__ & ~new_new_n477__;
  assign new_new_n3391__ = ~new_new_n302__ & ~new_new_n441__;
  assign new_new_n3392__ = ~new_new_n694__ & ~new_new_n950__;
  assign new_new_n3393__ = ~new_new_n508__ & ~new_new_n1212__;
  assign new_new_n3394__ = ~new_new_n260__ & ~new_new_n606__;
  assign new_new_n3395__ = new_new_n3392__ & new_new_n3394__;
  assign new_new_n3396__ = new_new_n3393__ & new_new_n3395__;
  assign new_new_n3397__ = ~new_new_n473__ & ~new_new_n1343__;
  assign new_new_n3398__ = ~new_new_n749__ & ~new_new_n945__;
  assign new_new_n3399__ = ~new_new_n222__ & ~new_new_n940__;
  assign new_new_n3400__ = ~new_new_n232__ & new_new_n3399__;
  assign new_new_n3401__ = new_new_n3391__ & new_new_n3397__;
  assign new_new_n3402__ = new_new_n3400__ & new_new_n3401__;
  assign new_new_n3403__ = ~new_new_n373__ & new_new_n1097__;
  assign new_new_n3404__ = new_new_n3385__ & new_new_n3390__;
  assign new_new_n3405__ = new_new_n3398__ & new_new_n3404__;
  assign new_new_n3406__ = new_new_n3402__ & new_new_n3403__;
  assign new_new_n3407__ = new_new_n1338__ & ~new_new_n1539__;
  assign new_new_n3408__ = new_new_n2709__ & new_new_n3022__;
  assign new_new_n3409__ = new_new_n3407__ & new_new_n3408__;
  assign new_new_n3410__ = new_new_n3405__ & new_new_n3406__;
  assign new_new_n3411__ = new_new_n3389__ & new_new_n3396__;
  assign new_new_n3412__ = new_new_n3410__ & new_new_n3411__;
  assign new_new_n3413__ = new_new_n3409__ & new_new_n3412__;
  assign new_new_n3414__ = ~new_new_n374__ & ~new_new_n843__;
  assign new_new_n3415__ = ~new_new_n103__ & ~new_new_n729__;
  assign new_new_n3416__ = ~new_new_n438__ & ~new_new_n828__;
  assign new_new_n3417__ = ~new_new_n439__ & new_new_n3416__;
  assign new_new_n3418__ = ~new_new_n937__ & ~new_new_n2170__;
  assign new_new_n3419__ = ~new_new_n136__ & ~new_new_n196__;
  assign new_new_n3420__ = ~new_new_n270__ & ~new_new_n300__;
  assign new_new_n3421__ = ~new_new_n160__ & ~new_new_n624__;
  assign new_new_n3422__ = ~new_new_n869__ & new_new_n3421__;
  assign new_new_n3423__ = new_new_n2425__ & new_new_n3415__;
  assign new_new_n3424__ = new_new_n3418__ & new_new_n3423__;
  assign new_new_n3425__ = ~new_new_n218__ & new_new_n3422__;
  assign new_new_n3426__ = new_new_n3419__ & new_new_n3420__;
  assign new_new_n3427__ = new_new_n3425__ & new_new_n3426__;
  assign new_new_n3428__ = new_new_n3417__ & new_new_n3424__;
  assign new_new_n3429__ = new_new_n3427__ & new_new_n3428__;
  assign new_new_n3430__ = ~new_new_n209__ & ~new_new_n634__;
  assign new_new_n3431__ = ~new_new_n101__ & ~new_new_n472__;
  assign new_new_n3432__ = ~new_new_n603__ & ~new_new_n656__;
  assign new_new_n3433__ = ~new_new_n671__ & ~new_new_n963__;
  assign new_new_n3434__ = new_new_n3432__ & new_new_n3433__;
  assign new_new_n3435__ = ~new_new_n348__ & new_new_n3431__;
  assign new_new_n3436__ = new_new_n3430__ & new_new_n3435__;
  assign new_new_n3437__ = new_new_n2769__ & new_new_n3434__;
  assign new_new_n3438__ = new_new_n3436__ & new_new_n3437__;
  assign new_new_n3439__ = ~new_new_n207__ & ~new_new_n425__;
  assign new_new_n3440__ = ~new_new_n249__ & ~new_new_n267__;
  assign new_new_n3441__ = ~new_new_n496__ & ~new_new_n632__;
  assign new_new_n3442__ = ~new_new_n637__ & ~new_new_n811__;
  assign new_new_n3443__ = ~new_new_n995__ & ~new_new_n1007__;
  assign new_new_n3444__ = ~new_new_n1372__ & new_new_n3443__;
  assign new_new_n3445__ = new_new_n3441__ & new_new_n3442__;
  assign new_new_n3446__ = ~new_new_n277__ & new_new_n3440__;
  assign new_new_n3447__ = ~new_new_n1003__ & new_new_n1709__;
  assign new_new_n3448__ = new_new_n3414__ & new_new_n3439__;
  assign new_new_n3449__ = new_new_n3447__ & new_new_n3448__;
  assign new_new_n3450__ = new_new_n340__ & new_new_n3446__;
  assign new_new_n3451__ = new_new_n3444__ & new_new_n3445__;
  assign new_new_n3452__ = ~new_new_n124__ & new_new_n2653__;
  assign new_new_n3453__ = new_new_n3451__ & new_new_n3452__;
  assign new_new_n3454__ = new_new_n3449__ & new_new_n3450__;
  assign new_new_n3455__ = new_new_n1608__ & new_new_n3454__;
  assign new_new_n3456__ = new_new_n3438__ & new_new_n3453__;
  assign new_new_n3457__ = new_new_n3455__ & new_new_n3456__;
  assign new_new_n3458__ = new_new_n3429__ & new_new_n3457__;
  assign new_new_n3459__ = new_new_n3384__ & new_new_n3458__;
  assign new_new_n3460__ = new_new_n3413__ & new_new_n3459__;
  assign new_new_n3461__ = new_new_n2886__ & new_new_n3460__;
  assign new_new_n3462__ = ~new_new_n3362__ & ~new_new_n3461__;
  assign new_new_n3463__ = new_new_n2960__ & ~new_new_n3462__;
  assign new_new_n3464__ = new_new_n2886__ & new_new_n3361__;
  assign new_new_n3465__ = ~new_new_n2961__ & ~new_new_n3464__;
  assign new_new_n3466__ = new_new_n3460__ & ~new_new_n3465__;
  assign new_new_n3467__ = ~new_new_n2887__ & ~new_new_n3463__;
  assign new_new_n3468__ = ~new_new_n3466__ & new_new_n3467__;
  assign new_new_n3469__ = ~new_new_n2739__ & ~new_new_n3468__;
  assign new_new_n3470__ = new_new_n2572__ & new_new_n2737__;
  assign new_new_n3471__ = ~new_new_n2638__ & ~new_new_n3470__;
  assign new_new_n3472__ = new_new_n2636__ & ~new_new_n3471__;
  assign new_new_n3473__ = ~new_new_n2573__ & ~new_new_n3472__;
  assign new_new_n3474__ = ~new_new_n3469__ & new_new_n3473__;
  assign new_new_n3475__ = new_new_n2313__ & ~new_new_n3474__;
  assign new_new_n3476__ = ~new_new_n2420__ & ~new_new_n3475__;
  assign new_new_n3477__ = new_new_n2130__ & new_new_n2224__;
  assign new_new_n3478__ = ~new_new_n3476__ & new_new_n3477__;
  assign new_new_n3479__ = ~new_new_n2423__ & ~new_new_n3478__;
  assign new_new_n3480__ = new_new_n1902__ & ~new_new_n3479__;
  assign new_new_n3481__ = ~new_new_n1824__ & ~new_new_n3480__;
  assign new_new_n3482__ = ~new_new_n213__ & ~new_new_n781__;
  assign new_new_n3483__ = ~new_new_n207__ & ~new_new_n950__;
  assign new_new_n3484__ = ~new_new_n675__ & ~new_new_n1094__;
  assign new_new_n3485__ = ~new_new_n271__ & ~new_new_n511__;
  assign new_new_n3486__ = ~new_new_n179__ & ~new_new_n495__;
  assign new_new_n3487__ = ~new_new_n168__ & ~new_new_n251__;
  assign new_new_n3488__ = ~new_new_n335__ & new_new_n3487__;
  assign new_new_n3489__ = new_new_n93__ & ~new_new_n321__;
  assign new_new_n3490__ = new_new_n3486__ & new_new_n3489__;
  assign new_new_n3491__ = new_new_n199__ & new_new_n3488__;
  assign new_new_n3492__ = new_new_n1078__ & new_new_n1340__;
  assign new_new_n3493__ = new_new_n2653__ & new_new_n3280__;
  assign new_new_n3494__ = new_new_n3492__ & new_new_n3493__;
  assign new_new_n3495__ = new_new_n3490__ & new_new_n3491__;
  assign new_new_n3496__ = new_new_n3494__ & new_new_n3495__;
  assign new_new_n3497__ = ~new_new_n940__ & new_new_n2099__;
  assign new_new_n3498__ = new_new_n2160__ & new_new_n3210__;
  assign new_new_n3499__ = new_new_n3483__ & new_new_n3485__;
  assign new_new_n3500__ = new_new_n3498__ & new_new_n3499__;
  assign new_new_n3501__ = new_new_n944__ & new_new_n3497__;
  assign new_new_n3502__ = new_new_n1114__ & new_new_n1471__;
  assign new_new_n3503__ = new_new_n1707__ & new_new_n2549__;
  assign new_new_n3504__ = new_new_n2710__ & new_new_n3484__;
  assign new_new_n3505__ = new_new_n3503__ & new_new_n3504__;
  assign new_new_n3506__ = new_new_n3501__ & new_new_n3502__;
  assign new_new_n3507__ = new_new_n1826__ & new_new_n3500__;
  assign new_new_n3508__ = new_new_n2700__ & new_new_n3507__;
  assign new_new_n3509__ = new_new_n3505__ & new_new_n3506__;
  assign new_new_n3510__ = new_new_n2757__ & new_new_n3509__;
  assign new_new_n3511__ = new_new_n3496__ & new_new_n3508__;
  assign new_new_n3512__ = new_new_n3510__ & new_new_n3511__;
  assign new_new_n3513__ = ~new_new_n280__ & ~new_new_n306__;
  assign new_new_n3514__ = ~new_new_n260__ & ~new_new_n284__;
  assign new_new_n3515__ = ~new_new_n843__ & ~new_new_n1398__;
  assign new_new_n3516__ = new_new_n3514__ & new_new_n3515__;
  assign new_new_n3517__ = ~new_new_n282__ & ~new_new_n875__;
  assign new_new_n3518__ = ~new_new_n390__ & new_new_n3517__;
  assign new_new_n3519__ = ~new_new_n588__ & ~new_new_n869__;
  assign new_new_n3520__ = new_new_n3518__ & new_new_n3519__;
  assign new_new_n3521__ = new_new_n3516__ & new_new_n3520__;
  assign new_new_n3522__ = ~new_new_n488__ & ~new_new_n884__;
  assign new_new_n3523__ = new_new_n1709__ & new_new_n3415__;
  assign new_new_n3524__ = new_new_n3522__ & new_new_n3523__;
  assign new_new_n3525__ = new_new_n2851__ & new_new_n3167__;
  assign new_new_n3526__ = new_new_n3185__ & new_new_n3482__;
  assign new_new_n3527__ = new_new_n3513__ & new_new_n3526__;
  assign new_new_n3528__ = new_new_n3524__ & new_new_n3525__;
  assign new_new_n3529__ = new_new_n1336__ & new_new_n2028__;
  assign new_new_n3530__ = new_new_n3528__ & new_new_n3529__;
  assign new_new_n3531__ = new_new_n3521__ & new_new_n3527__;
  assign new_new_n3532__ = new_new_n3530__ & new_new_n3531__;
  assign new_new_n3533__ = new_new_n1959__ & new_new_n3532__;
  assign new_new_n3534__ = new_new_n2538__ & new_new_n3533__;
  assign new_new_n3535__ = new_new_n3512__ & new_new_n3534__;
  assign new_new_n3536__ = ~new_new_n3481__ & new_new_n3535__;
  assign new_new_n3537__ = new_new_n1902__ & new_new_n3535__;
  assign new_new_n3538__ = new_new_n1824__ & ~new_new_n3479__;
  assign new_new_n3539__ = ~new_new_n3537__ & ~new_new_n3538__;
  assign new_new_n3540__ = new_new_n2130__ & ~new_new_n3539__;
  assign new_new_n3541__ = ~new_new_n1660__ & ~new_new_n1823__;
  assign new_new_n3542__ = new_new_n1902__ & ~new_new_n3541__;
  assign new_new_n3543__ = ~new_new_n3536__ & ~new_new_n3542__;
  assign new_new_n3544__ = ~new_new_n3540__ & new_new_n3543__;
  assign new_new_n3545__ = new_new_n1739__ & new_new_n3544__;
  assign new_new_n3546__ = ~new_new_n1738__ & ~new_new_n3545__;
  assign new_new_n3547__ = ~new_new_n1660__ & ~new_new_n3546__;
  assign new_new_n3548__ = ~new_new_n1556__ & new_new_n3544__;
  assign new_new_n3549__ = ~new_new_n1739__ & ~new_new_n3548__;
  assign new_new_n3550__ = ~new_new_n1737__ & ~new_new_n3549__;
  assign new_new_n3551__ = ~new_new_n1557__ & ~new_new_n3547__;
  assign new_new_n3552__ = ~new_new_n3550__ & new_new_n3551__;
  assign new_new_n3553__ = new_new_n1325__ & new_new_n3552__;
  assign new_new_n3554__ = ~new_new_n1207__ & ~new_new_n3553__;
  assign new_new_n3555__ = new_new_n1061__ & ~new_new_n1208__;
  assign new_new_n3556__ = ~new_new_n3554__ & new_new_n3555__;
  assign new_new_n3557__ = new_new_n1207__ & new_new_n3552__;
  assign new_new_n3558__ = new_new_n868__ & new_new_n1061__;
  assign new_new_n3559__ = ~new_new_n3557__ & ~new_new_n3558__;
  assign new_new_n3560__ = ~new_new_n332__ & new_new_n1448__;
  assign new_new_n3561__ = new_new_n428__ & ~new_new_n835__;
  assign new_new_n3562__ = new_new_n1827__ & new_new_n3561__;
  assign new_new_n3563__ = new_new_n3560__ & new_new_n3562__;
  assign new_new_n3564__ = ~new_new_n375__ & ~new_new_n816__;
  assign new_new_n3565__ = ~new_new_n126__ & ~new_new_n718__;
  assign new_new_n3566__ = new_new_n75__ & ~new_new_n3565__;
  assign new_new_n3567__ = ~new_new_n124__ & ~new_new_n1073__;
  assign new_new_n3568__ = ~new_new_n837__ & ~new_new_n1105__;
  assign new_new_n3569__ = ~new_new_n120__ & ~new_new_n996__;
  assign new_new_n3570__ = ~new_new_n300__ & new_new_n3569__;
  assign new_new_n3571__ = new_new_n1469__ & new_new_n2340__;
  assign new_new_n3572__ = ~new_new_n3566__ & new_new_n3571__;
  assign new_new_n3573__ = new_new_n1611__ & new_new_n3570__;
  assign new_new_n3574__ = new_new_n1707__ & new_new_n2384__;
  assign new_new_n3575__ = new_new_n3564__ & new_new_n3574__;
  assign new_new_n3576__ = new_new_n3572__ & new_new_n3573__;
  assign new_new_n3577__ = ~new_new_n1539__ & new_new_n3567__;
  assign new_new_n3578__ = new_new_n3568__ & new_new_n3577__;
  assign new_new_n3579__ = new_new_n3575__ & new_new_n3576__;
  assign new_new_n3580__ = new_new_n3578__ & new_new_n3579__;
  assign new_new_n3581__ = ~new_new_n168__ & ~new_new_n384__;
  assign new_new_n3582__ = ~new_new_n138__ & ~new_new_n937__;
  assign new_new_n3583__ = ~new_new_n302__ & ~new_new_n919__;
  assign new_new_n3584__ = new_new_n234__ & ~new_new_n355__;
  assign new_new_n3585__ = new_new_n941__ & ~new_new_n3584__;
  assign new_new_n3586__ = ~new_new_n209__ & ~new_new_n630__;
  assign new_new_n3587__ = ~new_new_n88__ & ~new_new_n246__;
  assign new_new_n3588__ = ~new_new_n588__ & ~new_new_n947__;
  assign new_new_n3589__ = ~new_new_n441__ & ~new_new_n698__;
  assign new_new_n3590__ = ~new_new_n380__ & new_new_n3589__;
  assign new_new_n3591__ = ~new_new_n483__ & new_new_n1106__;
  assign new_new_n3592__ = new_new_n1563__ & new_new_n3414__;
  assign new_new_n3593__ = new_new_n3587__ & new_new_n3592__;
  assign new_new_n3594__ = new_new_n3590__ & new_new_n3591__;
  assign new_new_n3595__ = new_new_n999__ & new_new_n1645__;
  assign new_new_n3596__ = new_new_n3076__ & new_new_n3484__;
  assign new_new_n3597__ = new_new_n3588__ & new_new_n3596__;
  assign new_new_n3598__ = new_new_n3594__ & new_new_n3595__;
  assign new_new_n3599__ = new_new_n3585__ & new_new_n3593__;
  assign new_new_n3600__ = new_new_n3586__ & new_new_n3599__;
  assign new_new_n3601__ = new_new_n3597__ & new_new_n3598__;
  assign new_new_n3602__ = new_new_n3600__ & new_new_n3601__;
  assign new_new_n3603__ = ~new_new_n631__ & ~new_new_n963__;
  assign new_new_n3604__ = new_new_n1449__ & new_new_n1942__;
  assign new_new_n3605__ = new_new_n3168__ & new_new_n3581__;
  assign new_new_n3606__ = new_new_n3582__ & new_new_n3605__;
  assign new_new_n3607__ = new_new_n3603__ & new_new_n3604__;
  assign new_new_n3608__ = new_new_n830__ & new_new_n2341__;
  assign new_new_n3609__ = new_new_n3583__ & new_new_n3608__;
  assign new_new_n3610__ = new_new_n3606__ & new_new_n3607__;
  assign new_new_n3611__ = new_new_n2089__ & new_new_n2893__;
  assign new_new_n3612__ = new_new_n3610__ & new_new_n3611__;
  assign new_new_n3613__ = new_new_n3609__ & new_new_n3612__;
  assign new_new_n3614__ = new_new_n3110__ & new_new_n3563__;
  assign new_new_n3615__ = new_new_n3613__ & new_new_n3614__;
  assign new_new_n3616__ = new_new_n3580__ & new_new_n3602__;
  assign new_new_n3617__ = new_new_n3615__ & new_new_n3616__;
  assign new_new_n3618__ = new_new_n763__ & new_new_n3617__;
  assign new_new_n3619__ = ~new_new_n3559__ & new_new_n3618__;
  assign new_new_n3620__ = new_new_n868__ & new_new_n1207__;
  assign new_new_n3621__ = ~new_new_n3556__ & ~new_new_n3620__;
  assign new_new_n3622__ = ~new_new_n3619__ & new_new_n3621__;
  assign new_new_n3623__ = new_new_n912__ & ~new_new_n3622__;
  assign new_new_n3624__ = new_new_n583__ & new_new_n691__;
  assign new_new_n3625__ = ~new_new_n438__ & ~new_new_n604__;
  assign new_new_n3626__ = ~new_new_n103__ & ~new_new_n138__;
  assign new_new_n3627__ = ~new_new_n600__ & new_new_n3626__;
  assign new_new_n3628__ = ~new_new_n286__ & ~new_new_n427__;
  assign new_new_n3629__ = new_new_n3625__ & new_new_n3628__;
  assign new_new_n3630__ = new_new_n1097__ & new_new_n3627__;
  assign new_new_n3631__ = new_new_n3629__ & new_new_n3630__;
  assign new_new_n3632__ = ~new_new_n246__ & ~new_new_n1070__;
  assign new_new_n3633__ = new_new_n256__ & ~new_new_n311__;
  assign new_new_n3634__ = new_new_n131__ & new_new_n830__;
  assign new_new_n3635__ = ~new_new_n232__ & ~new_new_n445__;
  assign new_new_n3636__ = ~new_new_n240__ & ~new_new_n284__;
  assign new_new_n3637__ = ~new_new_n222__ & new_new_n3636__;
  assign new_new_n3638__ = ~new_new_n950__ & ~new_new_n1113__;
  assign new_new_n3639__ = ~new_new_n585__ & ~new_new_n921__;
  assign new_new_n3640__ = ~new_new_n308__ & ~new_new_n935__;
  assign new_new_n3641__ = new_new_n163__ & ~new_new_n1129__;
  assign new_new_n3642__ = ~new_new_n842__ & ~new_new_n1212__;
  assign new_new_n3643__ = ~new_new_n202__ & ~new_new_n584__;
  assign new_new_n3644__ = ~new_new_n3641__ & new_new_n3643__;
  assign new_new_n3645__ = ~new_new_n439__ & new_new_n3642__;
  assign new_new_n3646__ = new_new_n3644__ & new_new_n3645__;
  assign new_new_n3647__ = new_new_n3640__ & new_new_n3646__;
  assign new_new_n3648__ = ~new_new_n242__ & new_new_n1709__;
  assign new_new_n3649__ = new_new_n2131__ & new_new_n3648__;
  assign new_new_n3650__ = ~new_new_n388__ & ~new_new_n624__;
  assign new_new_n3651__ = ~new_new_n380__ & new_new_n3650__;
  assign new_new_n3652__ = ~new_new_n635__ & new_new_n1106__;
  assign new_new_n3653__ = ~new_new_n1217__ & new_new_n1257__;
  assign new_new_n3654__ = new_new_n3638__ & new_new_n3653__;
  assign new_new_n3655__ = new_new_n3651__ & new_new_n3652__;
  assign new_new_n3656__ = new_new_n1848__ & new_new_n2098__;
  assign new_new_n3657__ = new_new_n3637__ & new_new_n3639__;
  assign new_new_n3658__ = new_new_n3656__ & new_new_n3657__;
  assign new_new_n3659__ = new_new_n3654__ & new_new_n3655__;
  assign new_new_n3660__ = new_new_n3649__ & new_new_n3659__;
  assign new_new_n3661__ = new_new_n3658__ & new_new_n3660__;
  assign new_new_n3662__ = new_new_n3647__ & new_new_n3661__;
  assign new_new_n3663__ = ~new_new_n375__ & ~new_new_n701__;
  assign new_new_n3664__ = ~new_new_n1009__ & new_new_n3663__;
  assign new_new_n3665__ = ~new_new_n1064__ & new_new_n1559__;
  assign new_new_n3666__ = new_new_n2267__ & new_new_n3665__;
  assign new_new_n3667__ = new_new_n3076__ & new_new_n3664__;
  assign new_new_n3668__ = new_new_n3666__ & new_new_n3667__;
  assign new_new_n3669__ = ~new_new_n480__ & ~new_new_n700__;
  assign new_new_n3670__ = ~new_new_n778__ & new_new_n3669__;
  assign new_new_n3671__ = ~new_new_n332__ & ~new_new_n939__;
  assign new_new_n3672__ = new_new_n1410__ & ~new_new_n1701__;
  assign new_new_n3673__ = ~new_new_n2329__ & new_new_n2642__;
  assign new_new_n3674__ = new_new_n3632__ & new_new_n3673__;
  assign new_new_n3675__ = new_new_n3671__ & new_new_n3672__;
  assign new_new_n3676__ = ~new_new_n546__ & new_new_n3670__;
  assign new_new_n3677__ = new_new_n1645__ & new_new_n1748__;
  assign new_new_n3678__ = new_new_n3635__ & new_new_n3677__;
  assign new_new_n3679__ = new_new_n3675__ & new_new_n3676__;
  assign new_new_n3680__ = new_new_n3634__ & new_new_n3674__;
  assign new_new_n3681__ = new_new_n3679__ & new_new_n3680__;
  assign new_new_n3682__ = new_new_n3633__ & new_new_n3678__;
  assign new_new_n3683__ = new_new_n3668__ & new_new_n3682__;
  assign new_new_n3684__ = new_new_n3681__ & new_new_n3683__;
  assign new_new_n3685__ = new_new_n3662__ & new_new_n3684__;
  assign new_new_n3686__ = ~new_new_n321__ & ~new_new_n874__;
  assign new_new_n3687__ = ~new_new_n96__ & ~new_new_n143__;
  assign new_new_n3688__ = ~new_new_n209__ & ~new_new_n1080__;
  assign new_new_n3689__ = ~new_new_n212__ & ~new_new_n1515__;
  assign new_new_n3690__ = ~new_new_n106__ & ~new_new_n634__;
  assign new_new_n3691__ = ~new_new_n715__ & ~new_new_n1081__;
  assign new_new_n3692__ = new_new_n3690__ & new_new_n3691__;
  assign new_new_n3693__ = ~new_new_n1507__ & new_new_n3688__;
  assign new_new_n3694__ = new_new_n3689__ & new_new_n3693__;
  assign new_new_n3695__ = ~new_new_n115__ & new_new_n3692__;
  assign new_new_n3696__ = new_new_n3686__ & new_new_n3687__;
  assign new_new_n3697__ = new_new_n3695__ & new_new_n3696__;
  assign new_new_n3698__ = new_new_n3694__ & new_new_n3697__;
  assign new_new_n3699__ = ~new_new_n473__ & new_new_n628__;
  assign new_new_n3700__ = ~new_new_n120__ & ~new_new_n124__;
  assign new_new_n3701__ = ~new_new_n101__ & ~new_new_n312__;
  assign new_new_n3702__ = ~new_new_n510__ & ~new_new_n811__;
  assign new_new_n3703__ = ~new_new_n826__ & ~new_new_n990__;
  assign new_new_n3704__ = new_new_n3702__ & new_new_n3703__;
  assign new_new_n3705__ = ~new_new_n150__ & new_new_n3701__;
  assign new_new_n3706__ = new_new_n2477__ & new_new_n3209__;
  assign new_new_n3707__ = new_new_n3705__ & new_new_n3706__;
  assign new_new_n3708__ = ~new_new_n373__ & new_new_n3704__;
  assign new_new_n3709__ = ~new_new_n630__ & new_new_n913__;
  assign new_new_n3710__ = new_new_n1341__ & new_new_n1970__;
  assign new_new_n3711__ = new_new_n3709__ & new_new_n3710__;
  assign new_new_n3712__ = new_new_n3707__ & new_new_n3708__;
  assign new_new_n3713__ = new_new_n347__ & new_new_n2755__;
  assign new_new_n3714__ = new_new_n3699__ & new_new_n3700__;
  assign new_new_n3715__ = new_new_n3713__ & new_new_n3714__;
  assign new_new_n3716__ = new_new_n3711__ & new_new_n3712__;
  assign new_new_n3717__ = new_new_n3631__ & new_new_n3716__;
  assign new_new_n3718__ = new_new_n3698__ & new_new_n3715__;
  assign new_new_n3719__ = new_new_n3717__ & new_new_n3718__;
  assign new_new_n3720__ = new_new_n3685__ & new_new_n3719__;
  assign new_new_n3721__ = new_new_n3624__ & new_new_n3720__;
  assign new_new_n3722__ = ~new_new_n3623__ & ~new_new_n3721__;
  assign new_new_n3723__ = new_new_n868__ & ~new_new_n3722__;
  assign new_new_n3724__ = ~new_new_n3622__ & new_new_n3624__;
  assign new_new_n3725__ = ~new_new_n912__ & ~new_new_n3724__;
  assign new_new_n3726__ = new_new_n3720__ & ~new_new_n3725__;
  assign new_new_n3727__ = new_new_n691__ & ~new_new_n910__;
  assign new_new_n3728__ = ~new_new_n583__ & new_new_n3727__;
  assign new_new_n3729__ = new_new_n583__ & ~new_new_n691__;
  assign new_new_n3730__ = new_new_n3622__ & new_new_n3729__;
  assign new_new_n3731__ = ~new_new_n3728__ & ~new_new_n3730__;
  assign new_new_n3732__ = ~new_new_n3720__ & ~new_new_n3731__;
  assign new_new_n3733__ = new_new_n3622__ & new_new_n3728__;
  assign new_new_n3734__ = ~new_new_n3720__ & new_new_n3729__;
  assign new_new_n3735__ = ~new_new_n3733__ & ~new_new_n3734__;
  assign new_new_n3736__ = ~new_new_n868__ & ~new_new_n3735__;
  assign new_new_n3737__ = new_new_n583__ & ~new_new_n911__;
  assign new_new_n3738__ = ~new_new_n3727__ & new_new_n3737__;
  assign new_new_n3739__ = ~new_new_n3723__ & ~new_new_n3738__;
  assign new_new_n3740__ = ~new_new_n3726__ & ~new_new_n3732__;
  assign new_new_n3741__ = ~new_new_n3736__ & new_new_n3740__;
  assign new_new_n3742__ = new_new_n3739__ & new_new_n3741__;
  assign new_new_n3743__ = ~new_new_n691__ & ~new_new_n3742__;
  assign new_new_n3744__ = new_new_n583__ & ~new_new_n3743__;
  assign new_new_n3745__ = pi24 & new_new_n430__;
  assign new_new_n3746__ = pi23 & ~new_new_n133__;
  assign new_new_n3747__ = new_new_n550__ & new_new_n3746__;
  assign new_new_n3748__ = ~new_new_n3745__ & ~new_new_n3747__;
  assign new_new_n3749__ = new_new_n126__ & ~new_new_n3748__;
  assign new_new_n3750__ = ~new_new_n86__ & new_new_n3015__;
  assign new_new_n3751__ = new_new_n594__ & new_new_n3750__;
  assign new_new_n3752__ = ~new_new_n585__ & ~new_new_n604__;
  assign new_new_n3753__ = ~new_new_n657__ & new_new_n3752__;
  assign new_new_n3754__ = ~new_new_n588__ & ~new_new_n3751__;
  assign new_new_n3755__ = new_new_n3753__ & new_new_n3754__;
  assign new_new_n3756__ = ~new_new_n3749__ & new_new_n3755__;
  assign new_new_n3757__ = new_new_n149__ & ~new_new_n550__;
  assign new_new_n3758__ = new_new_n126__ & new_new_n447__;
  assign new_new_n3759__ = new_new_n560__ & new_new_n3758__;
  assign new_new_n3760__ = ~new_new_n495__ & ~new_new_n3757__;
  assign new_new_n3761__ = ~new_new_n3759__ & new_new_n3760__;
  assign new_new_n3762__ = new_new_n471__ & new_new_n3761__;
  assign new_new_n3763__ = new_new_n3756__ & new_new_n3762__;
  assign new_new_n3764__ = new_new_n2753__ & new_new_n3763__;
  assign new_new_n3765__ = new_new_n2328__ & new_new_n3764__;
  assign new_new_n3766__ = ~new_new_n88__ & ~new_new_n1372__;
  assign new_new_n3767__ = new_new_n421__ & new_new_n3766__;
  assign new_new_n3768__ = new_new_n3765__ & new_new_n3767__;
  assign new_new_n3769__ = ~new_new_n3744__ & ~new_new_n3768__;
  assign new_new_n3770__ = pi29 & new_new_n3769__;
  assign new_new_n3771__ = new_new_n466__ & ~new_new_n3770__;
  assign new_new_n3772__ = pi31 & ~new_new_n3771__;
  assign new_new_n3773__ = ~new_new_n495__ & ~new_new_n732__;
  assign new_new_n3774__ = ~new_new_n302__ & ~new_new_n479__;
  assign new_new_n3775__ = ~new_new_n838__ & ~new_new_n1033__;
  assign new_new_n3776__ = ~new_new_n248__ & ~new_new_n657__;
  assign new_new_n3777__ = ~new_new_n778__ & new_new_n3776__;
  assign new_new_n3778__ = new_new_n314__ & ~new_new_n348__;
  assign new_new_n3779__ = ~new_new_n673__ & new_new_n745__;
  assign new_new_n3780__ = new_new_n784__ & new_new_n1077__;
  assign new_new_n3781__ = new_new_n3775__ & new_new_n3780__;
  assign new_new_n3782__ = new_new_n3778__ & new_new_n3779__;
  assign new_new_n3783__ = new_new_n3777__ & new_new_n3782__;
  assign new_new_n3784__ = new_new_n3774__ & new_new_n3781__;
  assign new_new_n3785__ = new_new_n3783__ & new_new_n3784__;
  assign new_new_n3786__ = ~new_new_n119__ & new_new_n3773__;
  assign new_new_n3787__ = new_new_n3785__ & new_new_n3786__;
  assign new_new_n3788__ = ~new_new_n658__ & ~new_new_n696__;
  assign new_new_n3789__ = new_new_n163__ & ~new_new_n310__;
  assign new_new_n3790__ = ~new_new_n192__ & ~new_new_n427__;
  assign new_new_n3791__ = ~new_new_n3789__ & new_new_n3790__;
  assign new_new_n3792__ = ~new_new_n306__ & ~new_new_n482__;
  assign new_new_n3793__ = ~new_new_n136__ & ~new_new_n845__;
  assign new_new_n3794__ = ~new_new_n179__ & ~new_new_n896__;
  assign new_new_n3795__ = ~new_new_n120__ & ~new_new_n700__;
  assign new_new_n3796__ = ~new_new_n591__ & new_new_n3795__;
  assign new_new_n3797__ = ~new_new_n675__ & ~new_new_n828__;
  assign new_new_n3798__ = new_new_n3794__ & new_new_n3797__;
  assign new_new_n3799__ = new_new_n1251__ & new_new_n3796__;
  assign new_new_n3800__ = new_new_n3096__ & new_new_n3792__;
  assign new_new_n3801__ = new_new_n3793__ & new_new_n3800__;
  assign new_new_n3802__ = new_new_n3798__ & new_new_n3799__;
  assign new_new_n3803__ = new_new_n3801__ & new_new_n3802__;
  assign new_new_n3804__ = ~new_new_n259__ & ~new_new_n511__;
  assign new_new_n3805__ = ~new_new_n103__ & ~new_new_n723__;
  assign new_new_n3806__ = ~new_new_n155__ & ~new_new_n238__;
  assign new_new_n3807__ = ~new_new_n942__ & ~new_new_n1094__;
  assign new_new_n3808__ = new_new_n2116__ & new_new_n3807__;
  assign new_new_n3809__ = new_new_n3804__ & new_new_n3805__;
  assign new_new_n3810__ = new_new_n3808__ & new_new_n3809__;
  assign new_new_n3811__ = new_new_n628__ & new_new_n962__;
  assign new_new_n3812__ = new_new_n2653__ & new_new_n2778__;
  assign new_new_n3813__ = new_new_n3788__ & new_new_n3806__;
  assign new_new_n3814__ = new_new_n3812__ & new_new_n3813__;
  assign new_new_n3815__ = new_new_n3810__ & new_new_n3811__;
  assign new_new_n3816__ = new_new_n601__ & new_new_n2989__;
  assign new_new_n3817__ = new_new_n3791__ & new_new_n3816__;
  assign new_new_n3818__ = new_new_n3814__ & new_new_n3815__;
  assign new_new_n3819__ = new_new_n2381__ & new_new_n3818__;
  assign new_new_n3820__ = new_new_n1407__ & new_new_n3817__;
  assign new_new_n3821__ = new_new_n3803__ & new_new_n3820__;
  assign new_new_n3822__ = new_new_n3787__ & new_new_n3819__;
  assign new_new_n3823__ = new_new_n3821__ & new_new_n3822__;
  assign new_new_n3824__ = new_new_n1795__ & new_new_n3823__;
  assign new_new_n3825__ = ~pi26 & ~new_new_n141__;
  assign new_new_n3826__ = new_new_n446__ & new_new_n550__;
  assign new_new_n3827__ = ~new_new_n3825__ & ~new_new_n3826__;
  assign new_new_n3828__ = new_new_n97__ & ~new_new_n3827__;
  assign new_new_n3829__ = new_new_n165__ & ~new_new_n429__;
  assign new_new_n3830__ = ~new_new_n447__ & new_new_n3829__;
  assign new_new_n3831__ = ~new_new_n3828__ & ~new_new_n3830__;
  assign new_new_n3832__ = ~new_new_n476__ & ~new_new_n747__;
  assign new_new_n3833__ = ~new_new_n945__ & new_new_n3832__;
  assign new_new_n3834__ = new_new_n1627__ & new_new_n3833__;
  assign new_new_n3835__ = new_new_n651__ & new_new_n3834__;
  assign new_new_n3836__ = ~new_new_n200__ & ~new_new_n896__;
  assign new_new_n3837__ = ~new_new_n120__ & ~new_new_n724__;
  assign new_new_n3838__ = ~new_new_n776__ & new_new_n3837__;
  assign new_new_n3839__ = ~new_new_n198__ & ~new_new_n321__;
  assign new_new_n3840__ = new_new_n527__ & ~new_new_n541__;
  assign new_new_n3841__ = new_new_n659__ & new_new_n3836__;
  assign new_new_n3842__ = new_new_n3840__ & new_new_n3841__;
  assign new_new_n3843__ = new_new_n3838__ & new_new_n3839__;
  assign new_new_n3844__ = new_new_n1804__ & new_new_n3843__;
  assign new_new_n3845__ = new_new_n3831__ & new_new_n3842__;
  assign new_new_n3846__ = new_new_n3844__ & new_new_n3845__;
  assign new_new_n3847__ = new_new_n187__ & new_new_n3846__;
  assign new_new_n3848__ = new_new_n3835__ & new_new_n3847__;
  assign new_new_n3849__ = ~new_new_n3824__ & ~new_new_n3848__;
  assign new_new_n3850__ = new_new_n3824__ & new_new_n3848__;
  assign new_new_n3851__ = ~pi29 & ~new_new_n3850__;
  assign new_new_n3852__ = ~new_new_n3849__ & ~new_new_n3851__;
  assign new_new_n3853__ = ~new_new_n3772__ & new_new_n3852__;
  assign new_new_n3854__ = new_new_n3772__ & ~new_new_n3852__;
  assign new_new_n3855__ = ~new_new_n3853__ & ~new_new_n3854__;
  assign new_new_n3856__ = new_new_n210__ & ~new_new_n959__;
  assign new_new_n3857__ = ~new_new_n1035__ & new_new_n3856__;
  assign new_new_n3858__ = new_new_n628__ & new_new_n3857__;
  assign new_new_n3859__ = new_new_n3756__ & new_new_n3858__;
  assign new_new_n3860__ = ~new_new_n430__ & new_new_n2672__;
  assign new_new_n3861__ = ~pi27 & new_new_n125__;
  assign new_new_n3862__ = ~new_new_n3860__ & ~new_new_n3861__;
  assign new_new_n3863__ = pi28 & ~new_new_n3862__;
  assign new_new_n3864__ = new_new_n86__ & new_new_n191__;
  assign new_new_n3865__ = new_new_n78__ & new_new_n3014__;
  assign new_new_n3866__ = ~new_new_n3864__ & ~new_new_n3865__;
  assign new_new_n3867__ = pi24 & ~new_new_n3866__;
  assign new_new_n3868__ = ~new_new_n634__ & ~new_new_n670__;
  assign new_new_n3869__ = ~new_new_n1064__ & new_new_n3868__;
  assign new_new_n3870__ = new_new_n1847__ & new_new_n3869__;
  assign new_new_n3871__ = new_new_n1947__ & new_new_n2382__;
  assign new_new_n3872__ = new_new_n3870__ & new_new_n3871__;
  assign new_new_n3873__ = ~new_new_n3867__ & new_new_n3872__;
  assign new_new_n3874__ = new_new_n743__ & ~new_new_n3863__;
  assign new_new_n3875__ = new_new_n454__ & new_new_n3874__;
  assign new_new_n3876__ = new_new_n669__ & new_new_n3875__;
  assign new_new_n3877__ = new_new_n187__ & new_new_n3859__;
  assign new_new_n3878__ = new_new_n3873__ & new_new_n3877__;
  assign new_new_n3879__ = new_new_n575__ & new_new_n3876__;
  assign new_new_n3880__ = new_new_n825__ & new_new_n3879__;
  assign new_new_n3881__ = new_new_n3878__ & new_new_n3880__;
  assign new_new_n3882__ = ~new_new_n3855__ & new_new_n3881__;
  assign new_new_n3883__ = new_new_n3855__ & ~new_new_n3881__;
  assign new_new_n3884__ = ~new_new_n3882__ & ~new_new_n3883__;
  assign new_new_n3885__ = ~new_new_n3849__ & ~new_new_n3850__;
  assign new_new_n3886__ = ~pi29 & ~new_new_n3885__;
  assign new_new_n3887__ = pi29 & new_new_n3885__;
  assign new_new_n3888__ = ~new_new_n3886__ & ~new_new_n3887__;
  assign new_new_n3889__ = pi26 & pi27;
  assign new_new_n3890__ = new_new_n220__ & new_new_n3889__;
  assign new_new_n3891__ = ~new_new_n466__ & new_new_n3890__;
  assign new_new_n3892__ = ~pi29 & ~new_new_n3891__;
  assign new_new_n3893__ = ~new_new_n380__ & ~new_new_n749__;
  assign new_new_n3894__ = new_new_n440__ & ~new_new_n1007__;
  assign new_new_n3895__ = new_new_n2888__ & new_new_n3894__;
  assign new_new_n3896__ = ~new_new_n196__ & ~new_new_n249__;
  assign new_new_n3897__ = ~new_new_n990__ & new_new_n3896__;
  assign new_new_n3898__ = new_new_n710__ & ~new_new_n747__;
  assign new_new_n3899__ = new_new_n1154__ & new_new_n3898__;
  assign new_new_n3900__ = new_new_n184__ & new_new_n3897__;
  assign new_new_n3901__ = new_new_n3893__ & new_new_n3900__;
  assign new_new_n3902__ = new_new_n3899__ & new_new_n3901__;
  assign new_new_n3903__ = new_new_n3895__ & new_new_n3902__;
  assign new_new_n3904__ = ~new_new_n300__ & ~new_new_n427__;
  assign new_new_n3905__ = ~new_new_n212__ & ~new_new_n597__;
  assign new_new_n3906__ = ~new_new_n1176__ & new_new_n3905__;
  assign new_new_n3907__ = ~new_new_n373__ & new_new_n3906__;
  assign new_new_n3908__ = new_new_n2376__ & new_new_n3263__;
  assign new_new_n3909__ = new_new_n3904__ & new_new_n3908__;
  assign new_new_n3910__ = new_new_n3907__ & new_new_n3909__;
  assign new_new_n3911__ = ~new_new_n724__ & new_new_n948__;
  assign new_new_n3912__ = ~new_new_n258__ & new_new_n2116__;
  assign new_new_n3913__ = ~new_new_n120__ & ~new_new_n1167__;
  assign new_new_n3914__ = ~new_new_n312__ & ~new_new_n586__;
  assign new_new_n3915__ = ~new_new_n785__ & new_new_n3914__;
  assign new_new_n3916__ = ~new_new_n828__ & ~new_new_n1507__;
  assign new_new_n3917__ = new_new_n2679__ & new_new_n3916__;
  assign new_new_n3918__ = new_new_n2710__ & new_new_n3915__;
  assign new_new_n3919__ = new_new_n2913__ & new_new_n3484__;
  assign new_new_n3920__ = new_new_n3911__ & new_new_n3912__;
  assign new_new_n3921__ = new_new_n3913__ & new_new_n3920__;
  assign new_new_n3922__ = new_new_n3918__ & new_new_n3919__;
  assign new_new_n3923__ = new_new_n1152__ & new_new_n3917__;
  assign new_new_n3924__ = new_new_n2605__ & new_new_n3923__;
  assign new_new_n3925__ = new_new_n3921__ & new_new_n3922__;
  assign new_new_n3926__ = new_new_n3924__ & new_new_n3925__;
  assign new_new_n3927__ = new_new_n3910__ & new_new_n3926__;
  assign new_new_n3928__ = ~new_new_n473__ & ~new_new_n509__;
  assign new_new_n3929__ = ~new_new_n896__ & new_new_n3928__;
  assign new_new_n3930__ = ~new_new_n919__ & new_new_n3929__;
  assign new_new_n3931__ = ~new_new_n248__ & ~new_new_n591__;
  assign new_new_n3932__ = ~new_new_n130__ & ~new_new_n390__;
  assign new_new_n3933__ = new_new_n3931__ & new_new_n3932__;
  assign new_new_n3934__ = ~new_new_n425__ & ~new_new_n715__;
  assign new_new_n3935__ = ~new_new_n838__ & new_new_n3934__;
  assign new_new_n3936__ = ~new_new_n1003__ & new_new_n2001__;
  assign new_new_n3937__ = new_new_n3193__ & new_new_n3936__;
  assign new_new_n3938__ = new_new_n733__ & new_new_n3935__;
  assign new_new_n3939__ = new_new_n744__ & new_new_n2909__;
  assign new_new_n3940__ = new_new_n3588__ & new_new_n3939__;
  assign new_new_n3941__ = new_new_n3937__ & new_new_n3938__;
  assign new_new_n3942__ = new_new_n709__ & new_new_n3930__;
  assign new_new_n3943__ = new_new_n3933__ & new_new_n3942__;
  assign new_new_n3944__ = new_new_n3940__ & new_new_n3941__;
  assign new_new_n3945__ = new_new_n3943__ & new_new_n3944__;
  assign new_new_n3946__ = new_new_n3903__ & new_new_n3945__;
  assign new_new_n3947__ = new_new_n3310__ & new_new_n3946__;
  assign new_new_n3948__ = new_new_n3927__ & new_new_n3947__;
  assign new_new_n3949__ = ~pi26 & ~new_new_n3948__;
  assign new_new_n3950__ = pi26 & new_new_n3948__;
  assign new_new_n3951__ = ~new_new_n308__ & ~new_new_n480__;
  assign new_new_n3952__ = ~new_new_n1176__ & new_new_n3951__;
  assign new_new_n3953__ = ~new_new_n380__ & ~new_new_n1217__;
  assign new_new_n3954__ = new_new_n3952__ & new_new_n3953__;
  assign new_new_n3955__ = new_new_n2499__ & new_new_n3954__;
  assign new_new_n3956__ = ~new_new_n168__ & ~new_new_n719__;
  assign new_new_n3957__ = ~new_new_n717__ & ~new_new_n1372__;
  assign new_new_n3958__ = ~new_new_n940__ & ~new_new_n942__;
  assign new_new_n3959__ = ~new_new_n247__ & ~new_new_n479__;
  assign new_new_n3960__ = ~new_new_n383__ & ~new_new_n586__;
  assign new_new_n3961__ = ~new_new_n1031__ & new_new_n3960__;
  assign new_new_n3962__ = new_new_n2768__ & new_new_n3957__;
  assign new_new_n3963__ = new_new_n3958__ & new_new_n3962__;
  assign new_new_n3964__ = new_new_n3419__ & new_new_n3961__;
  assign new_new_n3965__ = new_new_n3963__ & new_new_n3964__;
  assign new_new_n3966__ = new_new_n3959__ & new_new_n3965__;
  assign new_new_n3967__ = ~new_new_n253__ & ~new_new_n1343__;
  assign new_new_n3968__ = ~new_new_n472__ & ~new_new_n510__;
  assign new_new_n3969__ = ~new_new_n476__ & ~new_new_n635__;
  assign new_new_n3970__ = ~new_new_n138__ & ~new_new_n315__;
  assign new_new_n3971__ = ~new_new_n332__ & new_new_n3970__;
  assign new_new_n3972__ = ~new_new_n747__ & new_new_n779__;
  assign new_new_n3973__ = new_new_n3967__ & new_new_n3968__;
  assign new_new_n3974__ = new_new_n3972__ & new_new_n3973__;
  assign new_new_n3975__ = new_new_n2289__ & new_new_n3971__;
  assign new_new_n3976__ = new_new_n3956__ & new_new_n3969__;
  assign new_new_n3977__ = new_new_n3975__ & new_new_n3976__;
  assign new_new_n3978__ = new_new_n2028__ & new_new_n3974__;
  assign new_new_n3979__ = new_new_n3977__ & new_new_n3978__;
  assign new_new_n3980__ = new_new_n3955__ & new_new_n3979__;
  assign new_new_n3981__ = new_new_n3966__ & new_new_n3980__;
  assign new_new_n3982__ = ~new_new_n316__ & ~new_new_n489__;
  assign new_new_n3983__ = ~new_new_n252__ & ~new_new_n637__;
  assign new_new_n3984__ = ~new_new_n851__ & new_new_n3983__;
  assign new_new_n3985__ = ~new_new_n143__ & ~new_new_n258__;
  assign new_new_n3986__ = ~new_new_n276__ & new_new_n3985__;
  assign new_new_n3987__ = new_new_n3984__ & new_new_n3986__;
  assign new_new_n3988__ = new_new_n3982__ & new_new_n3987__;
  assign new_new_n3989__ = ~new_new_n298__ & ~new_new_n884__;
  assign new_new_n3990__ = new_new_n100__ & ~new_new_n3565__;
  assign new_new_n3991__ = ~new_new_n212__ & ~new_new_n309__;
  assign new_new_n3992__ = ~new_new_n1081__ & new_new_n3991__;
  assign new_new_n3993__ = ~new_new_n306__ & ~new_new_n894__;
  assign new_new_n3994__ = new_new_n1211__ & new_new_n3636__;
  assign new_new_n3995__ = new_new_n3993__ & new_new_n3994__;
  assign new_new_n3996__ = new_new_n1720__ & new_new_n3992__;
  assign new_new_n3997__ = ~new_new_n439__ & new_new_n2770__;
  assign new_new_n3998__ = new_new_n3996__ & new_new_n3997__;
  assign new_new_n3999__ = new_new_n3995__ & new_new_n3998__;
  assign new_new_n4000__ = ~new_new_n776__ & ~new_new_n2170__;
  assign new_new_n4001__ = ~new_new_n222__ & ~new_new_n588__;
  assign new_new_n4002__ = ~new_new_n379__ & ~new_new_n995__;
  assign new_new_n4003__ = ~new_new_n346__ & new_new_n4002__;
  assign new_new_n4004__ = ~new_new_n919__ & ~new_new_n2697__;
  assign new_new_n4005__ = new_new_n3179__ & new_new_n3430__;
  assign new_new_n4006__ = ~new_new_n3990__ & new_new_n4000__;
  assign new_new_n4007__ = new_new_n4005__ & new_new_n4006__;
  assign new_new_n4008__ = new_new_n4003__ & new_new_n4004__;
  assign new_new_n4009__ = ~new_new_n115__ & new_new_n484__;
  assign new_new_n4010__ = new_new_n830__ & new_new_n3989__;
  assign new_new_n4011__ = new_new_n4001__ & new_new_n4010__;
  assign new_new_n4012__ = new_new_n2688__ & new_new_n4009__;
  assign new_new_n4013__ = new_new_n4007__ & new_new_n4008__;
  assign new_new_n4014__ = new_new_n4012__ & new_new_n4013__;
  assign new_new_n4015__ = new_new_n4011__ & new_new_n4014__;
  assign new_new_n4016__ = new_new_n3988__ & new_new_n3999__;
  assign new_new_n4017__ = new_new_n4015__ & new_new_n4016__;
  assign new_new_n4018__ = new_new_n1992__ & new_new_n4017__;
  assign new_new_n4019__ = new_new_n3981__ & new_new_n4018__;
  assign new_new_n4020__ = ~new_new_n3950__ & ~new_new_n4019__;
  assign new_new_n4021__ = ~new_new_n3949__ & ~new_new_n4020__;
  assign new_new_n4022__ = pi30 & ~new_new_n691__;
  assign new_new_n4023__ = ~new_new_n583__ & new_new_n765__;
  assign new_new_n4024__ = ~new_new_n4022__ & ~new_new_n4023__;
  assign new_new_n4025__ = ~pi31 & ~new_new_n4024__;
  assign new_new_n4026__ = ~pi30 & new_new_n583__;
  assign new_new_n4027__ = ~new_new_n161__ & new_new_n691__;
  assign new_new_n4028__ = ~new_new_n4026__ & ~new_new_n4027__;
  assign new_new_n4029__ = ~new_new_n910__ & ~new_new_n3720__;
  assign new_new_n4030__ = ~new_new_n868__ & ~new_new_n3622__;
  assign new_new_n4031__ = new_new_n868__ & new_new_n3622__;
  assign new_new_n4032__ = ~new_new_n4030__ & ~new_new_n4031__;
  assign new_new_n4033__ = new_new_n868__ & new_new_n3720__;
  assign new_new_n4034__ = ~new_new_n868__ & ~new_new_n3720__;
  assign new_new_n4035__ = ~new_new_n4033__ & ~new_new_n4034__;
  assign new_new_n4036__ = new_new_n4032__ & new_new_n4035__;
  assign new_new_n4037__ = new_new_n910__ & new_new_n3720__;
  assign new_new_n4038__ = ~new_new_n4029__ & ~new_new_n4037__;
  assign new_new_n4039__ = ~new_new_n4036__ & new_new_n4038__;
  assign new_new_n4040__ = new_new_n691__ & ~new_new_n4039__;
  assign new_new_n4041__ = ~new_new_n691__ & new_new_n4039__;
  assign new_new_n4042__ = ~new_new_n4040__ & ~new_new_n4041__;
  assign new_new_n4043__ = pi29 & new_new_n3624__;
  assign new_new_n4044__ = ~new_new_n4042__ & new_new_n4043__;
  assign new_new_n4045__ = ~new_new_n4028__ & ~new_new_n4044__;
  assign new_new_n4046__ = ~new_new_n910__ & ~new_new_n4045__;
  assign new_new_n4047__ = ~new_new_n125__ & new_new_n691__;
  assign new_new_n4048__ = new_new_n691__ & new_new_n910__;
  assign new_new_n4049__ = ~new_new_n4039__ & ~new_new_n4048__;
  assign new_new_n4050__ = ~new_new_n583__ & ~new_new_n4047__;
  assign new_new_n4051__ = ~new_new_n4049__ & new_new_n4050__;
  assign new_new_n4052__ = new_new_n583__ & new_new_n910__;
  assign new_new_n4053__ = ~new_new_n4039__ & new_new_n4052__;
  assign new_new_n4054__ = ~new_new_n71__ & ~new_new_n4053__;
  assign new_new_n4055__ = ~new_new_n691__ & ~new_new_n4054__;
  assign new_new_n4056__ = ~new_new_n4051__ & ~new_new_n4055__;
  assign new_new_n4057__ = ~new_new_n4046__ & new_new_n4056__;
  assign new_new_n4058__ = pi31 & ~new_new_n4057__;
  assign new_new_n4059__ = ~new_new_n4025__ & ~new_new_n4058__;
  assign new_new_n4060__ = new_new_n3824__ & ~new_new_n4059__;
  assign new_new_n4061__ = new_new_n4021__ & new_new_n4060__;
  assign new_new_n4062__ = ~new_new_n246__ & ~new_new_n776__;
  assign new_new_n4063__ = ~new_new_n284__ & ~new_new_n510__;
  assign new_new_n4064__ = ~new_new_n963__ & ~new_new_n1372__;
  assign new_new_n4065__ = new_new_n4063__ & new_new_n4064__;
  assign new_new_n4066__ = ~new_new_n166__ & ~new_new_n202__;
  assign new_new_n4067__ = ~new_new_n884__ & new_new_n1333__;
  assign new_new_n4068__ = new_new_n2943__ & new_new_n4062__;
  assign new_new_n4069__ = new_new_n4067__ & new_new_n4068__;
  assign new_new_n4070__ = new_new_n4065__ & new_new_n4066__;
  assign new_new_n4071__ = ~new_new_n1486__ & new_new_n4070__;
  assign new_new_n4072__ = new_new_n4069__ & new_new_n4071__;
  assign new_new_n4073__ = ~new_new_n138__ & ~new_new_n894__;
  assign new_new_n4074__ = ~new_new_n585__ & ~new_new_n1008__;
  assign new_new_n4075__ = ~new_new_n196__ & ~new_new_n374__;
  assign new_new_n4076__ = ~new_new_n729__ & ~new_new_n875__;
  assign new_new_n4077__ = new_new_n4075__ & new_new_n4076__;
  assign new_new_n4078__ = new_new_n131__ & ~new_new_n150__;
  assign new_new_n4079__ = ~new_new_n266__ & ~new_new_n781__;
  assign new_new_n4080__ = ~new_new_n1151__ & new_new_n1177__;
  assign new_new_n4081__ = new_new_n1371__ & new_new_n4080__;
  assign new_new_n4082__ = new_new_n4078__ & new_new_n4079__;
  assign new_new_n4083__ = ~new_new_n676__ & new_new_n4077__;
  assign new_new_n4084__ = new_new_n941__ & new_new_n4073__;
  assign new_new_n4085__ = new_new_n4074__ & new_new_n4084__;
  assign new_new_n4086__ = new_new_n4082__ & new_new_n4083__;
  assign new_new_n4087__ = new_new_n1745__ & new_new_n4081__;
  assign new_new_n4088__ = new_new_n4086__ & new_new_n4087__;
  assign new_new_n4089__ = new_new_n4085__ & new_new_n4088__;
  assign new_new_n4090__ = ~new_new_n348__ & ~new_new_n837__;
  assign new_new_n4091__ = ~new_new_n218__ & ~new_new_n315__;
  assign new_new_n4092__ = ~new_new_n329__ & ~new_new_n1003__;
  assign new_new_n4093__ = ~new_new_n511__ & ~new_new_n604__;
  assign new_new_n4094__ = ~new_new_n634__ & ~new_new_n717__;
  assign new_new_n4095__ = new_new_n4093__ & new_new_n4094__;
  assign new_new_n4096__ = ~new_new_n1064__ & new_new_n1423__;
  assign new_new_n4097__ = new_new_n4095__ & new_new_n4096__;
  assign new_new_n4098__ = new_new_n1331__ & new_new_n2265__;
  assign new_new_n4099__ = new_new_n3793__ & new_new_n4092__;
  assign new_new_n4100__ = new_new_n4098__ & new_new_n4099__;
  assign new_new_n4101__ = new_new_n1384__ & new_new_n4097__;
  assign new_new_n4102__ = new_new_n4090__ & new_new_n4091__;
  assign new_new_n4103__ = new_new_n4101__ & new_new_n4102__;
  assign new_new_n4104__ = new_new_n3396__ & new_new_n4100__;
  assign new_new_n4105__ = new_new_n4103__ & new_new_n4104__;
  assign new_new_n4106__ = new_new_n2704__ & new_new_n2830__;
  assign new_new_n4107__ = new_new_n4105__ & new_new_n4106__;
  assign new_new_n4108__ = ~new_new_n302__ & ~new_new_n1217__;
  assign new_new_n4109__ = ~new_new_n351__ & ~new_new_n480__;
  assign new_new_n4110__ = ~new_new_n826__ & ~new_new_n995__;
  assign new_new_n4111__ = new_new_n4109__ & new_new_n4110__;
  assign new_new_n4112__ = ~new_new_n566__ & new_new_n1284__;
  assign new_new_n4113__ = new_new_n1511__ & new_new_n4112__;
  assign new_new_n4114__ = new_new_n233__ & new_new_n4111__;
  assign new_new_n4115__ = new_new_n387__ & new_new_n1078__;
  assign new_new_n4116__ = new_new_n1097__ & new_new_n1473__;
  assign new_new_n4117__ = ~new_new_n2403__ & new_new_n4108__;
  assign new_new_n4118__ = new_new_n4116__ & new_new_n4117__;
  assign new_new_n4119__ = new_new_n4114__ & new_new_n4115__;
  assign new_new_n4120__ = new_new_n4113__ & new_new_n4119__;
  assign new_new_n4121__ = new_new_n927__ & new_new_n4118__;
  assign new_new_n4122__ = new_new_n4120__ & new_new_n4121__;
  assign new_new_n4123__ = new_new_n4072__ & new_new_n4122__;
  assign new_new_n4124__ = new_new_n4089__ & new_new_n4123__;
  assign new_new_n4125__ = new_new_n4107__ & new_new_n4124__;
  assign new_new_n4126__ = new_new_n4021__ & ~new_new_n4125__;
  assign new_new_n4127__ = new_new_n3824__ & ~new_new_n4021__;
  assign new_new_n4128__ = ~new_new_n3824__ & new_new_n4021__;
  assign new_new_n4129__ = ~new_new_n4127__ & ~new_new_n4128__;
  assign new_new_n4130__ = ~new_new_n4126__ & ~new_new_n4129__;
  assign new_new_n4131__ = new_new_n4059__ & new_new_n4130__;
  assign new_new_n4132__ = ~new_new_n4021__ & ~new_new_n4059__;
  assign new_new_n4133__ = ~new_new_n3824__ & ~new_new_n4132__;
  assign new_new_n4134__ = ~new_new_n4060__ & ~new_new_n4125__;
  assign new_new_n4135__ = ~new_new_n4133__ & new_new_n4134__;
  assign new_new_n4136__ = ~new_new_n4061__ & ~new_new_n4131__;
  assign new_new_n4137__ = ~new_new_n4135__ & new_new_n4136__;
  assign new_new_n4138__ = new_new_n3892__ & ~new_new_n4137__;
  assign new_new_n4139__ = new_new_n691__ & new_new_n3742__;
  assign new_new_n4140__ = ~new_new_n583__ & ~new_new_n4139__;
  assign new_new_n4141__ = ~new_new_n3744__ & ~new_new_n4140__;
  assign new_new_n4142__ = ~new_new_n3768__ & ~new_new_n4141__;
  assign new_new_n4143__ = new_new_n3768__ & new_new_n4141__;
  assign new_new_n4144__ = ~new_new_n4142__ & ~new_new_n4143__;
  assign new_new_n4145__ = pi31 & new_new_n4144__;
  assign new_new_n4146__ = new_new_n125__ & ~new_new_n4145__;
  assign new_new_n4147__ = pi31 & ~new_new_n71__;
  assign new_new_n4148__ = ~pi29 & ~pi31;
  assign new_new_n4149__ = ~new_new_n4147__ & ~new_new_n4148__;
  assign new_new_n4150__ = ~new_new_n583__ & new_new_n4149__;
  assign new_new_n4151__ = pi31 & ~new_new_n691__;
  assign new_new_n4152__ = pi29 & ~new_new_n4151__;
  assign new_new_n4153__ = pi30 & ~new_new_n4152__;
  assign new_new_n4154__ = ~new_new_n4144__ & new_new_n4153__;
  assign new_new_n4155__ = ~new_new_n4150__ & ~new_new_n4154__;
  assign new_new_n4156__ = ~new_new_n4146__ & new_new_n4155__;
  assign new_new_n4157__ = ~new_new_n3824__ & new_new_n4132__;
  assign new_new_n4158__ = new_new_n3824__ & ~new_new_n4132__;
  assign new_new_n4159__ = ~new_new_n4157__ & ~new_new_n4158__;
  assign new_new_n4160__ = ~new_new_n4125__ & ~new_new_n4159__;
  assign new_new_n4161__ = new_new_n4021__ & ~new_new_n4059__;
  assign new_new_n4162__ = new_new_n4125__ & ~new_new_n4129__;
  assign new_new_n4163__ = ~new_new_n4161__ & new_new_n4162__;
  assign new_new_n4164__ = ~new_new_n3892__ & ~new_new_n4163__;
  assign new_new_n4165__ = ~new_new_n4160__ & new_new_n4164__;
  assign new_new_n4166__ = new_new_n4156__ & ~new_new_n4165__;
  assign new_new_n4167__ = ~new_new_n4138__ & ~new_new_n4166__;
  assign new_new_n4168__ = new_new_n3768__ & ~new_new_n4140__;
  assign new_new_n4169__ = ~new_new_n3769__ & ~new_new_n4168__;
  assign new_new_n4170__ = new_new_n466__ & ~new_new_n4169__;
  assign new_new_n4171__ = ~new_new_n466__ & new_new_n4169__;
  assign new_new_n4172__ = ~new_new_n4170__ & ~new_new_n4171__;
  assign new_new_n4173__ = new_new_n125__ & ~new_new_n4172__;
  assign new_new_n4174__ = pi30 & ~new_new_n583__;
  assign new_new_n4175__ = new_new_n3768__ & ~new_new_n4174__;
  assign new_new_n4176__ = pi31 & ~new_new_n4175__;
  assign new_new_n4177__ = ~new_new_n4173__ & new_new_n4176__;
  assign new_new_n4178__ = ~new_new_n4167__ & ~new_new_n4177__;
  assign new_new_n4179__ = new_new_n3888__ & new_new_n4178__;
  assign new_new_n4180__ = ~new_new_n3892__ & new_new_n4156__;
  assign new_new_n4181__ = ~new_new_n4021__ & new_new_n4125__;
  assign new_new_n4182__ = new_new_n4180__ & new_new_n4181__;
  assign new_new_n4183__ = new_new_n3892__ & ~new_new_n4156__;
  assign new_new_n4184__ = new_new_n4059__ & new_new_n4183__;
  assign new_new_n4185__ = new_new_n4021__ & new_new_n4180__;
  assign new_new_n4186__ = ~new_new_n4184__ & ~new_new_n4185__;
  assign new_new_n4187__ = ~new_new_n4125__ & ~new_new_n4186__;
  assign new_new_n4188__ = new_new_n4161__ & new_new_n4183__;
  assign new_new_n4189__ = ~new_new_n4182__ & ~new_new_n4188__;
  assign new_new_n4190__ = ~new_new_n4187__ & new_new_n4189__;
  assign new_new_n4191__ = new_new_n3824__ & ~new_new_n4190__;
  assign new_new_n4192__ = ~new_new_n4180__ & ~new_new_n4183__;
  assign new_new_n4193__ = ~new_new_n4125__ & new_new_n4132__;
  assign new_new_n4194__ = new_new_n4021__ & new_new_n4125__;
  assign new_new_n4195__ = new_new_n4059__ & new_new_n4194__;
  assign new_new_n4196__ = ~new_new_n4193__ & ~new_new_n4195__;
  assign new_new_n4197__ = ~new_new_n3824__ & new_new_n4196__;
  assign new_new_n4198__ = new_new_n3824__ & ~new_new_n4196__;
  assign new_new_n4199__ = new_new_n4192__ & ~new_new_n4197__;
  assign new_new_n4200__ = ~new_new_n4198__ & new_new_n4199__;
  assign new_new_n4201__ = new_new_n4125__ & new_new_n4128__;
  assign new_new_n4202__ = new_new_n4059__ & new_new_n4201__;
  assign new_new_n4203__ = ~new_new_n4127__ & ~new_new_n4193__;
  assign new_new_n4204__ = ~new_new_n4060__ & ~new_new_n4203__;
  assign new_new_n4205__ = ~new_new_n4192__ & ~new_new_n4202__;
  assign new_new_n4206__ = ~new_new_n4204__ & new_new_n4205__;
  assign new_new_n4207__ = ~new_new_n4200__ & ~new_new_n4206__;
  assign new_new_n4208__ = ~new_new_n4191__ & ~new_new_n4207__;
  assign new_new_n4209__ = ~pi26 & ~pi27;
  assign new_new_n4210__ = pi28 & ~new_new_n4209__;
  assign new_new_n4211__ = ~pi28 & ~new_new_n3889__;
  assign new_new_n4212__ = ~new_new_n4210__ & ~new_new_n4211__;
  assign new_new_n4213__ = ~new_new_n691__ & new_new_n4212__;
  assign new_new_n4214__ = ~new_new_n3889__ & ~new_new_n4209__;
  assign new_new_n4215__ = ~new_new_n220__ & ~new_new_n236__;
  assign new_new_n4216__ = new_new_n583__ & new_new_n4215__;
  assign new_new_n4217__ = new_new_n4214__ & ~new_new_n4216__;
  assign new_new_n4218__ = new_new_n3742__ & new_new_n4217__;
  assign new_new_n4219__ = ~new_new_n4213__ & ~new_new_n4218__;
  assign new_new_n4220__ = ~pi29 & ~new_new_n4219__;
  assign new_new_n4221__ = ~pi28 & new_new_n4209__;
  assign new_new_n4222__ = ~new_new_n910__ & new_new_n4221__;
  assign new_new_n4223__ = pi29 & ~new_new_n4222__;
  assign new_new_n4224__ = new_new_n66__ & ~new_new_n910__;
  assign new_new_n4225__ = ~new_new_n4223__ & ~new_new_n4224__;
  assign new_new_n4226__ = new_new_n4219__ & ~new_new_n4225__;
  assign new_new_n4227__ = ~new_new_n4220__ & ~new_new_n4226__;
  assign new_new_n4228__ = ~new_new_n835__ & ~new_new_n1033__;
  assign new_new_n4229__ = ~new_new_n631__ & new_new_n1332__;
  assign new_new_n4230__ = ~new_new_n259__ & ~new_new_n321__;
  assign new_new_n4231__ = ~new_new_n996__ & ~new_new_n1081__;
  assign new_new_n4232__ = ~new_new_n921__ & ~new_new_n1070__;
  assign new_new_n4233__ = ~new_new_n306__ & ~new_new_n723__;
  assign new_new_n4234__ = new_new_n167__ & new_new_n347__;
  assign new_new_n4235__ = ~new_new_n566__ & new_new_n3484__;
  assign new_new_n4236__ = ~new_new_n380__ & ~new_new_n933__;
  assign new_new_n4237__ = ~new_new_n150__ & new_new_n3806__;
  assign new_new_n4238__ = new_new_n4236__ & new_new_n4237__;
  assign new_new_n4239__ = new_new_n2701__ & new_new_n4238__;
  assign new_new_n4240__ = new_new_n3279__ & new_new_n4239__;
  assign new_new_n4241__ = ~new_new_n604__ & ~new_new_n1515__;
  assign new_new_n4242__ = ~new_new_n329__ & new_new_n4241__;
  assign new_new_n4243__ = ~new_new_n382__ & ~new_new_n871__;
  assign new_new_n4244__ = ~new_new_n993__ & new_new_n4243__;
  assign new_new_n4245__ = new_new_n722__ & new_new_n4242__;
  assign new_new_n4246__ = new_new_n4233__ & new_new_n4245__;
  assign new_new_n4247__ = new_new_n2791__ & new_new_n4244__;
  assign new_new_n4248__ = new_new_n3261__ & new_new_n4235__;
  assign new_new_n4249__ = new_new_n4247__ & new_new_n4248__;
  assign new_new_n4250__ = new_new_n4234__ & new_new_n4246__;
  assign new_new_n4251__ = new_new_n4249__ & new_new_n4250__;
  assign new_new_n4252__ = new_new_n4240__ & new_new_n4251__;
  assign new_new_n4253__ = ~new_new_n312__ & ~new_new_n637__;
  assign new_new_n4254__ = ~new_new_n242__ & ~new_new_n250__;
  assign new_new_n4255__ = ~new_new_n327__ & ~new_new_n1291__;
  assign new_new_n4256__ = new_new_n4254__ & new_new_n4255__;
  assign new_new_n4257__ = ~new_new_n202__ & new_new_n4253__;
  assign new_new_n4258__ = new_new_n4256__ & new_new_n4257__;
  assign new_new_n4259__ = new_new_n2168__ & new_new_n4258__;
  assign new_new_n4260__ = ~new_new_n717__ & ~new_new_n1109__;
  assign new_new_n4261__ = ~new_new_n1113__ & ~new_new_n2170__;
  assign new_new_n4262__ = new_new_n4260__ & new_new_n4261__;
  assign new_new_n4263__ = ~new_new_n274__ & ~new_new_n1166__;
  assign new_new_n4264__ = new_new_n1284__ & new_new_n4231__;
  assign new_new_n4265__ = new_new_n4263__ & new_new_n4264__;
  assign new_new_n4266__ = new_new_n1145__ & new_new_n4262__;
  assign new_new_n4267__ = new_new_n4228__ & new_new_n4229__;
  assign new_new_n4268__ = new_new_n4230__ & new_new_n4232__;
  assign new_new_n4269__ = new_new_n4267__ & new_new_n4268__;
  assign new_new_n4270__ = new_new_n4265__ & new_new_n4266__;
  assign new_new_n4271__ = new_new_n3317__ & new_new_n4270__;
  assign new_new_n4272__ = new_new_n4259__ & new_new_n4269__;
  assign new_new_n4273__ = new_new_n4271__ & new_new_n4272__;
  assign new_new_n4274__ = new_new_n1676__ & new_new_n4273__;
  assign new_new_n4275__ = new_new_n3413__ & new_new_n4274__;
  assign new_new_n4276__ = new_new_n4252__ & new_new_n4275__;
  assign new_new_n4277__ = new_new_n71__ & new_new_n3618__;
  assign new_new_n4278__ = ~new_new_n1061__ & new_new_n1325__;
  assign new_new_n4279__ = ~new_new_n3552__ & new_new_n4278__;
  assign new_new_n4280__ = new_new_n1061__ & new_new_n3618__;
  assign new_new_n4281__ = new_new_n1061__ & new_new_n1325__;
  assign new_new_n4282__ = ~new_new_n3618__ & ~new_new_n4281__;
  assign new_new_n4283__ = ~new_new_n4280__ & ~new_new_n4282__;
  assign new_new_n4284__ = new_new_n3552__ & new_new_n4283__;
  assign new_new_n4285__ = ~new_new_n4279__ & ~new_new_n4284__;
  assign new_new_n4286__ = ~new_new_n161__ & ~new_new_n4285__;
  assign new_new_n4287__ = new_new_n1061__ & ~new_new_n3552__;
  assign new_new_n4288__ = new_new_n3618__ & ~new_new_n4287__;
  assign new_new_n4289__ = new_new_n1061__ & ~new_new_n3618__;
  assign new_new_n4290__ = ~new_new_n4288__ & ~new_new_n4289__;
  assign new_new_n4291__ = ~new_new_n161__ & ~new_new_n4290__;
  assign new_new_n4292__ = ~new_new_n1325__ & ~new_new_n4291__;
  assign new_new_n4293__ = new_new_n4147__ & ~new_new_n4286__;
  assign new_new_n4294__ = ~new_new_n4292__ & new_new_n4293__;
  assign new_new_n4295__ = new_new_n161__ & new_new_n3618__;
  assign new_new_n4296__ = ~new_new_n161__ & new_new_n1061__;
  assign new_new_n4297__ = ~new_new_n71__ & ~new_new_n4295__;
  assign new_new_n4298__ = ~new_new_n4296__ & new_new_n4297__;
  assign new_new_n4299__ = ~pi31 & ~new_new_n4298__;
  assign new_new_n4300__ = ~new_new_n4277__ & ~new_new_n4299__;
  assign new_new_n4301__ = ~new_new_n4294__ & new_new_n4300__;
  assign new_new_n4302__ = new_new_n4276__ & ~new_new_n4301__;
  assign new_new_n4303__ = ~new_new_n240__ & ~new_new_n344__;
  assign new_new_n4304__ = ~new_new_n119__ & ~new_new_n164__;
  assign new_new_n4305__ = ~new_new_n327__ & new_new_n4304__;
  assign new_new_n4306__ = ~new_new_n721__ & ~new_new_n919__;
  assign new_new_n4307__ = ~new_new_n959__ & new_new_n1170__;
  assign new_new_n4308__ = ~new_new_n1506__ & new_new_n4307__;
  assign new_new_n4309__ = new_new_n4305__ & new_new_n4306__;
  assign new_new_n4310__ = new_new_n2455__ & new_new_n4309__;
  assign new_new_n4311__ = new_new_n3568__ & new_new_n4308__;
  assign new_new_n4312__ = new_new_n4303__ & new_new_n4311__;
  assign new_new_n4313__ = new_new_n4310__ & new_new_n4312__;
  assign new_new_n4314__ = ~new_new_n309__ & ~new_new_n383__;
  assign new_new_n4315__ = ~new_new_n95__ & ~new_new_n237__;
  assign new_new_n4316__ = new_new_n163__ & ~new_new_n4315__;
  assign new_new_n4317__ = ~new_new_n701__ & ~new_new_n875__;
  assign new_new_n4318__ = ~new_new_n143__ & new_new_n4317__;
  assign new_new_n4319__ = ~new_new_n192__ & ~new_new_n277__;
  assign new_new_n4320__ = ~new_new_n4316__ & new_new_n4319__;
  assign new_new_n4321__ = new_new_n4318__ & new_new_n4320__;
  assign new_new_n4322__ = ~new_new_n939__ & ~new_new_n2170__;
  assign new_new_n4323__ = ~new_new_n160__ & ~new_new_n284__;
  assign new_new_n4324__ = ~new_new_n1515__ & new_new_n4323__;
  assign new_new_n4325__ = new_new_n210__ & ~new_new_n258__;
  assign new_new_n4326__ = ~new_new_n675__ & ~new_new_n1073__;
  assign new_new_n4327__ = new_new_n1332__ & new_new_n1740__;
  assign new_new_n4328__ = new_new_n4314__ & new_new_n4327__;
  assign new_new_n4329__ = new_new_n4325__ & new_new_n4326__;
  assign new_new_n4330__ = new_new_n1065__ & new_new_n4324__;
  assign new_new_n4331__ = new_new_n1341__ & new_new_n1840__;
  assign new_new_n4332__ = new_new_n2335__ & new_new_n2427__;
  assign new_new_n4333__ = new_new_n4230__ & new_new_n4322__;
  assign new_new_n4334__ = new_new_n4332__ & new_new_n4333__;
  assign new_new_n4335__ = new_new_n4330__ & new_new_n4331__;
  assign new_new_n4336__ = new_new_n4328__ & new_new_n4329__;
  assign new_new_n4337__ = new_new_n3140__ & new_new_n4336__;
  assign new_new_n4338__ = new_new_n4334__ & new_new_n4335__;
  assign new_new_n4339__ = new_new_n4321__ & new_new_n4338__;
  assign new_new_n4340__ = new_new_n4337__ & new_new_n4339__;
  assign new_new_n4341__ = ~new_new_n809__ & new_new_n2653__;
  assign new_new_n4342__ = ~new_new_n963__ & ~new_new_n1162__;
  assign new_new_n4343__ = ~new_new_n476__ & ~new_new_n717__;
  assign new_new_n4344__ = ~new_new_n82__ & ~new_new_n509__;
  assign new_new_n4345__ = ~new_new_n724__ & new_new_n4344__;
  assign new_new_n4346__ = ~new_new_n306__ & ~new_new_n346__;
  assign new_new_n4347__ = ~new_new_n816__ & ~new_new_n874__;
  assign new_new_n4348__ = new_new_n2267__ & new_new_n4343__;
  assign new_new_n4349__ = new_new_n4347__ & new_new_n4348__;
  assign new_new_n4350__ = new_new_n4345__ & new_new_n4346__;
  assign new_new_n4351__ = new_new_n4349__ & new_new_n4350__;
  assign new_new_n4352__ = new_new_n1112__ & new_new_n4351__;
  assign new_new_n4353__ = new_new_n1569__ & new_new_n4352__;
  assign new_new_n4354__ = ~new_new_n101__ & ~new_new_n250__;
  assign new_new_n4355__ = ~new_new_n1003__ & new_new_n4354__;
  assign new_new_n4356__ = new_new_n1263__ & new_new_n1424__;
  assign new_new_n4357__ = new_new_n4342__ & new_new_n4356__;
  assign new_new_n4358__ = ~new_new_n254__ & new_new_n4355__;
  assign new_new_n4359__ = new_new_n3385__ & new_new_n3956__;
  assign new_new_n4360__ = new_new_n4358__ & new_new_n4359__;
  assign new_new_n4361__ = new_new_n4341__ & new_new_n4357__;
  assign new_new_n4362__ = new_new_n4360__ & new_new_n4361__;
  assign new_new_n4363__ = new_new_n1999__ & new_new_n4362__;
  assign new_new_n4364__ = new_new_n4353__ & new_new_n4363__;
  assign new_new_n4365__ = ~new_new_n488__ & ~new_new_n811__;
  assign new_new_n4366__ = ~new_new_n251__ & ~new_new_n783__;
  assign new_new_n4367__ = ~new_new_n843__ & new_new_n4366__;
  assign new_new_n4368__ = ~new_new_n255__ & ~new_new_n266__;
  assign new_new_n4369__ = ~new_new_n894__ & new_new_n4368__;
  assign new_new_n4370__ = new_new_n1679__ & new_new_n4367__;
  assign new_new_n4371__ = new_new_n4108__ & new_new_n4365__;
  assign new_new_n4372__ = new_new_n4370__ & new_new_n4371__;
  assign new_new_n4373__ = new_new_n4369__ & new_new_n4372__;
  assign new_new_n4374__ = ~new_new_n603__ & ~new_new_n785__;
  assign new_new_n4375__ = ~new_new_n1151__ & new_new_n4374__;
  assign new_new_n4376__ = new_new_n1449__ & new_new_n3486__;
  assign new_new_n4377__ = new_new_n4375__ & new_new_n4376__;
  assign new_new_n4378__ = new_new_n775__ & ~new_new_n1486__;
  assign new_new_n4379__ = new_new_n3365__ & new_new_n4378__;
  assign new_new_n4380__ = new_new_n4377__ & new_new_n4379__;
  assign new_new_n4381__ = new_new_n3631__ & new_new_n4380__;
  assign new_new_n4382__ = new_new_n4373__ & new_new_n4381__;
  assign new_new_n4383__ = new_new_n4313__ & new_new_n4382__;
  assign new_new_n4384__ = new_new_n4340__ & new_new_n4364__;
  assign new_new_n4385__ = new_new_n4383__ & new_new_n4384__;
  assign new_new_n4386__ = ~pi20 & ~new_new_n4385__;
  assign new_new_n4387__ = pi20 & new_new_n4385__;
  assign new_new_n4388__ = new_new_n1230__ & new_new_n2850__;
  assign new_new_n4389__ = ~new_new_n700__ & ~new_new_n828__;
  assign new_new_n4390__ = ~new_new_n232__ & ~new_new_n1113__;
  assign new_new_n4391__ = ~new_new_n597__ & ~new_new_n842__;
  assign new_new_n4392__ = ~new_new_n519__ & new_new_n4391__;
  assign new_new_n4393__ = ~new_new_n226__ & ~new_new_n335__;
  assign new_new_n4394__ = new_new_n180__ & ~new_new_n1880__;
  assign new_new_n4395__ = ~new_new_n92__ & ~new_new_n811__;
  assign new_new_n4396__ = ~new_new_n942__ & new_new_n4395__;
  assign new_new_n4397__ = new_new_n2822__ & ~new_new_n4394__;
  assign new_new_n4398__ = new_new_n4396__ & new_new_n4397__;
  assign new_new_n4399__ = ~new_new_n586__ & ~new_new_n637__;
  assign new_new_n4400__ = ~new_new_n723__ & ~new_new_n1109__;
  assign new_new_n4401__ = new_new_n4399__ & new_new_n4400__;
  assign new_new_n4402__ = ~new_new_n380__ & new_new_n2160__;
  assign new_new_n4403__ = new_new_n4401__ & new_new_n4402__;
  assign new_new_n4404__ = new_new_n167__ & new_new_n387__;
  assign new_new_n4405__ = new_new_n1032__ & new_new_n3012__;
  assign new_new_n4406__ = new_new_n3027__ & new_new_n3912__;
  assign new_new_n4407__ = new_new_n4393__ & new_new_n4406__;
  assign new_new_n4408__ = new_new_n4404__ & new_new_n4405__;
  assign new_new_n4409__ = new_new_n440__ & new_new_n4403__;
  assign new_new_n4410__ = new_new_n4398__ & new_new_n4409__;
  assign new_new_n4411__ = new_new_n4407__ & new_new_n4408__;
  assign new_new_n4412__ = new_new_n4410__ & new_new_n4411__;
  assign new_new_n4413__ = ~new_new_n510__ & ~new_new_n1003__;
  assign new_new_n4414__ = ~new_new_n196__ & ~new_new_n603__;
  assign new_new_n4415__ = ~new_new_n101__ & ~new_new_n634__;
  assign new_new_n4416__ = ~new_new_n656__ & ~new_new_n2170__;
  assign new_new_n4417__ = new_new_n4415__ & new_new_n4416__;
  assign new_new_n4418__ = ~new_new_n350__ & ~new_new_n835__;
  assign new_new_n4419__ = new_new_n3392__ & new_new_n3957__;
  assign new_new_n4420__ = new_new_n4414__ & new_new_n4419__;
  assign new_new_n4421__ = new_new_n4417__ & new_new_n4418__;
  assign new_new_n4422__ = new_new_n4413__ & new_new_n4421__;
  assign new_new_n4423__ = new_new_n4420__ & new_new_n4422__;
  assign new_new_n4424__ = ~new_new_n213__ & ~new_new_n282__;
  assign new_new_n4425__ = ~new_new_n379__ & new_new_n4424__;
  assign new_new_n4426__ = ~new_new_n198__ & ~new_new_n266__;
  assign new_new_n4427__ = new_new_n1177__ & new_new_n3179__;
  assign new_new_n4428__ = new_new_n4426__ & new_new_n4427__;
  assign new_new_n4429__ = new_new_n354__ & new_new_n4425__;
  assign new_new_n4430__ = new_new_n1340__ & new_new_n1481__;
  assign new_new_n4431__ = new_new_n2334__ & new_new_n4430__;
  assign new_new_n4432__ = new_new_n4428__ & new_new_n4429__;
  assign new_new_n4433__ = new_new_n2764__ & new_new_n4432__;
  assign new_new_n4434__ = new_new_n4431__ & new_new_n4433__;
  assign new_new_n4435__ = new_new_n2554__ & new_new_n4423__;
  assign new_new_n4436__ = new_new_n4434__ & new_new_n4435__;
  assign new_new_n4437__ = ~new_new_n82__ & ~new_new_n246__;
  assign new_new_n4438__ = ~new_new_n302__ & new_new_n4437__;
  assign new_new_n4439__ = ~new_new_n507__ & new_new_n3688__;
  assign new_new_n4440__ = new_new_n4438__ & new_new_n4439__;
  assign new_new_n4441__ = ~new_new_n218__ & ~new_new_n344__;
  assign new_new_n4442__ = new_new_n4389__ & new_new_n4390__;
  assign new_new_n4443__ = new_new_n4441__ & new_new_n4442__;
  assign new_new_n4444__ = new_new_n2028__ & new_new_n4440__;
  assign new_new_n4445__ = new_new_n3640__ & new_new_n4388__;
  assign new_new_n4446__ = new_new_n4392__ & new_new_n4445__;
  assign new_new_n4447__ = new_new_n4443__ & new_new_n4444__;
  assign new_new_n4448__ = new_new_n1879__ & new_new_n4447__;
  assign new_new_n4449__ = new_new_n1916__ & new_new_n4446__;
  assign new_new_n4450__ = new_new_n4448__ & new_new_n4449__;
  assign new_new_n4451__ = new_new_n4412__ & new_new_n4450__;
  assign new_new_n4452__ = new_new_n4436__ & new_new_n4451__;
  assign new_new_n4453__ = ~new_new_n4387__ & ~new_new_n4452__;
  assign new_new_n4454__ = ~new_new_n4386__ & ~new_new_n4453__;
  assign new_new_n4455__ = new_new_n4302__ & new_new_n4454__;
  assign new_new_n4456__ = ~new_new_n4276__ & new_new_n4301__;
  assign new_new_n4457__ = ~new_new_n4454__ & new_new_n4456__;
  assign new_new_n4458__ = ~new_new_n1151__ & ~new_new_n1515__;
  assign new_new_n4459__ = ~new_new_n384__ & ~new_new_n772__;
  assign new_new_n4460__ = ~new_new_n313__ & ~new_new_n1081__;
  assign new_new_n4461__ = ~new_new_n884__ & new_new_n4460__;
  assign new_new_n4462__ = new_new_n4459__ & new_new_n4461__;
  assign new_new_n4463__ = new_new_n4458__ & new_new_n4462__;
  assign new_new_n4464__ = new_new_n1255__ & new_new_n4463__;
  assign new_new_n4465__ = ~new_new_n92__ & ~new_new_n778__;
  assign new_new_n4466__ = ~new_new_n511__ & ~new_new_n637__;
  assign new_new_n4467__ = ~new_new_n933__ & ~new_new_n1398__;
  assign new_new_n4468__ = new_new_n4466__ & new_new_n4467__;
  assign new_new_n4469__ = ~new_new_n226__ & ~new_new_n719__;
  assign new_new_n4470__ = ~new_new_n2645__ & new_new_n3582__;
  assign new_new_n4471__ = new_new_n4465__ & new_new_n4470__;
  assign new_new_n4472__ = new_new_n4468__ & new_new_n4469__;
  assign new_new_n4473__ = new_new_n3282__ & new_new_n3686__;
  assign new_new_n4474__ = new_new_n4472__ & new_new_n4473__;
  assign new_new_n4475__ = new_new_n1160__ & new_new_n4471__;
  assign new_new_n4476__ = new_new_n4474__ & new_new_n4475__;
  assign new_new_n4477__ = ~new_new_n148__ & ~new_new_n894__;
  assign new_new_n4478__ = ~new_new_n300__ & ~new_new_n344__;
  assign new_new_n4479__ = ~new_new_n91__ & ~new_new_n163__;
  assign new_new_n4480__ = ~new_new_n202__ & ~new_new_n718__;
  assign new_new_n4481__ = ~new_new_n878__ & new_new_n4480__;
  assign new_new_n4482__ = ~new_new_n4479__ & ~new_new_n4481__;
  assign new_new_n4483__ = ~new_new_n82__ & ~new_new_n729__;
  assign new_new_n4484__ = ~new_new_n189__ & new_new_n4483__;
  assign new_new_n4485__ = new_new_n3439__ & new_new_n4484__;
  assign new_new_n4486__ = ~new_new_n4482__ & new_new_n4485__;
  assign new_new_n4487__ = ~new_new_n213__ & ~new_new_n996__;
  assign new_new_n4488__ = ~new_new_n155__ & new_new_n4487__;
  assign new_new_n4489__ = ~new_new_n939__ & new_new_n3836__;
  assign new_new_n4490__ = new_new_n4488__ & new_new_n4489__;
  assign new_new_n4491__ = new_new_n1920__ & new_new_n4477__;
  assign new_new_n4492__ = new_new_n4490__ & new_new_n4491__;
  assign new_new_n4493__ = new_new_n4478__ & new_new_n4492__;
  assign new_new_n4494__ = new_new_n3192__ & new_new_n4493__;
  assign new_new_n4495__ = new_new_n4464__ & new_new_n4476__;
  assign new_new_n4496__ = new_new_n4486__ & new_new_n4495__;
  assign new_new_n4497__ = new_new_n4494__ & new_new_n4496__;
  assign new_new_n4498__ = ~new_new_n482__ & ~new_new_n1210__;
  assign new_new_n4499__ = ~new_new_n380__ & new_new_n4498__;
  assign new_new_n4500__ = ~new_new_n1009__ & ~new_new_n1035__;
  assign new_new_n4501__ = new_new_n4499__ & new_new_n4500__;
  assign new_new_n4502__ = ~new_new_n935__ & new_new_n4501__;
  assign new_new_n4503__ = ~new_new_n1539__ & new_new_n4502__;
  assign new_new_n4504__ = ~new_new_n350__ & ~new_new_n676__;
  assign new_new_n4505__ = ~new_new_n316__ & ~new_new_n508__;
  assign new_new_n4506__ = ~new_new_n229__ & ~new_new_n242__;
  assign new_new_n4507__ = ~new_new_n1007__ & new_new_n4506__;
  assign new_new_n4508__ = ~new_new_n483__ & ~new_new_n1073__;
  assign new_new_n4509__ = new_new_n4507__ & new_new_n4508__;
  assign new_new_n4510__ = ~new_new_n208__ & ~new_new_n379__;
  assign new_new_n4511__ = ~new_new_n950__ & new_new_n4510__;
  assign new_new_n4512__ = new_new_n121__ & new_new_n1597__;
  assign new_new_n4513__ = new_new_n2116__ & new_new_n3968__;
  assign new_new_n4514__ = new_new_n4512__ & new_new_n4513__;
  assign new_new_n4515__ = new_new_n744__ & new_new_n4511__;
  assign new_new_n4516__ = new_new_n1905__ & new_new_n4515__;
  assign new_new_n4517__ = new_new_n2478__ & new_new_n4514__;
  assign new_new_n4518__ = new_new_n4504__ & new_new_n4505__;
  assign new_new_n4519__ = new_new_n4509__ & new_new_n4518__;
  assign new_new_n4520__ = new_new_n4516__ & new_new_n4517__;
  assign new_new_n4521__ = new_new_n4519__ & new_new_n4520__;
  assign new_new_n4522__ = new_new_n2514__ & new_new_n4503__;
  assign new_new_n4523__ = new_new_n4521__ & new_new_n4522__;
  assign new_new_n4524__ = new_new_n4497__ & new_new_n4523__;
  assign new_new_n4525__ = ~new_new_n4457__ & ~new_new_n4524__;
  assign new_new_n4526__ = ~new_new_n4455__ & ~new_new_n4525__;
  assign new_new_n4527__ = new_new_n71__ & new_new_n1207__;
  assign new_new_n4528__ = ~new_new_n1061__ & new_new_n3620__;
  assign new_new_n4529__ = ~new_new_n3552__ & new_new_n4528__;
  assign new_new_n4530__ = new_new_n1208__ & ~new_new_n3618__;
  assign new_new_n4531__ = ~new_new_n4529__ & ~new_new_n4530__;
  assign new_new_n4532__ = ~new_new_n1325__ & ~new_new_n4531__;
  assign new_new_n4533__ = new_new_n1208__ & ~new_new_n3552__;
  assign new_new_n4534__ = ~new_new_n4528__ & ~new_new_n4533__;
  assign new_new_n4535__ = ~new_new_n3618__ & ~new_new_n4534__;
  assign new_new_n4536__ = ~new_new_n868__ & ~new_new_n3618__;
  assign new_new_n4537__ = ~new_new_n1208__ & ~new_new_n3620__;
  assign new_new_n4538__ = new_new_n868__ & ~new_new_n4281__;
  assign new_new_n4539__ = ~new_new_n4536__ & new_new_n4537__;
  assign new_new_n4540__ = ~new_new_n4538__ & new_new_n4539__;
  assign new_new_n4541__ = new_new_n3552__ & new_new_n4540__;
  assign new_new_n4542__ = ~new_new_n1207__ & ~new_new_n3618__;
  assign new_new_n4543__ = new_new_n1061__ & ~new_new_n4542__;
  assign new_new_n4544__ = new_new_n4537__ & new_new_n4543__;
  assign new_new_n4545__ = ~new_new_n4541__ & ~new_new_n4544__;
  assign new_new_n4546__ = ~new_new_n4532__ & new_new_n4545__;
  assign new_new_n4547__ = ~new_new_n4535__ & new_new_n4546__;
  assign new_new_n4548__ = ~new_new_n1061__ & ~new_new_n1207__;
  assign new_new_n4549__ = ~new_new_n868__ & new_new_n4548__;
  assign new_new_n4550__ = new_new_n4547__ & ~new_new_n4549__;
  assign new_new_n4551__ = new_new_n765__ & new_new_n4550__;
  assign new_new_n4552__ = new_new_n161__ & new_new_n1061__;
  assign new_new_n4553__ = ~new_new_n4551__ & ~new_new_n4552__;
  assign new_new_n4554__ = pi31 & ~new_new_n4553__;
  assign new_new_n4555__ = new_new_n161__ & new_new_n1207__;
  assign new_new_n4556__ = ~new_new_n161__ & new_new_n868__;
  assign new_new_n4557__ = ~new_new_n71__ & ~new_new_n4555__;
  assign new_new_n4558__ = ~new_new_n4556__ & new_new_n4557__;
  assign new_new_n4559__ = ~pi31 & ~new_new_n4558__;
  assign new_new_n4560__ = ~new_new_n4527__ & ~new_new_n4559__;
  assign new_new_n4561__ = ~new_new_n4554__ & new_new_n4560__;
  assign new_new_n4562__ = ~new_new_n4526__ & ~new_new_n4561__;
  assign new_new_n4563__ = new_new_n4526__ & new_new_n4561__;
  assign new_new_n4564__ = ~new_new_n101__ & ~new_new_n776__;
  assign new_new_n4565__ = ~new_new_n607__ & ~new_new_n631__;
  assign new_new_n4566__ = ~new_new_n127__ & ~new_new_n480__;
  assign new_new_n4567__ = ~new_new_n246__ & ~new_new_n271__;
  assign new_new_n4568__ = ~new_new_n509__ & ~new_new_n1033__;
  assign new_new_n4569__ = new_new_n4567__ & new_new_n4568__;
  assign new_new_n4570__ = new_new_n1994__ & new_new_n4566__;
  assign new_new_n4571__ = new_new_n3792__ & new_new_n4569__;
  assign new_new_n4572__ = new_new_n4570__ & new_new_n4571__;
  assign new_new_n4573__ = new_new_n592__ & ~new_new_n945__;
  assign new_new_n4574__ = new_new_n78__ & new_new_n371__;
  assign new_new_n4575__ = ~new_new_n374__ & ~new_new_n637__;
  assign new_new_n4576__ = new_new_n2962__ & new_new_n4575__;
  assign new_new_n4577__ = ~new_new_n624__ & ~new_new_n772__;
  assign new_new_n4578__ = ~new_new_n213__ & ~new_new_n253__;
  assign new_new_n4579__ = ~new_new_n315__ & ~new_new_n510__;
  assign new_new_n4580__ = ~new_new_n729__ & ~new_new_n2170__;
  assign new_new_n4581__ = ~new_new_n4574__ & new_new_n4580__;
  assign new_new_n4582__ = new_new_n4578__ & new_new_n4579__;
  assign new_new_n4583__ = ~new_new_n183__ & ~new_new_n566__;
  assign new_new_n4584__ = ~new_new_n894__ & new_new_n1373__;
  assign new_new_n4585__ = ~new_new_n1701__ & new_new_n4577__;
  assign new_new_n4586__ = new_new_n4584__ & new_new_n4585__;
  assign new_new_n4587__ = new_new_n4582__ & new_new_n4583__;
  assign new_new_n4588__ = new_new_n4581__ & new_new_n4587__;
  assign new_new_n4589__ = new_new_n771__ & new_new_n4586__;
  assign new_new_n4590__ = ~new_new_n1539__ & new_new_n2641__;
  assign new_new_n4591__ = new_new_n4573__ & new_new_n4576__;
  assign new_new_n4592__ = new_new_n4590__ & new_new_n4591__;
  assign new_new_n4593__ = new_new_n4588__ & new_new_n4589__;
  assign new_new_n4594__ = new_new_n4592__ & new_new_n4593__;
  assign new_new_n4595__ = ~new_new_n209__ & ~new_new_n260__;
  assign new_new_n4596__ = ~new_new_n143__ & new_new_n944__;
  assign new_new_n4597__ = ~new_new_n350__ & ~new_new_n732__;
  assign new_new_n4598__ = ~new_new_n717__ & ~new_new_n815__;
  assign new_new_n4599__ = new_new_n4597__ & new_new_n4598__;
  assign new_new_n4600__ = new_new_n4596__ & new_new_n4599__;
  assign new_new_n4601__ = ~new_new_n218__ & ~new_new_n508__;
  assign new_new_n4602__ = ~new_new_n846__ & ~new_new_n1094__;
  assign new_new_n4603__ = ~new_new_n1176__ & new_new_n4602__;
  assign new_new_n4604__ = ~new_new_n869__ & ~new_new_n1217__;
  assign new_new_n4605__ = new_new_n1368__ & new_new_n1639__;
  assign new_new_n4606__ = new_new_n4595__ & new_new_n4605__;
  assign new_new_n4607__ = new_new_n4603__ & new_new_n4604__;
  assign new_new_n4608__ = new_new_n3280__ & new_new_n4607__;
  assign new_new_n4609__ = new_new_n1627__ & new_new_n4606__;
  assign new_new_n4610__ = new_new_n2092__ & new_new_n4601__;
  assign new_new_n4611__ = new_new_n4609__ & new_new_n4610__;
  assign new_new_n4612__ = new_new_n957__ & new_new_n4608__;
  assign new_new_n4613__ = new_new_n4600__ & new_new_n4612__;
  assign new_new_n4614__ = new_new_n1928__ & new_new_n4611__;
  assign new_new_n4615__ = new_new_n3895__ & new_new_n4614__;
  assign new_new_n4616__ = new_new_n4594__ & new_new_n4613__;
  assign new_new_n4617__ = new_new_n4615__ & new_new_n4616__;
  assign new_new_n4618__ = ~new_new_n82__ & ~new_new_n267__;
  assign new_new_n4619__ = ~new_new_n302__ & new_new_n4618__;
  assign new_new_n4620__ = ~new_new_n332__ & ~new_new_n348__;
  assign new_new_n4621__ = ~new_new_n673__ & new_new_n3258__;
  assign new_new_n4622__ = new_new_n3804__ & new_new_n4621__;
  assign new_new_n4623__ = new_new_n4619__ & new_new_n4620__;
  assign new_new_n4624__ = new_new_n885__ & new_new_n941__;
  assign new_new_n4625__ = new_new_n984__ & new_new_n1885__;
  assign new_new_n4626__ = new_new_n4624__ & new_new_n4625__;
  assign new_new_n4627__ = new_new_n4622__ & new_new_n4623__;
  assign new_new_n4628__ = new_new_n4626__ & new_new_n4627__;
  assign new_new_n4629__ = ~new_new_n96__ & ~new_new_n207__;
  assign new_new_n4630__ = ~new_new_n698__ & ~new_new_n838__;
  assign new_new_n4631__ = ~new_new_n933__ & new_new_n4630__;
  assign new_new_n4632__ = ~new_new_n255__ & new_new_n4629__;
  assign new_new_n4633__ = new_new_n3128__ & new_new_n4314__;
  assign new_new_n4634__ = new_new_n4564__ & new_new_n4633__;
  assign new_new_n4635__ = new_new_n4631__ & new_new_n4632__;
  assign new_new_n4636__ = new_new_n2197__ & new_new_n2336__;
  assign new_new_n4637__ = new_new_n3284__ & new_new_n4636__;
  assign new_new_n4638__ = new_new_n4634__ & new_new_n4635__;
  assign new_new_n4639__ = new_new_n1883__ & new_new_n4565__;
  assign new_new_n4640__ = new_new_n4638__ & new_new_n4639__;
  assign new_new_n4641__ = new_new_n4572__ & new_new_n4637__;
  assign new_new_n4642__ = new_new_n4640__ & new_new_n4641__;
  assign new_new_n4643__ = new_new_n4628__ & new_new_n4642__;
  assign new_new_n4644__ = new_new_n4617__ & new_new_n4643__;
  assign new_new_n4645__ = new_new_n4524__ & new_new_n4644__;
  assign new_new_n4646__ = ~new_new_n4524__ & ~new_new_n4644__;
  assign new_new_n4647__ = ~pi23 & ~new_new_n4645__;
  assign new_new_n4648__ = ~new_new_n4646__ & ~new_new_n4647__;
  assign new_new_n4649__ = ~new_new_n4645__ & new_new_n4648__;
  assign new_new_n4650__ = pi23 & ~new_new_n4649__;
  assign new_new_n4651__ = ~new_new_n4646__ & new_new_n4647__;
  assign new_new_n4652__ = ~new_new_n4650__ & ~new_new_n4651__;
  assign new_new_n4653__ = ~new_new_n4563__ & ~new_new_n4652__;
  assign new_new_n4654__ = ~new_new_n4562__ & ~new_new_n4653__;
  assign new_new_n4655__ = new_new_n4227__ & ~new_new_n4654__;
  assign new_new_n4656__ = new_new_n765__ & ~new_new_n3720__;
  assign new_new_n4657__ = new_new_n161__ & ~new_new_n868__;
  assign new_new_n4658__ = ~new_new_n4656__ & ~new_new_n4657__;
  assign new_new_n4659__ = ~pi31 & ~new_new_n4658__;
  assign new_new_n4660__ = new_new_n3622__ & ~new_new_n3720__;
  assign new_new_n4661__ = ~new_new_n3622__ & new_new_n3720__;
  assign new_new_n4662__ = ~new_new_n4660__ & ~new_new_n4661__;
  assign new_new_n4663__ = new_new_n3622__ & ~new_new_n3662__;
  assign new_new_n4664__ = new_new_n765__ & ~new_new_n868__;
  assign new_new_n4665__ = ~new_new_n4663__ & new_new_n4664__;
  assign new_new_n4666__ = new_new_n4662__ & new_new_n4665__;
  assign new_new_n4667__ = ~new_new_n71__ & new_new_n4662__;
  assign new_new_n4668__ = new_new_n4556__ & ~new_new_n4667__;
  assign new_new_n4669__ = pi31 & ~new_new_n4555__;
  assign new_new_n4670__ = ~new_new_n4666__ & new_new_n4669__;
  assign new_new_n4671__ = ~new_new_n4668__ & new_new_n4670__;
  assign new_new_n4672__ = ~new_new_n4659__ & ~new_new_n4671__;
  assign new_new_n4673__ = new_new_n4019__ & ~new_new_n4672__;
  assign new_new_n4674__ = ~new_new_n4648__ & new_new_n4673__;
  assign new_new_n4675__ = ~new_new_n4655__ & new_new_n4674__;
  assign new_new_n4676__ = ~new_new_n4227__ & new_new_n4654__;
  assign new_new_n4677__ = ~new_new_n4019__ & new_new_n4672__;
  assign new_new_n4678__ = ~new_new_n4648__ & ~new_new_n4677__;
  assign new_new_n4679__ = ~new_new_n4673__ & ~new_new_n4678__;
  assign new_new_n4680__ = ~new_new_n4676__ & new_new_n4679__;
  assign new_new_n4681__ = new_new_n4648__ & new_new_n4677__;
  assign new_new_n4682__ = ~new_new_n4655__ & ~new_new_n4681__;
  assign new_new_n4683__ = new_new_n4680__ & ~new_new_n4682__;
  assign new_new_n4684__ = ~new_new_n4030__ & ~new_new_n4660__;
  assign new_new_n4685__ = new_new_n765__ & ~new_new_n4684__;
  assign new_new_n4686__ = ~new_new_n4033__ & ~new_new_n4685__;
  assign new_new_n4687__ = new_new_n910__ & ~new_new_n4686__;
  assign new_new_n4688__ = ~new_new_n3622__ & new_new_n4029__;
  assign new_new_n4689__ = ~new_new_n161__ & ~new_new_n4688__;
  assign new_new_n4690__ = ~new_new_n71__ & new_new_n868__;
  assign new_new_n4691__ = ~new_new_n4689__ & new_new_n4690__;
  assign new_new_n4692__ = ~new_new_n868__ & ~new_new_n910__;
  assign new_new_n4693__ = new_new_n3622__ & new_new_n4692__;
  assign new_new_n4694__ = ~new_new_n71__ & ~new_new_n4693__;
  assign new_new_n4695__ = ~new_new_n161__ & new_new_n3720__;
  assign new_new_n4696__ = ~new_new_n4694__ & new_new_n4695__;
  assign new_new_n4697__ = ~new_new_n4691__ & ~new_new_n4696__;
  assign new_new_n4698__ = ~new_new_n4687__ & new_new_n4697__;
  assign new_new_n4699__ = pi31 & ~new_new_n4698__;
  assign new_new_n4700__ = new_new_n161__ & ~new_new_n3720__;
  assign new_new_n4701__ = new_new_n765__ & ~new_new_n910__;
  assign new_new_n4702__ = ~pi31 & ~new_new_n4700__;
  assign new_new_n4703__ = ~new_new_n4701__ & new_new_n4702__;
  assign new_new_n4704__ = ~new_new_n4699__ & ~new_new_n4703__;
  assign new_new_n4705__ = new_new_n201__ & ~new_new_n333__;
  assign new_new_n4706__ = ~new_new_n250__ & ~new_new_n476__;
  assign new_new_n4707__ = ~new_new_n950__ & new_new_n4706__;
  assign new_new_n4708__ = ~new_new_n348__ & new_new_n3141__;
  assign new_new_n4709__ = new_new_n3179__ & new_new_n3391__;
  assign new_new_n4710__ = ~new_new_n4705__ & new_new_n4709__;
  assign new_new_n4711__ = new_new_n4707__ & new_new_n4708__;
  assign new_new_n4712__ = ~new_new_n1105__ & new_new_n1884__;
  assign new_new_n4713__ = new_new_n4711__ & new_new_n4712__;
  assign new_new_n4714__ = new_new_n4710__ & new_new_n4713__;
  assign new_new_n4715__ = new_new_n1498__ & new_new_n4714__;
  assign new_new_n4716__ = ~new_new_n591__ & ~new_new_n1081__;
  assign new_new_n4717__ = ~new_new_n329__ & new_new_n3702__;
  assign new_new_n4718__ = ~new_new_n1217__ & new_new_n4717__;
  assign new_new_n4719__ = new_new_n4716__ & new_new_n4718__;
  assign new_new_n4720__ = ~new_new_n308__ & ~new_new_n388__;
  assign new_new_n4721__ = ~new_new_n315__ & ~new_new_n379__;
  assign new_new_n4722__ = ~new_new_n637__ & ~new_new_n772__;
  assign new_new_n4723__ = new_new_n4721__ & new_new_n4722__;
  assign new_new_n4724__ = new_new_n4720__ & new_new_n4723__;
  assign new_new_n4725__ = new_new_n2469__ & new_new_n3138__;
  assign new_new_n4726__ = new_new_n4724__ & new_new_n4725__;
  assign new_new_n4727__ = ~new_new_n106__ & ~new_new_n632__;
  assign new_new_n4728__ = ~new_new_n246__ & ~new_new_n723__;
  assign new_new_n4729__ = ~new_new_n332__ & ~new_new_n783__;
  assign new_new_n4730__ = ~new_new_n76__ & ~new_new_n700__;
  assign new_new_n4731__ = ~new_new_n251__ & ~new_new_n890__;
  assign new_new_n4732__ = ~new_new_n183__ & ~new_new_n1162__;
  assign new_new_n4733__ = ~new_new_n438__ & ~new_new_n778__;
  assign new_new_n4734__ = ~new_new_n339__ & new_new_n4733__;
  assign new_new_n4735__ = new_new_n386__ & ~new_new_n588__;
  assign new_new_n4736__ = new_new_n3020__ & new_new_n4735__;
  assign new_new_n4737__ = new_new_n1645__ & new_new_n4734__;
  assign new_new_n4738__ = new_new_n2962__ & new_new_n3390__;
  assign new_new_n4739__ = new_new_n4732__ & new_new_n4738__;
  assign new_new_n4740__ = new_new_n4736__ & new_new_n4737__;
  assign new_new_n4741__ = new_new_n4739__ & new_new_n4740__;
  assign new_new_n4742__ = new_new_n2865__ & new_new_n4741__;
  assign new_new_n4743__ = ~new_new_n282__ & ~new_new_n676__;
  assign new_new_n4744__ = ~new_new_n597__ & ~new_new_n829__;
  assign new_new_n4745__ = ~new_new_n875__ & new_new_n4744__;
  assign new_new_n4746__ = ~new_new_n871__ & ~new_new_n878__;
  assign new_new_n4747__ = ~new_new_n1151__ & new_new_n2468__;
  assign new_new_n4748__ = new_new_n2576__ & ~new_new_n3566__;
  assign new_new_n4749__ = new_new_n4727__ & new_new_n4728__;
  assign new_new_n4750__ = new_new_n4730__ & new_new_n4731__;
  assign new_new_n4751__ = new_new_n4749__ & new_new_n4750__;
  assign new_new_n4752__ = new_new_n4747__ & new_new_n4748__;
  assign new_new_n4753__ = new_new_n4745__ & new_new_n4746__;
  assign new_new_n4754__ = ~new_new_n630__ & new_new_n743__;
  assign new_new_n4755__ = new_new_n1841__ & new_new_n2145__;
  assign new_new_n4756__ = new_new_n2258__ & new_new_n4729__;
  assign new_new_n4757__ = new_new_n4755__ & new_new_n4756__;
  assign new_new_n4758__ = new_new_n4753__ & new_new_n4754__;
  assign new_new_n4759__ = new_new_n4751__ & new_new_n4752__;
  assign new_new_n4760__ = new_new_n1974__ & new_new_n4743__;
  assign new_new_n4761__ = new_new_n4759__ & new_new_n4760__;
  assign new_new_n4762__ = new_new_n4757__ & new_new_n4758__;
  assign new_new_n4763__ = new_new_n4719__ & new_new_n4726__;
  assign new_new_n4764__ = new_new_n4762__ & new_new_n4763__;
  assign new_new_n4765__ = new_new_n4761__ & new_new_n4764__;
  assign new_new_n4766__ = new_new_n4742__ & new_new_n4765__;
  assign new_new_n4767__ = new_new_n4715__ & new_new_n4766__;
  assign new_new_n4768__ = new_new_n4704__ & ~new_new_n4767__;
  assign new_new_n4769__ = ~new_new_n4704__ & new_new_n4767__;
  assign new_new_n4770__ = ~new_new_n4768__ & ~new_new_n4769__;
  assign new_new_n4771__ = new_new_n4019__ & new_new_n4770__;
  assign new_new_n4772__ = ~new_new_n4019__ & ~new_new_n4770__;
  assign new_new_n4773__ = ~new_new_n4771__ & ~new_new_n4772__;
  assign new_new_n4774__ = ~new_new_n4683__ & new_new_n4773__;
  assign new_new_n4775__ = new_new_n4676__ & ~new_new_n4679__;
  assign new_new_n4776__ = ~new_new_n4675__ & ~new_new_n4775__;
  assign new_new_n4777__ = ~new_new_n4774__ & new_new_n4776__;
  assign new_new_n4778__ = pi25 & ~new_new_n466__;
  assign new_new_n4779__ = ~pi26 & ~new_new_n4778__;
  assign new_new_n4780__ = ~new_new_n74__ & ~new_new_n99__;
  assign new_new_n4781__ = ~new_new_n466__ & new_new_n4780__;
  assign new_new_n4782__ = ~new_new_n4779__ & ~new_new_n4781__;
  assign new_new_n4783__ = ~new_new_n4168__ & ~new_new_n4778__;
  assign new_new_n4784__ = ~pi26 & new_new_n4168__;
  assign new_new_n4785__ = ~new_new_n104__ & ~new_new_n4783__;
  assign new_new_n4786__ = ~new_new_n4784__ & new_new_n4785__;
  assign new_new_n4787__ = ~new_new_n4782__ & ~new_new_n4786__;
  assign new_new_n4788__ = ~new_new_n4655__ & ~new_new_n4679__;
  assign new_new_n4789__ = ~new_new_n4680__ & ~new_new_n4788__;
  assign new_new_n4790__ = ~new_new_n4655__ & ~new_new_n4676__;
  assign new_new_n4791__ = ~new_new_n4674__ & ~new_new_n4681__;
  assign new_new_n4792__ = new_new_n4790__ & new_new_n4791__;
  assign new_new_n4793__ = ~new_new_n4773__ & ~new_new_n4789__;
  assign new_new_n4794__ = ~new_new_n4792__ & new_new_n4793__;
  assign new_new_n4795__ = new_new_n4655__ & new_new_n4677__;
  assign new_new_n4796__ = ~new_new_n4672__ & new_new_n4676__;
  assign new_new_n4797__ = new_new_n4019__ & new_new_n4796__;
  assign new_new_n4798__ = new_new_n4672__ & ~new_new_n4676__;
  assign new_new_n4799__ = ~new_new_n4019__ & new_new_n4798__;
  assign new_new_n4800__ = new_new_n4655__ & ~new_new_n4673__;
  assign new_new_n4801__ = new_new_n4648__ & ~new_new_n4800__;
  assign new_new_n4802__ = ~new_new_n4799__ & new_new_n4801__;
  assign new_new_n4803__ = new_new_n4019__ & ~new_new_n4655__;
  assign new_new_n4804__ = ~new_new_n4798__ & new_new_n4803__;
  assign new_new_n4805__ = ~new_new_n4648__ & ~new_new_n4796__;
  assign new_new_n4806__ = ~new_new_n4804__ & new_new_n4805__;
  assign new_new_n4807__ = ~new_new_n4802__ & ~new_new_n4806__;
  assign new_new_n4808__ = new_new_n4773__ & ~new_new_n4795__;
  assign new_new_n4809__ = ~new_new_n4797__ & new_new_n4808__;
  assign new_new_n4810__ = ~new_new_n4807__ & new_new_n4809__;
  assign new_new_n4811__ = ~new_new_n4794__ & ~new_new_n4810__;
  assign new_new_n4812__ = ~new_new_n4787__ & new_new_n4811__;
  assign new_new_n4813__ = new_new_n4214__ & ~new_new_n4215__;
  assign new_new_n4814__ = ~new_new_n4144__ & new_new_n4813__;
  assign new_new_n4815__ = new_new_n4214__ & new_new_n4215__;
  assign new_new_n4816__ = ~new_new_n3768__ & new_new_n4815__;
  assign new_new_n4817__ = new_new_n236__ & new_new_n4209__;
  assign new_new_n4818__ = ~new_new_n3890__ & ~new_new_n4817__;
  assign new_new_n4819__ = ~new_new_n691__ & ~new_new_n4818__;
  assign new_new_n4820__ = ~new_new_n583__ & new_new_n4212__;
  assign new_new_n4821__ = ~new_new_n4816__ & ~new_new_n4819__;
  assign new_new_n4822__ = ~new_new_n4820__ & new_new_n4821__;
  assign new_new_n4823__ = ~new_new_n4814__ & new_new_n4822__;
  assign new_new_n4824__ = pi29 & ~new_new_n4823__;
  assign new_new_n4825__ = pi28 & new_new_n4214__;
  assign new_new_n4826__ = ~pi29 & new_new_n4822__;
  assign new_new_n4827__ = ~new_new_n4825__ & new_new_n4826__;
  assign new_new_n4828__ = new_new_n4811__ & ~new_new_n4827__;
  assign new_new_n4829__ = new_new_n4787__ & ~new_new_n4828__;
  assign new_new_n4830__ = new_new_n4144__ & new_new_n4826__;
  assign new_new_n4831__ = ~new_new_n4824__ & ~new_new_n4830__;
  assign new_new_n4832__ = ~new_new_n4829__ & new_new_n4831__;
  assign new_new_n4833__ = ~new_new_n4812__ & ~new_new_n4832__;
  assign new_new_n4834__ = ~new_new_n3768__ & new_new_n4212__;
  assign new_new_n4835__ = ~new_new_n583__ & ~new_new_n4818__;
  assign new_new_n4836__ = ~new_new_n466__ & new_new_n4815__;
  assign new_new_n4837__ = ~new_new_n4834__ & ~new_new_n4835__;
  assign new_new_n4838__ = ~new_new_n4836__ & new_new_n4837__;
  assign new_new_n4839__ = pi29 & ~new_new_n4838__;
  assign new_new_n4840__ = new_new_n4172__ & new_new_n4214__;
  assign new_new_n4841__ = pi29 & ~new_new_n4840__;
  assign new_new_n4842__ = ~new_new_n4825__ & new_new_n4838__;
  assign new_new_n4843__ = ~new_new_n4841__ & new_new_n4842__;
  assign new_new_n4844__ = ~new_new_n4839__ & ~new_new_n4843__;
  assign new_new_n4845__ = new_new_n4833__ & ~new_new_n4844__;
  assign new_new_n4846__ = ~new_new_n3949__ & ~new_new_n3950__;
  assign new_new_n4847__ = ~new_new_n4019__ & ~new_new_n4846__;
  assign new_new_n4848__ = ~new_new_n4034__ & ~new_new_n4660__;
  assign new_new_n4849__ = new_new_n691__ & ~new_new_n4848__;
  assign new_new_n4850__ = ~new_new_n691__ & new_new_n3720__;
  assign new_new_n4851__ = ~pi30 & new_new_n4850__;
  assign new_new_n4852__ = ~new_new_n4849__ & ~new_new_n4851__;
  assign new_new_n4853__ = new_new_n910__ & ~new_new_n4852__;
  assign new_new_n4854__ = ~new_new_n691__ & new_new_n4036__;
  assign new_new_n4855__ = ~pi30 & ~new_new_n4854__;
  assign new_new_n4856__ = ~new_new_n3720__ & ~new_new_n4855__;
  assign new_new_n4857__ = ~new_new_n4853__ & ~new_new_n4856__;
  assign new_new_n4858__ = pi29 & ~new_new_n4857__;
  assign new_new_n4859__ = ~pi29 & new_new_n4850__;
  assign new_new_n4860__ = ~new_new_n4849__ & ~new_new_n4859__;
  assign new_new_n4861__ = new_new_n910__ & ~new_new_n4860__;
  assign new_new_n4862__ = ~new_new_n691__ & ~new_new_n3720__;
  assign new_new_n4863__ = new_new_n4036__ & new_new_n4862__;
  assign new_new_n4864__ = ~new_new_n4861__ & ~new_new_n4863__;
  assign new_new_n4865__ = pi30 & ~new_new_n4864__;
  assign new_new_n4866__ = new_new_n691__ & new_new_n3720__;
  assign new_new_n4867__ = ~new_new_n4036__ & new_new_n4866__;
  assign new_new_n4868__ = ~new_new_n4854__ & ~new_new_n4867__;
  assign new_new_n4869__ = ~new_new_n161__ & ~new_new_n4868__;
  assign new_new_n4870__ = ~new_new_n71__ & ~new_new_n4862__;
  assign new_new_n4871__ = ~new_new_n4869__ & new_new_n4870__;
  assign new_new_n4872__ = ~new_new_n910__ & ~new_new_n4871__;
  assign new_new_n4873__ = ~new_new_n4858__ & ~new_new_n4865__;
  assign new_new_n4874__ = ~new_new_n4872__ & new_new_n4873__;
  assign new_new_n4875__ = pi31 & ~new_new_n4874__;
  assign new_new_n4876__ = ~pi31 & ~new_new_n71__;
  assign new_new_n4877__ = ~new_new_n4027__ & new_new_n4876__;
  assign new_new_n4878__ = ~new_new_n4048__ & new_new_n4877__;
  assign new_new_n4879__ = ~new_new_n4875__ & ~new_new_n4878__;
  assign new_new_n4880__ = ~new_new_n4768__ & new_new_n4879__;
  assign new_new_n4881__ = new_new_n4847__ & ~new_new_n4880__;
  assign new_new_n4882__ = new_new_n4019__ & new_new_n4846__;
  assign new_new_n4883__ = new_new_n4019__ & ~new_new_n4769__;
  assign new_new_n4884__ = ~new_new_n4768__ & ~new_new_n4882__;
  assign new_new_n4885__ = ~new_new_n4883__ & new_new_n4884__;
  assign new_new_n4886__ = ~new_new_n4769__ & new_new_n4882__;
  assign new_new_n4887__ = new_new_n4879__ & ~new_new_n4886__;
  assign new_new_n4888__ = ~new_new_n4885__ & ~new_new_n4887__;
  assign new_new_n4889__ = ~new_new_n4881__ & ~new_new_n4888__;
  assign new_new_n4890__ = new_new_n4768__ & ~new_new_n4879__;
  assign new_new_n4891__ = ~new_new_n4889__ & ~new_new_n4890__;
  assign new_new_n4892__ = new_new_n4847__ & ~new_new_n4891__;
  assign new_new_n4893__ = ~new_new_n4879__ & new_new_n4886__;
  assign new_new_n4894__ = ~new_new_n4889__ & ~new_new_n4893__;
  assign new_new_n4895__ = new_new_n4879__ & new_new_n4885__;
  assign new_new_n4896__ = ~new_new_n4894__ & ~new_new_n4895__;
  assign new_new_n4897__ = ~new_new_n4892__ & ~new_new_n4896__;
  assign new_new_n4898__ = ~pi25 & ~new_new_n110__;
  assign new_new_n4899__ = pi26 & new_new_n4898__;
  assign new_new_n4900__ = ~new_new_n504__ & ~new_new_n4899__;
  assign new_new_n4901__ = new_new_n4172__ & ~new_new_n4900__;
  assign new_new_n4902__ = ~new_new_n466__ & new_new_n3311__;
  assign new_new_n4903__ = new_new_n873__ & ~new_new_n3768__;
  assign new_new_n4904__ = ~new_new_n4902__ & ~new_new_n4903__;
  assign new_new_n4905__ = ~new_new_n4901__ & new_new_n4904__;
  assign new_new_n4906__ = new_new_n303__ & ~new_new_n583__;
  assign new_new_n4907__ = pi26 & ~new_new_n4906__;
  assign new_new_n4908__ = new_new_n145__ & ~new_new_n583__;
  assign new_new_n4909__ = ~pi26 & ~new_new_n4908__;
  assign new_new_n4910__ = pi23 & ~new_new_n4909__;
  assign new_new_n4911__ = ~new_new_n4907__ & ~new_new_n4910__;
  assign new_new_n4912__ = new_new_n4905__ & ~new_new_n4911__;
  assign new_new_n4913__ = ~pi26 & ~new_new_n4905__;
  assign new_new_n4914__ = ~new_new_n4912__ & ~new_new_n4913__;
  assign new_new_n4915__ = ~new_new_n1061__ & new_new_n3553__;
  assign new_new_n4916__ = ~new_new_n4287__ & ~new_new_n4915__;
  assign new_new_n4917__ = ~new_new_n3618__ & ~new_new_n4916__;
  assign new_new_n4918__ = ~new_new_n1325__ & ~new_new_n3552__;
  assign new_new_n4919__ = ~new_new_n3553__ & ~new_new_n4918__;
  assign new_new_n4920__ = ~new_new_n1148__ & ~new_new_n3552__;
  assign new_new_n4921__ = new_new_n4919__ & ~new_new_n4920__;
  assign new_new_n4922__ = new_new_n1061__ & new_new_n4921__;
  assign new_new_n4923__ = ~new_new_n1061__ & ~new_new_n4918__;
  assign new_new_n4924__ = new_new_n4288__ & ~new_new_n4923__;
  assign new_new_n4925__ = ~new_new_n4922__ & ~new_new_n4924__;
  assign new_new_n4926__ = ~new_new_n4917__ & new_new_n4925__;
  assign new_new_n4927__ = new_new_n1061__ & ~new_new_n4926__;
  assign new_new_n4928__ = new_new_n3618__ & new_new_n4925__;
  assign new_new_n4929__ = new_new_n765__ & ~new_new_n4928__;
  assign new_new_n4930__ = ~new_new_n4927__ & new_new_n4929__;
  assign new_new_n4931__ = ~new_new_n4280__ & ~new_new_n4930__;
  assign new_new_n4932__ = new_new_n1207__ & ~new_new_n4931__;
  assign new_new_n4933__ = new_new_n4548__ & new_new_n4926__;
  assign new_new_n4934__ = ~new_new_n161__ & ~new_new_n4933__;
  assign new_new_n4935__ = ~new_new_n71__ & new_new_n3618__;
  assign new_new_n4936__ = ~new_new_n4934__ & new_new_n4935__;
  assign new_new_n4937__ = new_new_n4542__ & ~new_new_n4926__;
  assign new_new_n4938__ = ~new_new_n71__ & ~new_new_n4937__;
  assign new_new_n4939__ = new_new_n4296__ & ~new_new_n4938__;
  assign new_new_n4940__ = pi31 & ~new_new_n4936__;
  assign new_new_n4941__ = ~new_new_n4939__ & new_new_n4940__;
  assign new_new_n4942__ = ~new_new_n4932__ & new_new_n4941__;
  assign new_new_n4943__ = ~new_new_n71__ & ~new_new_n1207__;
  assign new_new_n4944__ = ~new_new_n161__ & ~new_new_n4943__;
  assign new_new_n4945__ = ~pi31 & ~new_new_n4552__;
  assign new_new_n4946__ = ~new_new_n4944__ & new_new_n4945__;
  assign new_new_n4947__ = ~new_new_n4942__ & ~new_new_n4946__;
  assign new_new_n4948__ = ~new_new_n729__ & ~new_new_n1515__;
  assign new_new_n4949__ = ~new_new_n280__ & ~new_new_n724__;
  assign new_new_n4950__ = ~new_new_n222__ & ~new_new_n630__;
  assign new_new_n4951__ = ~new_new_n511__ & ~new_new_n656__;
  assign new_new_n4952__ = ~new_new_n942__ & new_new_n4951__;
  assign new_new_n4953__ = new_new_n4948__ & new_new_n4952__;
  assign new_new_n4954__ = new_new_n4949__ & new_new_n4953__;
  assign new_new_n4955__ = new_new_n4950__ & new_new_n4954__;
  assign new_new_n4956__ = ~new_new_n441__ & ~new_new_n700__;
  assign new_new_n4957__ = ~new_new_n202__ & new_new_n4956__;
  assign new_new_n4958__ = ~new_new_n961__ & new_new_n4957__;
  assign new_new_n4959__ = ~new_new_n218__ & new_new_n4958__;
  assign new_new_n4960__ = ~new_new_n148__ & ~new_new_n781__;
  assign new_new_n4961__ = ~new_new_n1265__ & new_new_n4960__;
  assign new_new_n4962__ = ~new_new_n1105__ & new_new_n4961__;
  assign new_new_n4963__ = new_new_n131__ & new_new_n1742__;
  assign new_new_n4964__ = ~new_new_n103__ & ~new_new_n476__;
  assign new_new_n4965__ = ~new_new_n693__ & ~new_new_n990__;
  assign new_new_n4966__ = new_new_n4964__ & new_new_n4965__;
  assign new_new_n4967__ = ~new_new_n721__ & new_new_n1106__;
  assign new_new_n4968__ = new_new_n3632__ & new_new_n4967__;
  assign new_new_n4969__ = new_new_n307__ & new_new_n4966__;
  assign new_new_n4970__ = ~new_new_n439__ & new_new_n1840__;
  assign new_new_n4971__ = new_new_n2866__ & new_new_n4963__;
  assign new_new_n4972__ = new_new_n4970__ & new_new_n4971__;
  assign new_new_n4973__ = new_new_n4968__ & new_new_n4969__;
  assign new_new_n4974__ = new_new_n1006__ & new_new_n4973__;
  assign new_new_n4975__ = new_new_n4959__ & new_new_n4972__;
  assign new_new_n4976__ = new_new_n4962__ & new_new_n4975__;
  assign new_new_n4977__ = new_new_n4955__ & new_new_n4974__;
  assign new_new_n4978__ = new_new_n4976__ & new_new_n4977__;
  assign new_new_n4979__ = ~new_new_n258__ & ~new_new_n382__;
  assign new_new_n4980__ = ~new_new_n658__ & ~new_new_n2170__;
  assign new_new_n4981__ = ~new_new_n263__ & ~new_new_n346__;
  assign new_new_n4982__ = ~new_new_n226__ & ~new_new_n783__;
  assign new_new_n4983__ = ~new_new_n1008__ & new_new_n4980__;
  assign new_new_n4984__ = new_new_n4982__ & new_new_n4983__;
  assign new_new_n4985__ = new_new_n4979__ & new_new_n4981__;
  assign new_new_n4986__ = new_new_n4984__ & new_new_n4985__;
  assign new_new_n4987__ = new_new_n1961__ & new_new_n2454__;
  assign new_new_n4988__ = ~new_new_n254__ & ~new_new_n322__;
  assign new_new_n4989__ = ~new_new_n101__ & ~new_new_n488__;
  assign new_new_n4990__ = ~new_new_n196__ & ~new_new_n480__;
  assign new_new_n4991__ = ~new_new_n995__ & new_new_n4990__;
  assign new_new_n4992__ = ~new_new_n255__ & new_new_n4991__;
  assign new_new_n4993__ = new_new_n4989__ & new_new_n4992__;
  assign new_new_n4994__ = new_new_n4988__ & new_new_n4993__;
  assign new_new_n4995__ = new_new_n1213__ & new_new_n1424__;
  assign new_new_n4996__ = ~new_new_n106__ & ~new_new_n267__;
  assign new_new_n4997__ = ~new_new_n749__ & new_new_n4996__;
  assign new_new_n4998__ = ~new_new_n150__ & ~new_new_n1073__;
  assign new_new_n4999__ = new_new_n4997__ & new_new_n4998__;
  assign new_new_n5000__ = ~new_new_n115__ & new_new_n1679__;
  assign new_new_n5001__ = new_new_n4995__ & new_new_n5000__;
  assign new_new_n5002__ = new_new_n3281__ & new_new_n4999__;
  assign new_new_n5003__ = new_new_n4743__ & new_new_n4987__;
  assign new_new_n5004__ = new_new_n5002__ & new_new_n5003__;
  assign new_new_n5005__ = new_new_n4986__ & new_new_n5001__;
  assign new_new_n5006__ = new_new_n5004__ & new_new_n5005__;
  assign new_new_n5007__ = new_new_n4994__ & new_new_n5006__;
  assign new_new_n5008__ = ~new_new_n92__ & ~new_new_n772__;
  assign new_new_n5009__ = ~new_new_n270__ & new_new_n5008__;
  assign new_new_n5010__ = new_new_n1332__ & new_new_n1830__;
  assign new_new_n5011__ = new_new_n5009__ & new_new_n5010__;
  assign new_new_n5012__ = new_new_n1306__ & new_new_n1775__;
  assign new_new_n5013__ = new_new_n3773__ & new_new_n5012__;
  assign new_new_n5014__ = new_new_n378__ & new_new_n5011__;
  assign new_new_n5015__ = new_new_n5013__ & new_new_n5014__;
  assign new_new_n5016__ = new_new_n1262__ & new_new_n2430__;
  assign new_new_n5017__ = new_new_n5015__ & new_new_n5016__;
  assign new_new_n5018__ = new_new_n2802__ & new_new_n5017__;
  assign new_new_n5019__ = new_new_n4978__ & new_new_n5018__;
  assign new_new_n5020__ = new_new_n5007__ & new_new_n5019__;
  assign new_new_n5021__ = ~pi31 & new_new_n765__;
  assign new_new_n5022__ = ~new_new_n1325__ & new_new_n5021__;
  assign new_new_n5023__ = new_new_n161__ & ~new_new_n1466__;
  assign new_new_n5024__ = new_new_n1466__ & ~new_new_n1556__;
  assign new_new_n5025__ = ~new_new_n1466__ & new_new_n1556__;
  assign new_new_n5026__ = ~new_new_n5024__ & ~new_new_n5025__;
  assign new_new_n5027__ = new_new_n1325__ & new_new_n5026__;
  assign new_new_n5028__ = ~new_new_n1325__ & new_new_n5024__;
  assign new_new_n5029__ = ~new_new_n3544__ & new_new_n5028__;
  assign new_new_n5030__ = new_new_n1325__ & ~new_new_n1466__;
  assign new_new_n5031__ = new_new_n1737__ & new_new_n5030__;
  assign new_new_n5032__ = ~new_new_n5029__ & ~new_new_n5031__;
  assign new_new_n5033__ = new_new_n1660__ & ~new_new_n5032__;
  assign new_new_n5034__ = new_new_n1467__ & ~new_new_n1737__;
  assign new_new_n5035__ = new_new_n1556__ & new_new_n1739__;
  assign new_new_n5036__ = new_new_n3544__ & new_new_n5035__;
  assign new_new_n5037__ = ~new_new_n5034__ & ~new_new_n5036__;
  assign new_new_n5038__ = ~new_new_n1660__ & ~new_new_n5037__;
  assign new_new_n5039__ = ~new_new_n3544__ & new_new_n5030__;
  assign new_new_n5040__ = ~new_new_n5028__ & ~new_new_n5039__;
  assign new_new_n5041__ = new_new_n1737__ & ~new_new_n5040__;
  assign new_new_n5042__ = new_new_n1467__ & new_new_n3544__;
  assign new_new_n5043__ = ~new_new_n5035__ & ~new_new_n5042__;
  assign new_new_n5044__ = ~new_new_n1737__ & ~new_new_n5043__;
  assign new_new_n5045__ = ~new_new_n5027__ & ~new_new_n5033__;
  assign new_new_n5046__ = ~new_new_n5038__ & ~new_new_n5041__;
  assign new_new_n5047__ = ~new_new_n5044__ & new_new_n5046__;
  assign new_new_n5048__ = new_new_n5045__ & new_new_n5047__;
  assign new_new_n5049__ = new_new_n765__ & new_new_n5048__;
  assign new_new_n5050__ = ~new_new_n5023__ & ~new_new_n5049__;
  assign new_new_n5051__ = pi31 & ~new_new_n5050__;
  assign new_new_n5052__ = ~pi31 & ~new_new_n161__;
  assign new_new_n5053__ = ~new_new_n4147__ & ~new_new_n5052__;
  assign new_new_n5054__ = ~new_new_n1556__ & new_new_n5053__;
  assign new_new_n5055__ = ~new_new_n5022__ & ~new_new_n5054__;
  assign new_new_n5056__ = ~new_new_n5051__ & new_new_n5055__;
  assign new_new_n5057__ = ~new_new_n5020__ & ~new_new_n5056__;
  assign new_new_n5058__ = ~new_new_n1325__ & new_new_n5053__;
  assign new_new_n5059__ = pi31 & new_new_n161__;
  assign new_new_n5060__ = ~new_new_n1556__ & new_new_n5059__;
  assign new_new_n5061__ = ~new_new_n3618__ & new_new_n4921__;
  assign new_new_n5062__ = pi31 & new_new_n5061__;
  assign new_new_n5063__ = pi31 & new_new_n4921__;
  assign new_new_n5064__ = new_new_n3618__ & ~new_new_n5063__;
  assign new_new_n5065__ = new_new_n765__ & ~new_new_n5062__;
  assign new_new_n5066__ = ~new_new_n5064__ & new_new_n5065__;
  assign new_new_n5067__ = ~new_new_n5058__ & ~new_new_n5060__;
  assign new_new_n5068__ = ~new_new_n5066__ & new_new_n5067__;
  assign new_new_n5069__ = new_new_n5057__ & ~new_new_n5068__;
  assign new_new_n5070__ = new_new_n5020__ & new_new_n5056__;
  assign new_new_n5071__ = ~new_new_n4386__ & ~new_new_n4387__;
  assign new_new_n5072__ = new_new_n5070__ & ~new_new_n5071__;
  assign new_new_n5073__ = ~new_new_n5070__ & new_new_n5071__;
  assign new_new_n5074__ = new_new_n5068__ & ~new_new_n5073__;
  assign new_new_n5075__ = new_new_n4452__ & ~new_new_n5072__;
  assign new_new_n5076__ = ~new_new_n5074__ & new_new_n5075__;
  assign new_new_n5077__ = ~new_new_n5057__ & new_new_n5068__;
  assign new_new_n5078__ = ~new_new_n4452__ & ~new_new_n5071__;
  assign new_new_n5079__ = ~new_new_n5077__ & new_new_n5078__;
  assign new_new_n5080__ = ~new_new_n5069__ & ~new_new_n5076__;
  assign new_new_n5081__ = ~new_new_n5079__ & new_new_n5080__;
  assign new_new_n5082__ = ~new_new_n4302__ & ~new_new_n4456__;
  assign new_new_n5083__ = new_new_n4454__ & new_new_n5082__;
  assign new_new_n5084__ = ~new_new_n4454__ & ~new_new_n5082__;
  assign new_new_n5085__ = ~new_new_n5083__ & ~new_new_n5084__;
  assign new_new_n5086__ = new_new_n5081__ & ~new_new_n5085__;
  assign new_new_n5087__ = ~new_new_n5081__ & new_new_n5085__;
  assign new_new_n5088__ = ~new_new_n868__ & new_new_n4212__;
  assign new_new_n5089__ = ~new_new_n4032__ & ~new_new_n4215__;
  assign new_new_n5090__ = new_new_n3720__ & ~new_new_n5089__;
  assign new_new_n5091__ = ~new_new_n3720__ & new_new_n5089__;
  assign new_new_n5092__ = new_new_n4214__ & ~new_new_n5090__;
  assign new_new_n5093__ = ~new_new_n5091__ & new_new_n5092__;
  assign new_new_n5094__ = ~new_new_n5088__ & ~new_new_n5093__;
  assign new_new_n5095__ = new_new_n67__ & ~new_new_n1207__;
  assign new_new_n5096__ = pi29 & ~new_new_n5095__;
  assign new_new_n5097__ = new_new_n65__ & ~new_new_n1207__;
  assign new_new_n5098__ = ~pi29 & ~new_new_n5097__;
  assign new_new_n5099__ = pi26 & ~new_new_n5098__;
  assign new_new_n5100__ = ~new_new_n5096__ & ~new_new_n5099__;
  assign new_new_n5101__ = new_new_n5094__ & ~new_new_n5100__;
  assign new_new_n5102__ = ~pi29 & ~new_new_n5094__;
  assign new_new_n5103__ = ~new_new_n5101__ & ~new_new_n5102__;
  assign new_new_n5104__ = ~new_new_n5087__ & new_new_n5103__;
  assign new_new_n5105__ = ~new_new_n5086__ & ~new_new_n5104__;
  assign new_new_n5106__ = ~new_new_n4947__ & new_new_n5105__;
  assign new_new_n5107__ = new_new_n4947__ & ~new_new_n5105__;
  assign new_new_n5108__ = ~new_new_n5106__ & ~new_new_n5107__;
  assign new_new_n5109__ = ~new_new_n4455__ & ~new_new_n4457__;
  assign new_new_n5110__ = new_new_n4524__ & ~new_new_n5109__;
  assign new_new_n5111__ = ~new_new_n4524__ & new_new_n5109__;
  assign new_new_n5112__ = ~new_new_n5110__ & ~new_new_n5111__;
  assign new_new_n5113__ = new_new_n5108__ & new_new_n5112__;
  assign new_new_n5114__ = ~new_new_n5108__ & ~new_new_n5112__;
  assign new_new_n5115__ = ~new_new_n5113__ & ~new_new_n5114__;
  assign new_new_n5116__ = ~new_new_n910__ & ~new_new_n4036__;
  assign new_new_n5117__ = pi29 & new_new_n5116__;
  assign new_new_n5118__ = ~new_new_n868__ & ~new_new_n4818__;
  assign new_new_n5119__ = ~new_new_n3720__ & new_new_n4212__;
  assign new_new_n5120__ = ~new_new_n5118__ & ~new_new_n5119__;
  assign new_new_n5121__ = new_new_n910__ & new_new_n4036__;
  assign new_new_n5122__ = ~pi28 & new_new_n5120__;
  assign new_new_n5123__ = new_new_n5121__ & new_new_n5122__;
  assign new_new_n5124__ = ~new_new_n5117__ & ~new_new_n5123__;
  assign new_new_n5125__ = new_new_n4214__ & ~new_new_n5124__;
  assign new_new_n5126__ = ~pi29 & new_new_n4214__;
  assign new_new_n5127__ = ~new_new_n910__ & new_new_n4036__;
  assign new_new_n5128__ = pi28 & new_new_n5127__;
  assign new_new_n5129__ = new_new_n910__ & ~new_new_n4036__;
  assign new_new_n5130__ = new_new_n5126__ & ~new_new_n5129__;
  assign new_new_n5131__ = ~new_new_n5128__ & new_new_n5130__;
  assign new_new_n5132__ = ~pi29 & ~new_new_n5120__;
  assign new_new_n5133__ = pi29 & new_new_n5120__;
  assign new_new_n5134__ = ~new_new_n5132__ & ~new_new_n5133__;
  assign new_new_n5135__ = ~new_new_n5131__ & new_new_n5134__;
  assign new_new_n5136__ = ~new_new_n5125__ & ~new_new_n5135__;
  assign new_new_n5137__ = new_new_n5115__ & ~new_new_n5136__;
  assign new_new_n5138__ = ~new_new_n5115__ & new_new_n5136__;
  assign new_new_n5139__ = ~new_new_n4144__ & ~new_new_n4900__;
  assign new_new_n5140__ = new_new_n3311__ & ~new_new_n3768__;
  assign new_new_n5141__ = ~new_new_n333__ & ~new_new_n691__;
  assign new_new_n5142__ = ~new_new_n583__ & new_new_n873__;
  assign new_new_n5143__ = ~new_new_n5140__ & ~new_new_n5141__;
  assign new_new_n5144__ = ~new_new_n5142__ & new_new_n5143__;
  assign new_new_n5145__ = ~new_new_n5139__ & new_new_n5144__;
  assign new_new_n5146__ = pi26 & ~new_new_n5145__;
  assign new_new_n5147__ = ~pi26 & new_new_n5145__;
  assign new_new_n5148__ = ~new_new_n5146__ & ~new_new_n5147__;
  assign new_new_n5149__ = ~new_new_n5138__ & ~new_new_n5148__;
  assign new_new_n5150__ = ~new_new_n5137__ & ~new_new_n5149__;
  assign new_new_n5151__ = new_new_n4914__ & ~new_new_n5150__;
  assign new_new_n5152__ = ~new_new_n4914__ & new_new_n5150__;
  assign new_new_n5153__ = ~new_new_n5107__ & ~new_new_n5112__;
  assign new_new_n5154__ = ~new_new_n5106__ & ~new_new_n5153__;
  assign new_new_n5155__ = ~new_new_n3720__ & ~new_new_n4818__;
  assign new_new_n5156__ = ~new_new_n691__ & new_new_n4815__;
  assign new_new_n5157__ = ~new_new_n910__ & new_new_n4212__;
  assign new_new_n5158__ = ~new_new_n5155__ & ~new_new_n5156__;
  assign new_new_n5159__ = ~new_new_n5157__ & new_new_n5158__;
  assign new_new_n5160__ = new_new_n4042__ & new_new_n4214__;
  assign new_new_n5161__ = pi29 & ~new_new_n5160__;
  assign new_new_n5162__ = new_new_n4042__ & new_new_n4825__;
  assign new_new_n5163__ = ~new_new_n5161__ & ~new_new_n5162__;
  assign new_new_n5164__ = new_new_n5159__ & ~new_new_n5163__;
  assign new_new_n5165__ = ~pi29 & ~new_new_n5159__;
  assign new_new_n5166__ = ~new_new_n5164__ & ~new_new_n5165__;
  assign new_new_n5167__ = ~new_new_n4562__ & ~new_new_n4563__;
  assign new_new_n5168__ = ~new_new_n4652__ & new_new_n5167__;
  assign new_new_n5169__ = new_new_n4652__ & ~new_new_n5167__;
  assign new_new_n5170__ = ~new_new_n5168__ & ~new_new_n5169__;
  assign new_new_n5171__ = new_new_n5166__ & ~new_new_n5170__;
  assign new_new_n5172__ = ~new_new_n5166__ & new_new_n5170__;
  assign new_new_n5173__ = ~new_new_n5171__ & ~new_new_n5172__;
  assign new_new_n5174__ = new_new_n5154__ & new_new_n5173__;
  assign new_new_n5175__ = ~new_new_n5154__ & ~new_new_n5173__;
  assign new_new_n5176__ = ~new_new_n5174__ & ~new_new_n5175__;
  assign new_new_n5177__ = ~new_new_n5152__ & ~new_new_n5176__;
  assign new_new_n5178__ = ~new_new_n5151__ & ~new_new_n5177__;
  assign new_new_n5179__ = ~pi20 & ~pi21;
  assign new_new_n5180__ = pi22 & ~new_new_n5179__;
  assign new_new_n5181__ = pi20 & pi21;
  assign new_new_n5182__ = ~pi22 & ~new_new_n5181__;
  assign new_new_n5183__ = ~new_new_n5180__ & ~new_new_n5182__;
  assign new_new_n5184__ = ~new_new_n3768__ & new_new_n5183__;
  assign new_new_n5185__ = ~pi21 & ~pi22;
  assign new_new_n5186__ = ~pi20 & new_new_n5185__;
  assign new_new_n5187__ = pi23 & ~new_new_n5186__;
  assign new_new_n5188__ = pi21 & pi22;
  assign new_new_n5189__ = pi20 & new_new_n5188__;
  assign new_new_n5190__ = ~pi23 & ~new_new_n5189__;
  assign new_new_n5191__ = ~new_new_n5187__ & ~new_new_n5190__;
  assign new_new_n5192__ = ~new_new_n583__ & new_new_n5191__;
  assign new_new_n5193__ = ~new_new_n5184__ & ~new_new_n5192__;
  assign new_new_n5194__ = ~new_new_n466__ & ~new_new_n4169__;
  assign new_new_n5195__ = ~new_new_n5179__ & ~new_new_n5181__;
  assign new_new_n5196__ = new_new_n5194__ & new_new_n5195__;
  assign new_new_n5197__ = new_new_n5193__ & ~new_new_n5196__;
  assign new_new_n5198__ = pi23 & ~new_new_n5197__;
  assign new_new_n5199__ = ~new_new_n4170__ & new_new_n5195__;
  assign new_new_n5200__ = pi23 & ~new_new_n5199__;
  assign new_new_n5201__ = ~pi22 & ~new_new_n466__;
  assign new_new_n5202__ = pi22 & new_new_n4172__;
  assign new_new_n5203__ = ~new_new_n5201__ & ~new_new_n5202__;
  assign new_new_n5204__ = new_new_n5199__ & ~new_new_n5203__;
  assign new_new_n5205__ = new_new_n5193__ & ~new_new_n5200__;
  assign new_new_n5206__ = ~new_new_n5204__ & new_new_n5205__;
  assign new_new_n5207__ = ~new_new_n5198__ & ~new_new_n5206__;
  assign new_new_n5208__ = ~new_new_n910__ & new_new_n5191__;
  assign new_new_n5209__ = ~new_new_n691__ & new_new_n5183__;
  assign new_new_n5210__ = ~pi22 & ~pi23;
  assign new_new_n5211__ = pi22 & pi23;
  assign new_new_n5212__ = ~new_new_n5210__ & ~new_new_n5211__;
  assign new_new_n5213__ = new_new_n5195__ & ~new_new_n5212__;
  assign new_new_n5214__ = ~new_new_n583__ & new_new_n5213__;
  assign new_new_n5215__ = new_new_n5195__ & new_new_n5212__;
  assign new_new_n5216__ = new_new_n3742__ & new_new_n5215__;
  assign new_new_n5217__ = ~new_new_n5209__ & ~new_new_n5214__;
  assign new_new_n5218__ = ~new_new_n5208__ & new_new_n5217__;
  assign new_new_n5219__ = ~new_new_n5216__ & new_new_n5218__;
  assign new_new_n5220__ = new_new_n4542__ & ~new_new_n4921__;
  assign new_new_n5221__ = ~new_new_n1061__ & new_new_n1207__;
  assign new_new_n5222__ = new_new_n3618__ & new_new_n5221__;
  assign new_new_n5223__ = ~new_new_n5220__ & ~new_new_n5222__;
  assign new_new_n5224__ = new_new_n3552__ & ~new_new_n5223__;
  assign new_new_n5225__ = new_new_n1207__ & new_new_n1325__;
  assign new_new_n5226__ = new_new_n3618__ & new_new_n5225__;
  assign new_new_n5227__ = ~new_new_n4542__ & ~new_new_n5226__;
  assign new_new_n5228__ = ~new_new_n1061__ & ~new_new_n5227__;
  assign new_new_n5229__ = ~new_new_n1207__ & new_new_n3618__;
  assign new_new_n5230__ = ~new_new_n4923__ & new_new_n5229__;
  assign new_new_n5231__ = new_new_n1207__ & new_new_n4289__;
  assign new_new_n5232__ = ~new_new_n3553__ & new_new_n5231__;
  assign new_new_n5233__ = ~new_new_n5228__ & ~new_new_n5232__;
  assign new_new_n5234__ = ~new_new_n5230__ & new_new_n5233__;
  assign new_new_n5235__ = ~new_new_n5224__ & new_new_n5234__;
  assign new_new_n5236__ = ~new_new_n4900__ & ~new_new_n5235__;
  assign new_new_n5237__ = new_new_n873__ & ~new_new_n1061__;
  assign new_new_n5238__ = ~new_new_n333__ & ~new_new_n3618__;
  assign new_new_n5239__ = ~new_new_n1207__ & new_new_n3311__;
  assign new_new_n5240__ = ~new_new_n5237__ & ~new_new_n5238__;
  assign new_new_n5241__ = ~new_new_n5239__ & new_new_n5240__;
  assign new_new_n5242__ = ~new_new_n5236__ & new_new_n5241__;
  assign new_new_n5243__ = pi26 & ~new_new_n5242__;
  assign new_new_n5244__ = ~pi26 & new_new_n5242__;
  assign new_new_n5245__ = ~new_new_n5243__ & ~new_new_n5244__;
  assign new_new_n5246__ = new_new_n765__ & ~new_new_n1660__;
  assign new_new_n5247__ = new_new_n161__ & ~new_new_n1902__;
  assign new_new_n5248__ = ~new_new_n5246__ & ~new_new_n5247__;
  assign new_new_n5249__ = ~pi31 & ~new_new_n5248__;
  assign new_new_n5250__ = ~pi29 & new_new_n1902__;
  assign new_new_n5251__ = ~pi30 & new_new_n5250__;
  assign new_new_n5252__ = ~new_new_n1902__ & new_new_n3541__;
  assign new_new_n5253__ = new_new_n1823__ & ~new_new_n3535__;
  assign new_new_n5254__ = ~new_new_n1660__ & new_new_n5253__;
  assign new_new_n5255__ = new_new_n1660__ & ~new_new_n1823__;
  assign new_new_n5256__ = new_new_n1902__ & new_new_n5255__;
  assign new_new_n5257__ = new_new_n3479__ & new_new_n5256__;
  assign new_new_n5258__ = ~new_new_n5254__ & ~new_new_n5257__;
  assign new_new_n5259__ = ~new_new_n2130__ & ~new_new_n5258__;
  assign new_new_n5260__ = new_new_n1824__ & ~new_new_n1902__;
  assign new_new_n5261__ = new_new_n2130__ & new_new_n5260__;
  assign new_new_n5262__ = new_new_n3535__ & new_new_n3541__;
  assign new_new_n5263__ = ~new_new_n5261__ & ~new_new_n5262__;
  assign new_new_n5264__ = ~new_new_n3479__ & ~new_new_n5263__;
  assign new_new_n5265__ = new_new_n2130__ & new_new_n3541__;
  assign new_new_n5266__ = ~new_new_n5260__ & ~new_new_n5265__;
  assign new_new_n5267__ = new_new_n3535__ & ~new_new_n5266__;
  assign new_new_n5268__ = ~new_new_n1823__ & ~new_new_n3535__;
  assign new_new_n5269__ = new_new_n1660__ & ~new_new_n5268__;
  assign new_new_n5270__ = new_new_n3542__ & ~new_new_n5269__;
  assign new_new_n5271__ = ~new_new_n5267__ & ~new_new_n5270__;
  assign new_new_n5272__ = ~new_new_n5264__ & new_new_n5271__;
  assign new_new_n5273__ = ~new_new_n5259__ & new_new_n5272__;
  assign new_new_n5274__ = ~new_new_n5252__ & new_new_n5273__;
  assign new_new_n5275__ = new_new_n765__ & new_new_n5274__;
  assign new_new_n5276__ = pi30 & new_new_n1823__;
  assign new_new_n5277__ = pi29 & new_new_n5276__;
  assign new_new_n5278__ = pi31 & ~new_new_n5251__;
  assign new_new_n5279__ = ~new_new_n5277__ & new_new_n5278__;
  assign new_new_n5280__ = ~new_new_n5275__ & new_new_n5279__;
  assign new_new_n5281__ = ~new_new_n5249__ & ~new_new_n5280__;
  assign new_new_n5282__ = ~new_new_n274__ & ~new_new_n2170__;
  assign new_new_n5283__ = ~new_new_n1033__ & ~new_new_n2344__;
  assign new_new_n5284__ = ~new_new_n935__ & new_new_n5283__;
  assign new_new_n5285__ = new_new_n5282__ & new_new_n5284__;
  assign new_new_n5286__ = new_new_n3774__ & new_new_n5285__;
  assign new_new_n5287__ = ~new_new_n76__ & ~new_new_n637__;
  assign new_new_n5288__ = ~new_new_n270__ & ~new_new_n308__;
  assign new_new_n5289__ = ~new_new_n606__ & new_new_n5287__;
  assign new_new_n5290__ = new_new_n5288__ & new_new_n5289__;
  assign new_new_n5291__ = ~new_new_n344__ & new_new_n1447__;
  assign new_new_n5292__ = new_new_n2758__ & new_new_n3139__;
  assign new_new_n5293__ = new_new_n4092__ & new_new_n5292__;
  assign new_new_n5294__ = new_new_n5290__ & new_new_n5291__;
  assign new_new_n5295__ = new_new_n709__ & new_new_n3567__;
  assign new_new_n5296__ = new_new_n3699__ & new_new_n5295__;
  assign new_new_n5297__ = new_new_n5293__ & new_new_n5294__;
  assign new_new_n5298__ = new_new_n3389__ & new_new_n5297__;
  assign new_new_n5299__ = new_new_n4994__ & new_new_n5296__;
  assign new_new_n5300__ = new_new_n5298__ & new_new_n5299__;
  assign new_new_n5301__ = ~new_new_n838__ & ~new_new_n961__;
  assign new_new_n5302__ = ~new_new_n717__ & ~new_new_n828__;
  assign new_new_n5303__ = ~new_new_n438__ & ~new_new_n952__;
  assign new_new_n5304__ = ~new_new_n300__ & ~new_new_n921__;
  assign new_new_n5305__ = ~new_new_n1632__ & new_new_n5304__;
  assign new_new_n5306__ = new_new_n3367__ & new_new_n5301__;
  assign new_new_n5307__ = new_new_n5302__ & new_new_n5303__;
  assign new_new_n5308__ = new_new_n5306__ & new_new_n5307__;
  assign new_new_n5309__ = new_new_n1752__ & new_new_n5305__;
  assign new_new_n5310__ = new_new_n5308__ & new_new_n5309__;
  assign new_new_n5311__ = ~new_new_n82__ & ~new_new_n313__;
  assign new_new_n5312__ = ~new_new_n249__ & ~new_new_n316__;
  assign new_new_n5313__ = ~new_new_n350__ & ~new_new_n602__;
  assign new_new_n5314__ = ~new_new_n160__ & ~new_new_n588__;
  assign new_new_n5315__ = ~new_new_n947__ & new_new_n5314__;
  assign new_new_n5316__ = ~new_new_n698__ & ~new_new_n701__;
  assign new_new_n5317__ = ~new_new_n724__ & new_new_n5316__;
  assign new_new_n5318__ = ~new_new_n919__ & new_new_n1909__;
  assign new_new_n5319__ = new_new_n2174__ & new_new_n5318__;
  assign new_new_n5320__ = new_new_n5313__ & new_new_n5317__;
  assign new_new_n5321__ = new_new_n5319__ & new_new_n5320__;
  assign new_new_n5322__ = new_new_n1598__ & new_new_n5312__;
  assign new_new_n5323__ = new_new_n5315__ & new_new_n5322__;
  assign new_new_n5324__ = new_new_n5321__ & new_new_n5323__;
  assign new_new_n5325__ = new_new_n241__ & ~new_new_n1165__;
  assign new_new_n5326__ = ~new_new_n130__ & ~new_new_n179__;
  assign new_new_n5327__ = ~new_new_n222__ & ~new_new_n1113__;
  assign new_new_n5328__ = new_new_n5326__ & new_new_n5327__;
  assign new_new_n5329__ = new_new_n1505__ & new_new_n3587__;
  assign new_new_n5330__ = ~new_new_n5325__ & new_new_n5329__;
  assign new_new_n5331__ = new_new_n1230__ & new_new_n5328__;
  assign new_new_n5332__ = new_new_n1994__ & new_new_n1995__;
  assign new_new_n5333__ = new_new_n3642__ & new_new_n5332__;
  assign new_new_n5334__ = new_new_n5330__ & new_new_n5331__;
  assign new_new_n5335__ = new_new_n5333__ & new_new_n5334__;
  assign new_new_n5336__ = new_new_n3698__ & new_new_n5335__;
  assign new_new_n5337__ = new_new_n5324__ & new_new_n5336__;
  assign new_new_n5338__ = ~new_new_n164__ & ~new_new_n482__;
  assign new_new_n5339__ = ~new_new_n1291__ & new_new_n5338__;
  assign new_new_n5340__ = ~new_new_n150__ & ~new_new_n311__;
  assign new_new_n5341__ = new_new_n1368__ & new_new_n3204__;
  assign new_new_n5342__ = new_new_n5311__ & new_new_n5341__;
  assign new_new_n5343__ = new_new_n5339__ & new_new_n5340__;
  assign new_new_n5344__ = ~new_new_n439__ & new_new_n830__;
  assign new_new_n5345__ = ~new_new_n837__ & new_new_n2581__;
  assign new_new_n5346__ = new_new_n3276__ & new_new_n3482__;
  assign new_new_n5347__ = new_new_n3484__ & new_new_n5346__;
  assign new_new_n5348__ = new_new_n5344__ & new_new_n5345__;
  assign new_new_n5349__ = new_new_n5342__ & new_new_n5343__;
  assign new_new_n5350__ = new_new_n5348__ & new_new_n5349__;
  assign new_new_n5351__ = new_new_n5347__ & new_new_n5350__;
  assign new_new_n5352__ = new_new_n5286__ & new_new_n5310__;
  assign new_new_n5353__ = new_new_n5351__ & new_new_n5352__;
  assign new_new_n5354__ = new_new_n5300__ & new_new_n5353__;
  assign new_new_n5355__ = new_new_n5337__ & new_new_n5354__;
  assign new_new_n5356__ = ~pi14 & ~new_new_n5355__;
  assign new_new_n5357__ = pi14 & new_new_n5355__;
  assign new_new_n5358__ = ~new_new_n308__ & ~new_new_n1372__;
  assign new_new_n5359__ = ~new_new_n207__ & ~new_new_n271__;
  assign new_new_n5360__ = ~new_new_n155__ & new_new_n5359__;
  assign new_new_n5361__ = ~new_new_n489__ & new_new_n1946__;
  assign new_new_n5362__ = new_new_n5358__ & new_new_n5361__;
  assign new_new_n5363__ = new_new_n5360__ & new_new_n5362__;
  assign new_new_n5364__ = new_new_n2641__ & new_new_n5363__;
  assign new_new_n5365__ = ~new_new_n835__ & ~new_new_n845__;
  assign new_new_n5366__ = ~new_new_n332__ & ~new_new_n675__;
  assign new_new_n5367__ = ~new_new_n200__ & ~new_new_n283__;
  assign new_new_n5368__ = ~new_new_n309__ & ~new_new_n656__;
  assign new_new_n5369__ = new_new_n5367__ & new_new_n5368__;
  assign new_new_n5370__ = ~new_new_n192__ & ~new_new_n270__;
  assign new_new_n5371__ = new_new_n5369__ & new_new_n5370__;
  assign new_new_n5372__ = ~new_new_n373__ & new_new_n2161__;
  assign new_new_n5373__ = new_new_n5365__ & new_new_n5366__;
  assign new_new_n5374__ = new_new_n5372__ & new_new_n5373__;
  assign new_new_n5375__ = new_new_n4504__ & new_new_n5371__;
  assign new_new_n5376__ = new_new_n4950__ & new_new_n5375__;
  assign new_new_n5377__ = new_new_n5374__ & new_new_n5376__;
  assign new_new_n5378__ = ~new_new_n351__ & ~new_new_n700__;
  assign new_new_n5379__ = ~new_new_n276__ & ~new_new_n624__;
  assign new_new_n5380__ = ~new_new_n250__ & ~new_new_n869__;
  assign new_new_n5381__ = new_new_n5378__ & new_new_n5380__;
  assign new_new_n5382__ = new_new_n5379__ & new_new_n5381__;
  assign new_new_n5383__ = ~new_new_n940__ & ~new_new_n947__;
  assign new_new_n5384__ = ~new_new_n183__ & new_new_n3206__;
  assign new_new_n5385__ = new_new_n2027__ & new_new_n2708__;
  assign new_new_n5386__ = new_new_n3056__ & new_new_n5385__;
  assign new_new_n5387__ = new_new_n3098__ & new_new_n5386__;
  assign new_new_n5388__ = new_new_n5384__ & new_new_n5387__;
  assign new_new_n5389__ = new_new_n133__ & new_new_n424__;
  assign new_new_n5390__ = ~new_new_n221__ & ~new_new_n224__;
  assign new_new_n5391__ = ~new_new_n217__ & new_new_n5390__;
  assign new_new_n5392__ = new_new_n118__ & ~new_new_n5391__;
  assign new_new_n5393__ = ~new_new_n248__ & ~new_new_n875__;
  assign new_new_n5394__ = new_new_n2340__ & new_new_n5393__;
  assign new_new_n5395__ = ~new_new_n5389__ & new_new_n5394__;
  assign new_new_n5396__ = ~new_new_n5392__ & new_new_n5395__;
  assign new_new_n5397__ = ~new_new_n843__ & ~new_new_n1212__;
  assign new_new_n5398__ = ~new_new_n202__ & new_new_n2477__;
  assign new_new_n5399__ = ~new_new_n226__ & ~new_new_n477__;
  assign new_new_n5400__ = new_new_n1366__ & new_new_n5383__;
  assign new_new_n5401__ = new_new_n5397__ & new_new_n5400__;
  assign new_new_n5402__ = new_new_n5398__ & new_new_n5399__;
  assign new_new_n5403__ = new_new_n1074__ & new_new_n1253__;
  assign new_new_n5404__ = new_new_n2919__ & new_new_n5403__;
  assign new_new_n5405__ = new_new_n5401__ & new_new_n5402__;
  assign new_new_n5406__ = new_new_n2028__ & new_new_n5405__;
  assign new_new_n5407__ = new_new_n5382__ & new_new_n5404__;
  assign new_new_n5408__ = new_new_n5396__ & new_new_n5407__;
  assign new_new_n5409__ = new_new_n5388__ & new_new_n5406__;
  assign new_new_n5410__ = new_new_n5408__ & new_new_n5409__;
  assign new_new_n5411__ = ~new_new_n1398__ & ~new_new_n1507__;
  assign new_new_n5412__ = ~new_new_n344__ & new_new_n5411__;
  assign new_new_n5413__ = ~new_new_n127__ & ~new_new_n1162__;
  assign new_new_n5414__ = ~new_new_n168__ & ~new_new_n496__;
  assign new_new_n5415__ = new_new_n5413__ & new_new_n5414__;
  assign new_new_n5416__ = ~new_new_n119__ & ~new_new_n208__;
  assign new_new_n5417__ = ~new_new_n259__ & new_new_n5416__;
  assign new_new_n5418__ = new_new_n605__ & new_new_n2314__;
  assign new_new_n5419__ = new_new_n5311__ & new_new_n5418__;
  assign new_new_n5420__ = ~new_new_n607__ & new_new_n5417__;
  assign new_new_n5421__ = new_new_n965__ & new_new_n3913__;
  assign new_new_n5422__ = new_new_n5415__ & new_new_n5421__;
  assign new_new_n5423__ = new_new_n5419__ & new_new_n5420__;
  assign new_new_n5424__ = ~new_new_n1539__ & new_new_n2989__;
  assign new_new_n5425__ = new_new_n4090__ & new_new_n5412__;
  assign new_new_n5426__ = new_new_n5424__ & new_new_n5425__;
  assign new_new_n5427__ = new_new_n5422__ & new_new_n5423__;
  assign new_new_n5428__ = new_new_n1068__ & new_new_n5427__;
  assign new_new_n5429__ = new_new_n5426__ & new_new_n5428__;
  assign new_new_n5430__ = ~new_new_n658__ & ~new_new_n853__;
  assign new_new_n5431__ = ~new_new_n232__ & ~new_new_n721__;
  assign new_new_n5432__ = ~new_new_n150__ & ~new_new_n479__;
  assign new_new_n5433__ = ~new_new_n724__ & ~new_new_n729__;
  assign new_new_n5434__ = ~new_new_n772__ & ~new_new_n995__;
  assign new_new_n5435__ = new_new_n5433__ & new_new_n5434__;
  assign new_new_n5436__ = ~new_new_n588__ & ~new_new_n602__;
  assign new_new_n5437__ = ~new_new_n842__ & ~new_new_n993__;
  assign new_new_n5438__ = new_new_n2078__ & ~new_new_n2329__;
  assign new_new_n5439__ = new_new_n5430__ & new_new_n5438__;
  assign new_new_n5440__ = new_new_n5436__ & new_new_n5437__;
  assign new_new_n5441__ = new_new_n381__ & new_new_n5435__;
  assign new_new_n5442__ = new_new_n674__ & new_new_n5431__;
  assign new_new_n5443__ = new_new_n5441__ & new_new_n5442__;
  assign new_new_n5444__ = new_new_n5439__ & new_new_n5440__;
  assign new_new_n5445__ = new_new_n440__ & new_new_n5432__;
  assign new_new_n5446__ = new_new_n5444__ & new_new_n5445__;
  assign new_new_n5447__ = new_new_n5443__ & new_new_n5446__;
  assign new_new_n5448__ = new_new_n5364__ & new_new_n5447__;
  assign new_new_n5449__ = new_new_n5377__ & new_new_n5448__;
  assign new_new_n5450__ = new_new_n5410__ & new_new_n5429__;
  assign new_new_n5451__ = new_new_n5449__ & new_new_n5450__;
  assign new_new_n5452__ = ~new_new_n5357__ & ~new_new_n5451__;
  assign new_new_n5453__ = ~new_new_n5356__ & ~new_new_n5452__;
  assign new_new_n5454__ = ~new_new_n5281__ & ~new_new_n5453__;
  assign new_new_n5455__ = new_new_n5281__ & new_new_n5453__;
  assign new_new_n5456__ = ~new_new_n5454__ & ~new_new_n5455__;
  assign new_new_n5457__ = ~new_new_n317__ & ~new_new_n842__;
  assign new_new_n5458__ = ~new_new_n477__ & ~new_new_n871__;
  assign new_new_n5459__ = ~new_new_n168__ & ~new_new_n772__;
  assign new_new_n5460__ = ~new_new_n130__ & ~new_new_n259__;
  assign new_new_n5461__ = ~new_new_n309__ & ~new_new_n1070__;
  assign new_new_n5462__ = new_new_n5460__ & new_new_n5461__;
  assign new_new_n5463__ = ~new_new_n263__ & new_new_n1960__;
  assign new_new_n5464__ = ~new_new_n5325__ & new_new_n5459__;
  assign new_new_n5465__ = new_new_n5463__ & new_new_n5464__;
  assign new_new_n5466__ = new_new_n744__ & new_new_n5462__;
  assign new_new_n5467__ = new_new_n5457__ & new_new_n5458__;
  assign new_new_n5468__ = new_new_n5466__ & new_new_n5467__;
  assign new_new_n5469__ = new_new_n891__ & new_new_n5465__;
  assign new_new_n5470__ = new_new_n1369__ & new_new_n5469__;
  assign new_new_n5471__ = new_new_n2584__ & new_new_n5468__;
  assign new_new_n5472__ = new_new_n5470__ & new_new_n5471__;
  assign new_new_n5473__ = ~new_new_n82__ & ~new_new_n482__;
  assign new_new_n5474__ = ~new_new_n277__ & ~new_new_n439__;
  assign new_new_n5475__ = ~new_new_n283__ & ~new_new_n603__;
  assign new_new_n5476__ = ~new_new_n657__ & new_new_n5475__;
  assign new_new_n5477__ = ~new_new_n148__ & new_new_n3184__;
  assign new_new_n5478__ = new_new_n3418__ & new_new_n5473__;
  assign new_new_n5479__ = new_new_n5477__ & new_new_n5478__;
  assign new_new_n5480__ = new_new_n167__ & new_new_n5476__;
  assign new_new_n5481__ = new_new_n2505__ & new_new_n5480__;
  assign new_new_n5482__ = new_new_n1267__ & new_new_n5479__;
  assign new_new_n5483__ = new_new_n1662__ & new_new_n2989__;
  assign new_new_n5484__ = new_new_n5474__ & new_new_n5483__;
  assign new_new_n5485__ = new_new_n5481__ & new_new_n5482__;
  assign new_new_n5486__ = new_new_n2973__ & new_new_n3374__;
  assign new_new_n5487__ = new_new_n5485__ & new_new_n5486__;
  assign new_new_n5488__ = new_new_n5388__ & new_new_n5484__;
  assign new_new_n5489__ = new_new_n5487__ & new_new_n5488__;
  assign new_new_n5490__ = new_new_n5472__ & new_new_n5489__;
  assign new_new_n5491__ = new_new_n4107__ & new_new_n5490__;
  assign new_new_n5492__ = ~new_new_n5456__ & new_new_n5491__;
  assign new_new_n5493__ = new_new_n5456__ & ~new_new_n5491__;
  assign new_new_n5494__ = ~new_new_n5492__ & ~new_new_n5493__;
  assign new_new_n5495__ = new_new_n3479__ & ~new_new_n3535__;
  assign new_new_n5496__ = ~new_new_n3479__ & new_new_n3535__;
  assign new_new_n5497__ = ~new_new_n5495__ & ~new_new_n5496__;
  assign new_new_n5498__ = new_new_n2130__ & ~new_new_n3479__;
  assign new_new_n5499__ = ~new_new_n2130__ & ~new_new_n2423__;
  assign new_new_n5500__ = ~new_new_n5498__ & ~new_new_n5499__;
  assign new_new_n5501__ = new_new_n5497__ & ~new_new_n5500__;
  assign new_new_n5502__ = new_new_n1902__ & new_new_n5501__;
  assign new_new_n5503__ = ~pi30 & ~new_new_n5502__;
  assign new_new_n5504__ = new_new_n3535__ & ~new_new_n5503__;
  assign new_new_n5505__ = new_new_n3535__ & ~new_new_n5501__;
  assign new_new_n5506__ = ~pi30 & new_new_n1902__;
  assign new_new_n5507__ = ~new_new_n5505__ & ~new_new_n5506__;
  assign new_new_n5508__ = ~new_new_n1823__ & ~new_new_n3537__;
  assign new_new_n5509__ = ~new_new_n5507__ & new_new_n5508__;
  assign new_new_n5510__ = ~new_new_n5504__ & ~new_new_n5509__;
  assign new_new_n5511__ = pi29 & ~new_new_n5510__;
  assign new_new_n5512__ = ~new_new_n1902__ & ~new_new_n5501__;
  assign new_new_n5513__ = ~new_new_n5502__ & ~new_new_n5512__;
  assign new_new_n5514__ = ~new_new_n161__ & ~new_new_n5505__;
  assign new_new_n5515__ = ~new_new_n5513__ & new_new_n5514__;
  assign new_new_n5516__ = ~new_new_n71__ & ~new_new_n3537__;
  assign new_new_n5517__ = ~new_new_n5515__ & new_new_n5516__;
  assign new_new_n5518__ = new_new_n1823__ & ~new_new_n5517__;
  assign new_new_n5519__ = new_new_n5250__ & new_new_n5268__;
  assign new_new_n5520__ = new_new_n1823__ & ~new_new_n5501__;
  assign new_new_n5521__ = new_new_n3535__ & ~new_new_n5520__;
  assign new_new_n5522__ = ~new_new_n5513__ & new_new_n5521__;
  assign new_new_n5523__ = ~new_new_n5519__ & ~new_new_n5522__;
  assign new_new_n5524__ = pi30 & ~new_new_n5523__;
  assign new_new_n5525__ = pi31 & ~new_new_n5511__;
  assign new_new_n5526__ = ~new_new_n5518__ & ~new_new_n5524__;
  assign new_new_n5527__ = new_new_n5525__ & new_new_n5526__;
  assign new_new_n5528__ = ~new_new_n71__ & ~new_new_n1902__;
  assign new_new_n5529__ = ~new_new_n161__ & ~new_new_n5528__;
  assign new_new_n5530__ = ~pi31 & ~new_new_n5277__;
  assign new_new_n5531__ = ~new_new_n5529__ & new_new_n5530__;
  assign new_new_n5532__ = ~new_new_n5527__ & ~new_new_n5531__;
  assign new_new_n5533__ = ~new_new_n3535__ & ~new_new_n5276__;
  assign new_new_n5534__ = pi30 & ~new_new_n5495__;
  assign new_new_n5535__ = ~new_new_n5533__ & ~new_new_n5534__;
  assign new_new_n5536__ = ~new_new_n1823__ & new_new_n3535__;
  assign new_new_n5537__ = new_new_n3479__ & ~new_new_n5536__;
  assign new_new_n5538__ = ~new_new_n3479__ & ~new_new_n5276__;
  assign new_new_n5539__ = ~new_new_n2130__ & ~new_new_n5537__;
  assign new_new_n5540__ = ~new_new_n5538__ & new_new_n5539__;
  assign new_new_n5541__ = ~new_new_n5535__ & ~new_new_n5540__;
  assign new_new_n5542__ = ~pi29 & ~new_new_n5541__;
  assign new_new_n5543__ = new_new_n1823__ & new_new_n3535__;
  assign new_new_n5544__ = ~new_new_n71__ & new_new_n5268__;
  assign new_new_n5545__ = ~new_new_n3479__ & new_new_n5544__;
  assign new_new_n5546__ = ~new_new_n161__ & ~new_new_n5543__;
  assign new_new_n5547__ = ~new_new_n5545__ & new_new_n5546__;
  assign new_new_n5548__ = new_new_n2130__ & ~new_new_n5547__;
  assign new_new_n5549__ = ~new_new_n3479__ & ~new_new_n5543__;
  assign new_new_n5550__ = ~new_new_n2130__ & new_new_n5536__;
  assign new_new_n5551__ = pi29 & new_new_n5253__;
  assign new_new_n5552__ = ~new_new_n5550__ & ~new_new_n5551__;
  assign new_new_n5553__ = new_new_n3479__ & new_new_n5552__;
  assign new_new_n5554__ = ~pi30 & ~new_new_n5549__;
  assign new_new_n5555__ = ~new_new_n5553__ & new_new_n5554__;
  assign new_new_n5556__ = pi31 & ~new_new_n5548__;
  assign new_new_n5557__ = ~new_new_n5555__ & new_new_n5556__;
  assign new_new_n5558__ = ~new_new_n5542__ & new_new_n5557__;
  assign new_new_n5559__ = new_new_n765__ & ~new_new_n1823__;
  assign new_new_n5560__ = new_new_n161__ & ~new_new_n3535__;
  assign new_new_n5561__ = ~new_new_n5559__ & ~new_new_n5560__;
  assign new_new_n5562__ = ~pi31 & ~new_new_n5561__;
  assign new_new_n5563__ = ~new_new_n5558__ & ~new_new_n5562__;
  assign new_new_n5564__ = ~new_new_n183__ & new_new_n1509__;
  assign new_new_n5565__ = new_new_n936__ & new_new_n5564__;
  assign new_new_n5566__ = ~new_new_n270__ & ~new_new_n1151__;
  assign new_new_n5567__ = ~new_new_n277__ & ~new_new_n1109__;
  assign new_new_n5568__ = ~new_new_n496__ & ~new_new_n607__;
  assign new_new_n5569__ = new_new_n5567__ & new_new_n5568__;
  assign new_new_n5570__ = ~new_new_n160__ & ~new_new_n335__;
  assign new_new_n5571__ = new_new_n386__ & new_new_n5570__;
  assign new_new_n5572__ = ~new_new_n871__ & ~new_new_n993__;
  assign new_new_n5573__ = ~new_new_n1035__ & new_new_n3430__;
  assign new_new_n5574__ = new_new_n4465__ & new_new_n5573__;
  assign new_new_n5575__ = new_new_n5571__ & new_new_n5572__;
  assign new_new_n5576__ = ~new_new_n316__ & new_new_n2131__;
  assign new_new_n5577__ = new_new_n5566__ & new_new_n5576__;
  assign new_new_n5578__ = new_new_n5574__ & new_new_n5575__;
  assign new_new_n5579__ = new_new_n1704__ & new_new_n2764__;
  assign new_new_n5580__ = new_new_n5578__ & new_new_n5579__;
  assign new_new_n5581__ = new_new_n5565__ & new_new_n5577__;
  assign new_new_n5582__ = new_new_n5569__ & new_new_n5581__;
  assign new_new_n5583__ = new_new_n3563__ & new_new_n5580__;
  assign new_new_n5584__ = new_new_n5582__ & new_new_n5583__;
  assign new_new_n5585__ = ~new_new_n252__ & ~new_new_n597__;
  assign new_new_n5586__ = ~new_new_n1372__ & new_new_n5585__;
  assign new_new_n5587__ = ~new_new_n382__ & new_new_n5586__;
  assign new_new_n5588__ = new_new_n1340__ & new_new_n1471__;
  assign new_new_n5589__ = new_new_n5587__ & new_new_n5588__;
  assign new_new_n5590__ = new_new_n153__ & ~new_new_n1129__;
  assign new_new_n5591__ = ~new_new_n896__ & ~new_new_n995__;
  assign new_new_n5592__ = ~new_new_n842__ & new_new_n5591__;
  assign new_new_n5593__ = new_new_n2619__ & new_new_n5592__;
  assign new_new_n5594__ = ~new_new_n96__ & ~new_new_n196__;
  assign new_new_n5595__ = ~new_new_n656__ & ~new_new_n723__;
  assign new_new_n5596__ = new_new_n5594__ & new_new_n5595__;
  assign new_new_n5597__ = ~new_new_n1008__ & new_new_n2479__;
  assign new_new_n5598__ = ~new_new_n5590__ & new_new_n5597__;
  assign new_new_n5599__ = new_new_n1705__ & new_new_n5596__;
  assign new_new_n5600__ = new_new_n3893__ & new_new_n3989__;
  assign new_new_n5601__ = new_new_n5599__ & new_new_n5600__;
  assign new_new_n5602__ = new_new_n1001__ & new_new_n5598__;
  assign new_new_n5603__ = new_new_n2031__ & new_new_n4388__;
  assign new_new_n5604__ = new_new_n5593__ & new_new_n5603__;
  assign new_new_n5605__ = new_new_n5601__ & new_new_n5602__;
  assign new_new_n5606__ = new_new_n4726__ & new_new_n5605__;
  assign new_new_n5607__ = new_new_n5604__ & new_new_n5606__;
  assign new_new_n5608__ = ~new_new_n816__ & new_new_n5607__;
  assign new_new_n5609__ = ~new_new_n600__ & ~new_new_n768__;
  assign new_new_n5610__ = ~new_new_n202__ & new_new_n5609__;
  assign new_new_n5611__ = ~new_new_n1167__ & new_new_n5610__;
  assign new_new_n5612__ = ~new_new_n254__ & new_new_n5611__;
  assign new_new_n5613__ = ~new_new_n120__ & ~new_new_n511__;
  assign new_new_n5614__ = ~new_new_n694__ & ~new_new_n1176__;
  assign new_new_n5615__ = new_new_n5613__ & new_new_n5614__;
  assign new_new_n5616__ = ~new_new_n1166__ & new_new_n3415__;
  assign new_new_n5617__ = new_new_n5615__ & new_new_n5616__;
  assign new_new_n5618__ = ~new_new_n115__ & ~new_new_n439__;
  assign new_new_n5619__ = ~new_new_n809__ & new_new_n5618__;
  assign new_new_n5620__ = new_new_n3023__ & new_new_n5617__;
  assign new_new_n5621__ = new_new_n5619__ & new_new_n5620__;
  assign new_new_n5622__ = new_new_n5612__ & new_new_n5621__;
  assign new_new_n5623__ = new_new_n1154__ & ~new_new_n1217__;
  assign new_new_n5624__ = ~new_new_n138__ & ~new_new_n247__;
  assign new_new_n5625__ = ~new_new_n843__ & ~new_new_n963__;
  assign new_new_n5626__ = new_new_n5624__ & new_new_n5625__;
  assign new_new_n5627__ = ~new_new_n329__ & ~new_new_n675__;
  assign new_new_n5628__ = new_new_n2160__ & new_new_n2873__;
  assign new_new_n5629__ = new_new_n5626__ & new_new_n5627__;
  assign new_new_n5630__ = new_new_n1063__ & new_new_n1153__;
  assign new_new_n5631__ = new_new_n5623__ & new_new_n5630__;
  assign new_new_n5632__ = new_new_n5628__ & new_new_n5629__;
  assign new_new_n5633__ = new_new_n5631__ & new_new_n5632__;
  assign new_new_n5634__ = new_new_n841__ & new_new_n5589__;
  assign new_new_n5635__ = new_new_n5633__ & new_new_n5634__;
  assign new_new_n5636__ = new_new_n5622__ & new_new_n5635__;
  assign new_new_n5637__ = new_new_n5584__ & new_new_n5636__;
  assign new_new_n5638__ = new_new_n5608__ & new_new_n5637__;
  assign new_new_n5639__ = ~new_new_n5563__ & ~new_new_n5638__;
  assign new_new_n5640__ = ~new_new_n5356__ & ~new_new_n5357__;
  assign new_new_n5641__ = new_new_n5563__ & new_new_n5638__;
  assign new_new_n5642__ = ~new_new_n5640__ & new_new_n5641__;
  assign new_new_n5643__ = new_new_n5451__ & ~new_new_n5642__;
  assign new_new_n5644__ = ~new_new_n5639__ & ~new_new_n5643__;
  assign new_new_n5645__ = ~new_new_n5532__ & ~new_new_n5644__;
  assign new_new_n5646__ = new_new_n5640__ & ~new_new_n5641__;
  assign new_new_n5647__ = new_new_n5643__ & new_new_n5646__;
  assign new_new_n5648__ = new_new_n5532__ & ~new_new_n5639__;
  assign new_new_n5649__ = ~new_new_n5451__ & ~new_new_n5640__;
  assign new_new_n5650__ = ~new_new_n5648__ & new_new_n5649__;
  assign new_new_n5651__ = ~new_new_n5645__ & ~new_new_n5647__;
  assign new_new_n5652__ = ~new_new_n5650__ & new_new_n5651__;
  assign new_new_n5653__ = new_new_n5494__ & new_new_n5652__;
  assign new_new_n5654__ = ~new_new_n5494__ & ~new_new_n5652__;
  assign new_new_n5655__ = ~new_new_n1556__ & new_new_n4815__;
  assign new_new_n5656__ = ~new_new_n1737__ & ~new_new_n4818__;
  assign new_new_n5657__ = ~new_new_n1466__ & new_new_n4212__;
  assign new_new_n5658__ = ~new_new_n1660__ & ~new_new_n1737__;
  assign new_new_n5659__ = new_new_n1660__ & new_new_n1737__;
  assign new_new_n5660__ = ~new_new_n5658__ & ~new_new_n5659__;
  assign new_new_n5661__ = new_new_n1737__ & new_new_n3544__;
  assign new_new_n5662__ = ~new_new_n1737__ & ~new_new_n3544__;
  assign new_new_n5663__ = ~new_new_n5661__ & ~new_new_n5662__;
  assign new_new_n5664__ = new_new_n5660__ & ~new_new_n5663__;
  assign new_new_n5665__ = new_new_n1466__ & new_new_n5664__;
  assign new_new_n5666__ = new_new_n3544__ & new_new_n5660__;
  assign new_new_n5667__ = new_new_n1737__ & ~new_new_n5666__;
  assign new_new_n5668__ = ~new_new_n5665__ & ~new_new_n5667__;
  assign new_new_n5669__ = new_new_n5026__ & new_new_n5668__;
  assign new_new_n5670__ = ~new_new_n5026__ & ~new_new_n5668__;
  assign new_new_n5671__ = ~new_new_n5669__ & ~new_new_n5670__;
  assign new_new_n5672__ = new_new_n4813__ & ~new_new_n5671__;
  assign new_new_n5673__ = ~new_new_n5655__ & ~new_new_n5656__;
  assign new_new_n5674__ = ~new_new_n5657__ & new_new_n5673__;
  assign new_new_n5675__ = ~new_new_n5672__ & new_new_n5674__;
  assign new_new_n5676__ = pi29 & ~new_new_n5675__;
  assign new_new_n5677__ = ~pi29 & new_new_n5675__;
  assign new_new_n5678__ = ~new_new_n5676__ & ~new_new_n5677__;
  assign new_new_n5679__ = ~new_new_n5654__ & ~new_new_n5678__;
  assign new_new_n5680__ = ~new_new_n5653__ & ~new_new_n5679__;
  assign new_new_n5681__ = ~new_new_n5245__ & ~new_new_n5680__;
  assign new_new_n5682__ = new_new_n5245__ & new_new_n5680__;
  assign new_new_n5683__ = new_new_n161__ & ~new_new_n1660__;
  assign new_new_n5684__ = new_new_n765__ & ~new_new_n1737__;
  assign new_new_n5685__ = ~new_new_n5683__ & ~new_new_n5684__;
  assign new_new_n5686__ = ~pi31 & ~new_new_n5685__;
  assign new_new_n5687__ = ~new_new_n3544__ & ~new_new_n5660__;
  assign new_new_n5688__ = ~new_new_n5666__ & ~new_new_n5687__;
  assign new_new_n5689__ = new_new_n765__ & new_new_n5688__;
  assign new_new_n5690__ = new_new_n71__ & ~new_new_n1660__;
  assign new_new_n5691__ = ~new_new_n5247__ & ~new_new_n5690__;
  assign new_new_n5692__ = ~new_new_n5689__ & new_new_n5691__;
  assign new_new_n5693__ = pi31 & ~new_new_n5692__;
  assign new_new_n5694__ = ~new_new_n5686__ & ~new_new_n5693__;
  assign new_new_n5695__ = ~new_new_n353__ & ~new_new_n781__;
  assign new_new_n5696__ = ~new_new_n884__ & new_new_n5695__;
  assign new_new_n5697__ = ~new_new_n652__ & new_new_n5696__;
  assign new_new_n5698__ = ~new_new_n747__ & ~new_new_n851__;
  assign new_new_n5699__ = ~new_new_n383__ & ~new_new_n656__;
  assign new_new_n5700__ = new_new_n239__ & ~new_new_n276__;
  assign new_new_n5701__ = ~new_new_n1003__ & new_new_n1263__;
  assign new_new_n5702__ = new_new_n1711__ & new_new_n2340__;
  assign new_new_n5703__ = new_new_n2404__ & new_new_n5699__;
  assign new_new_n5704__ = new_new_n5702__ & new_new_n5703__;
  assign new_new_n5705__ = new_new_n5700__ & new_new_n5701__;
  assign new_new_n5706__ = new_new_n5458__ & new_new_n5566__;
  assign new_new_n5707__ = new_new_n5698__ & new_new_n5706__;
  assign new_new_n5708__ = new_new_n5704__ & new_new_n5705__;
  assign new_new_n5709__ = new_new_n932__ & new_new_n5708__;
  assign new_new_n5710__ = new_new_n5697__ & new_new_n5707__;
  assign new_new_n5711__ = new_new_n5709__ & new_new_n5710__;
  assign new_new_n5712__ = new_new_n2777__ & new_new_n5711__;
  assign new_new_n5713__ = new_new_n621__ & new_new_n3089__;
  assign new_new_n5714__ = new_new_n5712__ & new_new_n5713__;
  assign new_new_n5715__ = new_new_n3662__ & new_new_n5714__;
  assign new_new_n5716__ = new_new_n5455__ & new_new_n5491__;
  assign new_new_n5717__ = new_new_n5454__ & ~new_new_n5491__;
  assign new_new_n5718__ = ~new_new_n5716__ & ~new_new_n5717__;
  assign new_new_n5719__ = new_new_n5715__ & ~new_new_n5718__;
  assign new_new_n5720__ = ~new_new_n5715__ & new_new_n5718__;
  assign new_new_n5721__ = ~new_new_n5719__ & ~new_new_n5720__;
  assign new_new_n5722__ = ~new_new_n5694__ & ~new_new_n5721__;
  assign new_new_n5723__ = new_new_n5694__ & new_new_n5721__;
  assign new_new_n5724__ = ~new_new_n5722__ & ~new_new_n5723__;
  assign new_new_n5725__ = ~new_new_n1325__ & new_new_n4815__;
  assign new_new_n5726__ = ~new_new_n1466__ & ~new_new_n4818__;
  assign new_new_n5727__ = ~new_new_n1556__ & new_new_n4212__;
  assign new_new_n5728__ = ~new_new_n5725__ & ~new_new_n5726__;
  assign new_new_n5729__ = ~new_new_n5727__ & new_new_n5728__;
  assign new_new_n5730__ = new_new_n4214__ & new_new_n5048__;
  assign new_new_n5731__ = ~pi29 & ~new_new_n5730__;
  assign new_new_n5732__ = ~pi28 & new_new_n4214__;
  assign new_new_n5733__ = new_new_n5048__ & new_new_n5732__;
  assign new_new_n5734__ = ~new_new_n5731__ & ~new_new_n5733__;
  assign new_new_n5735__ = new_new_n5729__ & ~new_new_n5734__;
  assign new_new_n5736__ = pi29 & ~new_new_n5729__;
  assign new_new_n5737__ = ~new_new_n5735__ & ~new_new_n5736__;
  assign new_new_n5738__ = ~new_new_n5724__ & new_new_n5737__;
  assign new_new_n5739__ = new_new_n5724__ & ~new_new_n5737__;
  assign new_new_n5740__ = ~new_new_n5738__ & ~new_new_n5739__;
  assign new_new_n5741__ = ~new_new_n5682__ & new_new_n5740__;
  assign new_new_n5742__ = ~new_new_n5681__ & ~new_new_n5741__;
  assign new_new_n5743__ = ~new_new_n1325__ & new_new_n4212__;
  assign new_new_n5744__ = ~new_new_n1556__ & ~new_new_n4818__;
  assign new_new_n5745__ = ~new_new_n5743__ & ~new_new_n5744__;
  assign new_new_n5746__ = new_new_n3618__ & ~new_new_n4921__;
  assign new_new_n5747__ = new_new_n4214__ & ~new_new_n5746__;
  assign new_new_n5748__ = pi29 & ~new_new_n5747__;
  assign new_new_n5749__ = ~pi28 & new_new_n3618__;
  assign new_new_n5750__ = pi28 & ~new_new_n3618__;
  assign new_new_n5751__ = new_new_n4214__ & ~new_new_n5749__;
  assign new_new_n5752__ = ~new_new_n5750__ & new_new_n5751__;
  assign new_new_n5753__ = new_new_n4921__ & new_new_n5752__;
  assign new_new_n5754__ = ~new_new_n5748__ & ~new_new_n5753__;
  assign new_new_n5755__ = new_new_n5745__ & ~new_new_n5754__;
  assign new_new_n5756__ = ~new_new_n3618__ & ~new_new_n4921__;
  assign new_new_n5757__ = new_new_n4214__ & new_new_n5756__;
  assign new_new_n5758__ = new_new_n5745__ & ~new_new_n5757__;
  assign new_new_n5759__ = ~pi29 & ~new_new_n5758__;
  assign new_new_n5760__ = ~new_new_n5755__ & ~new_new_n5759__;
  assign new_new_n5761__ = ~new_new_n5491__ & ~new_new_n5715__;
  assign new_new_n5762__ = ~new_new_n5455__ & ~new_new_n5761__;
  assign new_new_n5763__ = new_new_n161__ & ~new_new_n1737__;
  assign new_new_n5764__ = new_new_n765__ & ~new_new_n1466__;
  assign new_new_n5765__ = ~new_new_n5763__ & ~new_new_n5764__;
  assign new_new_n5766__ = ~pi31 & ~new_new_n5765__;
  assign new_new_n5767__ = new_new_n71__ & new_new_n1737__;
  assign new_new_n5768__ = new_new_n1466__ & new_new_n3544__;
  assign new_new_n5769__ = ~new_new_n1737__ & new_new_n5768__;
  assign new_new_n5770__ = ~new_new_n1466__ & ~new_new_n5661__;
  assign new_new_n5771__ = ~new_new_n1660__ & ~new_new_n5768__;
  assign new_new_n5772__ = ~new_new_n5770__ & new_new_n5771__;
  assign new_new_n5773__ = ~new_new_n5769__ & ~new_new_n5772__;
  assign new_new_n5774__ = ~new_new_n161__ & ~new_new_n5773__;
  assign new_new_n5775__ = ~new_new_n1466__ & new_new_n5662__;
  assign new_new_n5776__ = new_new_n1466__ & new_new_n1737__;
  assign new_new_n5777__ = ~new_new_n161__ & ~new_new_n5776__;
  assign new_new_n5778__ = ~new_new_n5775__ & new_new_n5777__;
  assign new_new_n5779__ = new_new_n1660__ & ~new_new_n5778__;
  assign new_new_n5780__ = ~new_new_n5774__ & ~new_new_n5779__;
  assign new_new_n5781__ = ~new_new_n71__ & ~new_new_n5780__;
  assign new_new_n5782__ = pi31 & ~new_new_n5767__;
  assign new_new_n5783__ = ~new_new_n5781__ & new_new_n5782__;
  assign new_new_n5784__ = ~new_new_n5766__ & ~new_new_n5783__;
  assign new_new_n5785__ = ~new_new_n150__ & ~new_new_n382__;
  assign new_new_n5786__ = ~pi23 & ~new_new_n162__;
  assign new_new_n5787__ = pi23 & ~new_new_n85__;
  assign new_new_n5788__ = ~new_new_n333__ & ~new_new_n5786__;
  assign new_new_n5789__ = ~new_new_n5787__ & new_new_n5788__;
  assign new_new_n5790__ = ~new_new_n719__ & ~new_new_n875__;
  assign new_new_n5791__ = ~new_new_n5789__ & new_new_n5790__;
  assign new_new_n5792__ = ~new_new_n108__ & ~new_new_n388__;
  assign new_new_n5793__ = ~new_new_n1151__ & new_new_n5792__;
  assign new_new_n5794__ = new_new_n481__ & new_new_n5793__;
  assign new_new_n5795__ = new_new_n1850__ & new_new_n5794__;
  assign new_new_n5796__ = ~new_new_n284__ & ~new_new_n312__;
  assign new_new_n5797__ = ~new_new_n313__ & ~new_new_n671__;
  assign new_new_n5798__ = ~new_new_n783__ & new_new_n5797__;
  assign new_new_n5799__ = ~new_new_n286__ & new_new_n5796__;
  assign new_new_n5800__ = ~new_new_n842__ & new_new_n1740__;
  assign new_new_n5801__ = new_new_n5799__ & new_new_n5800__;
  assign new_new_n5802__ = new_new_n1499__ & new_new_n5798__;
  assign new_new_n5803__ = new_new_n1645__ & new_new_n1828__;
  assign new_new_n5804__ = new_new_n2316__ & new_new_n3363__;
  assign new_new_n5805__ = new_new_n5785__ & new_new_n5804__;
  assign new_new_n5806__ = new_new_n5802__ & new_new_n5803__;
  assign new_new_n5807__ = new_new_n2700__ & new_new_n5801__;
  assign new_new_n5808__ = new_new_n5791__ & new_new_n5807__;
  assign new_new_n5809__ = new_new_n5805__ & new_new_n5806__;
  assign new_new_n5810__ = new_new_n4234__ & new_new_n5809__;
  assign new_new_n5811__ = new_new_n5795__ & new_new_n5808__;
  assign new_new_n5812__ = new_new_n5810__ & new_new_n5811__;
  assign new_new_n5813__ = ~new_new_n383__ & ~new_new_n482__;
  assign new_new_n5814__ = ~new_new_n277__ & new_new_n5813__;
  assign new_new_n5815__ = ~new_new_n721__ & new_new_n5814__;
  assign new_new_n5816__ = new_new_n118__ & ~new_new_n1880__;
  assign new_new_n5817__ = ~new_new_n947__ & ~new_new_n1291__;
  assign new_new_n5818__ = ~new_new_n207__ & ~new_new_n700__;
  assign new_new_n5819__ = ~new_new_n890__ & new_new_n5818__;
  assign new_new_n5820__ = ~new_new_n189__ & ~new_new_n1003__;
  assign new_new_n5821__ = new_new_n1366__ & ~new_new_n1632__;
  assign new_new_n5822__ = ~new_new_n5816__ & new_new_n5817__;
  assign new_new_n5823__ = new_new_n5821__ & new_new_n5822__;
  assign new_new_n5824__ = new_new_n5819__ & new_new_n5820__;
  assign new_new_n5825__ = ~new_new_n218__ & ~new_new_n546__;
  assign new_new_n5826__ = new_new_n1707__ & new_new_n1971__;
  assign new_new_n5827__ = new_new_n5314__ & new_new_n5826__;
  assign new_new_n5828__ = new_new_n5824__ & new_new_n5825__;
  assign new_new_n5829__ = new_new_n985__ & new_new_n5823__;
  assign new_new_n5830__ = new_new_n5815__ & new_new_n5829__;
  assign new_new_n5831__ = new_new_n5827__ & new_new_n5828__;
  assign new_new_n5832__ = new_new_n5830__ & new_new_n5831__;
  assign new_new_n5833__ = new_new_n5812__ & new_new_n5832__;
  assign new_new_n5834__ = new_new_n1141__ & new_new_n5833__;
  assign new_new_n5835__ = new_new_n3102__ & new_new_n5834__;
  assign new_new_n5836__ = ~pi17 & ~new_new_n5835__;
  assign new_new_n5837__ = pi17 & new_new_n5834__;
  assign new_new_n5838__ = new_new_n3102__ & new_new_n5837__;
  assign new_new_n5839__ = ~new_new_n5836__ & ~new_new_n5838__;
  assign new_new_n5840__ = new_new_n5784__ & ~new_new_n5839__;
  assign new_new_n5841__ = ~new_new_n5784__ & new_new_n5839__;
  assign new_new_n5842__ = ~new_new_n5840__ & ~new_new_n5841__;
  assign new_new_n5843__ = new_new_n5491__ & new_new_n5715__;
  assign new_new_n5844__ = ~new_new_n5454__ & ~new_new_n5843__;
  assign new_new_n5845__ = ~new_new_n5762__ & ~new_new_n5844__;
  assign new_new_n5846__ = new_new_n5842__ & new_new_n5845__;
  assign new_new_n5847__ = ~new_new_n5715__ & new_new_n5717__;
  assign new_new_n5848__ = new_new_n5455__ & new_new_n5843__;
  assign new_new_n5849__ = ~new_new_n5847__ & ~new_new_n5848__;
  assign new_new_n5850__ = ~new_new_n5842__ & new_new_n5849__;
  assign new_new_n5851__ = ~new_new_n5846__ & ~new_new_n5850__;
  assign new_new_n5852__ = new_new_n5760__ & new_new_n5851__;
  assign new_new_n5853__ = ~new_new_n5760__ & ~new_new_n5851__;
  assign new_new_n5854__ = ~new_new_n5852__ & ~new_new_n5853__;
  assign new_new_n5855__ = ~new_new_n5723__ & new_new_n5737__;
  assign new_new_n5856__ = ~new_new_n5722__ & ~new_new_n5855__;
  assign new_new_n5857__ = new_new_n5854__ & ~new_new_n5856__;
  assign new_new_n5858__ = ~new_new_n5854__ & new_new_n5856__;
  assign new_new_n5859__ = ~new_new_n5857__ & ~new_new_n5858__;
  assign new_new_n5860__ = ~new_new_n5742__ & ~new_new_n5859__;
  assign new_new_n5861__ = ~new_new_n4550__ & ~new_new_n4900__;
  assign new_new_n5862__ = ~new_new_n868__ & new_new_n3311__;
  assign new_new_n5863__ = ~new_new_n333__ & ~new_new_n1061__;
  assign new_new_n5864__ = new_new_n873__ & ~new_new_n1207__;
  assign new_new_n5865__ = ~new_new_n5862__ & ~new_new_n5863__;
  assign new_new_n5866__ = ~new_new_n5864__ & new_new_n5865__;
  assign new_new_n5867__ = ~new_new_n5861__ & new_new_n5866__;
  assign new_new_n5868__ = pi26 & ~new_new_n5867__;
  assign new_new_n5869__ = ~pi26 & new_new_n5867__;
  assign new_new_n5870__ = ~new_new_n5868__ & ~new_new_n5869__;
  assign new_new_n5871__ = new_new_n5742__ & new_new_n5859__;
  assign new_new_n5872__ = ~new_new_n5870__ & ~new_new_n5871__;
  assign new_new_n5873__ = ~new_new_n5860__ & ~new_new_n5872__;
  assign new_new_n5874__ = new_new_n1466__ & ~new_new_n5664__;
  assign new_new_n5875__ = ~new_new_n1466__ & new_new_n5664__;
  assign new_new_n5876__ = new_new_n1737__ & ~new_new_n5875__;
  assign new_new_n5877__ = new_new_n765__ & ~new_new_n5874__;
  assign new_new_n5878__ = ~new_new_n5876__ & new_new_n5877__;
  assign new_new_n5879__ = ~new_new_n5776__ & ~new_new_n5878__;
  assign new_new_n5880__ = new_new_n1556__ & ~new_new_n5879__;
  assign new_new_n5881__ = ~new_new_n1466__ & ~new_new_n5664__;
  assign new_new_n5882__ = ~new_new_n1556__ & new_new_n5881__;
  assign new_new_n5883__ = ~new_new_n161__ & ~new_new_n5882__;
  assign new_new_n5884__ = ~new_new_n71__ & new_new_n1737__;
  assign new_new_n5885__ = ~new_new_n5883__ & new_new_n5884__;
  assign new_new_n5886__ = new_new_n1738__ & ~new_new_n5664__;
  assign new_new_n5887__ = ~new_new_n71__ & ~new_new_n5886__;
  assign new_new_n5888__ = ~new_new_n161__ & new_new_n1466__;
  assign new_new_n5889__ = ~new_new_n5887__ & new_new_n5888__;
  assign new_new_n5890__ = pi31 & ~new_new_n5889__;
  assign new_new_n5891__ = ~new_new_n5885__ & new_new_n5890__;
  assign new_new_n5892__ = ~new_new_n5880__ & new_new_n5891__;
  assign new_new_n5893__ = new_new_n765__ & ~new_new_n1556__;
  assign new_new_n5894__ = ~new_new_n5023__ & ~new_new_n5893__;
  assign new_new_n5895__ = ~pi31 & ~new_new_n5894__;
  assign new_new_n5896__ = ~new_new_n5892__ & ~new_new_n5895__;
  assign new_new_n5897__ = ~new_new_n3618__ & new_new_n4212__;
  assign new_new_n5898__ = ~new_new_n1061__ & new_new_n4815__;
  assign new_new_n5899__ = ~new_new_n1325__ & ~new_new_n4818__;
  assign new_new_n5900__ = ~new_new_n5897__ & ~new_new_n5898__;
  assign new_new_n5901__ = ~new_new_n5899__ & new_new_n5900__;
  assign new_new_n5902__ = new_new_n4214__ & new_new_n4926__;
  assign new_new_n5903__ = ~pi29 & ~new_new_n5902__;
  assign new_new_n5904__ = new_new_n4926__ & new_new_n5732__;
  assign new_new_n5905__ = ~new_new_n5903__ & ~new_new_n5904__;
  assign new_new_n5906__ = new_new_n5901__ & ~new_new_n5905__;
  assign new_new_n5907__ = pi29 & ~new_new_n5901__;
  assign new_new_n5908__ = ~new_new_n5906__ & ~new_new_n5907__;
  assign new_new_n5909__ = ~new_new_n5896__ & new_new_n5908__;
  assign new_new_n5910__ = new_new_n5896__ & ~new_new_n5908__;
  assign new_new_n5911__ = ~new_new_n5909__ & ~new_new_n5910__;
  assign new_new_n5912__ = ~new_new_n5852__ & ~new_new_n5856__;
  assign new_new_n5913__ = ~new_new_n5853__ & ~new_new_n5912__;
  assign new_new_n5914__ = ~new_new_n333__ & ~new_new_n1207__;
  assign new_new_n5915__ = new_new_n3311__ & ~new_new_n3720__;
  assign new_new_n5916__ = ~new_new_n868__ & new_new_n873__;
  assign new_new_n5917__ = ~new_new_n5914__ & ~new_new_n5915__;
  assign new_new_n5918__ = ~new_new_n5916__ & new_new_n5917__;
  assign new_new_n5919__ = ~new_new_n4033__ & ~new_new_n5918__;
  assign new_new_n5920__ = ~new_new_n3622__ & new_new_n4035__;
  assign new_new_n5921__ = new_new_n3622__ & new_new_n4034__;
  assign new_new_n5922__ = ~new_new_n5920__ & ~new_new_n5921__;
  assign new_new_n5923__ = ~new_new_n4900__ & ~new_new_n5922__;
  assign new_new_n5924__ = ~new_new_n5919__ & ~new_new_n5923__;
  assign new_new_n5925__ = pi26 & ~new_new_n5924__;
  assign new_new_n5926__ = new_new_n3622__ & ~new_new_n4035__;
  assign new_new_n5927__ = ~new_new_n5920__ & ~new_new_n5926__;
  assign new_new_n5928__ = ~new_new_n4900__ & ~new_new_n5927__;
  assign new_new_n5929__ = ~pi26 & new_new_n5918__;
  assign new_new_n5930__ = ~new_new_n5928__ & new_new_n5929__;
  assign new_new_n5931__ = ~new_new_n5925__ & ~new_new_n5930__;
  assign new_new_n5932__ = ~new_new_n5784__ & ~new_new_n5848__;
  assign new_new_n5933__ = ~new_new_n5847__ & ~new_new_n5932__;
  assign new_new_n5934__ = ~new_new_n5839__ & ~new_new_n5933__;
  assign new_new_n5935__ = new_new_n5715__ & ~new_new_n5836__;
  assign new_new_n5936__ = ~new_new_n5838__ & new_new_n5935__;
  assign new_new_n5937__ = new_new_n5717__ & ~new_new_n5784__;
  assign new_new_n5938__ = ~new_new_n5936__ & ~new_new_n5937__;
  assign new_new_n5939__ = new_new_n5716__ & new_new_n5784__;
  assign new_new_n5940__ = ~new_new_n5938__ & ~new_new_n5939__;
  assign new_new_n5941__ = ~new_new_n5934__ & ~new_new_n5940__;
  assign new_new_n5942__ = ~new_new_n5837__ & ~new_new_n5935__;
  assign new_new_n5943__ = new_new_n4452__ & ~new_new_n5942__;
  assign new_new_n5944__ = ~new_new_n4452__ & new_new_n5942__;
  assign new_new_n5945__ = ~new_new_n5943__ & ~new_new_n5944__;
  assign new_new_n5946__ = new_new_n5941__ & ~new_new_n5945__;
  assign new_new_n5947__ = ~new_new_n5941__ & new_new_n5945__;
  assign new_new_n5948__ = ~new_new_n5946__ & ~new_new_n5947__;
  assign new_new_n5949__ = new_new_n5931__ & new_new_n5948__;
  assign new_new_n5950__ = ~new_new_n5931__ & ~new_new_n5948__;
  assign new_new_n5951__ = ~new_new_n5949__ & ~new_new_n5950__;
  assign new_new_n5952__ = new_new_n5913__ & ~new_new_n5951__;
  assign new_new_n5953__ = ~new_new_n5913__ & new_new_n5951__;
  assign new_new_n5954__ = ~new_new_n5952__ & ~new_new_n5953__;
  assign new_new_n5955__ = new_new_n5911__ & new_new_n5954__;
  assign new_new_n5956__ = ~new_new_n5911__ & ~new_new_n5954__;
  assign new_new_n5957__ = ~new_new_n5955__ & ~new_new_n5956__;
  assign new_new_n5958__ = ~new_new_n5873__ & new_new_n5957__;
  assign new_new_n5959__ = new_new_n5873__ & ~new_new_n5957__;
  assign new_new_n5960__ = ~new_new_n5958__ & ~new_new_n5959__;
  assign new_new_n5961__ = pi23 & ~new_new_n5960__;
  assign new_new_n5962__ = ~pi23 & new_new_n5960__;
  assign new_new_n5963__ = ~new_new_n5961__ & ~new_new_n5962__;
  assign new_new_n5964__ = new_new_n5219__ & new_new_n5963__;
  assign new_new_n5965__ = ~new_new_n5219__ & ~new_new_n5963__;
  assign new_new_n5966__ = ~new_new_n5964__ & ~new_new_n5965__;
  assign new_new_n5967__ = ~new_new_n868__ & new_new_n5213__;
  assign new_new_n5968__ = ~new_new_n1061__ & new_new_n5191__;
  assign new_new_n5969__ = ~new_new_n1207__ & new_new_n5183__;
  assign new_new_n5970__ = ~new_new_n5967__ & ~new_new_n5968__;
  assign new_new_n5971__ = ~new_new_n5969__ & new_new_n5970__;
  assign new_new_n5972__ = ~new_new_n4550__ & new_new_n5195__;
  assign new_new_n5973__ = ~pi23 & ~new_new_n5972__;
  assign new_new_n5974__ = ~pi22 & new_new_n5195__;
  assign new_new_n5975__ = ~new_new_n4550__ & new_new_n5974__;
  assign new_new_n5976__ = ~new_new_n5973__ & ~new_new_n5975__;
  assign new_new_n5977__ = new_new_n5971__ & ~new_new_n5976__;
  assign new_new_n5978__ = pi23 & ~new_new_n5971__;
  assign new_new_n5979__ = ~new_new_n5977__ & ~new_new_n5978__;
  assign new_new_n5980__ = new_new_n3311__ & ~new_new_n3618__;
  assign new_new_n5981__ = ~new_new_n3618__ & ~new_new_n4919__;
  assign new_new_n5982__ = new_new_n3618__ & ~new_new_n4918__;
  assign new_new_n5983__ = ~new_new_n3553__ & new_new_n5982__;
  assign new_new_n5984__ = ~new_new_n5981__ & ~new_new_n5983__;
  assign new_new_n5985__ = ~new_new_n4900__ & ~new_new_n5984__;
  assign new_new_n5986__ = new_new_n873__ & ~new_new_n1325__;
  assign new_new_n5987__ = ~new_new_n333__ & ~new_new_n1556__;
  assign new_new_n5988__ = ~new_new_n5980__ & ~new_new_n5986__;
  assign new_new_n5989__ = ~new_new_n5987__ & new_new_n5988__;
  assign new_new_n5990__ = ~new_new_n5985__ & new_new_n5989__;
  assign new_new_n5991__ = pi26 & ~new_new_n5990__;
  assign new_new_n5992__ = ~pi26 & new_new_n5990__;
  assign new_new_n5993__ = ~new_new_n5991__ & ~new_new_n5992__;
  assign new_new_n5994__ = ~new_new_n1823__ & ~new_new_n4818__;
  assign new_new_n5995__ = ~new_new_n1902__ & new_new_n4212__;
  assign new_new_n5996__ = new_new_n4813__ & ~new_new_n5274__;
  assign new_new_n5997__ = ~new_new_n5994__ & ~new_new_n5995__;
  assign new_new_n5998__ = ~new_new_n5996__ & new_new_n5997__;
  assign new_new_n5999__ = ~new_new_n1660__ & new_new_n4214__;
  assign new_new_n6000__ = pi29 & ~new_new_n5999__;
  assign new_new_n6001__ = ~new_new_n1660__ & new_new_n5732__;
  assign new_new_n6002__ = ~new_new_n6000__ & ~new_new_n6001__;
  assign new_new_n6003__ = new_new_n5998__ & ~new_new_n6002__;
  assign new_new_n6004__ = ~pi29 & ~new_new_n5998__;
  assign new_new_n6005__ = ~new_new_n6003__ & ~new_new_n6004__;
  assign new_new_n6006__ = new_new_n161__ & ~new_new_n2024__;
  assign new_new_n6007__ = new_new_n765__ & ~new_new_n2130__;
  assign new_new_n6008__ = ~new_new_n6006__ & ~new_new_n6007__;
  assign new_new_n6009__ = ~pi31 & ~new_new_n6008__;
  assign new_new_n6010__ = new_new_n71__ & ~new_new_n2024__;
  assign new_new_n6011__ = new_new_n161__ & ~new_new_n2224__;
  assign new_new_n6012__ = new_new_n2225__ & new_new_n2420__;
  assign new_new_n6013__ = ~new_new_n2024__ & new_new_n2224__;
  assign new_new_n6014__ = new_new_n2130__ & new_new_n6013__;
  assign new_new_n6015__ = ~new_new_n3474__ & new_new_n6014__;
  assign new_new_n6016__ = ~new_new_n6012__ & ~new_new_n6015__;
  assign new_new_n6017__ = new_new_n2313__ & ~new_new_n6016__;
  assign new_new_n6018__ = ~new_new_n2130__ & new_new_n2224__;
  assign new_new_n6019__ = ~new_new_n2420__ & new_new_n6018__;
  assign new_new_n6020__ = new_new_n2024__ & ~new_new_n2224__;
  assign new_new_n6021__ = new_new_n2130__ & new_new_n6020__;
  assign new_new_n6022__ = ~new_new_n2313__ & new_new_n6021__;
  assign new_new_n6023__ = ~new_new_n6019__ & ~new_new_n6022__;
  assign new_new_n6024__ = new_new_n3474__ & ~new_new_n6023__;
  assign new_new_n6025__ = ~new_new_n2313__ & new_new_n6018__;
  assign new_new_n6026__ = ~new_new_n6021__ & ~new_new_n6025__;
  assign new_new_n6027__ = ~new_new_n2420__ & ~new_new_n6026__;
  assign new_new_n6028__ = new_new_n2224__ & new_new_n2420__;
  assign new_new_n6029__ = new_new_n2130__ & ~new_new_n6028__;
  assign new_new_n6030__ = ~new_new_n2024__ & ~new_new_n6018__;
  assign new_new_n6031__ = ~new_new_n6029__ & new_new_n6030__;
  assign new_new_n6032__ = ~new_new_n6027__ & ~new_new_n6031__;
  assign new_new_n6033__ = ~new_new_n6024__ & new_new_n6032__;
  assign new_new_n6034__ = ~new_new_n6017__ & new_new_n6033__;
  assign new_new_n6035__ = new_new_n2024__ & new_new_n6018__;
  assign new_new_n6036__ = new_new_n6034__ & ~new_new_n6035__;
  assign new_new_n6037__ = new_new_n765__ & ~new_new_n6036__;
  assign new_new_n6038__ = ~new_new_n6010__ & ~new_new_n6011__;
  assign new_new_n6039__ = ~new_new_n6037__ & new_new_n6038__;
  assign new_new_n6040__ = pi31 & ~new_new_n6039__;
  assign new_new_n6041__ = ~new_new_n6009__ & ~new_new_n6040__;
  assign new_new_n6042__ = new_new_n2420__ & new_new_n3474__;
  assign new_new_n6043__ = ~new_new_n3475__ & ~new_new_n6042__;
  assign new_new_n6044__ = new_new_n765__ & new_new_n6043__;
  assign new_new_n6045__ = ~new_new_n2421__ & ~new_new_n6044__;
  assign new_new_n6046__ = new_new_n2224__ & ~new_new_n6045__;
  assign new_new_n6047__ = ~new_new_n2224__ & ~new_new_n2420__;
  assign new_new_n6048__ = ~new_new_n3474__ & new_new_n6047__;
  assign new_new_n6049__ = ~new_new_n161__ & ~new_new_n6048__;
  assign new_new_n6050__ = ~new_new_n71__ & new_new_n2313__;
  assign new_new_n6051__ = ~new_new_n6049__ & new_new_n6050__;
  assign new_new_n6052__ = ~new_new_n2313__ & new_new_n3474__;
  assign new_new_n6053__ = ~new_new_n2224__ & new_new_n6052__;
  assign new_new_n6054__ = ~new_new_n71__ & ~new_new_n6053__;
  assign new_new_n6055__ = ~new_new_n161__ & new_new_n2420__;
  assign new_new_n6056__ = ~new_new_n6054__ & new_new_n6055__;
  assign new_new_n6057__ = pi31 & ~new_new_n6051__;
  assign new_new_n6058__ = ~new_new_n6056__ & new_new_n6057__;
  assign new_new_n6059__ = ~new_new_n6046__ & new_new_n6058__;
  assign new_new_n6060__ = new_new_n765__ & ~new_new_n2224__;
  assign new_new_n6061__ = new_new_n161__ & ~new_new_n2420__;
  assign new_new_n6062__ = ~new_new_n6060__ & ~new_new_n6061__;
  assign new_new_n6063__ = ~pi31 & ~new_new_n6062__;
  assign new_new_n6064__ = ~new_new_n6059__ & ~new_new_n6063__;
  assign new_new_n6065__ = ~new_new_n383__ & ~new_new_n1035__;
  assign new_new_n6066__ = ~new_new_n346__ & ~new_new_n768__;
  assign new_new_n6067__ = ~new_new_n749__ & ~new_new_n937__;
  assign new_new_n6068__ = new_new_n3211__ & new_new_n6067__;
  assign new_new_n6069__ = new_new_n2025__ & new_new_n6068__;
  assign new_new_n6070__ = ~new_new_n249__ & ~new_new_n427__;
  assign new_new_n6071__ = ~new_new_n160__ & ~new_new_n248__;
  assign new_new_n6072__ = ~new_new_n438__ & ~new_new_n853__;
  assign new_new_n6073__ = new_new_n6071__ & new_new_n6072__;
  assign new_new_n6074__ = ~new_new_n136__ & new_new_n4304__;
  assign new_new_n6075__ = ~new_new_n143__ & new_new_n695__;
  assign new_new_n6076__ = ~new_new_n1009__ & new_new_n6075__;
  assign new_new_n6077__ = new_new_n6073__ & new_new_n6074__;
  assign new_new_n6078__ = new_new_n6065__ & new_new_n6066__;
  assign new_new_n6079__ = new_new_n6070__ & new_new_n6078__;
  assign new_new_n6080__ = new_new_n6076__ & new_new_n6077__;
  assign new_new_n6081__ = new_new_n2478__ & new_new_n6080__;
  assign new_new_n6082__ = new_new_n1962__ & new_new_n6079__;
  assign new_new_n6083__ = new_new_n6069__ & new_new_n6082__;
  assign new_new_n6084__ = new_new_n2140__ & new_new_n6081__;
  assign new_new_n6085__ = new_new_n4486__ & new_new_n6084__;
  assign new_new_n6086__ = new_new_n6083__ & new_new_n6085__;
  assign new_new_n6087__ = new_new_n1446__ & new_new_n2195__;
  assign new_new_n6088__ = new_new_n6086__ & new_new_n6087__;
  assign new_new_n6089__ = ~new_new_n6064__ & ~new_new_n6088__;
  assign new_new_n6090__ = ~new_new_n103__ & ~new_new_n479__;
  assign new_new_n6091__ = ~new_new_n240__ & ~new_new_n843__;
  assign new_new_n6092__ = ~new_new_n1031__ & new_new_n6091__;
  assign new_new_n6093__ = ~new_new_n266__ & ~new_new_n1308__;
  assign new_new_n6094__ = new_new_n1922__ & new_new_n4231__;
  assign new_new_n6095__ = new_new_n6093__ & new_new_n6094__;
  assign new_new_n6096__ = new_new_n3416__ & new_new_n6092__;
  assign new_new_n6097__ = new_new_n5314__ & new_new_n5379__;
  assign new_new_n6098__ = new_new_n6096__ & new_new_n6097__;
  assign new_new_n6099__ = new_new_n2028__ & new_new_n6095__;
  assign new_new_n6100__ = new_new_n6090__ & new_new_n6099__;
  assign new_new_n6101__ = new_new_n6098__ & new_new_n6100__;
  assign new_new_n6102__ = ~new_new_n213__ & ~new_new_n332__;
  assign new_new_n6103__ = new_new_n2768__ & new_new_n6102__;
  assign new_new_n6104__ = new_new_n2331__ & new_new_n6070__;
  assign new_new_n6105__ = new_new_n6103__ & new_new_n6104__;
  assign new_new_n6106__ = ~new_new_n164__ & ~new_new_n222__;
  assign new_new_n6107__ = ~new_new_n251__ & ~new_new_n267__;
  assign new_new_n6108__ = ~new_new_n351__ & ~new_new_n694__;
  assign new_new_n6109__ = ~new_new_n1094__ & ~new_new_n1398__;
  assign new_new_n6110__ = new_new_n6108__ & new_new_n6109__;
  assign new_new_n6111__ = new_new_n6106__ & new_new_n6107__;
  assign new_new_n6112__ = ~new_new_n835__ & new_new_n4314__;
  assign new_new_n6113__ = new_new_n6111__ & new_new_n6112__;
  assign new_new_n6114__ = ~new_new_n218__ & new_new_n6110__;
  assign new_new_n6115__ = new_new_n876__ & new_new_n2259__;
  assign new_new_n6116__ = new_new_n2993__ & new_new_n6115__;
  assign new_new_n6117__ = new_new_n6113__ & new_new_n6114__;
  assign new_new_n6118__ = new_new_n709__ & ~new_new_n1539__;
  assign new_new_n6119__ = new_new_n6117__ & new_new_n6118__;
  assign new_new_n6120__ = new_new_n6105__ & new_new_n6116__;
  assign new_new_n6121__ = new_new_n6119__ & new_new_n6120__;
  assign new_new_n6122__ = ~new_new_n675__ & ~new_new_n1507__;
  assign new_new_n6123__ = ~new_new_n327__ & ~new_new_n701__;
  assign new_new_n6124__ = ~new_new_n255__ & ~new_new_n851__;
  assign new_new_n6125__ = ~new_new_n189__ & new_new_n1470__;
  assign new_new_n6126__ = ~new_new_n1568__ & new_new_n6123__;
  assign new_new_n6127__ = new_new_n6125__ & new_new_n6126__;
  assign new_new_n6128__ = new_new_n1339__ & new_new_n2469__;
  assign new_new_n6129__ = new_new_n2909__ & new_new_n3793__;
  assign new_new_n6130__ = new_new_n6122__ & new_new_n6124__;
  assign new_new_n6131__ = new_new_n6129__ & new_new_n6130__;
  assign new_new_n6132__ = new_new_n6127__ & new_new_n6128__;
  assign new_new_n6133__ = new_new_n6131__ & new_new_n6132__;
  assign new_new_n6134__ = new_new_n2181__ & new_new_n6133__;
  assign new_new_n6135__ = new_new_n5364__ & new_new_n6134__;
  assign new_new_n6136__ = new_new_n6101__ & new_new_n6121__;
  assign new_new_n6137__ = new_new_n6135__ & new_new_n6136__;
  assign new_new_n6138__ = new_new_n983__ & new_new_n6137__;
  assign new_new_n6139__ = ~new_new_n6089__ & ~new_new_n6138__;
  assign new_new_n6140__ = new_new_n6064__ & new_new_n6088__;
  assign new_new_n6141__ = new_new_n6138__ & ~new_new_n6140__;
  assign new_new_n6142__ = ~new_new_n160__ & ~new_new_n329__;
  assign new_new_n6143__ = ~new_new_n947__ & new_new_n2160__;
  assign new_new_n6144__ = ~new_new_n222__ & ~new_new_n1064__;
  assign new_new_n6145__ = ~new_new_n607__ & new_new_n6144__;
  assign new_new_n6146__ = new_new_n6142__ & new_new_n6143__;
  assign new_new_n6147__ = new_new_n6145__ & new_new_n6146__;
  assign new_new_n6148__ = new_new_n1250__ & new_new_n6147__;
  assign new_new_n6149__ = ~new_new_n1007__ & ~new_new_n1094__;
  assign new_new_n6150__ = ~new_new_n179__ & ~new_new_n996__;
  assign new_new_n6151__ = ~new_new_n380__ & new_new_n6150__;
  assign new_new_n6152__ = ~new_new_n721__ & new_new_n1709__;
  assign new_new_n6153__ = new_new_n6151__ & new_new_n6152__;
  assign new_new_n6154__ = new_new_n1037__ & new_new_n6153__;
  assign new_new_n6155__ = ~new_new_n959__ & ~new_new_n1176__;
  assign new_new_n6156__ = ~new_new_n82__ & ~new_new_n182__;
  assign new_new_n6157__ = ~new_new_n692__ & ~new_new_n723__;
  assign new_new_n6158__ = new_new_n6156__ & new_new_n6157__;
  assign new_new_n6159__ = ~new_new_n317__ & ~new_new_n566__;
  assign new_new_n6160__ = ~new_new_n945__ & new_new_n6159__;
  assign new_new_n6161__ = new_new_n1778__ & new_new_n6158__;
  assign new_new_n6162__ = new_new_n2196__ & new_new_n2758__;
  assign new_new_n6163__ = new_new_n6161__ & new_new_n6162__;
  assign new_new_n6164__ = new_new_n6160__ & new_new_n6163__;
  assign new_new_n6165__ = ~new_new_n248__ & ~new_new_n251__;
  assign new_new_n6166__ = ~new_new_n309__ & ~new_new_n476__;
  assign new_new_n6167__ = ~new_new_n496__ & ~new_new_n701__;
  assign new_new_n6168__ = new_new_n6166__ & new_new_n6167__;
  assign new_new_n6169__ = ~new_new_n1701__ & new_new_n6165__;
  assign new_new_n6170__ = new_new_n1742__ & new_new_n2158__;
  assign new_new_n6171__ = new_new_n6149__ & new_new_n6170__;
  assign new_new_n6172__ = new_new_n6168__ & new_new_n6169__;
  assign new_new_n6173__ = new_new_n743__ & ~new_new_n1486__;
  assign new_new_n6174__ = new_new_n1840__ & new_new_n6155__;
  assign new_new_n6175__ = new_new_n6173__ & new_new_n6174__;
  assign new_new_n6176__ = new_new_n6171__ & new_new_n6172__;
  assign new_new_n6177__ = new_new_n378__ & new_new_n3417__;
  assign new_new_n6178__ = new_new_n6176__ & new_new_n6177__;
  assign new_new_n6179__ = new_new_n6154__ & new_new_n6175__;
  assign new_new_n6180__ = new_new_n6178__ & new_new_n6179__;
  assign new_new_n6181__ = new_new_n6164__ & new_new_n6180__;
  assign new_new_n6182__ = ~new_new_n298__ & ~new_new_n875__;
  assign new_new_n6183__ = ~new_new_n286__ & ~new_new_n1003__;
  assign new_new_n6184__ = new_new_n87__ & ~new_new_n1165__;
  assign new_new_n6185__ = ~new_new_n937__ & ~new_new_n940__;
  assign new_new_n6186__ = ~new_new_n259__ & ~new_new_n312__;
  assign new_new_n6187__ = ~new_new_n388__ & ~new_new_n473__;
  assign new_new_n6188__ = ~new_new_n320__ & new_new_n6187__;
  assign new_new_n6189__ = ~new_new_n588__ & new_new_n6091__;
  assign new_new_n6190__ = new_new_n6185__ & new_new_n6186__;
  assign new_new_n6191__ = new_new_n6189__ & new_new_n6190__;
  assign new_new_n6192__ = ~new_new_n218__ & new_new_n6188__;
  assign new_new_n6193__ = ~new_new_n809__ & new_new_n1330__;
  assign new_new_n6194__ = new_new_n6192__ & new_new_n6193__;
  assign new_new_n6195__ = new_new_n6191__ & new_new_n6194__;
  assign new_new_n6196__ = ~new_new_n168__ & ~new_new_n510__;
  assign new_new_n6197__ = ~new_new_n1167__ & new_new_n6196__;
  assign new_new_n6198__ = new_new_n6182__ & ~new_new_n6184__;
  assign new_new_n6199__ = new_new_n6197__ & new_new_n6198__;
  assign new_new_n6200__ = new_new_n484__ & new_new_n1000__;
  assign new_new_n6201__ = new_new_n1078__ & new_new_n2770__;
  assign new_new_n6202__ = new_new_n6183__ & new_new_n6201__;
  assign new_new_n6203__ = new_new_n6199__ & new_new_n6200__;
  assign new_new_n6204__ = new_new_n3700__ & new_new_n6203__;
  assign new_new_n6205__ = new_new_n4962__ & new_new_n6202__;
  assign new_new_n6206__ = new_new_n6204__ & new_new_n6205__;
  assign new_new_n6207__ = new_new_n6148__ & new_new_n6195__;
  assign new_new_n6208__ = new_new_n6206__ & new_new_n6207__;
  assign new_new_n6209__ = new_new_n5007__ & new_new_n6208__;
  assign new_new_n6210__ = new_new_n6181__ & new_new_n6209__;
  assign new_new_n6211__ = ~new_new_n483__ & ~new_new_n1080__;
  assign new_new_n6212__ = ~new_new_n108__ & ~new_new_n933__;
  assign new_new_n6213__ = ~new_new_n940__ & ~new_new_n1113__;
  assign new_new_n6214__ = new_new_n6212__ & new_new_n6213__;
  assign new_new_n6215__ = ~new_new_n591__ & ~new_new_n719__;
  assign new_new_n6216__ = new_new_n779__ & ~new_new_n2697__;
  assign new_new_n6217__ = new_new_n2970__ & new_new_n3258__;
  assign new_new_n6218__ = new_new_n4314__ & new_new_n5358__;
  assign new_new_n6219__ = new_new_n6217__ & new_new_n6218__;
  assign new_new_n6220__ = new_new_n6215__ & new_new_n6216__;
  assign new_new_n6221__ = ~new_new_n344__ & new_new_n6214__;
  assign new_new_n6222__ = ~new_new_n630__ & new_new_n1468__;
  assign new_new_n6223__ = new_new_n2316__ & new_new_n6211__;
  assign new_new_n6224__ = new_new_n6222__ & new_new_n6223__;
  assign new_new_n6225__ = new_new_n6220__ & new_new_n6221__;
  assign new_new_n6226__ = new_new_n6219__ & new_new_n6225__;
  assign new_new_n6227__ = new_new_n6224__ & new_new_n6226__;
  assign new_new_n6228__ = new_new_n5286__ & new_new_n6227__;
  assign new_new_n6229__ = ~new_new_n811__ & ~new_new_n871__;
  assign new_new_n6230__ = ~new_new_n1003__ & new_new_n4564__;
  assign new_new_n6231__ = new_new_n6229__ & new_new_n6230__;
  assign new_new_n6232__ = ~new_new_n316__ & new_new_n6231__;
  assign new_new_n6233__ = ~new_new_n652__ & new_new_n6232__;
  assign new_new_n6234__ = ~new_new_n785__ & ~new_new_n851__;
  assign new_new_n6235__ = ~new_new_n226__ & ~new_new_n495__;
  assign new_new_n6236__ = ~new_new_n1070__ & new_new_n2707__;
  assign new_new_n6237__ = new_new_n3181__ & new_new_n6236__;
  assign new_new_n6238__ = new_new_n5301__ & new_new_n6235__;
  assign new_new_n6239__ = new_new_n6237__ & new_new_n6238__;
  assign new_new_n6240__ = ~new_new_n196__ & ~new_new_n240__;
  assign new_new_n6241__ = ~new_new_n283__ & ~new_new_n438__;
  assign new_new_n6242__ = ~new_new_n473__ & ~new_new_n990__;
  assign new_new_n6243__ = new_new_n6241__ & new_new_n6242__;
  assign new_new_n6244__ = ~new_new_n266__ & ~new_new_n277__;
  assign new_new_n6245__ = new_new_n2585__ & new_new_n6240__;
  assign new_new_n6246__ = new_new_n6244__ & new_new_n6245__;
  assign new_new_n6247__ = new_new_n6243__ & new_new_n6246__;
  assign new_new_n6248__ = ~new_new_n166__ & ~new_new_n729__;
  assign new_new_n6249__ = ~new_new_n106__ & ~new_new_n260__;
  assign new_new_n6250__ = ~new_new_n183__ & new_new_n6249__;
  assign new_new_n6251__ = ~new_new_n878__ & new_new_n6250__;
  assign new_new_n6252__ = new_new_n2266__ & new_new_n6248__;
  assign new_new_n6253__ = new_new_n6251__ & new_new_n6252__;
  assign new_new_n6254__ = ~new_new_n1539__ & new_new_n2796__;
  assign new_new_n6255__ = new_new_n6253__ & new_new_n6254__;
  assign new_new_n6256__ = ~new_new_n632__ & new_new_n1747__;
  assign new_new_n6257__ = ~new_new_n92__ & ~new_new_n119__;
  assign new_new_n6258__ = ~new_new_n335__ & ~new_new_n509__;
  assign new_new_n6259__ = ~new_new_n1212__ & ~new_new_n1343__;
  assign new_new_n6260__ = new_new_n6258__ & new_new_n6259__;
  assign new_new_n6261__ = ~new_new_n675__ & new_new_n6257__;
  assign new_new_n6262__ = ~new_new_n835__ & new_new_n3483__;
  assign new_new_n6263__ = new_new_n6261__ & new_new_n6262__;
  assign new_new_n6264__ = ~new_new_n676__ & new_new_n6260__;
  assign new_new_n6265__ = new_new_n2639__ & new_new_n6155__;
  assign new_new_n6266__ = new_new_n6264__ & new_new_n6265__;
  assign new_new_n6267__ = new_new_n6256__ & new_new_n6263__;
  assign new_new_n6268__ = new_new_n6266__ & new_new_n6267__;
  assign new_new_n6269__ = new_new_n1610__ & new_new_n6247__;
  assign new_new_n6270__ = new_new_n6268__ & new_new_n6269__;
  assign new_new_n6271__ = new_new_n6255__ & new_new_n6270__;
  assign new_new_n6272__ = ~new_new_n189__ & ~new_new_n222__;
  assign new_new_n6273__ = ~new_new_n322__ & new_new_n6234__;
  assign new_new_n6274__ = new_new_n6272__ & new_new_n6273__;
  assign new_new_n6275__ = ~new_new_n508__ & new_new_n1037__;
  assign new_new_n6276__ = new_new_n1296__ & new_new_n1630__;
  assign new_new_n6277__ = new_new_n2507__ & new_new_n3322__;
  assign new_new_n6278__ = new_new_n6276__ & new_new_n6277__;
  assign new_new_n6279__ = new_new_n6274__ & new_new_n6275__;
  assign new_new_n6280__ = new_new_n2264__ & new_new_n6279__;
  assign new_new_n6281__ = new_new_n6239__ & new_new_n6278__;
  assign new_new_n6282__ = new_new_n6280__ & new_new_n6281__;
  assign new_new_n6283__ = new_new_n3873__ & new_new_n6233__;
  assign new_new_n6284__ = new_new_n6282__ & new_new_n6283__;
  assign new_new_n6285__ = new_new_n6228__ & new_new_n6284__;
  assign new_new_n6286__ = new_new_n6271__ & new_new_n6285__;
  assign new_new_n6287__ = ~new_new_n6210__ & ~new_new_n6286__;
  assign new_new_n6288__ = new_new_n6210__ & new_new_n6286__;
  assign new_new_n6289__ = ~pi08 & ~new_new_n6288__;
  assign new_new_n6290__ = ~new_new_n6287__ & ~new_new_n6289__;
  assign new_new_n6291__ = ~new_new_n6141__ & new_new_n6290__;
  assign new_new_n6292__ = ~new_new_n6139__ & ~new_new_n6291__;
  assign new_new_n6293__ = new_new_n6041__ & ~new_new_n6292__;
  assign new_new_n6294__ = ~new_new_n6041__ & new_new_n6292__;
  assign new_new_n6295__ = new_new_n830__ & new_new_n6101__;
  assign new_new_n6296__ = ~new_new_n106__ & ~new_new_n308__;
  assign new_new_n6297__ = ~new_new_n274__ & ~new_new_n675__;
  assign new_new_n6298__ = new_new_n6296__ & new_new_n6297__;
  assign new_new_n6299__ = ~new_new_n309__ & ~new_new_n746__;
  assign new_new_n6300__ = ~new_new_n1210__ & new_new_n6299__;
  assign new_new_n6301__ = new_new_n3205__ & new_new_n6300__;
  assign new_new_n6302__ = ~new_new_n935__ & ~new_new_n1486__;
  assign new_new_n6303__ = new_new_n5785__ & new_new_n6302__;
  assign new_new_n6304__ = new_new_n6298__ & new_new_n6301__;
  assign new_new_n6305__ = new_new_n6303__ & new_new_n6304__;
  assign new_new_n6306__ = ~new_new_n179__ & ~new_new_n388__;
  assign new_new_n6307__ = ~new_new_n724__ & new_new_n6306__;
  assign new_new_n6308__ = ~new_new_n255__ & ~new_new_n322__;
  assign new_new_n6309__ = ~new_new_n945__ & ~new_new_n1632__;
  assign new_new_n6310__ = new_new_n2093__ & ~new_new_n2697__;
  assign new_new_n6311__ = new_new_n6309__ & new_new_n6310__;
  assign new_new_n6312__ = new_new_n6307__ & new_new_n6308__;
  assign new_new_n6313__ = new_new_n2226__ & new_new_n3969__;
  assign new_new_n6314__ = new_new_n6312__ & new_new_n6313__;
  assign new_new_n6315__ = new_new_n4505__ & new_new_n6311__;
  assign new_new_n6316__ = new_new_n6314__ & new_new_n6315__;
  assign new_new_n6317__ = new_new_n1521__ & new_new_n2343__;
  assign new_new_n6318__ = new_new_n6316__ & new_new_n6317__;
  assign new_new_n6319__ = new_new_n6305__ & new_new_n6318__;
  assign new_new_n6320__ = ~new_new_n251__ & ~new_new_n947__;
  assign new_new_n6321__ = ~new_new_n657__ & ~new_new_n829__;
  assign new_new_n6322__ = ~new_new_n260__ & ~new_new_n871__;
  assign new_new_n6323__ = ~new_new_n482__ & ~new_new_n495__;
  assign new_new_n6324__ = ~new_new_n270__ & ~new_new_n473__;
  assign new_new_n6325__ = ~new_new_n329__ & ~new_new_n602__;
  assign new_new_n6326__ = ~new_new_n869__ & new_new_n1095__;
  assign new_new_n6327__ = new_new_n4566__ & new_new_n6320__;
  assign new_new_n6328__ = new_new_n6321__ & new_new_n6323__;
  assign new_new_n6329__ = new_new_n6327__ & new_new_n6328__;
  assign new_new_n6330__ = new_new_n6325__ & new_new_n6326__;
  assign new_new_n6331__ = new_new_n984__ & new_new_n6324__;
  assign new_new_n6332__ = new_new_n1209__ & new_new_n1599__;
  assign new_new_n6333__ = new_new_n2424__ & new_new_n6322__;
  assign new_new_n6334__ = new_new_n6332__ & new_new_n6333__;
  assign new_new_n6335__ = new_new_n6330__ & new_new_n6331__;
  assign new_new_n6336__ = new_new_n116__ & new_new_n6329__;
  assign new_new_n6337__ = new_new_n3791__ & new_new_n6336__;
  assign new_new_n6338__ = new_new_n6334__ & new_new_n6335__;
  assign new_new_n6339__ = new_new_n6337__ & new_new_n6338__;
  assign new_new_n6340__ = new_new_n4423__ & new_new_n4476__;
  assign new_new_n6341__ = new_new_n6339__ & new_new_n6340__;
  assign new_new_n6342__ = new_new_n6295__ & new_new_n6341__;
  assign new_new_n6343__ = new_new_n6319__ & new_new_n6342__;
  assign new_new_n6344__ = new_new_n6138__ & new_new_n6343__;
  assign new_new_n6345__ = ~new_new_n6138__ & ~new_new_n6343__;
  assign new_new_n6346__ = ~pi11 & ~new_new_n6344__;
  assign new_new_n6347__ = ~new_new_n6345__ & ~new_new_n6346__;
  assign new_new_n6348__ = ~new_new_n6344__ & new_new_n6347__;
  assign new_new_n6349__ = ~new_new_n6345__ & new_new_n6346__;
  assign new_new_n6350__ = ~pi11 & ~new_new_n6349__;
  assign new_new_n6351__ = ~new_new_n6348__ & ~new_new_n6350__;
  assign new_new_n6352__ = ~new_new_n6294__ & new_new_n6351__;
  assign new_new_n6353__ = ~new_new_n6293__ & ~new_new_n6352__;
  assign new_new_n6354__ = ~new_new_n6005__ & new_new_n6353__;
  assign new_new_n6355__ = new_new_n765__ & ~new_new_n3535__;
  assign new_new_n6356__ = new_new_n161__ & ~new_new_n2130__;
  assign new_new_n6357__ = ~new_new_n6355__ & ~new_new_n6356__;
  assign new_new_n6358__ = ~pi31 & ~new_new_n6357__;
  assign new_new_n6359__ = ~new_new_n71__ & new_new_n5497__;
  assign new_new_n6360__ = new_new_n2130__ & ~new_new_n6359__;
  assign new_new_n6361__ = new_new_n3479__ & ~new_new_n3496__;
  assign new_new_n6362__ = new_new_n2130__ & ~new_new_n6361__;
  assign new_new_n6363__ = new_new_n6359__ & ~new_new_n6362__;
  assign new_new_n6364__ = ~new_new_n161__ & ~new_new_n6360__;
  assign new_new_n6365__ = ~new_new_n6363__ & new_new_n6364__;
  assign new_new_n6366__ = ~new_new_n6006__ & ~new_new_n6365__;
  assign new_new_n6367__ = pi31 & ~new_new_n6366__;
  assign new_new_n6368__ = ~new_new_n6358__ & ~new_new_n6367__;
  assign new_new_n6369__ = ~new_new_n6347__ & ~new_new_n6368__;
  assign new_new_n6370__ = new_new_n6354__ & new_new_n6369__;
  assign new_new_n6371__ = ~new_new_n5639__ & ~new_new_n5641__;
  assign new_new_n6372__ = new_new_n6005__ & ~new_new_n6353__;
  assign new_new_n6373__ = new_new_n5451__ & new_new_n6372__;
  assign new_new_n6374__ = ~new_new_n6347__ & ~new_new_n6373__;
  assign new_new_n6375__ = new_new_n6368__ & ~new_new_n6374__;
  assign new_new_n6376__ = ~new_new_n5451__ & ~new_new_n6372__;
  assign new_new_n6377__ = ~new_new_n6375__ & new_new_n6376__;
  assign new_new_n6378__ = new_new_n6347__ & new_new_n6368__;
  assign new_new_n6379__ = new_new_n5451__ & new_new_n6378__;
  assign new_new_n6380__ = new_new_n6354__ & ~new_new_n6379__;
  assign new_new_n6381__ = ~new_new_n6368__ & new_new_n6374__;
  assign new_new_n6382__ = ~new_new_n6380__ & ~new_new_n6381__;
  assign new_new_n6383__ = ~new_new_n6377__ & new_new_n6382__;
  assign new_new_n6384__ = new_new_n6371__ & ~new_new_n6383__;
  assign new_new_n6385__ = new_new_n6372__ & new_new_n6378__;
  assign new_new_n6386__ = new_new_n5451__ & ~new_new_n6371__;
  assign new_new_n6387__ = ~new_new_n6385__ & new_new_n6386__;
  assign new_new_n6388__ = ~new_new_n6370__ & ~new_new_n6387__;
  assign new_new_n6389__ = ~new_new_n6384__ & new_new_n6388__;
  assign new_new_n6390__ = ~new_new_n5355__ & ~new_new_n5532__;
  assign new_new_n6391__ = new_new_n5355__ & new_new_n5532__;
  assign new_new_n6392__ = ~new_new_n6390__ & ~new_new_n6391__;
  assign new_new_n6393__ = new_new_n5451__ & new_new_n5641__;
  assign new_new_n6394__ = ~new_new_n5451__ & new_new_n5639__;
  assign new_new_n6395__ = ~new_new_n6393__ & ~new_new_n6394__;
  assign new_new_n6396__ = pi14 & ~new_new_n6395__;
  assign new_new_n6397__ = ~pi14 & new_new_n6395__;
  assign new_new_n6398__ = ~new_new_n6396__ & ~new_new_n6397__;
  assign new_new_n6399__ = ~new_new_n6392__ & new_new_n6398__;
  assign new_new_n6400__ = new_new_n5324__ & new_new_n6391__;
  assign new_new_n6401__ = ~new_new_n6390__ & ~new_new_n6398__;
  assign new_new_n6402__ = ~new_new_n6400__ & new_new_n6401__;
  assign new_new_n6403__ = ~new_new_n6399__ & ~new_new_n6402__;
  assign new_new_n6404__ = new_new_n6389__ & new_new_n6403__;
  assign new_new_n6405__ = ~new_new_n6389__ & ~new_new_n6403__;
  assign new_new_n6406__ = ~new_new_n6404__ & ~new_new_n6405__;
  assign new_new_n6407__ = ~new_new_n1660__ & ~new_new_n4818__;
  assign new_new_n6408__ = ~new_new_n1737__ & new_new_n4212__;
  assign new_new_n6409__ = ~new_new_n1466__ & new_new_n4815__;
  assign new_new_n6410__ = ~new_new_n5665__ & ~new_new_n5881__;
  assign new_new_n6411__ = new_new_n4813__ & ~new_new_n6410__;
  assign new_new_n6412__ = ~new_new_n6407__ & ~new_new_n6408__;
  assign new_new_n6413__ = ~new_new_n6409__ & new_new_n6412__;
  assign new_new_n6414__ = ~new_new_n6411__ & new_new_n6413__;
  assign new_new_n6415__ = pi29 & ~new_new_n6414__;
  assign new_new_n6416__ = ~pi29 & new_new_n6414__;
  assign new_new_n6417__ = ~new_new_n6415__ & ~new_new_n6416__;
  assign new_new_n6418__ = new_new_n6406__ & new_new_n6417__;
  assign new_new_n6419__ = ~new_new_n6406__ & ~new_new_n6417__;
  assign new_new_n6420__ = ~new_new_n6418__ & ~new_new_n6419__;
  assign new_new_n6421__ = new_new_n5993__ & new_new_n6420__;
  assign new_new_n6422__ = ~new_new_n5993__ & ~new_new_n6420__;
  assign new_new_n6423__ = ~new_new_n6421__ & ~new_new_n6422__;
  assign new_new_n6424__ = ~new_new_n4900__ & new_new_n5048__;
  assign new_new_n6425__ = ~new_new_n333__ & ~new_new_n1466__;
  assign new_new_n6426__ = new_new_n873__ & ~new_new_n1556__;
  assign new_new_n6427__ = ~new_new_n6425__ & ~new_new_n6426__;
  assign new_new_n6428__ = ~new_new_n6424__ & new_new_n6427__;
  assign new_new_n6429__ = pi26 & ~new_new_n6428__;
  assign new_new_n6430__ = new_new_n512__ & ~new_new_n1325__;
  assign new_new_n6431__ = new_new_n801__ & ~new_new_n1325__;
  assign new_new_n6432__ = ~pi26 & ~new_new_n6431__;
  assign new_new_n6433__ = ~new_new_n6430__ & ~new_new_n6432__;
  assign new_new_n6434__ = new_new_n6428__ & ~new_new_n6433__;
  assign new_new_n6435__ = ~new_new_n6429__ & ~new_new_n6434__;
  assign new_new_n6436__ = ~new_new_n6354__ & ~new_new_n6372__;
  assign new_new_n6437__ = ~new_new_n5451__ & ~new_new_n6378__;
  assign new_new_n6438__ = ~new_new_n6369__ & ~new_new_n6437__;
  assign new_new_n6439__ = ~new_new_n6371__ & ~new_new_n6438__;
  assign new_new_n6440__ = new_new_n6371__ & new_new_n6438__;
  assign new_new_n6441__ = new_new_n6436__ & ~new_new_n6439__;
  assign new_new_n6442__ = ~new_new_n6440__ & new_new_n6441__;
  assign new_new_n6443__ = new_new_n6353__ & ~new_new_n6371__;
  assign new_new_n6444__ = ~new_new_n6353__ & new_new_n6371__;
  assign new_new_n6445__ = ~new_new_n6443__ & ~new_new_n6444__;
  assign new_new_n6446__ = ~new_new_n6005__ & new_new_n6371__;
  assign new_new_n6447__ = new_new_n6379__ & ~new_new_n6446__;
  assign new_new_n6448__ = ~new_new_n6445__ & new_new_n6447__;
  assign new_new_n6449__ = ~new_new_n5451__ & new_new_n6369__;
  assign new_new_n6450__ = new_new_n6005__ & ~new_new_n6371__;
  assign new_new_n6451__ = new_new_n6449__ & ~new_new_n6450__;
  assign new_new_n6452__ = ~new_new_n6445__ & new_new_n6451__;
  assign new_new_n6453__ = ~new_new_n6379__ & ~new_new_n6449__;
  assign new_new_n6454__ = ~new_new_n6436__ & new_new_n6453__;
  assign new_new_n6455__ = new_new_n6445__ & new_new_n6454__;
  assign new_new_n6456__ = ~new_new_n6448__ & ~new_new_n6452__;
  assign new_new_n6457__ = ~new_new_n6455__ & new_new_n6456__;
  assign new_new_n6458__ = ~new_new_n6442__ & new_new_n6457__;
  assign new_new_n6459__ = new_new_n6435__ & new_new_n6458__;
  assign new_new_n6460__ = ~new_new_n6435__ & ~new_new_n6458__;
  assign new_new_n6461__ = ~new_new_n1660__ & new_new_n4212__;
  assign new_new_n6462__ = ~new_new_n1737__ & new_new_n4815__;
  assign new_new_n6463__ = ~new_new_n1902__ & ~new_new_n4818__;
  assign new_new_n6464__ = ~new_new_n6461__ & ~new_new_n6462__;
  assign new_new_n6465__ = ~new_new_n6463__ & new_new_n6464__;
  assign new_new_n6466__ = new_new_n4813__ & new_new_n5688__;
  assign new_new_n6467__ = new_new_n6465__ & ~new_new_n6466__;
  assign new_new_n6468__ = ~pi29 & ~new_new_n6467__;
  assign new_new_n6469__ = pi29 & new_new_n6467__;
  assign new_new_n6470__ = ~new_new_n6468__ & ~new_new_n6469__;
  assign new_new_n6471__ = ~new_new_n6460__ & ~new_new_n6470__;
  assign new_new_n6472__ = ~new_new_n6459__ & ~new_new_n6471__;
  assign new_new_n6473__ = new_new_n6423__ & ~new_new_n6472__;
  assign new_new_n6474__ = ~new_new_n6423__ & new_new_n6472__;
  assign new_new_n6475__ = ~new_new_n6473__ & ~new_new_n6474__;
  assign new_new_n6476__ = ~new_new_n5979__ & ~new_new_n6475__;
  assign new_new_n6477__ = new_new_n5979__ & new_new_n6475__;
  assign new_new_n6478__ = ~new_new_n3535__ & ~new_new_n4818__;
  assign new_new_n6479__ = ~new_new_n1902__ & new_new_n4815__;
  assign new_new_n6480__ = ~new_new_n1823__ & new_new_n4212__;
  assign new_new_n6481__ = ~new_new_n6478__ & ~new_new_n6479__;
  assign new_new_n6482__ = ~new_new_n6480__ & new_new_n6481__;
  assign new_new_n6483__ = ~new_new_n5268__ & ~new_new_n5543__;
  assign new_new_n6484__ = ~new_new_n5501__ & new_new_n6483__;
  assign new_new_n6485__ = ~new_new_n1902__ & ~new_new_n6484__;
  assign new_new_n6486__ = new_new_n1902__ & new_new_n6484__;
  assign new_new_n6487__ = ~new_new_n6485__ & ~new_new_n6486__;
  assign new_new_n6488__ = new_new_n4214__ & ~new_new_n6487__;
  assign new_new_n6489__ = ~pi29 & ~new_new_n6488__;
  assign new_new_n6490__ = new_new_n5732__ & ~new_new_n6487__;
  assign new_new_n6491__ = ~new_new_n6489__ & ~new_new_n6490__;
  assign new_new_n6492__ = new_new_n6482__ & ~new_new_n6491__;
  assign new_new_n6493__ = pi29 & ~new_new_n6482__;
  assign new_new_n6494__ = ~new_new_n6492__ & ~new_new_n6493__;
  assign new_new_n6495__ = ~new_new_n6293__ & ~new_new_n6294__;
  assign new_new_n6496__ = new_new_n6351__ & new_new_n6495__;
  assign new_new_n6497__ = ~new_new_n6351__ & ~new_new_n6495__;
  assign new_new_n6498__ = ~new_new_n6496__ & ~new_new_n6497__;
  assign new_new_n6499__ = ~new_new_n6494__ & new_new_n6498__;
  assign new_new_n6500__ = new_new_n6494__ & ~new_new_n6498__;
  assign new_new_n6501__ = ~new_new_n6064__ & new_new_n6138__;
  assign new_new_n6502__ = new_new_n6064__ & ~new_new_n6138__;
  assign new_new_n6503__ = ~new_new_n6501__ & ~new_new_n6502__;
  assign new_new_n6504__ = new_new_n6088__ & ~new_new_n6503__;
  assign new_new_n6505__ = ~new_new_n6089__ & ~new_new_n6140__;
  assign new_new_n6506__ = ~new_new_n6290__ & ~new_new_n6501__;
  assign new_new_n6507__ = ~new_new_n6505__ & new_new_n6506__;
  assign new_new_n6508__ = new_new_n6290__ & ~new_new_n6502__;
  assign new_new_n6509__ = new_new_n6505__ & new_new_n6508__;
  assign new_new_n6510__ = ~new_new_n6504__ & ~new_new_n6507__;
  assign new_new_n6511__ = ~new_new_n6509__ & new_new_n6510__;
  assign new_new_n6512__ = new_new_n2420__ & ~new_new_n6052__;
  assign new_new_n6513__ = new_new_n2224__ & ~new_new_n3475__;
  assign new_new_n6514__ = new_new_n765__ & ~new_new_n6512__;
  assign new_new_n6515__ = ~new_new_n6513__ & new_new_n6514__;
  assign new_new_n6516__ = ~new_new_n6028__ & ~new_new_n6515__;
  assign new_new_n6517__ = new_new_n2024__ & ~new_new_n6516__;
  assign new_new_n6518__ = ~new_new_n2421__ & ~new_new_n6043__;
  assign new_new_n6519__ = new_new_n2224__ & ~new_new_n6518__;
  assign new_new_n6520__ = ~new_new_n2224__ & new_new_n6518__;
  assign new_new_n6521__ = ~new_new_n6519__ & ~new_new_n6520__;
  assign new_new_n6522__ = ~new_new_n2024__ & ~new_new_n2420__;
  assign new_new_n6523__ = ~new_new_n6521__ & new_new_n6522__;
  assign new_new_n6524__ = ~new_new_n71__ & ~new_new_n6523__;
  assign new_new_n6525__ = ~new_new_n161__ & new_new_n2224__;
  assign new_new_n6526__ = ~new_new_n6524__ & new_new_n6525__;
  assign new_new_n6527__ = ~new_new_n2024__ & ~new_new_n2224__;
  assign new_new_n6528__ = ~new_new_n6518__ & new_new_n6527__;
  assign new_new_n6529__ = ~new_new_n161__ & ~new_new_n6528__;
  assign new_new_n6530__ = ~new_new_n71__ & new_new_n2420__;
  assign new_new_n6531__ = ~new_new_n6529__ & new_new_n6530__;
  assign new_new_n6532__ = ~new_new_n6517__ & ~new_new_n6531__;
  assign new_new_n6533__ = ~new_new_n6526__ & new_new_n6532__;
  assign new_new_n6534__ = pi31 & ~new_new_n6533__;
  assign new_new_n6535__ = new_new_n765__ & ~new_new_n2024__;
  assign new_new_n6536__ = ~pi31 & ~new_new_n6011__;
  assign new_new_n6537__ = ~new_new_n6535__ & new_new_n6536__;
  assign new_new_n6538__ = ~new_new_n6534__ & ~new_new_n6537__;
  assign new_new_n6539__ = ~new_new_n6511__ & ~new_new_n6538__;
  assign new_new_n6540__ = new_new_n6511__ & new_new_n6538__;
  assign new_new_n6541__ = ~new_new_n2130__ & ~new_new_n4818__;
  assign new_new_n6542__ = ~new_new_n3535__ & new_new_n4212__;
  assign new_new_n6543__ = ~new_new_n6541__ & ~new_new_n6542__;
  assign new_new_n6544__ = new_new_n4214__ & ~new_new_n5520__;
  assign new_new_n6545__ = pi29 & ~new_new_n6544__;
  assign new_new_n6546__ = ~pi28 & new_new_n1823__;
  assign new_new_n6547__ = pi28 & ~new_new_n1823__;
  assign new_new_n6548__ = new_new_n4214__ & ~new_new_n6546__;
  assign new_new_n6549__ = ~new_new_n6547__ & new_new_n6548__;
  assign new_new_n6550__ = new_new_n5501__ & new_new_n6549__;
  assign new_new_n6551__ = ~new_new_n6545__ & ~new_new_n6550__;
  assign new_new_n6552__ = new_new_n6543__ & ~new_new_n6551__;
  assign new_new_n6553__ = ~new_new_n1823__ & ~new_new_n5501__;
  assign new_new_n6554__ = new_new_n4214__ & new_new_n6553__;
  assign new_new_n6555__ = new_new_n6543__ & ~new_new_n6554__;
  assign new_new_n6556__ = ~pi29 & ~new_new_n6555__;
  assign new_new_n6557__ = ~new_new_n6552__ & ~new_new_n6556__;
  assign new_new_n6558__ = ~new_new_n6540__ & new_new_n6557__;
  assign new_new_n6559__ = ~new_new_n6539__ & ~new_new_n6558__;
  assign new_new_n6560__ = ~new_new_n6500__ & ~new_new_n6559__;
  assign new_new_n6561__ = ~new_new_n6499__ & ~new_new_n6560__;
  assign new_new_n6562__ = ~new_new_n6369__ & ~new_new_n6378__;
  assign new_new_n6563__ = new_new_n6436__ & ~new_new_n6562__;
  assign new_new_n6564__ = ~new_new_n6436__ & new_new_n6562__;
  assign new_new_n6565__ = ~new_new_n6563__ & ~new_new_n6564__;
  assign new_new_n6566__ = new_new_n5451__ & new_new_n6565__;
  assign new_new_n6567__ = ~new_new_n5451__ & ~new_new_n6565__;
  assign new_new_n6568__ = ~new_new_n6566__ & ~new_new_n6567__;
  assign new_new_n6569__ = ~new_new_n1556__ & new_new_n3311__;
  assign new_new_n6570__ = ~new_new_n333__ & ~new_new_n1737__;
  assign new_new_n6571__ = new_new_n873__ & ~new_new_n1466__;
  assign new_new_n6572__ = ~new_new_n4900__ & ~new_new_n5671__;
  assign new_new_n6573__ = ~new_new_n6569__ & ~new_new_n6570__;
  assign new_new_n6574__ = ~new_new_n6571__ & new_new_n6573__;
  assign new_new_n6575__ = ~new_new_n6572__ & new_new_n6574__;
  assign new_new_n6576__ = pi26 & ~new_new_n6575__;
  assign new_new_n6577__ = ~pi26 & new_new_n6575__;
  assign new_new_n6578__ = ~new_new_n6576__ & ~new_new_n6577__;
  assign new_new_n6579__ = new_new_n6568__ & new_new_n6578__;
  assign new_new_n6580__ = ~new_new_n6568__ & ~new_new_n6578__;
  assign new_new_n6581__ = ~new_new_n6579__ & ~new_new_n6580__;
  assign new_new_n6582__ = ~new_new_n6561__ & ~new_new_n6581__;
  assign new_new_n6583__ = new_new_n6568__ & ~new_new_n6578__;
  assign new_new_n6584__ = ~new_new_n6582__ & ~new_new_n6583__;
  assign new_new_n6585__ = ~new_new_n1207__ & new_new_n5213__;
  assign new_new_n6586__ = ~new_new_n3618__ & new_new_n5191__;
  assign new_new_n6587__ = ~new_new_n1061__ & new_new_n5183__;
  assign new_new_n6588__ = ~new_new_n6585__ & ~new_new_n6586__;
  assign new_new_n6589__ = ~new_new_n6587__ & new_new_n6588__;
  assign new_new_n6590__ = new_new_n5195__ & ~new_new_n5235__;
  assign new_new_n6591__ = ~pi23 & ~new_new_n6590__;
  assign new_new_n6592__ = ~new_new_n5235__ & new_new_n5974__;
  assign new_new_n6593__ = ~new_new_n6591__ & ~new_new_n6592__;
  assign new_new_n6594__ = new_new_n6589__ & ~new_new_n6593__;
  assign new_new_n6595__ = pi23 & ~new_new_n6589__;
  assign new_new_n6596__ = ~new_new_n6594__ & ~new_new_n6595__;
  assign new_new_n6597__ = new_new_n6584__ & new_new_n6596__;
  assign new_new_n6598__ = ~new_new_n6584__ & ~new_new_n6596__;
  assign new_new_n6599__ = new_new_n4214__ & new_new_n5688__;
  assign new_new_n6600__ = pi28 & ~new_new_n6458__;
  assign new_new_n6601__ = ~pi28 & new_new_n6458__;
  assign new_new_n6602__ = ~new_new_n6600__ & ~new_new_n6601__;
  assign new_new_n6603__ = new_new_n6599__ & ~new_new_n6602__;
  assign new_new_n6604__ = ~pi29 & ~new_new_n6458__;
  assign new_new_n6605__ = pi29 & new_new_n6458__;
  assign new_new_n6606__ = ~new_new_n6604__ & ~new_new_n6605__;
  assign new_new_n6607__ = ~new_new_n6599__ & new_new_n6606__;
  assign new_new_n6608__ = ~new_new_n6603__ & ~new_new_n6607__;
  assign new_new_n6609__ = new_new_n6465__ & ~new_new_n6608__;
  assign new_new_n6610__ = ~new_new_n6465__ & ~new_new_n6606__;
  assign new_new_n6611__ = ~new_new_n6609__ & ~new_new_n6610__;
  assign new_new_n6612__ = new_new_n6435__ & ~new_new_n6611__;
  assign new_new_n6613__ = ~new_new_n6435__ & new_new_n6611__;
  assign new_new_n6614__ = ~new_new_n6612__ & ~new_new_n6613__;
  assign new_new_n6615__ = ~new_new_n6598__ & new_new_n6614__;
  assign new_new_n6616__ = ~new_new_n6597__ & ~new_new_n6615__;
  assign new_new_n6617__ = ~new_new_n6477__ & new_new_n6616__;
  assign new_new_n6618__ = ~new_new_n6476__ & ~new_new_n6617__;
  assign new_new_n6619__ = pi17 & pi18;
  assign new_new_n6620__ = pi19 & ~pi20;
  assign new_new_n6621__ = new_new_n6619__ & new_new_n6620__;
  assign new_new_n6622__ = ~pi17 & ~pi18;
  assign new_new_n6623__ = ~pi19 & new_new_n6622__;
  assign new_new_n6624__ = pi20 & new_new_n6623__;
  assign new_new_n6625__ = ~new_new_n6621__ & ~new_new_n6624__;
  assign new_new_n6626__ = ~new_new_n910__ & ~new_new_n6625__;
  assign new_new_n6627__ = pi19 & ~new_new_n6622__;
  assign new_new_n6628__ = ~pi19 & ~new_new_n6619__;
  assign new_new_n6629__ = ~new_new_n6627__ & ~new_new_n6628__;
  assign new_new_n6630__ = ~new_new_n691__ & new_new_n6629__;
  assign new_new_n6631__ = ~new_new_n6619__ & ~new_new_n6622__;
  assign new_new_n6632__ = ~pi19 & pi20;
  assign new_new_n6633__ = ~new_new_n6620__ & ~new_new_n6632__;
  assign new_new_n6634__ = new_new_n6631__ & new_new_n6633__;
  assign new_new_n6635__ = ~new_new_n583__ & new_new_n6634__;
  assign new_new_n6636__ = ~new_new_n6630__ & ~new_new_n6635__;
  assign new_new_n6637__ = ~new_new_n6626__ & new_new_n6636__;
  assign new_new_n6638__ = new_new_n3742__ & new_new_n6631__;
  assign new_new_n6639__ = pi20 & ~new_new_n6638__;
  assign new_new_n6640__ = pi19 & new_new_n6631__;
  assign new_new_n6641__ = new_new_n3742__ & new_new_n6640__;
  assign new_new_n6642__ = ~new_new_n6639__ & ~new_new_n6641__;
  assign new_new_n6643__ = new_new_n6637__ & ~new_new_n6642__;
  assign new_new_n6644__ = ~pi20 & ~new_new_n6637__;
  assign new_new_n6645__ = ~new_new_n6643__ & ~new_new_n6644__;
  assign new_new_n6646__ = new_new_n6618__ & ~new_new_n6645__;
  assign new_new_n6647__ = ~new_new_n6618__ & new_new_n6645__;
  assign new_new_n6648__ = ~new_new_n6646__ & ~new_new_n6647__;
  assign new_new_n6649__ = new_new_n873__ & ~new_new_n3618__;
  assign new_new_n6650__ = ~new_new_n1061__ & new_new_n3311__;
  assign new_new_n6651__ = ~new_new_n333__ & ~new_new_n1325__;
  assign new_new_n6652__ = ~new_new_n6649__ & ~new_new_n6650__;
  assign new_new_n6653__ = ~new_new_n6651__ & new_new_n6652__;
  assign new_new_n6654__ = pi26 & ~new_new_n6653__;
  assign new_new_n6655__ = new_new_n4898__ & new_new_n4926__;
  assign new_new_n6656__ = new_new_n801__ & new_new_n4926__;
  assign new_new_n6657__ = ~pi26 & ~new_new_n6656__;
  assign new_new_n6658__ = ~new_new_n6655__ & ~new_new_n6657__;
  assign new_new_n6659__ = new_new_n6653__ & ~new_new_n6658__;
  assign new_new_n6660__ = ~new_new_n6654__ & ~new_new_n6659__;
  assign new_new_n6661__ = ~new_new_n6405__ & ~new_new_n6417__;
  assign new_new_n6662__ = ~new_new_n6404__ & ~new_new_n6661__;
  assign new_new_n6663__ = ~new_new_n5653__ & ~new_new_n5654__;
  assign new_new_n6664__ = new_new_n5678__ & new_new_n6663__;
  assign new_new_n6665__ = ~new_new_n5678__ & ~new_new_n6663__;
  assign new_new_n6666__ = ~new_new_n6664__ & ~new_new_n6665__;
  assign new_new_n6667__ = ~new_new_n6662__ & ~new_new_n6666__;
  assign new_new_n6668__ = new_new_n6662__ & new_new_n6666__;
  assign new_new_n6669__ = ~new_new_n6667__ & ~new_new_n6668__;
  assign new_new_n6670__ = new_new_n6660__ & ~new_new_n6669__;
  assign new_new_n6671__ = ~new_new_n6660__ & new_new_n6669__;
  assign new_new_n6672__ = ~new_new_n6670__ & ~new_new_n6671__;
  assign new_new_n6673__ = ~new_new_n868__ & new_new_n5183__;
  assign new_new_n6674__ = ~new_new_n4032__ & new_new_n5212__;
  assign new_new_n6675__ = new_new_n3720__ & ~new_new_n6674__;
  assign new_new_n6676__ = ~new_new_n3720__ & new_new_n6674__;
  assign new_new_n6677__ = new_new_n5195__ & ~new_new_n6675__;
  assign new_new_n6678__ = ~new_new_n6676__ & new_new_n6677__;
  assign new_new_n6679__ = ~new_new_n6673__ & ~new_new_n6678__;
  assign new_new_n6680__ = ~new_new_n1207__ & new_new_n5185__;
  assign new_new_n6681__ = pi23 & ~new_new_n6680__;
  assign new_new_n6682__ = ~new_new_n1207__ & new_new_n5188__;
  assign new_new_n6683__ = ~pi23 & ~new_new_n6682__;
  assign new_new_n6684__ = pi20 & ~new_new_n6683__;
  assign new_new_n6685__ = ~new_new_n6681__ & ~new_new_n6684__;
  assign new_new_n6686__ = new_new_n6679__ & ~new_new_n6685__;
  assign new_new_n6687__ = ~pi23 & ~new_new_n6679__;
  assign new_new_n6688__ = ~new_new_n6686__ & ~new_new_n6687__;
  assign new_new_n6689__ = ~new_new_n6421__ & new_new_n6472__;
  assign new_new_n6690__ = ~new_new_n6422__ & ~new_new_n6689__;
  assign new_new_n6691__ = ~new_new_n6688__ & new_new_n6690__;
  assign new_new_n6692__ = new_new_n6688__ & ~new_new_n6690__;
  assign new_new_n6693__ = ~new_new_n6691__ & ~new_new_n6692__;
  assign new_new_n6694__ = new_new_n6672__ & new_new_n6693__;
  assign new_new_n6695__ = ~new_new_n6672__ & ~new_new_n6693__;
  assign new_new_n6696__ = ~new_new_n6694__ & ~new_new_n6695__;
  assign new_new_n6697__ = new_new_n6648__ & ~new_new_n6696__;
  assign new_new_n6698__ = ~new_new_n6648__ & new_new_n6696__;
  assign new_new_n6699__ = ~new_new_n6697__ & ~new_new_n6698__;
  assign new_new_n6700__ = ~new_new_n6476__ & ~new_new_n6477__;
  assign new_new_n6701__ = ~new_new_n6616__ & new_new_n6700__;
  assign new_new_n6702__ = new_new_n6616__ & ~new_new_n6700__;
  assign new_new_n6703__ = ~new_new_n6701__ & ~new_new_n6702__;
  assign new_new_n6704__ = ~new_new_n3720__ & new_new_n6629__;
  assign new_new_n6705__ = ~new_new_n868__ & ~new_new_n6625__;
  assign new_new_n6706__ = ~new_new_n6704__ & ~new_new_n6705__;
  assign new_new_n6707__ = ~new_new_n5129__ & new_new_n6631__;
  assign new_new_n6708__ = pi20 & ~new_new_n6707__;
  assign new_new_n6709__ = ~pi19 & new_new_n910__;
  assign new_new_n6710__ = pi19 & ~new_new_n910__;
  assign new_new_n6711__ = new_new_n6631__ & ~new_new_n6709__;
  assign new_new_n6712__ = ~new_new_n6710__ & new_new_n6711__;
  assign new_new_n6713__ = new_new_n4036__ & new_new_n6712__;
  assign new_new_n6714__ = ~new_new_n6708__ & ~new_new_n6713__;
  assign new_new_n6715__ = new_new_n6706__ & ~new_new_n6714__;
  assign new_new_n6716__ = new_new_n5116__ & new_new_n6631__;
  assign new_new_n6717__ = new_new_n6706__ & ~new_new_n6716__;
  assign new_new_n6718__ = ~pi20 & ~new_new_n6717__;
  assign new_new_n6719__ = ~new_new_n6715__ & ~new_new_n6718__;
  assign new_new_n6720__ = new_new_n6561__ & new_new_n6581__;
  assign new_new_n6721__ = ~new_new_n6582__ & ~new_new_n6720__;
  assign new_new_n6722__ = ~new_new_n3618__ & new_new_n5183__;
  assign new_new_n6723__ = ~new_new_n1325__ & new_new_n5191__;
  assign new_new_n6724__ = ~new_new_n1061__ & new_new_n5213__;
  assign new_new_n6725__ = ~new_new_n6722__ & ~new_new_n6723__;
  assign new_new_n6726__ = ~new_new_n6724__ & new_new_n6725__;
  assign new_new_n6727__ = new_new_n4926__ & new_new_n5195__;
  assign new_new_n6728__ = ~pi23 & ~new_new_n6727__;
  assign new_new_n6729__ = new_new_n4926__ & new_new_n5974__;
  assign new_new_n6730__ = ~new_new_n6728__ & ~new_new_n6729__;
  assign new_new_n6731__ = new_new_n6726__ & ~new_new_n6730__;
  assign new_new_n6732__ = pi23 & ~new_new_n6726__;
  assign new_new_n6733__ = ~new_new_n6731__ & ~new_new_n6732__;
  assign new_new_n6734__ = new_new_n6721__ & ~new_new_n6733__;
  assign new_new_n6735__ = ~new_new_n6721__ & new_new_n6733__;
  assign new_new_n6736__ = ~new_new_n6499__ & ~new_new_n6500__;
  assign new_new_n6737__ = new_new_n6559__ & ~new_new_n6736__;
  assign new_new_n6738__ = ~new_new_n6559__ & new_new_n6736__;
  assign new_new_n6739__ = ~new_new_n6737__ & ~new_new_n6738__;
  assign new_new_n6740__ = new_new_n161__ & ~new_new_n2313__;
  assign new_new_n6741__ = new_new_n765__ & ~new_new_n2420__;
  assign new_new_n6742__ = ~new_new_n6740__ & ~new_new_n6741__;
  assign new_new_n6743__ = ~pi31 & ~new_new_n6742__;
  assign new_new_n6744__ = new_new_n161__ & ~new_new_n2572__;
  assign new_new_n6745__ = new_new_n71__ & ~new_new_n2313__;
  assign new_new_n6746__ = ~new_new_n6744__ & ~new_new_n6745__;
  assign new_new_n6747__ = pi31 & ~new_new_n6746__;
  assign new_new_n6748__ = ~new_new_n3475__ & ~new_new_n6052__;
  assign new_new_n6749__ = ~new_new_n2420__ & ~new_new_n6748__;
  assign new_new_n6750__ = new_new_n2420__ & new_new_n6748__;
  assign new_new_n6751__ = ~new_new_n6749__ & ~new_new_n6750__;
  assign new_new_n6752__ = ~pi31 & new_new_n2420__;
  assign new_new_n6753__ = new_new_n765__ & ~new_new_n6752__;
  assign new_new_n6754__ = ~new_new_n6751__ & new_new_n6753__;
  assign new_new_n6755__ = ~new_new_n6743__ & ~new_new_n6747__;
  assign new_new_n6756__ = ~new_new_n6754__ & new_new_n6755__;
  assign new_new_n6757__ = ~new_new_n247__ & ~new_new_n258__;
  assign new_new_n6758__ = ~new_new_n472__ & ~new_new_n482__;
  assign new_new_n6759__ = ~new_new_n88__ & ~new_new_n96__;
  assign new_new_n6760__ = ~new_new_n212__ & ~new_new_n249__;
  assign new_new_n6761__ = ~new_new_n312__ & ~new_new_n768__;
  assign new_new_n6762__ = new_new_n6760__ & new_new_n6761__;
  assign new_new_n6763__ = ~new_new_n732__ & new_new_n6759__;
  assign new_new_n6764__ = new_new_n2158__ & new_new_n6758__;
  assign new_new_n6765__ = new_new_n6763__ & new_new_n6764__;
  assign new_new_n6766__ = new_new_n849__ & new_new_n6762__;
  assign new_new_n6767__ = new_new_n1905__ & new_new_n3057__;
  assign new_new_n6768__ = new_new_n6757__ & new_new_n6767__;
  assign new_new_n6769__ = new_new_n6765__ & new_new_n6766__;
  assign new_new_n6770__ = new_new_n4596__ & new_new_n5384__;
  assign new_new_n6771__ = new_new_n6769__ & new_new_n6770__;
  assign new_new_n6772__ = new_new_n6768__ & new_new_n6771__;
  assign new_new_n6773__ = ~new_new_n76__ & ~new_new_n92__;
  assign new_new_n6774__ = ~new_new_n692__ & ~new_new_n933__;
  assign new_new_n6775__ = ~new_new_n1033__ & new_new_n6774__;
  assign new_new_n6776__ = ~new_new_n675__ & new_new_n6773__;
  assign new_new_n6777__ = ~new_new_n1166__ & new_new_n6185__;
  assign new_new_n6778__ = new_new_n6776__ & new_new_n6777__;
  assign new_new_n6779__ = ~new_new_n676__ & new_new_n6775__;
  assign new_new_n6780__ = new_new_n1253__ & new_new_n5695__;
  assign new_new_n6781__ = new_new_n6779__ & new_new_n6780__;
  assign new_new_n6782__ = new_new_n1803__ & new_new_n6778__;
  assign new_new_n6783__ = new_new_n2990__ & new_new_n6782__;
  assign new_new_n6784__ = new_new_n6154__ & new_new_n6781__;
  assign new_new_n6785__ = new_new_n6239__ & new_new_n6784__;
  assign new_new_n6786__ = new_new_n1353__ & new_new_n6783__;
  assign new_new_n6787__ = new_new_n6785__ & new_new_n6786__;
  assign new_new_n6788__ = new_new_n6772__ & new_new_n6787__;
  assign new_new_n6789__ = new_new_n4364__ & new_new_n6788__;
  assign new_new_n6790__ = ~new_new_n2497__ & new_new_n5053__;
  assign new_new_n6791__ = ~new_new_n2636__ & new_new_n5059__;
  assign new_new_n6792__ = ~pi31 & new_new_n2572__;
  assign new_new_n6793__ = new_new_n2737__ & ~new_new_n3468__;
  assign new_new_n6794__ = ~new_new_n2636__ & new_new_n6793__;
  assign new_new_n6795__ = ~new_new_n2737__ & new_new_n3468__;
  assign new_new_n6796__ = new_new_n2636__ & new_new_n6795__;
  assign new_new_n6797__ = ~new_new_n6794__ & ~new_new_n6796__;
  assign new_new_n6798__ = ~new_new_n2497__ & new_new_n2636__;
  assign new_new_n6799__ = new_new_n2497__ & ~new_new_n2636__;
  assign new_new_n6800__ = ~new_new_n6798__ & ~new_new_n6799__;
  assign new_new_n6801__ = new_new_n6797__ & ~new_new_n6800__;
  assign new_new_n6802__ = new_new_n2572__ & ~new_new_n6801__;
  assign new_new_n6803__ = ~new_new_n2572__ & new_new_n6801__;
  assign new_new_n6804__ = ~new_new_n6802__ & ~new_new_n6803__;
  assign new_new_n6805__ = pi31 & ~new_new_n6804__;
  assign new_new_n6806__ = new_new_n765__ & ~new_new_n6792__;
  assign new_new_n6807__ = ~new_new_n6805__ & new_new_n6806__;
  assign new_new_n6808__ = ~new_new_n6790__ & ~new_new_n6791__;
  assign new_new_n6809__ = ~new_new_n6807__ & new_new_n6808__;
  assign new_new_n6810__ = ~pi02 & ~pi05;
  assign new_new_n6811__ = pi02 & pi05;
  assign new_new_n6812__ = ~new_new_n229__ & ~new_new_n768__;
  assign new_new_n6813__ = ~new_new_n148__ & new_new_n6812__;
  assign new_new_n6814__ = ~new_new_n952__ & new_new_n1069__;
  assign new_new_n6815__ = new_new_n6813__ & new_new_n6814__;
  assign new_new_n6816__ = ~new_new_n837__ & new_new_n1401__;
  assign new_new_n6817__ = new_new_n6815__ & new_new_n6816__;
  assign new_new_n6818__ = ~new_new_n120__ & ~new_new_n267__;
  assign new_new_n6819__ = ~new_new_n335__ & ~new_new_n384__;
  assign new_new_n6820__ = ~new_new_n785__ & ~new_new_n950__;
  assign new_new_n6821__ = ~new_new_n1398__ & new_new_n6820__;
  assign new_new_n6822__ = new_new_n6818__ & new_new_n6819__;
  assign new_new_n6823__ = new_new_n672__ & ~new_new_n1073__;
  assign new_new_n6824__ = new_new_n2100__ & new_new_n6823__;
  assign new_new_n6825__ = new_new_n6821__ & new_new_n6822__;
  assign new_new_n6826__ = new_new_n1145__ & new_new_n4732__;
  assign new_new_n6827__ = new_new_n6825__ & new_new_n6826__;
  assign new_new_n6828__ = new_new_n1131__ & new_new_n6824__;
  assign new_new_n6829__ = ~new_new_n1539__ & new_new_n6828__;
  assign new_new_n6830__ = new_new_n1040__ & new_new_n6827__;
  assign new_new_n6831__ = new_new_n6817__ & new_new_n6830__;
  assign new_new_n6832__ = new_new_n1019__ & new_new_n6829__;
  assign new_new_n6833__ = new_new_n6831__ & new_new_n6832__;
  assign new_new_n6834__ = new_new_n3981__ & new_new_n6833__;
  assign new_new_n6835__ = new_new_n5337__ & new_new_n6834__;
  assign new_new_n6836__ = ~new_new_n6811__ & ~new_new_n6835__;
  assign new_new_n6837__ = ~new_new_n6810__ & ~new_new_n6836__;
  assign new_new_n6838__ = new_new_n6789__ & new_new_n6837__;
  assign new_new_n6839__ = new_new_n6809__ & new_new_n6838__;
  assign new_new_n6840__ = new_new_n6286__ & ~new_new_n6839__;
  assign new_new_n6841__ = ~new_new_n6789__ & ~new_new_n6809__;
  assign new_new_n6842__ = ~new_new_n6837__ & new_new_n6841__;
  assign new_new_n6843__ = ~new_new_n6840__ & ~new_new_n6842__;
  assign new_new_n6844__ = new_new_n6756__ & new_new_n6843__;
  assign new_new_n6845__ = ~new_new_n2130__ & new_new_n4212__;
  assign new_new_n6846__ = ~new_new_n3535__ & new_new_n4815__;
  assign new_new_n6847__ = ~new_new_n2024__ & ~new_new_n4818__;
  assign new_new_n6848__ = ~new_new_n6845__ & ~new_new_n6846__;
  assign new_new_n6849__ = ~new_new_n6847__ & new_new_n6848__;
  assign new_new_n6850__ = new_new_n3535__ & ~new_new_n5500__;
  assign new_new_n6851__ = ~new_new_n2097__ & new_new_n3479__;
  assign new_new_n6852__ = new_new_n5500__ & ~new_new_n6851__;
  assign new_new_n6853__ = ~new_new_n3535__ & new_new_n6852__;
  assign new_new_n6854__ = ~new_new_n6850__ & ~new_new_n6853__;
  assign new_new_n6855__ = new_new_n4214__ & new_new_n6854__;
  assign new_new_n6856__ = ~pi29 & ~new_new_n6855__;
  assign new_new_n6857__ = new_new_n5732__ & new_new_n6854__;
  assign new_new_n6858__ = ~new_new_n6856__ & ~new_new_n6857__;
  assign new_new_n6859__ = new_new_n6849__ & ~new_new_n6858__;
  assign new_new_n6860__ = pi29 & ~new_new_n6849__;
  assign new_new_n6861__ = ~new_new_n6859__ & ~new_new_n6860__;
  assign new_new_n6862__ = new_new_n6844__ & new_new_n6861__;
  assign new_new_n6863__ = ~new_new_n6844__ & ~new_new_n6861__;
  assign new_new_n6864__ = pi08 & ~new_new_n6863__;
  assign new_new_n6865__ = ~new_new_n6287__ & ~new_new_n6288__;
  assign new_new_n6866__ = ~new_new_n6756__ & ~new_new_n6843__;
  assign new_new_n6867__ = new_new_n6861__ & ~new_new_n6866__;
  assign new_new_n6868__ = ~pi08 & ~new_new_n6867__;
  assign new_new_n6869__ = ~new_new_n6864__ & new_new_n6865__;
  assign new_new_n6870__ = ~new_new_n6868__ & new_new_n6869__;
  assign new_new_n6871__ = pi08 & ~new_new_n6867__;
  assign new_new_n6872__ = ~pi08 & ~new_new_n6863__;
  assign new_new_n6873__ = ~new_new_n6865__ & ~new_new_n6871__;
  assign new_new_n6874__ = ~new_new_n6872__ & new_new_n6873__;
  assign new_new_n6875__ = ~new_new_n6861__ & new_new_n6866__;
  assign new_new_n6876__ = ~new_new_n6870__ & ~new_new_n6875__;
  assign new_new_n6877__ = ~new_new_n6874__ & new_new_n6876__;
  assign new_new_n6878__ = ~new_new_n6862__ & new_new_n6877__;
  assign new_new_n6879__ = new_new_n6290__ & new_new_n6503__;
  assign new_new_n6880__ = ~new_new_n6290__ & ~new_new_n6503__;
  assign new_new_n6881__ = ~new_new_n6879__ & ~new_new_n6880__;
  assign new_new_n6882__ = ~new_new_n6878__ & new_new_n6881__;
  assign new_new_n6883__ = ~new_new_n6861__ & new_new_n6877__;
  assign new_new_n6884__ = ~new_new_n6882__ & ~new_new_n6883__;
  assign new_new_n6885__ = ~new_new_n1737__ & new_new_n3311__;
  assign new_new_n6886__ = ~new_new_n333__ & ~new_new_n1902__;
  assign new_new_n6887__ = new_new_n873__ & ~new_new_n1660__;
  assign new_new_n6888__ = ~new_new_n4900__ & new_new_n5688__;
  assign new_new_n6889__ = ~new_new_n6885__ & ~new_new_n6886__;
  assign new_new_n6890__ = ~new_new_n6887__ & new_new_n6889__;
  assign new_new_n6891__ = ~new_new_n6888__ & new_new_n6890__;
  assign new_new_n6892__ = pi26 & ~new_new_n6891__;
  assign new_new_n6893__ = ~pi26 & new_new_n6891__;
  assign new_new_n6894__ = ~new_new_n6892__ & ~new_new_n6893__;
  assign new_new_n6895__ = ~new_new_n6884__ & ~new_new_n6894__;
  assign new_new_n6896__ = new_new_n6884__ & new_new_n6894__;
  assign new_new_n6897__ = ~new_new_n6539__ & ~new_new_n6540__;
  assign new_new_n6898__ = ~new_new_n6557__ & new_new_n6897__;
  assign new_new_n6899__ = new_new_n6557__ & ~new_new_n6897__;
  assign new_new_n6900__ = ~new_new_n6898__ & ~new_new_n6899__;
  assign new_new_n6901__ = ~new_new_n6896__ & ~new_new_n6900__;
  assign new_new_n6902__ = ~new_new_n6895__ & ~new_new_n6901__;
  assign new_new_n6903__ = new_new_n6739__ & ~new_new_n6902__;
  assign new_new_n6904__ = ~new_new_n6739__ & new_new_n6902__;
  assign new_new_n6905__ = ~new_new_n1466__ & new_new_n3311__;
  assign new_new_n6906__ = ~new_new_n333__ & ~new_new_n1660__;
  assign new_new_n6907__ = new_new_n873__ & ~new_new_n1737__;
  assign new_new_n6908__ = ~new_new_n6905__ & ~new_new_n6906__;
  assign new_new_n6909__ = ~new_new_n6907__ & new_new_n6908__;
  assign new_new_n6910__ = pi26 & ~new_new_n6909__;
  assign new_new_n6911__ = new_new_n4898__ & ~new_new_n6410__;
  assign new_new_n6912__ = new_new_n801__ & ~new_new_n6410__;
  assign new_new_n6913__ = ~pi26 & ~new_new_n6912__;
  assign new_new_n6914__ = ~new_new_n6911__ & ~new_new_n6913__;
  assign new_new_n6915__ = new_new_n6909__ & ~new_new_n6914__;
  assign new_new_n6916__ = ~new_new_n6910__ & ~new_new_n6915__;
  assign new_new_n6917__ = ~new_new_n6904__ & ~new_new_n6916__;
  assign new_new_n6918__ = ~new_new_n6903__ & ~new_new_n6917__;
  assign new_new_n6919__ = ~new_new_n6735__ & ~new_new_n6918__;
  assign new_new_n6920__ = ~new_new_n6734__ & ~new_new_n6919__;
  assign new_new_n6921__ = ~new_new_n6719__ & new_new_n6920__;
  assign new_new_n6922__ = new_new_n6719__ & ~new_new_n6920__;
  assign new_new_n6923__ = new_new_n6596__ & new_new_n6614__;
  assign new_new_n6924__ = ~new_new_n6596__ & ~new_new_n6614__;
  assign new_new_n6925__ = ~new_new_n6923__ & ~new_new_n6924__;
  assign new_new_n6926__ = ~new_new_n6584__ & new_new_n6925__;
  assign new_new_n6927__ = new_new_n6584__ & ~new_new_n6925__;
  assign new_new_n6928__ = ~new_new_n6926__ & ~new_new_n6927__;
  assign new_new_n6929__ = ~new_new_n6922__ & ~new_new_n6928__;
  assign new_new_n6930__ = ~new_new_n6921__ & ~new_new_n6929__;
  assign new_new_n6931__ = new_new_n6703__ & ~new_new_n6930__;
  assign new_new_n6932__ = ~new_new_n6703__ & new_new_n6930__;
  assign new_new_n6933__ = ~new_new_n910__ & new_new_n6629__;
  assign new_new_n6934__ = ~new_new_n3720__ & ~new_new_n6625__;
  assign new_new_n6935__ = ~new_new_n691__ & new_new_n6634__;
  assign new_new_n6936__ = new_new_n6631__ & ~new_new_n6633__;
  assign new_new_n6937__ = new_new_n4042__ & new_new_n6936__;
  assign new_new_n6938__ = ~new_new_n6934__ & ~new_new_n6935__;
  assign new_new_n6939__ = ~new_new_n6933__ & new_new_n6938__;
  assign new_new_n6940__ = ~new_new_n6937__ & new_new_n6939__;
  assign new_new_n6941__ = ~new_new_n6931__ & ~new_new_n6932__;
  assign new_new_n6942__ = pi20 & ~new_new_n6941__;
  assign new_new_n6943__ = ~pi20 & new_new_n6941__;
  assign new_new_n6944__ = ~new_new_n6942__ & ~new_new_n6943__;
  assign new_new_n6945__ = new_new_n6940__ & new_new_n6944__;
  assign new_new_n6946__ = ~new_new_n6940__ & ~new_new_n6944__;
  assign new_new_n6947__ = ~new_new_n6945__ & ~new_new_n6946__;
  assign new_new_n6948__ = ~new_new_n6932__ & ~new_new_n6947__;
  assign new_new_n6949__ = ~new_new_n6931__ & ~new_new_n6948__;
  assign new_new_n6950__ = ~new_new_n466__ & ~new_new_n4168__;
  assign new_new_n6951__ = new_new_n466__ & ~new_new_n3769__;
  assign new_new_n6952__ = ~new_new_n6950__ & ~new_new_n6951__;
  assign new_new_n6953__ = ~pi16 & ~pi17;
  assign new_new_n6954__ = pi16 & pi17;
  assign new_new_n6955__ = ~new_new_n6953__ & ~new_new_n6954__;
  assign new_new_n6956__ = ~pi14 & ~pi15;
  assign new_new_n6957__ = pi14 & pi15;
  assign new_new_n6958__ = ~new_new_n6956__ & ~new_new_n6957__;
  assign new_new_n6959__ = new_new_n6955__ & new_new_n6958__;
  assign new_new_n6960__ = new_new_n6952__ & new_new_n6959__;
  assign new_new_n6961__ = ~pi16 & new_new_n6956__;
  assign new_new_n6962__ = pi16 & new_new_n6957__;
  assign new_new_n6963__ = ~new_new_n6961__ & ~new_new_n6962__;
  assign new_new_n6964__ = new_new_n6955__ & ~new_new_n6963__;
  assign new_new_n6965__ = ~new_new_n3768__ & new_new_n6964__;
  assign new_new_n6966__ = pi16 & ~new_new_n6956__;
  assign new_new_n6967__ = ~pi16 & ~new_new_n6957__;
  assign new_new_n6968__ = ~new_new_n6966__ & ~new_new_n6967__;
  assign new_new_n6969__ = ~new_new_n466__ & new_new_n6968__;
  assign new_new_n6970__ = ~new_new_n6965__ & ~new_new_n6969__;
  assign new_new_n6971__ = ~new_new_n6960__ & new_new_n6970__;
  assign new_new_n6972__ = pi17 & ~new_new_n6971__;
  assign new_new_n6973__ = ~pi17 & new_new_n6971__;
  assign new_new_n6974__ = ~new_new_n6972__ & ~new_new_n6973__;
  assign new_new_n6975__ = new_new_n6949__ & new_new_n6974__;
  assign new_new_n6976__ = ~new_new_n6949__ & ~new_new_n6974__;
  assign new_new_n6977__ = ~new_new_n6975__ & ~new_new_n6976__;
  assign new_new_n6978__ = new_new_n6699__ & ~new_new_n6977__;
  assign new_new_n6979__ = ~new_new_n6949__ & new_new_n6974__;
  assign new_new_n6980__ = ~new_new_n6978__ & ~new_new_n6979__;
  assign new_new_n6981__ = ~pi11 & ~pi12;
  assign new_new_n6982__ = pi13 & ~new_new_n6981__;
  assign new_new_n6983__ = pi11 & pi12;
  assign new_new_n6984__ = ~pi13 & ~new_new_n6983__;
  assign new_new_n6985__ = ~new_new_n6982__ & ~new_new_n6984__;
  assign new_new_n6986__ = ~new_new_n583__ & new_new_n6985__;
  assign new_new_n6987__ = pi13 & new_new_n6983__;
  assign new_new_n6988__ = ~pi14 & ~new_new_n6987__;
  assign new_new_n6989__ = ~pi13 & new_new_n6981__;
  assign new_new_n6990__ = pi14 & ~new_new_n6989__;
  assign new_new_n6991__ = ~new_new_n6988__ & ~new_new_n6990__;
  assign new_new_n6992__ = ~new_new_n691__ & new_new_n6991__;
  assign new_new_n6993__ = ~new_new_n6986__ & ~new_new_n6992__;
  assign new_new_n6994__ = ~new_new_n6981__ & ~new_new_n6983__;
  assign new_new_n6995__ = new_new_n4142__ & new_new_n6994__;
  assign new_new_n6996__ = new_new_n6993__ & ~new_new_n6995__;
  assign new_new_n6997__ = ~pi14 & ~new_new_n6996__;
  assign new_new_n6998__ = pi13 & ~new_new_n3768__;
  assign new_new_n6999__ = ~pi13 & ~new_new_n4144__;
  assign new_new_n7000__ = new_new_n3768__ & ~new_new_n4141__;
  assign new_new_n7001__ = new_new_n6994__ & ~new_new_n7000__;
  assign new_new_n7002__ = ~new_new_n6998__ & new_new_n7001__;
  assign new_new_n7003__ = ~new_new_n6999__ & new_new_n7002__;
  assign new_new_n7004__ = pi14 & new_new_n6993__;
  assign new_new_n7005__ = ~new_new_n7001__ & new_new_n7004__;
  assign new_new_n7006__ = ~new_new_n6997__ & ~new_new_n7005__;
  assign new_new_n7007__ = ~new_new_n7003__ & new_new_n7006__;
  assign new_new_n7008__ = new_new_n4926__ & new_new_n6936__;
  assign new_new_n7009__ = ~new_new_n3618__ & new_new_n6629__;
  assign new_new_n7010__ = ~new_new_n1325__ & ~new_new_n6625__;
  assign new_new_n7011__ = ~new_new_n7009__ & ~new_new_n7010__;
  assign new_new_n7012__ = ~new_new_n7008__ & new_new_n7011__;
  assign new_new_n7013__ = ~new_new_n1061__ & new_new_n6631__;
  assign new_new_n7014__ = pi20 & ~new_new_n7013__;
  assign new_new_n7015__ = ~pi19 & new_new_n6631__;
  assign new_new_n7016__ = ~new_new_n1061__ & new_new_n7015__;
  assign new_new_n7017__ = ~new_new_n7014__ & ~new_new_n7016__;
  assign new_new_n7018__ = new_new_n7012__ & ~new_new_n7017__;
  assign new_new_n7019__ = ~pi20 & ~new_new_n7012__;
  assign new_new_n7020__ = ~new_new_n7018__ & ~new_new_n7019__;
  assign new_new_n7021__ = ~new_new_n4900__ & ~new_new_n6487__;
  assign new_new_n7022__ = ~new_new_n1902__ & new_new_n3311__;
  assign new_new_n7023__ = ~new_new_n333__ & ~new_new_n3535__;
  assign new_new_n7024__ = new_new_n873__ & ~new_new_n1823__;
  assign new_new_n7025__ = ~new_new_n7022__ & ~new_new_n7023__;
  assign new_new_n7026__ = ~new_new_n7024__ & new_new_n7025__;
  assign new_new_n7027__ = ~new_new_n7021__ & new_new_n7026__;
  assign new_new_n7028__ = pi26 & ~new_new_n7027__;
  assign new_new_n7029__ = ~pi26 & new_new_n7027__;
  assign new_new_n7030__ = ~new_new_n7028__ & ~new_new_n7029__;
  assign new_new_n7031__ = ~new_new_n2024__ & new_new_n4212__;
  assign new_new_n7032__ = ~new_new_n2130__ & new_new_n4815__;
  assign new_new_n7033__ = ~new_new_n2224__ & ~new_new_n4818__;
  assign new_new_n7034__ = ~new_new_n7031__ & ~new_new_n7032__;
  assign new_new_n7035__ = ~new_new_n7033__ & new_new_n7034__;
  assign new_new_n7036__ = new_new_n4214__ & ~new_new_n6036__;
  assign new_new_n7037__ = ~pi29 & ~new_new_n7036__;
  assign new_new_n7038__ = new_new_n5732__ & ~new_new_n6036__;
  assign new_new_n7039__ = ~new_new_n7037__ & ~new_new_n7038__;
  assign new_new_n7040__ = new_new_n7035__ & ~new_new_n7039__;
  assign new_new_n7041__ = pi29 & ~new_new_n7035__;
  assign new_new_n7042__ = ~new_new_n7040__ & ~new_new_n7041__;
  assign new_new_n7043__ = ~new_new_n2313__ & ~new_new_n4818__;
  assign new_new_n7044__ = ~new_new_n2224__ & new_new_n4815__;
  assign new_new_n7045__ = ~new_new_n2420__ & new_new_n4212__;
  assign new_new_n7046__ = ~new_new_n7043__ & ~new_new_n7044__;
  assign new_new_n7047__ = ~new_new_n7045__ & new_new_n7046__;
  assign new_new_n7048__ = new_new_n4214__ & new_new_n6521__;
  assign new_new_n7049__ = ~pi29 & ~new_new_n7048__;
  assign new_new_n7050__ = new_new_n5732__ & new_new_n6521__;
  assign new_new_n7051__ = ~new_new_n7049__ & ~new_new_n7050__;
  assign new_new_n7052__ = new_new_n7047__ & ~new_new_n7051__;
  assign new_new_n7053__ = pi29 & ~new_new_n7047__;
  assign new_new_n7054__ = ~new_new_n7052__ & ~new_new_n7053__;
  assign new_new_n7055__ = ~new_new_n2848__ & ~new_new_n3460__;
  assign new_new_n7056__ = ~new_new_n2848__ & new_new_n3361__;
  assign new_new_n7057__ = new_new_n2848__ & ~new_new_n3361__;
  assign new_new_n7058__ = ~new_new_n7056__ & ~new_new_n7057__;
  assign new_new_n7059__ = new_new_n2960__ & ~new_new_n3361__;
  assign new_new_n7060__ = ~new_new_n2960__ & new_new_n3361__;
  assign new_new_n7061__ = ~new_new_n3460__ & ~new_new_n7060__;
  assign new_new_n7062__ = ~new_new_n7059__ & ~new_new_n7061__;
  assign new_new_n7063__ = new_new_n7058__ & ~new_new_n7062__;
  assign new_new_n7064__ = ~new_new_n7058__ & new_new_n7062__;
  assign new_new_n7065__ = ~new_new_n7063__ & ~new_new_n7064__;
  assign new_new_n7066__ = new_new_n3460__ & new_new_n7065__;
  assign new_new_n7067__ = new_new_n2848__ & ~new_new_n7065__;
  assign new_new_n7068__ = ~new_new_n7066__ & ~new_new_n7067__;
  assign new_new_n7069__ = new_new_n765__ & ~new_new_n7068__;
  assign new_new_n7070__ = ~new_new_n7055__ & ~new_new_n7069__;
  assign new_new_n7071__ = ~new_new_n2886__ & ~new_new_n7070__;
  assign new_new_n7072__ = ~new_new_n71__ & ~new_new_n3460__;
  assign new_new_n7073__ = new_new_n2848__ & new_new_n2886__;
  assign new_new_n7074__ = new_new_n7065__ & new_new_n7073__;
  assign new_new_n7075__ = ~new_new_n161__ & ~new_new_n7074__;
  assign new_new_n7076__ = new_new_n7072__ & ~new_new_n7075__;
  assign new_new_n7077__ = new_new_n2886__ & ~new_new_n7065__;
  assign new_new_n7078__ = ~new_new_n71__ & ~new_new_n7077__;
  assign new_new_n7079__ = ~new_new_n161__ & ~new_new_n2848__;
  assign new_new_n7080__ = ~new_new_n7072__ & new_new_n7079__;
  assign new_new_n7081__ = ~new_new_n7078__ & new_new_n7080__;
  assign new_new_n7082__ = ~new_new_n7076__ & ~new_new_n7081__;
  assign new_new_n7083__ = ~new_new_n7071__ & new_new_n7082__;
  assign new_new_n7084__ = pi31 & ~new_new_n7083__;
  assign new_new_n7085__ = new_new_n161__ & new_new_n2848__;
  assign new_new_n7086__ = ~new_new_n71__ & ~new_new_n2886__;
  assign new_new_n7087__ = ~new_new_n161__ & ~new_new_n7086__;
  assign new_new_n7088__ = ~pi31 & ~new_new_n7085__;
  assign new_new_n7089__ = ~new_new_n7087__ & new_new_n7088__;
  assign new_new_n7090__ = ~new_new_n7084__ & ~new_new_n7089__;
  assign new_new_n7091__ = ~new_new_n277__ & ~new_new_n656__;
  assign new_new_n7092__ = new_new_n4392__ & new_new_n4465__;
  assign new_new_n7093__ = ~new_new_n247__ & ~new_new_n313__;
  assign new_new_n7094__ = ~new_new_n183__ & new_new_n7093__;
  assign new_new_n7095__ = new_new_n474__ & ~new_new_n488__;
  assign new_new_n7096__ = ~new_new_n959__ & new_new_n2176__;
  assign new_new_n7097__ = new_new_n7095__ & new_new_n7096__;
  assign new_new_n7098__ = new_new_n743__ & new_new_n7094__;
  assign new_new_n7099__ = new_new_n4995__ & new_new_n5302__;
  assign new_new_n7100__ = new_new_n7091__ & new_new_n7099__;
  assign new_new_n7101__ = new_new_n7097__ & new_new_n7098__;
  assign new_new_n7102__ = new_new_n985__ & new_new_n7101__;
  assign new_new_n7103__ = new_new_n957__ & new_new_n7100__;
  assign new_new_n7104__ = new_new_n5396__ & new_new_n7092__;
  assign new_new_n7105__ = new_new_n7103__ & new_new_n7104__;
  assign new_new_n7106__ = new_new_n3999__ & new_new_n7102__;
  assign new_new_n7107__ = new_new_n7105__ & new_new_n7106__;
  assign new_new_n7108__ = new_new_n3602__ & new_new_n7107__;
  assign new_new_n7109__ = new_new_n3237__ & new_new_n7108__;
  assign new_new_n7110__ = new_new_n7090__ & new_new_n7109__;
  assign new_new_n7111__ = ~new_new_n248__ & ~new_new_n630__;
  assign new_new_n7112__ = ~new_new_n327__ & ~new_new_n1033__;
  assign new_new_n7113__ = ~new_new_n346__ & new_new_n7112__;
  assign new_new_n7114__ = ~new_new_n1568__ & new_new_n2234__;
  assign new_new_n7115__ = new_new_n2425__ & new_new_n7114__;
  assign new_new_n7116__ = ~new_new_n124__ & new_new_n7113__;
  assign new_new_n7117__ = new_new_n567__ & new_new_n7116__;
  assign new_new_n7118__ = new_new_n985__ & new_new_n7115__;
  assign new_new_n7119__ = new_new_n1076__ & new_new_n3568__;
  assign new_new_n7120__ = new_new_n4987__ & new_new_n7111__;
  assign new_new_n7121__ = new_new_n7119__ & new_new_n7120__;
  assign new_new_n7122__ = new_new_n7117__ & new_new_n7118__;
  assign new_new_n7123__ = new_new_n7121__ & new_new_n7122__;
  assign new_new_n7124__ = new_new_n6233__ & new_new_n7123__;
  assign new_new_n7125__ = ~new_new_n260__ & ~new_new_n445__;
  assign new_new_n7126__ = ~new_new_n372__ & new_new_n7125__;
  assign new_new_n7127__ = ~new_new_n390__ & ~new_new_n632__;
  assign new_new_n7128__ = ~new_new_n696__ & ~new_new_n842__;
  assign new_new_n7129__ = new_new_n7127__ & new_new_n7128__;
  assign new_new_n7130__ = new_new_n1010__ & new_new_n7129__;
  assign new_new_n7131__ = ~new_new_n249__ & ~new_new_n425__;
  assign new_new_n7132__ = ~new_new_n937__ & new_new_n7131__;
  assign new_new_n7133__ = ~new_new_n150__ & new_new_n7132__;
  assign new_new_n7134__ = ~new_new_n607__ & new_new_n1875__;
  assign new_new_n7135__ = new_new_n3989__ & new_new_n7126__;
  assign new_new_n7136__ = new_new_n7134__ & new_new_n7135__;
  assign new_new_n7137__ = new_new_n3930__ & new_new_n7133__;
  assign new_new_n7138__ = new_new_n5474__ & new_new_n7137__;
  assign new_new_n7139__ = new_new_n7130__ & new_new_n7136__;
  assign new_new_n7140__ = new_new_n7138__ & new_new_n7139__;
  assign new_new_n7141__ = new_new_n3293__ & new_new_n3910__;
  assign new_new_n7142__ = new_new_n7140__ & new_new_n7141__;
  assign new_new_n7143__ = new_new_n3512__ & new_new_n7142__;
  assign new_new_n7144__ = new_new_n7124__ & new_new_n7143__;
  assign new_new_n7145__ = new_new_n7110__ & new_new_n7144__;
  assign new_new_n7146__ = pi02 & ~new_new_n7145__;
  assign new_new_n7147__ = ~new_new_n477__ & ~new_new_n630__;
  assign new_new_n7148__ = ~new_new_n138__ & ~new_new_n729__;
  assign new_new_n7149__ = ~new_new_n300__ & new_new_n7148__;
  assign new_new_n7150__ = ~new_new_n346__ & ~new_new_n696__;
  assign new_new_n7151__ = new_new_n1163__ & new_new_n7150__;
  assign new_new_n7152__ = new_new_n4477__ & new_new_n7149__;
  assign new_new_n7153__ = new_new_n7151__ & new_new_n7152__;
  assign new_new_n7154__ = new_new_n7147__ & new_new_n7153__;
  assign new_new_n7155__ = ~new_new_n252__ & ~new_new_n990__;
  assign new_new_n7156__ = ~new_new_n1033__ & new_new_n3397__;
  assign new_new_n7157__ = new_new_n7155__ & new_new_n7156__;
  assign new_new_n7158__ = new_new_n2643__ & new_new_n7157__;
  assign new_new_n7159__ = ~new_new_n251__ & ~new_new_n586__;
  assign new_new_n7160__ = ~new_new_n995__ & new_new_n7159__;
  assign new_new_n7161__ = ~new_new_n878__ & new_new_n4459__;
  assign new_new_n7162__ = new_new_n7160__ & new_new_n7161__;
  assign new_new_n7163__ = ~new_new_n519__ & new_new_n3989__;
  assign new_new_n7164__ = new_new_n6065__ & new_new_n7163__;
  assign new_new_n7165__ = new_new_n709__ & new_new_n7162__;
  assign new_new_n7166__ = new_new_n1076__ & new_new_n1861__;
  assign new_new_n7167__ = new_new_n6298__ & new_new_n7166__;
  assign new_new_n7168__ = new_new_n7164__ & new_new_n7165__;
  assign new_new_n7169__ = new_new_n7158__ & new_new_n7168__;
  assign new_new_n7170__ = new_new_n7154__ & new_new_n7167__;
  assign new_new_n7171__ = new_new_n7169__ & new_new_n7170__;
  assign new_new_n7172__ = new_new_n825__ & new_new_n2695__;
  assign new_new_n7173__ = new_new_n7171__ & new_new_n7172__;
  assign new_new_n7174__ = new_new_n2939__ & new_new_n7173__;
  assign new_new_n7175__ = ~new_new_n7146__ & new_new_n7174__;
  assign new_new_n7176__ = ~new_new_n7090__ & ~new_new_n7109__;
  assign new_new_n7177__ = ~new_new_n7144__ & new_new_n7176__;
  assign new_new_n7178__ = ~pi02 & ~new_new_n7177__;
  assign new_new_n7179__ = ~new_new_n7175__ & ~new_new_n7178__;
  assign new_new_n7180__ = ~new_new_n2737__ & new_new_n5059__;
  assign new_new_n7181__ = ~new_new_n2636__ & new_new_n5053__;
  assign new_new_n7182__ = pi31 & ~new_new_n6797__;
  assign new_new_n7183__ = new_new_n2497__ & ~new_new_n7182__;
  assign new_new_n7184__ = ~new_new_n2497__ & new_new_n7182__;
  assign new_new_n7185__ = new_new_n765__ & ~new_new_n7183__;
  assign new_new_n7186__ = ~new_new_n7184__ & new_new_n7185__;
  assign new_new_n7187__ = ~new_new_n7180__ & ~new_new_n7181__;
  assign new_new_n7188__ = ~new_new_n7186__ & new_new_n7187__;
  assign new_new_n7189__ = ~new_new_n7179__ & new_new_n7188__;
  assign new_new_n7190__ = new_new_n7179__ & ~new_new_n7188__;
  assign new_new_n7191__ = ~new_new_n6810__ & ~new_new_n6811__;
  assign new_new_n7192__ = new_new_n6835__ & ~new_new_n7191__;
  assign new_new_n7193__ = ~new_new_n6835__ & new_new_n7191__;
  assign new_new_n7194__ = ~new_new_n7192__ & ~new_new_n7193__;
  assign new_new_n7195__ = ~new_new_n7190__ & ~new_new_n7194__;
  assign new_new_n7196__ = ~new_new_n7189__ & ~new_new_n7195__;
  assign new_new_n7197__ = new_new_n7054__ & new_new_n7196__;
  assign new_new_n7198__ = new_new_n6809__ & ~new_new_n6837__;
  assign new_new_n7199__ = ~new_new_n6809__ & new_new_n6837__;
  assign new_new_n7200__ = ~new_new_n7198__ & ~new_new_n7199__;
  assign new_new_n7201__ = ~new_new_n6255__ & new_new_n7200__;
  assign new_new_n7202__ = ~new_new_n7054__ & ~new_new_n7196__;
  assign new_new_n7203__ = new_new_n6286__ & ~new_new_n7200__;
  assign new_new_n7204__ = ~new_new_n6286__ & new_new_n7200__;
  assign new_new_n7205__ = ~new_new_n7203__ & ~new_new_n7204__;
  assign new_new_n7206__ = ~new_new_n7201__ & new_new_n7205__;
  assign new_new_n7207__ = ~new_new_n7202__ & new_new_n7206__;
  assign new_new_n7208__ = ~new_new_n7197__ & ~new_new_n7207__;
  assign new_new_n7209__ = ~new_new_n2572__ & new_new_n5053__;
  assign new_new_n7210__ = ~new_new_n2497__ & new_new_n5059__;
  assign new_new_n7211__ = ~pi31 & new_new_n2313__;
  assign new_new_n7212__ = ~new_new_n2497__ & new_new_n2572__;
  assign new_new_n7213__ = new_new_n2313__ & new_new_n7212__;
  assign new_new_n7214__ = ~new_new_n2737__ & new_new_n7213__;
  assign new_new_n7215__ = ~new_new_n2313__ & new_new_n2497__;
  assign new_new_n7216__ = ~new_new_n2636__ & new_new_n7215__;
  assign new_new_n7217__ = ~new_new_n7214__ & ~new_new_n7216__;
  assign new_new_n7218__ = new_new_n3468__ & ~new_new_n7217__;
  assign new_new_n7219__ = new_new_n2498__ & new_new_n2636__;
  assign new_new_n7220__ = ~new_new_n2572__ & new_new_n2738__;
  assign new_new_n7221__ = ~new_new_n7219__ & ~new_new_n7220__;
  assign new_new_n7222__ = ~new_new_n3468__ & ~new_new_n7221__;
  assign new_new_n7223__ = new_new_n2498__ & new_new_n2737__;
  assign new_new_n7224__ = ~new_new_n2572__ & new_new_n2638__;
  assign new_new_n7225__ = ~new_new_n7223__ & ~new_new_n7224__;
  assign new_new_n7226__ = new_new_n2636__ & ~new_new_n7225__;
  assign new_new_n7227__ = ~new_new_n2737__ & new_new_n7215__;
  assign new_new_n7228__ = ~new_new_n7213__ & ~new_new_n7227__;
  assign new_new_n7229__ = ~new_new_n2636__ & ~new_new_n7228__;
  assign new_new_n7230__ = new_new_n2497__ & ~new_new_n2572__;
  assign new_new_n7231__ = ~new_new_n2313__ & ~new_new_n7212__;
  assign new_new_n7232__ = ~new_new_n7230__ & new_new_n7231__;
  assign new_new_n7233__ = ~new_new_n7226__ & ~new_new_n7232__;
  assign new_new_n7234__ = ~new_new_n7229__ & new_new_n7233__;
  assign new_new_n7235__ = ~new_new_n7218__ & new_new_n7234__;
  assign new_new_n7236__ = ~new_new_n7222__ & new_new_n7235__;
  assign new_new_n7237__ = pi31 & new_new_n7236__;
  assign new_new_n7238__ = new_new_n765__ & ~new_new_n7211__;
  assign new_new_n7239__ = ~new_new_n7237__ & new_new_n7238__;
  assign new_new_n7240__ = ~new_new_n7209__ & ~new_new_n7210__;
  assign new_new_n7241__ = ~new_new_n7239__ & new_new_n7240__;
  assign new_new_n7242__ = new_new_n7208__ & new_new_n7241__;
  assign new_new_n7243__ = ~new_new_n7208__ & ~new_new_n7241__;
  assign new_new_n7244__ = new_new_n6789__ & new_new_n6809__;
  assign new_new_n7245__ = ~new_new_n6841__ & ~new_new_n7244__;
  assign new_new_n7246__ = ~new_new_n6286__ & ~new_new_n7199__;
  assign new_new_n7247__ = ~new_new_n7245__ & new_new_n7246__;
  assign new_new_n7248__ = new_new_n6286__ & ~new_new_n7198__;
  assign new_new_n7249__ = new_new_n7245__ & new_new_n7248__;
  assign new_new_n7250__ = new_new_n6789__ & ~new_new_n7200__;
  assign new_new_n7251__ = ~new_new_n7247__ & ~new_new_n7249__;
  assign new_new_n7252__ = ~new_new_n7250__ & new_new_n7251__;
  assign new_new_n7253__ = ~new_new_n7243__ & ~new_new_n7252__;
  assign new_new_n7254__ = ~new_new_n7242__ & ~new_new_n7253__;
  assign new_new_n7255__ = ~new_new_n7042__ & ~new_new_n7254__;
  assign new_new_n7256__ = new_new_n7042__ & new_new_n7254__;
  assign new_new_n7257__ = ~new_new_n7255__ & ~new_new_n7256__;
  assign new_new_n7258__ = ~new_new_n6844__ & ~new_new_n6866__;
  assign new_new_n7259__ = pi08 & ~new_new_n7258__;
  assign new_new_n7260__ = ~pi08 & new_new_n7258__;
  assign new_new_n7261__ = ~new_new_n7259__ & ~new_new_n7260__;
  assign new_new_n7262__ = new_new_n6865__ & new_new_n7261__;
  assign new_new_n7263__ = ~new_new_n6865__ & ~new_new_n7261__;
  assign new_new_n7264__ = ~new_new_n7262__ & ~new_new_n7263__;
  assign new_new_n7265__ = new_new_n7257__ & ~new_new_n7264__;
  assign new_new_n7266__ = ~new_new_n7257__ & new_new_n7264__;
  assign new_new_n7267__ = ~new_new_n7265__ & ~new_new_n7266__;
  assign new_new_n7268__ = ~new_new_n333__ & ~new_new_n2130__;
  assign new_new_n7269__ = new_new_n873__ & ~new_new_n3535__;
  assign new_new_n7270__ = ~new_new_n1823__ & new_new_n3311__;
  assign new_new_n7271__ = ~new_new_n7268__ & ~new_new_n7269__;
  assign new_new_n7272__ = ~new_new_n7270__ & new_new_n7271__;
  assign new_new_n7273__ = ~new_new_n1823__ & new_new_n5501__;
  assign new_new_n7274__ = ~new_new_n5520__ & ~new_new_n7273__;
  assign new_new_n7275__ = new_new_n4898__ & new_new_n7274__;
  assign new_new_n7276__ = new_new_n801__ & new_new_n7274__;
  assign new_new_n7277__ = ~pi26 & ~new_new_n7276__;
  assign new_new_n7278__ = ~new_new_n7275__ & ~new_new_n7277__;
  assign new_new_n7279__ = new_new_n7272__ & ~new_new_n7278__;
  assign new_new_n7280__ = pi26 & ~new_new_n7272__;
  assign new_new_n7281__ = ~new_new_n7279__ & ~new_new_n7280__;
  assign new_new_n7282__ = ~new_new_n7242__ & ~new_new_n7243__;
  assign new_new_n7283__ = ~new_new_n7245__ & new_new_n7248__;
  assign new_new_n7284__ = new_new_n7245__ & new_new_n7246__;
  assign new_new_n7285__ = ~new_new_n6789__ & ~new_new_n7200__;
  assign new_new_n7286__ = ~new_new_n7283__ & ~new_new_n7284__;
  assign new_new_n7287__ = ~new_new_n7285__ & new_new_n7286__;
  assign new_new_n7288__ = ~new_new_n7282__ & ~new_new_n7287__;
  assign new_new_n7289__ = ~new_new_n7252__ & new_new_n7282__;
  assign new_new_n7290__ = ~new_new_n7288__ & ~new_new_n7289__;
  assign new_new_n7291__ = new_new_n7281__ & ~new_new_n7290__;
  assign new_new_n7292__ = ~new_new_n7281__ & new_new_n7290__;
  assign new_new_n7293__ = ~new_new_n2224__ & new_new_n4212__;
  assign new_new_n7294__ = ~new_new_n2420__ & ~new_new_n4818__;
  assign new_new_n7295__ = ~new_new_n2024__ & new_new_n4815__;
  assign new_new_n7296__ = new_new_n2024__ & new_new_n2224__;
  assign new_new_n7297__ = new_new_n6527__ & new_new_n6748__;
  assign new_new_n7298__ = ~new_new_n7296__ & ~new_new_n7297__;
  assign new_new_n7299__ = new_new_n2420__ & ~new_new_n7298__;
  assign new_new_n7300__ = new_new_n2420__ & new_new_n6527__;
  assign new_new_n7301__ = ~new_new_n3474__ & new_new_n7296__;
  assign new_new_n7302__ = ~new_new_n7300__ & ~new_new_n7301__;
  assign new_new_n7303__ = new_new_n2313__ & ~new_new_n7302__;
  assign new_new_n7304__ = new_new_n3474__ & new_new_n6013__;
  assign new_new_n7305__ = ~new_new_n6020__ & ~new_new_n7304__;
  assign new_new_n7306__ = ~new_new_n2420__ & ~new_new_n7305__;
  assign new_new_n7307__ = ~new_new_n2420__ & new_new_n6013__;
  assign new_new_n7308__ = new_new_n3474__ & new_new_n6020__;
  assign new_new_n7309__ = ~new_new_n7307__ & ~new_new_n7308__;
  assign new_new_n7310__ = ~new_new_n2313__ & ~new_new_n7309__;
  assign new_new_n7311__ = ~new_new_n7303__ & ~new_new_n7306__;
  assign new_new_n7312__ = ~new_new_n7310__ & new_new_n7311__;
  assign new_new_n7313__ = ~new_new_n7299__ & new_new_n7312__;
  assign new_new_n7314__ = new_new_n4813__ & new_new_n7313__;
  assign new_new_n7315__ = ~new_new_n7293__ & ~new_new_n7294__;
  assign new_new_n7316__ = ~new_new_n7295__ & new_new_n7315__;
  assign new_new_n7317__ = ~new_new_n7314__ & new_new_n7316__;
  assign new_new_n7318__ = pi29 & ~new_new_n7317__;
  assign new_new_n7319__ = ~pi29 & new_new_n7317__;
  assign new_new_n7320__ = ~new_new_n7318__ & ~new_new_n7319__;
  assign new_new_n7321__ = ~new_new_n7292__ & new_new_n7320__;
  assign new_new_n7322__ = ~new_new_n7291__ & ~new_new_n7321__;
  assign new_new_n7323__ = ~new_new_n7267__ & ~new_new_n7322__;
  assign new_new_n7324__ = new_new_n7267__ & new_new_n7322__;
  assign new_new_n7325__ = ~new_new_n7323__ & ~new_new_n7324__;
  assign new_new_n7326__ = new_new_n7030__ & ~new_new_n7325__;
  assign new_new_n7327__ = ~new_new_n7030__ & new_new_n7325__;
  assign new_new_n7328__ = ~new_new_n7326__ & ~new_new_n7327__;
  assign new_new_n7329__ = ~new_new_n4900__ & new_new_n6854__;
  assign new_new_n7330__ = ~new_new_n333__ & ~new_new_n2024__;
  assign new_new_n7331__ = new_new_n873__ & ~new_new_n2130__;
  assign new_new_n7332__ = ~new_new_n7330__ & ~new_new_n7331__;
  assign new_new_n7333__ = ~new_new_n7329__ & new_new_n7332__;
  assign new_new_n7334__ = ~pi26 & ~new_new_n7333__;
  assign new_new_n7335__ = ~new_new_n3535__ & new_new_n4898__;
  assign new_new_n7336__ = new_new_n801__ & ~new_new_n3535__;
  assign new_new_n7337__ = pi26 & ~new_new_n7336__;
  assign new_new_n7338__ = ~new_new_n7335__ & ~new_new_n7337__;
  assign new_new_n7339__ = new_new_n7333__ & ~new_new_n7338__;
  assign new_new_n7340__ = ~new_new_n7334__ & ~new_new_n7339__;
  assign new_new_n7341__ = ~new_new_n7197__ & new_new_n7207__;
  assign new_new_n7342__ = ~new_new_n7197__ & ~new_new_n7202__;
  assign new_new_n7343__ = ~new_new_n7205__ & ~new_new_n7342__;
  assign new_new_n7344__ = ~new_new_n7341__ & ~new_new_n7343__;
  assign new_new_n7345__ = ~new_new_n7146__ & ~new_new_n7178__;
  assign new_new_n7346__ = new_new_n7174__ & ~new_new_n7345__;
  assign new_new_n7347__ = ~new_new_n7174__ & new_new_n7345__;
  assign new_new_n7348__ = ~new_new_n7346__ & ~new_new_n7347__;
  assign new_new_n7349__ = new_new_n765__ & ~new_new_n2737__;
  assign new_new_n7350__ = new_new_n161__ & ~new_new_n2886__;
  assign new_new_n7351__ = ~new_new_n7349__ & ~new_new_n7350__;
  assign new_new_n7352__ = ~pi31 & ~new_new_n7351__;
  assign new_new_n7353__ = new_new_n71__ & new_new_n2886__;
  assign new_new_n7354__ = new_new_n2849__ & new_new_n3460__;
  assign new_new_n7355__ = ~new_new_n2886__ & new_new_n2961__;
  assign new_new_n7356__ = new_new_n3361__ & new_new_n7355__;
  assign new_new_n7357__ = ~new_new_n7354__ & ~new_new_n7356__;
  assign new_new_n7358__ = new_new_n2960__ & ~new_new_n7357__;
  assign new_new_n7359__ = ~new_new_n2848__ & ~new_new_n2886__;
  assign new_new_n7360__ = ~new_new_n7073__ & ~new_new_n7359__;
  assign new_new_n7361__ = ~new_new_n2737__ & ~new_new_n7360__;
  assign new_new_n7362__ = ~new_new_n2737__ & new_new_n2848__;
  assign new_new_n7363__ = ~new_new_n3460__ & new_new_n7362__;
  assign new_new_n7364__ = new_new_n2737__ & ~new_new_n2848__;
  assign new_new_n7365__ = new_new_n2886__ & new_new_n7364__;
  assign new_new_n7366__ = ~new_new_n3361__ & new_new_n7365__;
  assign new_new_n7367__ = ~new_new_n7363__ & ~new_new_n7366__;
  assign new_new_n7368__ = ~new_new_n2960__ & ~new_new_n7367__;
  assign new_new_n7369__ = new_new_n2849__ & new_new_n3361__;
  assign new_new_n7370__ = ~new_new_n7355__ & ~new_new_n7369__;
  assign new_new_n7371__ = new_new_n3460__ & ~new_new_n7370__;
  assign new_new_n7372__ = ~new_new_n3361__ & new_new_n7362__;
  assign new_new_n7373__ = ~new_new_n7365__ & ~new_new_n7372__;
  assign new_new_n7374__ = ~new_new_n3460__ & ~new_new_n7373__;
  assign new_new_n7375__ = ~new_new_n7358__ & ~new_new_n7361__;
  assign new_new_n7376__ = ~new_new_n7368__ & ~new_new_n7371__;
  assign new_new_n7377__ = ~new_new_n7374__ & new_new_n7376__;
  assign new_new_n7378__ = new_new_n7375__ & new_new_n7377__;
  assign new_new_n7379__ = new_new_n765__ & new_new_n7378__;
  assign new_new_n7380__ = pi31 & ~new_new_n7085__;
  assign new_new_n7381__ = ~new_new_n7353__ & new_new_n7380__;
  assign new_new_n7382__ = ~new_new_n7379__ & new_new_n7381__;
  assign new_new_n7383__ = ~new_new_n7352__ & ~new_new_n7382__;
  assign new_new_n7384__ = new_new_n161__ & ~new_new_n2960__;
  assign new_new_n7385__ = ~new_new_n161__ & new_new_n7072__;
  assign new_new_n7386__ = ~new_new_n7384__ & ~new_new_n7385__;
  assign new_new_n7387__ = ~pi31 & ~new_new_n7386__;
  assign new_new_n7388__ = ~new_new_n7059__ & ~new_new_n7060__;
  assign new_new_n7389__ = new_new_n3460__ & new_new_n7388__;
  assign new_new_n7390__ = ~new_new_n3460__ & ~new_new_n7388__;
  assign new_new_n7391__ = ~new_new_n7389__ & ~new_new_n7390__;
  assign new_new_n7392__ = new_new_n765__ & new_new_n7391__;
  assign new_new_n7393__ = new_new_n161__ & ~new_new_n3126__;
  assign new_new_n7394__ = new_new_n71__ & ~new_new_n2960__;
  assign new_new_n7395__ = ~new_new_n7393__ & ~new_new_n7394__;
  assign new_new_n7396__ = ~new_new_n7392__ & new_new_n7395__;
  assign new_new_n7397__ = pi31 & ~new_new_n7396__;
  assign new_new_n7398__ = ~new_new_n7387__ & ~new_new_n7397__;
  assign new_new_n7399__ = ~new_new_n671__ & ~new_new_n776__;
  assign new_new_n7400__ = ~new_new_n286__ & ~new_new_n896__;
  assign new_new_n7401__ = ~new_new_n329__ & ~new_new_n351__;
  assign new_new_n7402__ = ~new_new_n164__ & ~new_new_n242__;
  assign new_new_n7403__ = ~new_new_n315__ & ~new_new_n634__;
  assign new_new_n7404__ = ~new_new_n845__ & new_new_n7403__;
  assign new_new_n7405__ = new_new_n3581__ & new_new_n7402__;
  assign new_new_n7406__ = new_new_n3582__ & new_new_n5473__;
  assign new_new_n7407__ = new_new_n6320__ & new_new_n7406__;
  assign new_new_n7408__ = new_new_n7404__ & new_new_n7405__;
  assign new_new_n7409__ = ~new_new_n373__ & ~new_new_n607__;
  assign new_new_n7410__ = new_new_n1143__ & new_new_n7401__;
  assign new_new_n7411__ = new_new_n7409__ & new_new_n7410__;
  assign new_new_n7412__ = new_new_n7407__ & new_new_n7408__;
  assign new_new_n7413__ = new_new_n7411__ & new_new_n7412__;
  assign new_new_n7414__ = new_new_n669__ & new_new_n7413__;
  assign new_new_n7415__ = new_new_n5795__ & new_new_n7414__;
  assign new_new_n7416__ = ~new_new_n72__ & ~new_new_n224__;
  assign new_new_n7417__ = new_new_n142__ & ~new_new_n7416__;
  assign new_new_n7418__ = ~new_new_n247__ & ~new_new_n658__;
  assign new_new_n7419__ = ~new_new_n1081__ & new_new_n7418__;
  assign new_new_n7420__ = ~new_new_n192__ & new_new_n1213__;
  assign new_new_n7421__ = new_new_n7419__ & new_new_n7420__;
  assign new_new_n7422__ = ~new_new_n92__ & ~new_new_n441__;
  assign new_new_n7423__ = ~new_new_n1094__ & ~new_new_n3013__;
  assign new_new_n7424__ = new_new_n7422__ & new_new_n7423__;
  assign new_new_n7425__ = new_new_n1711__ & new_new_n1742__;
  assign new_new_n7426__ = new_new_n3968__ & new_new_n7399__;
  assign new_new_n7427__ = ~new_new_n7417__ & new_new_n7426__;
  assign new_new_n7428__ = new_new_n7424__ & new_new_n7425__;
  assign new_new_n7429__ = new_new_n1216__ & new_new_n2034__;
  assign new_new_n7430__ = new_new_n2331__ & new_new_n2619__;
  assign new_new_n7431__ = new_new_n3172__ & new_new_n7400__;
  assign new_new_n7432__ = new_new_n7430__ & new_new_n7431__;
  assign new_new_n7433__ = new_new_n7428__ & new_new_n7429__;
  assign new_new_n7434__ = new_new_n831__ & new_new_n7427__;
  assign new_new_n7435__ = new_new_n7421__ & new_new_n7434__;
  assign new_new_n7436__ = new_new_n7432__ & new_new_n7433__;
  assign new_new_n7437__ = new_new_n7435__ & new_new_n7436__;
  assign new_new_n7438__ = new_new_n6305__ & new_new_n7437__;
  assign new_new_n7439__ = new_new_n3580__ & new_new_n7438__;
  assign new_new_n7440__ = new_new_n7415__ & new_new_n7439__;
  assign new_new_n7441__ = ~new_new_n7398__ & ~new_new_n7440__;
  assign new_new_n7442__ = new_new_n7398__ & new_new_n7440__;
  assign new_new_n7443__ = new_new_n765__ & ~new_new_n2960__;
  assign new_new_n7444__ = ~new_new_n7393__ & ~new_new_n7443__;
  assign new_new_n7445__ = ~pi31 & ~new_new_n7444__;
  assign new_new_n7446__ = ~new_new_n3126__ & new_new_n3164__;
  assign new_new_n7447__ = new_new_n2960__ & new_new_n7446__;
  assign new_new_n7448__ = new_new_n3165__ & new_new_n3356__;
  assign new_new_n7449__ = ~new_new_n7447__ & ~new_new_n7448__;
  assign new_new_n7450__ = new_new_n3254__ & ~new_new_n7449__;
  assign new_new_n7451__ = ~new_new_n2960__ & new_new_n3164__;
  assign new_new_n7452__ = new_new_n2960__ & ~new_new_n3164__;
  assign new_new_n7453__ = ~new_new_n3254__ & new_new_n7452__;
  assign new_new_n7454__ = ~new_new_n7451__ & ~new_new_n7453__;
  assign new_new_n7455__ = new_new_n3126__ & ~new_new_n7454__;
  assign new_new_n7456__ = new_new_n3165__ & new_new_n3254__;
  assign new_new_n7457__ = ~new_new_n7447__ & ~new_new_n7456__;
  assign new_new_n7458__ = new_new_n3055__ & ~new_new_n7457__;
  assign new_new_n7459__ = ~new_new_n3254__ & new_new_n7451__;
  assign new_new_n7460__ = new_new_n3126__ & ~new_new_n3356__;
  assign new_new_n7461__ = new_new_n7452__ & new_new_n7460__;
  assign new_new_n7462__ = ~new_new_n7459__ & ~new_new_n7461__;
  assign new_new_n7463__ = ~new_new_n3055__ & ~new_new_n7462__;
  assign new_new_n7464__ = ~new_new_n3126__ & new_new_n3165__;
  assign new_new_n7465__ = ~new_new_n7450__ & ~new_new_n7464__;
  assign new_new_n7466__ = ~new_new_n7455__ & ~new_new_n7458__;
  assign new_new_n7467__ = ~new_new_n7463__ & new_new_n7466__;
  assign new_new_n7468__ = new_new_n7465__ & new_new_n7467__;
  assign new_new_n7469__ = new_new_n765__ & new_new_n7468__;
  assign new_new_n7470__ = new_new_n71__ & new_new_n3126__;
  assign new_new_n7471__ = new_new_n161__ & new_new_n3164__;
  assign new_new_n7472__ = pi31 & ~new_new_n7470__;
  assign new_new_n7473__ = ~new_new_n7471__ & new_new_n7472__;
  assign new_new_n7474__ = ~new_new_n7469__ & new_new_n7473__;
  assign new_new_n7475__ = ~new_new_n7445__ & ~new_new_n7474__;
  assign new_new_n7476__ = ~new_new_n327__ & ~new_new_n480__;
  assign new_new_n7477__ = ~new_new_n1372__ & new_new_n7476__;
  assign new_new_n7478__ = ~new_new_n150__ & ~new_new_n483__;
  assign new_new_n7479__ = ~new_new_n781__ & ~new_new_n1064__;
  assign new_new_n7480__ = new_new_n7478__ & new_new_n7479__;
  assign new_new_n7481__ = new_new_n2167__ & new_new_n7477__;
  assign new_new_n7482__ = new_new_n2550__ & new_new_n3277__;
  assign new_new_n7483__ = new_new_n7481__ & new_new_n7482__;
  assign new_new_n7484__ = new_new_n2144__ & new_new_n7480__;
  assign new_new_n7485__ = new_new_n3024__ & new_new_n3319__;
  assign new_new_n7486__ = new_new_n4573__ & new_new_n7485__;
  assign new_new_n7487__ = new_new_n7483__ & new_new_n7484__;
  assign new_new_n7488__ = new_new_n3633__ & new_new_n6069__;
  assign new_new_n7489__ = new_new_n7487__ & new_new_n7488__;
  assign new_new_n7490__ = new_new_n7486__ & new_new_n7489__;
  assign new_new_n7491__ = new_new_n1967__ & new_new_n2169__;
  assign new_new_n7492__ = new_new_n2574__ & new_new_n7491__;
  assign new_new_n7493__ = ~new_new_n120__ & ~new_new_n168__;
  assign new_new_n7494__ = ~new_new_n600__ & ~new_new_n1033__;
  assign new_new_n7495__ = new_new_n7493__ & new_new_n7494__;
  assign new_new_n7496__ = ~new_new_n258__ & new_new_n2822__;
  assign new_new_n7497__ = new_new_n7495__ & new_new_n7496__;
  assign new_new_n7498__ = new_new_n1664__ & new_new_n3588__;
  assign new_new_n7499__ = new_new_n4073__ & new_new_n7498__;
  assign new_new_n7500__ = new_new_n7497__ & new_new_n7499__;
  assign new_new_n7501__ = ~new_new_n164__ & ~new_new_n476__;
  assign new_new_n7502__ = ~new_new_n723__ & ~new_new_n1070__;
  assign new_new_n7503__ = new_new_n7501__ & new_new_n7502__;
  assign new_new_n7504__ = ~new_new_n372__ & ~new_new_n595__;
  assign new_new_n7505__ = ~new_new_n884__ & ~new_new_n952__;
  assign new_new_n7506__ = new_new_n7504__ & new_new_n7505__;
  assign new_new_n7507__ = new_new_n735__ & new_new_n7503__;
  assign new_new_n7508__ = new_new_n7506__ & new_new_n7507__;
  assign new_new_n7509__ = new_new_n394__ & new_new_n7508__;
  assign new_new_n7510__ = new_new_n3438__ & new_new_n7492__;
  assign new_new_n7511__ = new_new_n7509__ & new_new_n7510__;
  assign new_new_n7512__ = new_new_n7500__ & new_new_n7511__;
  assign new_new_n7513__ = new_new_n6271__ & new_new_n7512__;
  assign new_new_n7514__ = new_new_n7490__ & new_new_n7513__;
  assign new_new_n7515__ = ~new_new_n7475__ & ~new_new_n7514__;
  assign new_new_n7516__ = new_new_n7475__ & new_new_n7514__;
  assign new_new_n7517__ = ~new_new_n473__ & ~new_new_n585__;
  assign new_new_n7518__ = ~new_new_n248__ & ~new_new_n495__;
  assign new_new_n7519__ = ~new_new_n603__ & ~new_new_n671__;
  assign new_new_n7520__ = ~new_new_n1007__ & new_new_n7519__;
  assign new_new_n7521__ = ~new_new_n606__ & new_new_n7518__;
  assign new_new_n7522__ = new_new_n7520__ & new_new_n7521__;
  assign new_new_n7523__ = ~new_new_n477__ & ~new_new_n1113__;
  assign new_new_n7524__ = ~new_new_n259__ & ~new_new_n375__;
  assign new_new_n7525__ = ~new_new_n1372__ & new_new_n7524__;
  assign new_new_n7526__ = ~new_new_n136__ & ~new_new_n602__;
  assign new_new_n7527__ = new_new_n779__ & ~new_new_n1506__;
  assign new_new_n7528__ = new_new_n1830__ & new_new_n4731__;
  assign new_new_n7529__ = new_new_n6182__ & new_new_n7528__;
  assign new_new_n7530__ = new_new_n7526__ & new_new_n7527__;
  assign new_new_n7531__ = new_new_n1961__ & new_new_n7525__;
  assign new_new_n7532__ = new_new_n7523__ & new_new_n7531__;
  assign new_new_n7533__ = new_new_n7529__ & new_new_n7530__;
  assign new_new_n7534__ = new_new_n7532__ & new_new_n7533__;
  assign new_new_n7535__ = ~new_new_n260__ & ~new_new_n472__;
  assign new_new_n7536__ = ~new_new_n826__ & ~new_new_n896__;
  assign new_new_n7537__ = ~new_new_n1070__ & new_new_n7536__;
  assign new_new_n7538__ = ~new_new_n372__ & new_new_n7535__;
  assign new_new_n7539__ = new_new_n3179__ & new_new_n3805__;
  assign new_new_n7540__ = new_new_n7517__ & new_new_n7539__;
  assign new_new_n7541__ = new_new_n7537__ & new_new_n7538__;
  assign new_new_n7542__ = new_new_n628__ & new_new_n1331__;
  assign new_new_n7543__ = new_new_n1750__ & new_new_n4393__;
  assign new_new_n7544__ = new_new_n7542__ & new_new_n7543__;
  assign new_new_n7545__ = new_new_n7540__ & new_new_n7541__;
  assign new_new_n7546__ = new_new_n347__ & new_new_n2133__;
  assign new_new_n7547__ = new_new_n4576__ & new_new_n4988__;
  assign new_new_n7548__ = new_new_n7522__ & new_new_n7547__;
  assign new_new_n7549__ = new_new_n7545__ & new_new_n7546__;
  assign new_new_n7550__ = new_new_n7544__ & new_new_n7549__;
  assign new_new_n7551__ = new_new_n7534__ & new_new_n7548__;
  assign new_new_n7552__ = new_new_n7550__ & new_new_n7551__;
  assign new_new_n7553__ = new_new_n2788__ & new_new_n7552__;
  assign new_new_n7554__ = new_new_n2819__ & new_new_n7553__;
  assign new_new_n7555__ = new_new_n161__ & ~new_new_n3254__;
  assign new_new_n7556__ = new_new_n71__ & ~new_new_n3164__;
  assign new_new_n7557__ = ~new_new_n3126__ & new_new_n3358__;
  assign new_new_n7558__ = new_new_n3126__ & ~new_new_n3164__;
  assign new_new_n7559__ = ~new_new_n7446__ & ~new_new_n7558__;
  assign new_new_n7560__ = new_new_n3055__ & new_new_n3164__;
  assign new_new_n7561__ = ~new_new_n3254__ & ~new_new_n7560__;
  assign new_new_n7562__ = new_new_n7559__ & new_new_n7561__;
  assign new_new_n7563__ = new_new_n3254__ & ~new_new_n7460__;
  assign new_new_n7564__ = ~new_new_n7559__ & new_new_n7563__;
  assign new_new_n7565__ = ~new_new_n3164__ & ~new_new_n3254__;
  assign new_new_n7566__ = new_new_n3055__ & ~new_new_n7565__;
  assign new_new_n7567__ = ~new_new_n7559__ & new_new_n7566__;
  assign new_new_n7568__ = ~new_new_n7557__ & ~new_new_n7562__;
  assign new_new_n7569__ = ~new_new_n7564__ & ~new_new_n7567__;
  assign new_new_n7570__ = new_new_n7568__ & new_new_n7569__;
  assign new_new_n7571__ = new_new_n765__ & ~new_new_n7570__;
  assign new_new_n7572__ = ~new_new_n7555__ & ~new_new_n7556__;
  assign new_new_n7573__ = ~new_new_n7571__ & new_new_n7572__;
  assign new_new_n7574__ = pi31 & ~new_new_n7573__;
  assign new_new_n7575__ = ~new_new_n71__ & ~new_new_n3126__;
  assign new_new_n7576__ = ~new_new_n161__ & ~new_new_n7575__;
  assign new_new_n7577__ = ~pi31 & ~new_new_n7471__;
  assign new_new_n7578__ = ~new_new_n7576__ & new_new_n7577__;
  assign new_new_n7579__ = ~new_new_n7574__ & ~new_new_n7578__;
  assign new_new_n7580__ = ~new_new_n7554__ & ~new_new_n7579__;
  assign new_new_n7581__ = new_new_n7554__ & new_new_n7579__;
  assign new_new_n7582__ = new_new_n3164__ & new_new_n3356__;
  assign new_new_n7583__ = ~new_new_n3358__ & ~new_new_n7582__;
  assign new_new_n7584__ = ~new_new_n161__ & ~new_new_n7583__;
  assign new_new_n7585__ = ~new_new_n71__ & ~new_new_n7560__;
  assign new_new_n7586__ = ~new_new_n7584__ & new_new_n7585__;
  assign new_new_n7587__ = new_new_n3254__ & ~new_new_n7586__;
  assign new_new_n7588__ = new_new_n161__ & new_new_n3055__;
  assign new_new_n7589__ = new_new_n161__ & ~new_new_n3055__;
  assign new_new_n7590__ = ~new_new_n3254__ & ~new_new_n3357__;
  assign new_new_n7591__ = ~new_new_n7589__ & new_new_n7590__;
  assign new_new_n7592__ = new_new_n7585__ & new_new_n7591__;
  assign new_new_n7593__ = pi31 & ~new_new_n7588__;
  assign new_new_n7594__ = ~new_new_n7592__ & new_new_n7593__;
  assign new_new_n7595__ = ~new_new_n7587__ & new_new_n7594__;
  assign new_new_n7596__ = new_new_n765__ & ~new_new_n3164__;
  assign new_new_n7597__ = ~new_new_n7555__ & ~new_new_n7596__;
  assign new_new_n7598__ = ~pi31 & ~new_new_n7597__;
  assign new_new_n7599__ = ~new_new_n7595__ & ~new_new_n7598__;
  assign new_new_n7600__ = ~new_new_n283__ & ~new_new_n698__;
  assign new_new_n7601__ = ~new_new_n717__ & ~new_new_n940__;
  assign new_new_n7602__ = new_new_n7600__ & new_new_n7601__;
  assign new_new_n7603__ = ~new_new_n218__ & new_new_n7602__;
  assign new_new_n7604__ = new_new_n3076__ & new_new_n7603__;
  assign new_new_n7605__ = ~new_new_n271__ & ~new_new_n425__;
  assign new_new_n7606__ = ~new_new_n846__ & new_new_n7605__;
  assign new_new_n7607__ = ~new_new_n189__ & new_new_n7606__;
  assign new_new_n7608__ = ~new_new_n693__ & ~new_new_n995__;
  assign new_new_n7609__ = new_new_n3058__ & new_new_n7608__;
  assign new_new_n7610__ = new_new_n589__ & new_new_n7609__;
  assign new_new_n7611__ = new_new_n2183__ & new_new_n4232__;
  assign new_new_n7612__ = new_new_n7610__ & new_new_n7611__;
  assign new_new_n7613__ = new_new_n2990__ & new_new_n7612__;
  assign new_new_n7614__ = ~new_new_n101__ & ~new_new_n120__;
  assign new_new_n7615__ = ~new_new_n480__ & ~new_new_n632__;
  assign new_new_n7616__ = ~new_new_n724__ & ~new_new_n838__;
  assign new_new_n7617__ = ~new_new_n851__ & new_new_n7616__;
  assign new_new_n7618__ = new_new_n7614__ & new_new_n7615__;
  assign new_new_n7619__ = new_new_n1371__ & new_new_n1423__;
  assign new_new_n7620__ = new_new_n1741__ & new_new_n2942__;
  assign new_new_n7621__ = new_new_n7399__ & new_new_n7620__;
  assign new_new_n7622__ = new_new_n7618__ & new_new_n7619__;
  assign new_new_n7623__ = new_new_n1097__ & new_new_n7617__;
  assign new_new_n7624__ = new_new_n4074__ & new_new_n7623__;
  assign new_new_n7625__ = new_new_n7621__ & new_new_n7622__;
  assign new_new_n7626__ = new_new_n4303__ & new_new_n7607__;
  assign new_new_n7627__ = new_new_n7625__ & new_new_n7626__;
  assign new_new_n7628__ = new_new_n7624__ & new_new_n7627__;
  assign new_new_n7629__ = new_new_n7613__ & new_new_n7628__;
  assign new_new_n7630__ = ~new_new_n254__ & new_new_n1511__;
  assign new_new_n7631__ = ~new_new_n213__ & ~new_new_n1515__;
  assign new_new_n7632__ = ~new_new_n166__ & new_new_n7631__;
  assign new_new_n7633__ = ~new_new_n945__ & ~new_new_n1217__;
  assign new_new_n7634__ = new_new_n2287__ & new_new_n7633__;
  assign new_new_n7635__ = new_new_n4508__ & new_new_n7632__;
  assign new_new_n7636__ = new_new_n1975__ & new_new_n2324__;
  assign new_new_n7637__ = new_new_n7635__ & new_new_n7636__;
  assign new_new_n7638__ = new_new_n1627__ & new_new_n7634__;
  assign new_new_n7639__ = new_new_n7630__ & new_new_n7638__;
  assign new_new_n7640__ = new_new_n2173__ & new_new_n7637__;
  assign new_new_n7641__ = new_new_n7604__ & new_new_n7640__;
  assign new_new_n7642__ = new_new_n3178__ & new_new_n7639__;
  assign new_new_n7643__ = new_new_n7641__ & new_new_n7642__;
  assign new_new_n7644__ = new_new_n2061__ & new_new_n7643__;
  assign new_new_n7645__ = new_new_n7629__ & new_new_n7644__;
  assign new_new_n7646__ = ~new_new_n7599__ & ~new_new_n7645__;
  assign new_new_n7647__ = new_new_n7599__ & new_new_n7645__;
  assign new_new_n7648__ = ~new_new_n200__ & ~new_new_n604__;
  assign new_new_n7649__ = ~new_new_n693__ & new_new_n7648__;
  assign new_new_n7650__ = new_new_n1097__ & new_new_n7649__;
  assign new_new_n7651__ = ~new_new_n85__ & ~new_new_n594__;
  assign new_new_n7652__ = new_new_n272__ & ~new_new_n7651__;
  assign new_new_n7653__ = ~new_new_n348__ & new_new_n2182__;
  assign new_new_n7654__ = new_new_n2197__ & new_new_n7653__;
  assign new_new_n7655__ = new_new_n3076__ & ~new_new_n7652__;
  assign new_new_n7656__ = new_new_n7654__ & new_new_n7655__;
  assign new_new_n7657__ = ~new_new_n1105__ & new_new_n3274__;
  assign new_new_n7658__ = ~new_new_n837__ & ~new_new_n1515__;
  assign new_new_n7659__ = ~new_new_n120__ & ~new_new_n584__;
  assign new_new_n7660__ = ~new_new_n717__ & ~new_new_n1033__;
  assign new_new_n7661__ = new_new_n7659__ & new_new_n7660__;
  assign new_new_n7662__ = ~new_new_n871__ & ~new_new_n884__;
  assign new_new_n7663__ = new_new_n2500__ & new_new_n7662__;
  assign new_new_n7664__ = ~new_new_n373__ & new_new_n7661__;
  assign new_new_n7665__ = new_new_n962__ & new_new_n1143__;
  assign new_new_n7666__ = new_new_n1341__ & new_new_n7665__;
  assign new_new_n7667__ = new_new_n7663__ & new_new_n7664__;
  assign new_new_n7668__ = new_new_n7650__ & new_new_n7657__;
  assign new_new_n7669__ = new_new_n7658__ & new_new_n7668__;
  assign new_new_n7670__ = new_new_n7666__ & new_new_n7667__;
  assign new_new_n7671__ = new_new_n1569__ & new_new_n2343__;
  assign new_new_n7672__ = new_new_n7656__ & new_new_n7671__;
  assign new_new_n7673__ = new_new_n7669__ & new_new_n7670__;
  assign new_new_n7674__ = new_new_n2722__ & new_new_n7673__;
  assign new_new_n7675__ = new_new_n4594__ & new_new_n7672__;
  assign new_new_n7676__ = new_new_n7674__ & new_new_n7675__;
  assign new_new_n7677__ = new_new_n5812__ & new_new_n7676__;
  assign new_new_n7678__ = ~new_new_n3356__ & new_new_n5059__;
  assign new_new_n7679__ = ~new_new_n161__ & new_new_n3254__;
  assign new_new_n7680__ = new_new_n4876__ & ~new_new_n7679__;
  assign new_new_n7681__ = ~new_new_n3254__ & ~new_new_n3356__;
  assign new_new_n7682__ = new_new_n3254__ & new_new_n3356__;
  assign new_new_n7683__ = ~new_new_n161__ & new_new_n7682__;
  assign new_new_n7684__ = ~new_new_n71__ & ~new_new_n7681__;
  assign new_new_n7685__ = ~new_new_n7683__ & new_new_n7684__;
  assign new_new_n7686__ = pi31 & ~new_new_n7685__;
  assign new_new_n7687__ = ~new_new_n7680__ & ~new_new_n7686__;
  assign new_new_n7688__ = ~new_new_n3055__ & ~new_new_n7687__;
  assign new_new_n7689__ = new_new_n765__ & new_new_n3055__;
  assign new_new_n7690__ = ~new_new_n3254__ & new_new_n7689__;
  assign new_new_n7691__ = ~new_new_n7678__ & ~new_new_n7690__;
  assign new_new_n7692__ = ~new_new_n7688__ & new_new_n7691__;
  assign new_new_n7693__ = ~new_new_n7677__ & ~new_new_n7692__;
  assign new_new_n7694__ = ~new_new_n7647__ & new_new_n7693__;
  assign new_new_n7695__ = ~new_new_n7646__ & ~new_new_n7694__;
  assign new_new_n7696__ = ~new_new_n7581__ & ~new_new_n7695__;
  assign new_new_n7697__ = ~new_new_n7580__ & ~new_new_n7696__;
  assign new_new_n7698__ = ~new_new_n7516__ & ~new_new_n7697__;
  assign new_new_n7699__ = ~new_new_n7515__ & ~new_new_n7698__;
  assign new_new_n7700__ = ~new_new_n7442__ & ~new_new_n7699__;
  assign new_new_n7701__ = ~new_new_n7441__ & ~new_new_n7700__;
  assign new_new_n7702__ = new_new_n161__ & ~new_new_n3460__;
  assign new_new_n7703__ = new_new_n765__ & ~new_new_n2848__;
  assign new_new_n7704__ = ~new_new_n7702__ & ~new_new_n7703__;
  assign new_new_n7705__ = ~pi31 & ~new_new_n7704__;
  assign new_new_n7706__ = new_new_n71__ & new_new_n3460__;
  assign new_new_n7707__ = ~new_new_n3460__ & new_new_n7057__;
  assign new_new_n7708__ = ~new_new_n7055__ & new_new_n7058__;
  assign new_new_n7709__ = ~new_new_n2960__ & ~new_new_n7708__;
  assign new_new_n7710__ = new_new_n3361__ & new_new_n7055__;
  assign new_new_n7711__ = new_new_n2848__ & new_new_n3460__;
  assign new_new_n7712__ = ~new_new_n161__ & new_new_n2960__;
  assign new_new_n7713__ = ~new_new_n7711__ & new_new_n7712__;
  assign new_new_n7714__ = ~new_new_n7710__ & new_new_n7713__;
  assign new_new_n7715__ = ~new_new_n7709__ & ~new_new_n7714__;
  assign new_new_n7716__ = ~new_new_n7707__ & ~new_new_n7715__;
  assign new_new_n7717__ = ~new_new_n71__ & ~new_new_n7384__;
  assign new_new_n7718__ = ~new_new_n7716__ & new_new_n7717__;
  assign new_new_n7719__ = pi31 & ~new_new_n7706__;
  assign new_new_n7720__ = ~new_new_n7718__ & new_new_n7719__;
  assign new_new_n7721__ = ~new_new_n7705__ & ~new_new_n7720__;
  assign new_new_n7722__ = ~new_new_n7701__ & ~new_new_n7721__;
  assign new_new_n7723__ = new_new_n7701__ & new_new_n7721__;
  assign new_new_n7724__ = ~new_new_n585__ & ~new_new_n939__;
  assign new_new_n7725__ = ~new_new_n871__ & ~new_new_n1080__;
  assign new_new_n7726__ = ~new_new_n208__ & new_new_n6234__;
  assign new_new_n7727__ = new_new_n6248__ & new_new_n7726__;
  assign new_new_n7728__ = new_new_n303__ & new_new_n517__;
  assign new_new_n7729__ = ~new_new_n282__ & ~new_new_n656__;
  assign new_new_n7730__ = ~new_new_n332__ & new_new_n7729__;
  assign new_new_n7731__ = ~new_new_n353__ & ~new_new_n874__;
  assign new_new_n7732__ = ~new_new_n1167__ & new_new_n1740__;
  assign new_new_n7733__ = new_new_n2330__ & ~new_new_n7728__;
  assign new_new_n7734__ = new_new_n7732__ & new_new_n7733__;
  assign new_new_n7735__ = new_new_n7730__ & new_new_n7731__;
  assign new_new_n7736__ = new_new_n830__ & ~new_new_n935__;
  assign new_new_n7737__ = new_new_n5303__ & new_new_n6757__;
  assign new_new_n7738__ = new_new_n7736__ & new_new_n7737__;
  assign new_new_n7739__ = new_new_n7734__ & new_new_n7735__;
  assign new_new_n7740__ = new_new_n1704__ & new_new_n7739__;
  assign new_new_n7741__ = new_new_n5382__ & new_new_n7738__;
  assign new_new_n7742__ = new_new_n7740__ & new_new_n7741__;
  assign new_new_n7743__ = new_new_n2298__ & new_new_n7742__;
  assign new_new_n7744__ = ~new_new_n259__ & ~new_new_n496__;
  assign new_new_n7745__ = ~new_new_n671__ & new_new_n7744__;
  assign new_new_n7746__ = ~new_new_n346__ & new_new_n7745__;
  assign new_new_n7747__ = ~new_new_n586__ & ~new_new_n692__;
  assign new_new_n7748__ = ~new_new_n136__ & new_new_n7747__;
  assign new_new_n7749__ = ~new_new_n192__ & ~new_new_n595__;
  assign new_new_n7750__ = ~new_new_n1151__ & new_new_n1424__;
  assign new_new_n7751__ = ~new_new_n1506__ & ~new_new_n1921__;
  assign new_new_n7752__ = new_new_n7750__ & new_new_n7751__;
  assign new_new_n7753__ = new_new_n7748__ & new_new_n7749__;
  assign new_new_n7754__ = new_new_n2202__ & new_new_n2331__;
  assign new_new_n7755__ = new_new_n7724__ & new_new_n7725__;
  assign new_new_n7756__ = new_new_n7754__ & new_new_n7755__;
  assign new_new_n7757__ = new_new_n7752__ & new_new_n7753__;
  assign new_new_n7758__ = new_new_n985__ & new_new_n7727__;
  assign new_new_n7759__ = new_new_n7746__ & new_new_n7758__;
  assign new_new_n7760__ = new_new_n7756__ & new_new_n7757__;
  assign new_new_n7761__ = new_new_n7759__ & new_new_n7760__;
  assign new_new_n7762__ = new_new_n5324__ & new_new_n7761__;
  assign new_new_n7763__ = new_new_n5300__ & new_new_n7762__;
  assign new_new_n7764__ = new_new_n7743__ & new_new_n7763__;
  assign new_new_n7765__ = ~new_new_n7723__ & ~new_new_n7764__;
  assign new_new_n7766__ = ~new_new_n7722__ & ~new_new_n7765__;
  assign new_new_n7767__ = ~new_new_n2636__ & new_new_n4212__;
  assign new_new_n7768__ = ~new_new_n2497__ & new_new_n4815__;
  assign new_new_n7769__ = ~new_new_n2737__ & ~new_new_n4818__;
  assign new_new_n7770__ = ~new_new_n7767__ & ~new_new_n7768__;
  assign new_new_n7771__ = ~new_new_n7769__ & new_new_n7770__;
  assign new_new_n7772__ = ~new_new_n2497__ & new_new_n6797__;
  assign new_new_n7773__ = new_new_n2497__ & ~new_new_n6797__;
  assign new_new_n7774__ = ~new_new_n7772__ & ~new_new_n7773__;
  assign new_new_n7775__ = new_new_n4214__ & ~new_new_n7774__;
  assign new_new_n7776__ = ~pi29 & ~new_new_n7775__;
  assign new_new_n7777__ = new_new_n5732__ & ~new_new_n7774__;
  assign new_new_n7778__ = ~new_new_n7776__ & ~new_new_n7777__;
  assign new_new_n7779__ = new_new_n7771__ & ~new_new_n7778__;
  assign new_new_n7780__ = pi29 & ~new_new_n7771__;
  assign new_new_n7781__ = ~new_new_n7779__ & ~new_new_n7780__;
  assign new_new_n7782__ = new_new_n7766__ & ~new_new_n7781__;
  assign new_new_n7783__ = ~new_new_n7766__ & new_new_n7781__;
  assign new_new_n7784__ = new_new_n7090__ & ~new_new_n7144__;
  assign new_new_n7785__ = ~new_new_n7090__ & new_new_n7144__;
  assign new_new_n7786__ = ~new_new_n7784__ & ~new_new_n7785__;
  assign new_new_n7787__ = pi02 & new_new_n7786__;
  assign new_new_n7788__ = ~pi02 & ~new_new_n7786__;
  assign new_new_n7789__ = ~new_new_n7787__ & ~new_new_n7788__;
  assign new_new_n7790__ = ~new_new_n7783__ & new_new_n7789__;
  assign new_new_n7791__ = ~new_new_n7782__ & ~new_new_n7790__;
  assign new_new_n7792__ = new_new_n7383__ & ~new_new_n7791__;
  assign new_new_n7793__ = ~new_new_n7383__ & new_new_n7791__;
  assign new_new_n7794__ = ~new_new_n7110__ & ~new_new_n7176__;
  assign new_new_n7795__ = ~pi02 & ~new_new_n7785__;
  assign new_new_n7796__ = ~new_new_n7794__ & new_new_n7795__;
  assign new_new_n7797__ = pi02 & ~new_new_n7784__;
  assign new_new_n7798__ = new_new_n7794__ & new_new_n7797__;
  assign new_new_n7799__ = new_new_n7109__ & ~new_new_n7786__;
  assign new_new_n7800__ = ~new_new_n7796__ & ~new_new_n7798__;
  assign new_new_n7801__ = ~new_new_n7799__ & new_new_n7800__;
  assign new_new_n7802__ = ~new_new_n7793__ & ~new_new_n7801__;
  assign new_new_n7803__ = ~new_new_n7792__ & ~new_new_n7802__;
  assign new_new_n7804__ = ~new_new_n7348__ & ~new_new_n7803__;
  assign new_new_n7805__ = new_new_n7348__ & new_new_n7803__;
  assign new_new_n7806__ = new_new_n161__ & ~new_new_n2737__;
  assign new_new_n7807__ = new_new_n765__ & ~new_new_n2636__;
  assign new_new_n7808__ = ~new_new_n7806__ & ~new_new_n7807__;
  assign new_new_n7809__ = ~pi31 & ~new_new_n7808__;
  assign new_new_n7810__ = new_new_n71__ & ~new_new_n2737__;
  assign new_new_n7811__ = ~new_new_n6793__ & ~new_new_n6795__;
  assign new_new_n7812__ = ~new_new_n2636__ & ~new_new_n7811__;
  assign new_new_n7813__ = new_new_n2636__ & new_new_n7811__;
  assign new_new_n7814__ = ~new_new_n7812__ & ~new_new_n7813__;
  assign new_new_n7815__ = new_new_n765__ & ~new_new_n7814__;
  assign new_new_n7816__ = ~new_new_n7350__ & ~new_new_n7810__;
  assign new_new_n7817__ = ~new_new_n7815__ & new_new_n7816__;
  assign new_new_n7818__ = pi31 & ~new_new_n7817__;
  assign new_new_n7819__ = ~new_new_n7809__ & ~new_new_n7818__;
  assign new_new_n7820__ = ~new_new_n7805__ & new_new_n7819__;
  assign new_new_n7821__ = ~new_new_n7804__ & ~new_new_n7820__;
  assign new_new_n7822__ = new_new_n4813__ & ~new_new_n6751__;
  assign new_new_n7823__ = ~new_new_n2572__ & ~new_new_n4818__;
  assign new_new_n7824__ = ~new_new_n2420__ & new_new_n4815__;
  assign new_new_n7825__ = ~new_new_n2313__ & new_new_n4212__;
  assign new_new_n7826__ = ~new_new_n7823__ & ~new_new_n7824__;
  assign new_new_n7827__ = ~new_new_n7825__ & new_new_n7826__;
  assign new_new_n7828__ = ~new_new_n7822__ & new_new_n7827__;
  assign new_new_n7829__ = pi29 & ~new_new_n7828__;
  assign new_new_n7830__ = ~pi29 & new_new_n7828__;
  assign new_new_n7831__ = ~new_new_n7829__ & ~new_new_n7830__;
  assign new_new_n7832__ = ~new_new_n7189__ & ~new_new_n7190__;
  assign new_new_n7833__ = ~new_new_n7194__ & new_new_n7832__;
  assign new_new_n7834__ = new_new_n7194__ & ~new_new_n7832__;
  assign new_new_n7835__ = ~new_new_n7833__ & ~new_new_n7834__;
  assign new_new_n7836__ = ~new_new_n7831__ & new_new_n7835__;
  assign new_new_n7837__ = new_new_n7821__ & ~new_new_n7836__;
  assign new_new_n7838__ = new_new_n7831__ & ~new_new_n7835__;
  assign new_new_n7839__ = ~new_new_n7837__ & ~new_new_n7838__;
  assign new_new_n7840__ = new_new_n7344__ & ~new_new_n7839__;
  assign new_new_n7841__ = new_new_n7340__ & ~new_new_n7840__;
  assign new_new_n7842__ = ~new_new_n7344__ & new_new_n7839__;
  assign new_new_n7843__ = ~new_new_n7841__ & ~new_new_n7842__;
  assign new_new_n7844__ = ~new_new_n1660__ & new_new_n5183__;
  assign new_new_n7845__ = ~new_new_n1902__ & new_new_n5191__;
  assign new_new_n7846__ = ~new_new_n1737__ & new_new_n5213__;
  assign new_new_n7847__ = ~new_new_n7844__ & ~new_new_n7845__;
  assign new_new_n7848__ = ~new_new_n7846__ & new_new_n7847__;
  assign new_new_n7849__ = new_new_n5195__ & new_new_n5688__;
  assign new_new_n7850__ = ~pi23 & ~new_new_n7849__;
  assign new_new_n7851__ = new_new_n5688__ & new_new_n5974__;
  assign new_new_n7852__ = ~new_new_n7850__ & ~new_new_n7851__;
  assign new_new_n7853__ = new_new_n7848__ & ~new_new_n7852__;
  assign new_new_n7854__ = pi23 & ~new_new_n7848__;
  assign new_new_n7855__ = ~new_new_n7853__ & ~new_new_n7854__;
  assign new_new_n7856__ = ~new_new_n7843__ & ~new_new_n7855__;
  assign new_new_n7857__ = new_new_n7843__ & new_new_n7855__;
  assign new_new_n7858__ = ~pi29 & new_new_n7281__;
  assign new_new_n7859__ = pi29 & ~new_new_n7281__;
  assign new_new_n7860__ = ~new_new_n7858__ & ~new_new_n7859__;
  assign new_new_n7861__ = new_new_n7317__ & ~new_new_n7860__;
  assign new_new_n7862__ = ~new_new_n7317__ & new_new_n7860__;
  assign new_new_n7863__ = ~new_new_n7861__ & ~new_new_n7862__;
  assign new_new_n7864__ = new_new_n7290__ & new_new_n7863__;
  assign new_new_n7865__ = ~new_new_n7290__ & ~new_new_n7863__;
  assign new_new_n7866__ = ~new_new_n7864__ & ~new_new_n7865__;
  assign new_new_n7867__ = ~new_new_n7857__ & ~new_new_n7866__;
  assign new_new_n7868__ = ~new_new_n7856__ & ~new_new_n7867__;
  assign new_new_n7869__ = ~new_new_n7328__ & new_new_n7868__;
  assign new_new_n7870__ = new_new_n7328__ & ~new_new_n7868__;
  assign new_new_n7871__ = ~new_new_n1660__ & new_new_n5191__;
  assign new_new_n7872__ = ~new_new_n1466__ & new_new_n5213__;
  assign new_new_n7873__ = ~new_new_n1737__ & new_new_n5183__;
  assign new_new_n7874__ = ~new_new_n7871__ & ~new_new_n7872__;
  assign new_new_n7875__ = ~new_new_n7873__ & new_new_n7874__;
  assign new_new_n7876__ = new_new_n5195__ & ~new_new_n6410__;
  assign new_new_n7877__ = pi23 & ~new_new_n7876__;
  assign new_new_n7878__ = pi22 & new_new_n5195__;
  assign new_new_n7879__ = ~new_new_n6410__ & new_new_n7878__;
  assign new_new_n7880__ = ~new_new_n7877__ & ~new_new_n7879__;
  assign new_new_n7881__ = new_new_n7875__ & ~new_new_n7880__;
  assign new_new_n7882__ = ~pi23 & ~new_new_n7875__;
  assign new_new_n7883__ = ~new_new_n7881__ & ~new_new_n7882__;
  assign new_new_n7884__ = ~new_new_n7870__ & ~new_new_n7883__;
  assign new_new_n7885__ = ~new_new_n7869__ & ~new_new_n7884__;
  assign new_new_n7886__ = new_new_n7020__ & new_new_n7885__;
  assign new_new_n7887__ = ~new_new_n7020__ & ~new_new_n7885__;
  assign new_new_n7888__ = ~new_new_n7886__ & ~new_new_n7887__;
  assign new_new_n7889__ = new_new_n7030__ & ~new_new_n7324__;
  assign new_new_n7890__ = ~new_new_n7323__ & ~new_new_n7889__;
  assign new_new_n7891__ = new_new_n5215__ & ~new_new_n5671__;
  assign new_new_n7892__ = ~new_new_n1737__ & new_new_n5191__;
  assign new_new_n7893__ = ~new_new_n1466__ & new_new_n5183__;
  assign new_new_n7894__ = ~new_new_n7892__ & ~new_new_n7893__;
  assign new_new_n7895__ = ~new_new_n7891__ & new_new_n7894__;
  assign new_new_n7896__ = ~new_new_n1556__ & new_new_n5195__;
  assign new_new_n7897__ = pi23 & ~new_new_n7896__;
  assign new_new_n7898__ = ~new_new_n1556__ & new_new_n5974__;
  assign new_new_n7899__ = ~new_new_n7897__ & ~new_new_n7898__;
  assign new_new_n7900__ = new_new_n7895__ & ~new_new_n7899__;
  assign new_new_n7901__ = ~pi23 & ~new_new_n7895__;
  assign new_new_n7902__ = ~new_new_n7900__ & ~new_new_n7901__;
  assign new_new_n7903__ = new_new_n7890__ & new_new_n7902__;
  assign new_new_n7904__ = ~new_new_n7890__ & ~new_new_n7902__;
  assign new_new_n7905__ = ~new_new_n7903__ & ~new_new_n7904__;
  assign new_new_n7906__ = new_new_n6878__ & ~new_new_n6881__;
  assign new_new_n7907__ = ~new_new_n6882__ & ~new_new_n7906__;
  assign new_new_n7908__ = new_new_n873__ & ~new_new_n1902__;
  assign new_new_n7909__ = ~new_new_n1660__ & new_new_n3311__;
  assign new_new_n7910__ = ~new_new_n333__ & ~new_new_n1823__;
  assign new_new_n7911__ = ~new_new_n7908__ & ~new_new_n7909__;
  assign new_new_n7912__ = ~new_new_n7910__ & new_new_n7911__;
  assign new_new_n7913__ = pi26 & ~new_new_n7912__;
  assign new_new_n7914__ = new_new_n4898__ & ~new_new_n5274__;
  assign new_new_n7915__ = new_new_n801__ & ~new_new_n5274__;
  assign new_new_n7916__ = ~pi26 & ~new_new_n7915__;
  assign new_new_n7917__ = ~new_new_n7914__ & ~new_new_n7916__;
  assign new_new_n7918__ = new_new_n7912__ & ~new_new_n7917__;
  assign new_new_n7919__ = ~new_new_n7913__ & ~new_new_n7918__;
  assign new_new_n7920__ = ~new_new_n7256__ & ~new_new_n7264__;
  assign new_new_n7921__ = ~new_new_n7255__ & ~new_new_n7920__;
  assign new_new_n7922__ = ~new_new_n7919__ & ~new_new_n7921__;
  assign new_new_n7923__ = new_new_n7919__ & new_new_n7921__;
  assign new_new_n7924__ = ~new_new_n7922__ & ~new_new_n7923__;
  assign new_new_n7925__ = new_new_n7907__ & new_new_n7924__;
  assign new_new_n7926__ = ~new_new_n7907__ & ~new_new_n7924__;
  assign new_new_n7927__ = ~new_new_n7925__ & ~new_new_n7926__;
  assign new_new_n7928__ = ~new_new_n7905__ & new_new_n7927__;
  assign new_new_n7929__ = new_new_n7905__ & ~new_new_n7927__;
  assign new_new_n7930__ = ~new_new_n7928__ & ~new_new_n7929__;
  assign new_new_n7931__ = new_new_n7888__ & ~new_new_n7930__;
  assign new_new_n7932__ = ~new_new_n7888__ & new_new_n7930__;
  assign new_new_n7933__ = ~new_new_n7931__ & ~new_new_n7932__;
  assign new_new_n7934__ = ~new_new_n1207__ & new_new_n6964__;
  assign new_new_n7935__ = ~new_new_n6955__ & new_new_n6958__;
  assign new_new_n7936__ = ~new_new_n3720__ & new_new_n7935__;
  assign new_new_n7937__ = ~new_new_n868__ & new_new_n6968__;
  assign new_new_n7938__ = ~new_new_n7934__ & ~new_new_n7936__;
  assign new_new_n7939__ = ~new_new_n7937__ & new_new_n7938__;
  assign new_new_n7940__ = ~new_new_n5927__ & new_new_n6958__;
  assign new_new_n7941__ = pi17 & ~new_new_n7940__;
  assign new_new_n7942__ = pi16 & new_new_n6958__;
  assign new_new_n7943__ = ~new_new_n5927__ & new_new_n7942__;
  assign new_new_n7944__ = ~new_new_n7941__ & ~new_new_n7943__;
  assign new_new_n7945__ = new_new_n7939__ & ~new_new_n7944__;
  assign new_new_n7946__ = ~pi17 & ~new_new_n7939__;
  assign new_new_n7947__ = ~new_new_n7945__ & ~new_new_n7946__;
  assign new_new_n7948__ = ~new_new_n7933__ & ~new_new_n7947__;
  assign new_new_n7949__ = new_new_n7933__ & new_new_n7947__;
  assign new_new_n7950__ = ~new_new_n3618__ & new_new_n6634__;
  assign new_new_n7951__ = ~new_new_n1325__ & new_new_n6629__;
  assign new_new_n7952__ = ~new_new_n1556__ & ~new_new_n6625__;
  assign new_new_n7953__ = ~new_new_n7950__ & ~new_new_n7951__;
  assign new_new_n7954__ = ~new_new_n7952__ & new_new_n7953__;
  assign new_new_n7955__ = ~new_new_n5061__ & new_new_n6631__;
  assign new_new_n7956__ = ~new_new_n5746__ & new_new_n7955__;
  assign new_new_n7957__ = pi20 & ~new_new_n7956__;
  assign new_new_n7958__ = pi19 & new_new_n7956__;
  assign new_new_n7959__ = ~new_new_n7957__ & ~new_new_n7958__;
  assign new_new_n7960__ = new_new_n7954__ & ~new_new_n7959__;
  assign new_new_n7961__ = ~pi20 & ~new_new_n7954__;
  assign new_new_n7962__ = ~new_new_n7960__ & ~new_new_n7961__;
  assign new_new_n7963__ = new_new_n5215__ & ~new_new_n5274__;
  assign new_new_n7964__ = ~new_new_n1902__ & new_new_n5183__;
  assign new_new_n7965__ = ~new_new_n1660__ & new_new_n5213__;
  assign new_new_n7966__ = ~new_new_n1823__ & new_new_n5191__;
  assign new_new_n7967__ = ~new_new_n7964__ & ~new_new_n7965__;
  assign new_new_n7968__ = ~new_new_n7966__ & new_new_n7967__;
  assign new_new_n7969__ = ~new_new_n7963__ & new_new_n7968__;
  assign new_new_n7970__ = pi23 & ~new_new_n7969__;
  assign new_new_n7971__ = ~pi23 & new_new_n7969__;
  assign new_new_n7972__ = ~new_new_n7970__ & ~new_new_n7971__;
  assign new_new_n7973__ = ~new_new_n2572__ & new_new_n4212__;
  assign new_new_n7974__ = ~new_new_n2497__ & ~new_new_n4818__;
  assign new_new_n7975__ = ~new_new_n2313__ & new_new_n4815__;
  assign new_new_n7976__ = new_new_n4813__ & ~new_new_n7236__;
  assign new_new_n7977__ = ~new_new_n7973__ & ~new_new_n7974__;
  assign new_new_n7978__ = ~new_new_n7975__ & new_new_n7977__;
  assign new_new_n7979__ = ~new_new_n7976__ & new_new_n7978__;
  assign new_new_n7980__ = pi29 & ~new_new_n7979__;
  assign new_new_n7981__ = ~pi29 & new_new_n7979__;
  assign new_new_n7982__ = ~new_new_n7980__ & ~new_new_n7981__;
  assign new_new_n7983__ = ~new_new_n7804__ & ~new_new_n7805__;
  assign new_new_n7984__ = new_new_n7819__ & new_new_n7983__;
  assign new_new_n7985__ = ~new_new_n7819__ & ~new_new_n7983__;
  assign new_new_n7986__ = ~new_new_n7984__ & ~new_new_n7985__;
  assign new_new_n7987__ = ~new_new_n7982__ & new_new_n7986__;
  assign new_new_n7988__ = new_new_n7982__ & ~new_new_n7986__;
  assign new_new_n7989__ = new_new_n873__ & ~new_new_n2224__;
  assign new_new_n7990__ = ~new_new_n333__ & ~new_new_n2420__;
  assign new_new_n7991__ = ~new_new_n2024__ & new_new_n3311__;
  assign new_new_n7992__ = ~new_new_n4900__ & new_new_n7313__;
  assign new_new_n7993__ = ~new_new_n7989__ & ~new_new_n7990__;
  assign new_new_n7994__ = ~new_new_n7991__ & new_new_n7993__;
  assign new_new_n7995__ = ~new_new_n7992__ & new_new_n7994__;
  assign new_new_n7996__ = pi26 & ~new_new_n7995__;
  assign new_new_n7997__ = ~pi26 & new_new_n7995__;
  assign new_new_n7998__ = ~new_new_n7996__ & ~new_new_n7997__;
  assign new_new_n7999__ = ~new_new_n7988__ & ~new_new_n7998__;
  assign new_new_n8000__ = ~new_new_n7987__ & ~new_new_n7999__;
  assign new_new_n8001__ = ~new_new_n7836__ & ~new_new_n7838__;
  assign new_new_n8002__ = new_new_n7821__ & new_new_n8001__;
  assign new_new_n8003__ = ~new_new_n7821__ & ~new_new_n8001__;
  assign new_new_n8004__ = ~new_new_n8002__ & ~new_new_n8003__;
  assign new_new_n8005__ = ~new_new_n8000__ & ~new_new_n8004__;
  assign new_new_n8006__ = new_new_n8000__ & new_new_n8004__;
  assign new_new_n8007__ = ~new_new_n2130__ & new_new_n3311__;
  assign new_new_n8008__ = ~new_new_n333__ & ~new_new_n2224__;
  assign new_new_n8009__ = new_new_n873__ & ~new_new_n2024__;
  assign new_new_n8010__ = ~new_new_n4900__ & ~new_new_n6036__;
  assign new_new_n8011__ = ~new_new_n8007__ & ~new_new_n8008__;
  assign new_new_n8012__ = ~new_new_n8009__ & new_new_n8011__;
  assign new_new_n8013__ = ~new_new_n8010__ & new_new_n8012__;
  assign new_new_n8014__ = ~pi26 & ~new_new_n8013__;
  assign new_new_n8015__ = pi26 & new_new_n8013__;
  assign new_new_n8016__ = ~new_new_n8014__ & ~new_new_n8015__;
  assign new_new_n8017__ = ~new_new_n8006__ & new_new_n8016__;
  assign new_new_n8018__ = ~new_new_n8005__ & ~new_new_n8017__;
  assign new_new_n8019__ = new_new_n7972__ & new_new_n8018__;
  assign new_new_n8020__ = ~new_new_n7972__ & ~new_new_n8018__;
  assign new_new_n8021__ = ~new_new_n7840__ & ~new_new_n7842__;
  assign new_new_n8022__ = new_new_n7340__ & new_new_n8021__;
  assign new_new_n8023__ = ~new_new_n7340__ & ~new_new_n8021__;
  assign new_new_n8024__ = ~new_new_n8022__ & ~new_new_n8023__;
  assign new_new_n8025__ = ~new_new_n8020__ & ~new_new_n8024__;
  assign new_new_n8026__ = ~new_new_n8019__ & ~new_new_n8025__;
  assign new_new_n8027__ = ~new_new_n7317__ & new_new_n7843__;
  assign new_new_n8028__ = new_new_n7317__ & ~new_new_n7843__;
  assign new_new_n8029__ = ~new_new_n8027__ & ~new_new_n8028__;
  assign new_new_n8030__ = new_new_n7290__ & new_new_n8029__;
  assign new_new_n8031__ = ~new_new_n7290__ & ~new_new_n8029__;
  assign new_new_n8032__ = ~new_new_n8030__ & ~new_new_n8031__;
  assign new_new_n8033__ = new_new_n7860__ & ~new_new_n8032__;
  assign new_new_n8034__ = ~new_new_n7860__ & new_new_n8032__;
  assign new_new_n8035__ = ~new_new_n8033__ & ~new_new_n8034__;
  assign new_new_n8036__ = new_new_n7855__ & new_new_n8035__;
  assign new_new_n8037__ = ~new_new_n7855__ & ~new_new_n8035__;
  assign new_new_n8038__ = ~new_new_n8036__ & ~new_new_n8037__;
  assign new_new_n8039__ = ~new_new_n8026__ & ~new_new_n8038__;
  assign new_new_n8040__ = ~new_new_n1466__ & ~new_new_n6625__;
  assign new_new_n8041__ = ~new_new_n1556__ & new_new_n6629__;
  assign new_new_n8042__ = ~new_new_n1325__ & new_new_n6634__;
  assign new_new_n8043__ = new_new_n5048__ & new_new_n6936__;
  assign new_new_n8044__ = ~new_new_n8040__ & ~new_new_n8041__;
  assign new_new_n8045__ = ~new_new_n8042__ & new_new_n8044__;
  assign new_new_n8046__ = ~new_new_n8043__ & new_new_n8045__;
  assign new_new_n8047__ = ~pi20 & ~new_new_n8046__;
  assign new_new_n8048__ = pi20 & new_new_n8046__;
  assign new_new_n8049__ = ~new_new_n8047__ & ~new_new_n8048__;
  assign new_new_n8050__ = new_new_n8026__ & new_new_n8038__;
  assign new_new_n8051__ = ~new_new_n8049__ & ~new_new_n8050__;
  assign new_new_n8052__ = ~new_new_n8039__ & ~new_new_n8051__;
  assign new_new_n8053__ = ~new_new_n7962__ & ~new_new_n8052__;
  assign new_new_n8054__ = new_new_n7962__ & new_new_n8052__;
  assign new_new_n8055__ = ~new_new_n7869__ & ~new_new_n7870__;
  assign new_new_n8056__ = ~new_new_n7883__ & new_new_n8055__;
  assign new_new_n8057__ = new_new_n7883__ & ~new_new_n8055__;
  assign new_new_n8058__ = ~new_new_n8056__ & ~new_new_n8057__;
  assign new_new_n8059__ = ~new_new_n8054__ & new_new_n8058__;
  assign new_new_n8060__ = ~new_new_n8053__ & ~new_new_n8059__;
  assign new_new_n8061__ = ~new_new_n7949__ & ~new_new_n8060__;
  assign new_new_n8062__ = ~new_new_n7948__ & ~new_new_n8061__;
  assign new_new_n8063__ = ~new_new_n7007__ & ~new_new_n8062__;
  assign new_new_n8064__ = new_new_n7007__ & new_new_n8062__;
  assign new_new_n8065__ = ~new_new_n8063__ & ~new_new_n8064__;
  assign new_new_n8066__ = ~new_new_n3720__ & new_new_n6968__;
  assign new_new_n8067__ = ~new_new_n868__ & new_new_n6964__;
  assign new_new_n8068__ = ~new_new_n8066__ & ~new_new_n8067__;
  assign new_new_n8069__ = new_new_n5116__ & new_new_n6958__;
  assign new_new_n8070__ = new_new_n8068__ & ~new_new_n8069__;
  assign new_new_n8071__ = pi17 & ~new_new_n8070__;
  assign new_new_n8072__ = ~new_new_n5129__ & new_new_n6958__;
  assign new_new_n8073__ = ~pi17 & ~new_new_n8072__;
  assign new_new_n8074__ = pi16 & new_new_n910__;
  assign new_new_n8075__ = ~pi16 & ~new_new_n910__;
  assign new_new_n8076__ = new_new_n6958__ & ~new_new_n8074__;
  assign new_new_n8077__ = ~new_new_n8075__ & new_new_n8076__;
  assign new_new_n8078__ = new_new_n4036__ & new_new_n8077__;
  assign new_new_n8079__ = ~new_new_n8073__ & ~new_new_n8078__;
  assign new_new_n8080__ = new_new_n8068__ & ~new_new_n8079__;
  assign new_new_n8081__ = ~new_new_n8071__ & ~new_new_n8080__;
  assign new_new_n8082__ = ~new_new_n7886__ & ~new_new_n7931__;
  assign new_new_n8083__ = ~new_new_n1207__ & new_new_n6634__;
  assign new_new_n8084__ = ~new_new_n1061__ & new_new_n6629__;
  assign new_new_n8085__ = ~new_new_n3618__ & ~new_new_n6625__;
  assign new_new_n8086__ = ~new_new_n5235__ & new_new_n6936__;
  assign new_new_n8087__ = ~new_new_n8083__ & ~new_new_n8084__;
  assign new_new_n8088__ = ~new_new_n8085__ & new_new_n8087__;
  assign new_new_n8089__ = ~new_new_n8086__ & new_new_n8088__;
  assign new_new_n8090__ = ~pi20 & ~new_new_n8089__;
  assign new_new_n8091__ = pi20 & new_new_n8089__;
  assign new_new_n8092__ = ~new_new_n8090__ & ~new_new_n8091__;
  assign new_new_n8093__ = ~new_new_n1466__ & new_new_n5191__;
  assign new_new_n8094__ = ~new_new_n1556__ & new_new_n5183__;
  assign new_new_n8095__ = ~new_new_n1325__ & new_new_n5213__;
  assign new_new_n8096__ = new_new_n5048__ & new_new_n5215__;
  assign new_new_n8097__ = ~new_new_n8093__ & ~new_new_n8094__;
  assign new_new_n8098__ = ~new_new_n8095__ & new_new_n8097__;
  assign new_new_n8099__ = ~new_new_n8096__ & new_new_n8098__;
  assign new_new_n8100__ = ~pi23 & ~new_new_n8099__;
  assign new_new_n8101__ = pi23 & new_new_n8099__;
  assign new_new_n8102__ = ~new_new_n8100__ & ~new_new_n8101__;
  assign new_new_n8103__ = ~new_new_n6895__ & ~new_new_n6896__;
  assign new_new_n8104__ = ~new_new_n6900__ & new_new_n8103__;
  assign new_new_n8105__ = new_new_n6900__ & ~new_new_n8103__;
  assign new_new_n8106__ = ~new_new_n8104__ & ~new_new_n8105__;
  assign new_new_n8107__ = ~new_new_n8102__ & ~new_new_n8106__;
  assign new_new_n8108__ = new_new_n8102__ & new_new_n8106__;
  assign new_new_n8109__ = ~new_new_n8107__ & ~new_new_n8108__;
  assign new_new_n8110__ = new_new_n7907__ & ~new_new_n7923__;
  assign new_new_n8111__ = ~new_new_n7922__ & ~new_new_n8110__;
  assign new_new_n8112__ = new_new_n8109__ & new_new_n8111__;
  assign new_new_n8113__ = ~new_new_n8109__ & ~new_new_n8111__;
  assign new_new_n8114__ = ~new_new_n8112__ & ~new_new_n8113__;
  assign new_new_n8115__ = ~new_new_n7904__ & new_new_n7927__;
  assign new_new_n8116__ = ~new_new_n7903__ & ~new_new_n8115__;
  assign new_new_n8117__ = new_new_n8114__ & new_new_n8116__;
  assign new_new_n8118__ = ~new_new_n8114__ & ~new_new_n8116__;
  assign new_new_n8119__ = ~new_new_n8117__ & ~new_new_n8118__;
  assign new_new_n8120__ = ~new_new_n8092__ & new_new_n8119__;
  assign new_new_n8121__ = new_new_n8092__ & ~new_new_n8119__;
  assign new_new_n8122__ = ~new_new_n8120__ & ~new_new_n8121__;
  assign new_new_n8123__ = ~new_new_n8082__ & ~new_new_n8122__;
  assign new_new_n8124__ = new_new_n8082__ & new_new_n8122__;
  assign new_new_n8125__ = ~new_new_n8123__ & ~new_new_n8124__;
  assign new_new_n8126__ = new_new_n8081__ & new_new_n8125__;
  assign new_new_n8127__ = ~new_new_n8081__ & ~new_new_n8125__;
  assign new_new_n8128__ = ~new_new_n8126__ & ~new_new_n8127__;
  assign new_new_n8129__ = new_new_n8065__ & ~new_new_n8128__;
  assign new_new_n8130__ = ~new_new_n8065__ & new_new_n8128__;
  assign new_new_n8131__ = ~new_new_n8129__ & ~new_new_n8130__;
  assign new_new_n8132__ = ~new_new_n910__ & new_new_n6991__;
  assign new_new_n8133__ = ~new_new_n691__ & new_new_n6985__;
  assign new_new_n8134__ = ~new_new_n8132__ & ~new_new_n8133__;
  assign new_new_n8135__ = ~new_new_n583__ & new_new_n6994__;
  assign new_new_n8136__ = new_new_n3742__ & new_new_n8135__;
  assign new_new_n8137__ = new_new_n8134__ & ~new_new_n8136__;
  assign new_new_n8138__ = ~pi14 & ~new_new_n8137__;
  assign new_new_n8139__ = ~pi13 & new_new_n3742__;
  assign new_new_n8140__ = new_new_n583__ & ~new_new_n3742__;
  assign new_new_n8141__ = new_new_n6994__ & ~new_new_n8140__;
  assign new_new_n8142__ = pi13 & ~new_new_n583__;
  assign new_new_n8143__ = ~new_new_n8139__ & ~new_new_n8142__;
  assign new_new_n8144__ = new_new_n8141__ & new_new_n8143__;
  assign new_new_n8145__ = pi14 & new_new_n8134__;
  assign new_new_n8146__ = ~new_new_n8141__ & new_new_n8145__;
  assign new_new_n8147__ = ~new_new_n8138__ & ~new_new_n8144__;
  assign new_new_n8148__ = ~new_new_n8146__ & new_new_n8147__;
  assign new_new_n8149__ = ~new_new_n8039__ & ~new_new_n8050__;
  assign new_new_n8150__ = new_new_n8049__ & ~new_new_n8149__;
  assign new_new_n8151__ = ~new_new_n8049__ & new_new_n8149__;
  assign new_new_n8152__ = ~new_new_n8150__ & ~new_new_n8151__;
  assign new_new_n8153__ = ~new_new_n1207__ & new_new_n7935__;
  assign new_new_n8154__ = ~new_new_n3618__ & new_new_n6964__;
  assign new_new_n8155__ = ~new_new_n1061__ & new_new_n6968__;
  assign new_new_n8156__ = ~new_new_n8153__ & ~new_new_n8154__;
  assign new_new_n8157__ = ~new_new_n8155__ & new_new_n8156__;
  assign new_new_n8158__ = ~new_new_n5235__ & new_new_n6958__;
  assign new_new_n8159__ = ~pi17 & ~new_new_n8158__;
  assign new_new_n8160__ = ~pi16 & new_new_n6958__;
  assign new_new_n8161__ = ~new_new_n5235__ & new_new_n8160__;
  assign new_new_n8162__ = ~new_new_n8159__ & ~new_new_n8161__;
  assign new_new_n8163__ = new_new_n8157__ & ~new_new_n8162__;
  assign new_new_n8164__ = pi17 & ~new_new_n8157__;
  assign new_new_n8165__ = ~new_new_n8163__ & ~new_new_n8164__;
  assign new_new_n8166__ = ~new_new_n8152__ & ~new_new_n8165__;
  assign new_new_n8167__ = new_new_n8152__ & new_new_n8165__;
  assign new_new_n8168__ = ~new_new_n3535__ & new_new_n5183__;
  assign new_new_n8169__ = ~new_new_n2130__ & new_new_n5191__;
  assign new_new_n8170__ = ~new_new_n8168__ & ~new_new_n8169__;
  assign new_new_n8171__ = new_new_n5195__ & ~new_new_n5520__;
  assign new_new_n8172__ = pi23 & ~new_new_n8171__;
  assign new_new_n8173__ = ~pi22 & new_new_n1823__;
  assign new_new_n8174__ = pi22 & ~new_new_n1823__;
  assign new_new_n8175__ = new_new_n5195__ & ~new_new_n8173__;
  assign new_new_n8176__ = ~new_new_n8174__ & new_new_n8175__;
  assign new_new_n8177__ = new_new_n5501__ & new_new_n8176__;
  assign new_new_n8178__ = ~new_new_n8172__ & ~new_new_n8177__;
  assign new_new_n8179__ = new_new_n8170__ & ~new_new_n8178__;
  assign new_new_n8180__ = new_new_n5195__ & new_new_n6553__;
  assign new_new_n8181__ = new_new_n8170__ & ~new_new_n8180__;
  assign new_new_n8182__ = ~pi23 & ~new_new_n8181__;
  assign new_new_n8183__ = ~new_new_n8179__ & ~new_new_n8182__;
  assign new_new_n8184__ = ~new_new_n7987__ & ~new_new_n7988__;
  assign new_new_n8185__ = new_new_n7998__ & new_new_n8184__;
  assign new_new_n8186__ = ~new_new_n7998__ & ~new_new_n8184__;
  assign new_new_n8187__ = ~new_new_n8185__ & ~new_new_n8186__;
  assign new_new_n8188__ = new_new_n8183__ & ~new_new_n8187__;
  assign new_new_n8189__ = ~new_new_n8183__ & new_new_n8187__;
  assign new_new_n8190__ = ~new_new_n333__ & ~new_new_n2313__;
  assign new_new_n8191__ = ~new_new_n2224__ & new_new_n3311__;
  assign new_new_n8192__ = new_new_n873__ & ~new_new_n2420__;
  assign new_new_n8193__ = ~new_new_n4900__ & new_new_n6521__;
  assign new_new_n8194__ = ~new_new_n8190__ & ~new_new_n8191__;
  assign new_new_n8195__ = ~new_new_n8192__ & new_new_n8194__;
  assign new_new_n8196__ = ~new_new_n8193__ & new_new_n8195__;
  assign new_new_n8197__ = pi26 & ~new_new_n8196__;
  assign new_new_n8198__ = ~pi26 & new_new_n8196__;
  assign new_new_n8199__ = ~new_new_n8197__ & ~new_new_n8198__;
  assign new_new_n8200__ = ~new_new_n7792__ & ~new_new_n7793__;
  assign new_new_n8201__ = ~new_new_n7794__ & new_new_n7797__;
  assign new_new_n8202__ = new_new_n7794__ & new_new_n7795__;
  assign new_new_n8203__ = ~new_new_n7109__ & ~new_new_n7786__;
  assign new_new_n8204__ = ~new_new_n8201__ & ~new_new_n8202__;
  assign new_new_n8205__ = ~new_new_n8203__ & new_new_n8204__;
  assign new_new_n8206__ = new_new_n8200__ & ~new_new_n8205__;
  assign new_new_n8207__ = ~new_new_n7801__ & ~new_new_n8200__;
  assign new_new_n8208__ = ~new_new_n8206__ & ~new_new_n8207__;
  assign new_new_n8209__ = ~new_new_n8199__ & ~new_new_n8208__;
  assign new_new_n8210__ = new_new_n8199__ & new_new_n8208__;
  assign new_new_n8211__ = ~new_new_n2636__ & ~new_new_n4818__;
  assign new_new_n8212__ = ~new_new_n2497__ & new_new_n4212__;
  assign new_new_n8213__ = ~new_new_n2572__ & new_new_n4815__;
  assign new_new_n8214__ = ~new_new_n8211__ & ~new_new_n8212__;
  assign new_new_n8215__ = ~new_new_n8213__ & new_new_n8214__;
  assign new_new_n8216__ = new_new_n4214__ & new_new_n6804__;
  assign new_new_n8217__ = ~pi29 & ~new_new_n8216__;
  assign new_new_n8218__ = new_new_n5732__ & new_new_n6804__;
  assign new_new_n8219__ = ~new_new_n8217__ & ~new_new_n8218__;
  assign new_new_n8220__ = new_new_n8215__ & ~new_new_n8219__;
  assign new_new_n8221__ = pi29 & ~new_new_n8215__;
  assign new_new_n8222__ = ~new_new_n8220__ & ~new_new_n8221__;
  assign new_new_n8223__ = ~new_new_n8210__ & ~new_new_n8222__;
  assign new_new_n8224__ = ~new_new_n8209__ & ~new_new_n8223__;
  assign new_new_n8225__ = ~new_new_n8189__ & ~new_new_n8224__;
  assign new_new_n8226__ = ~new_new_n8188__ & ~new_new_n8225__;
  assign new_new_n8227__ = ~new_new_n8005__ & ~new_new_n8006__;
  assign new_new_n8228__ = ~new_new_n8016__ & new_new_n8227__;
  assign new_new_n8229__ = new_new_n8016__ & ~new_new_n8227__;
  assign new_new_n8230__ = ~new_new_n8228__ & ~new_new_n8229__;
  assign new_new_n8231__ = ~new_new_n8226__ & ~new_new_n8230__;
  assign new_new_n8232__ = new_new_n8226__ & new_new_n8230__;
  assign new_new_n8233__ = ~new_new_n1823__ & new_new_n5183__;
  assign new_new_n8234__ = ~new_new_n3535__ & new_new_n5191__;
  assign new_new_n8235__ = ~new_new_n1902__ & new_new_n5213__;
  assign new_new_n8236__ = new_new_n5215__ & ~new_new_n6487__;
  assign new_new_n8237__ = ~new_new_n8233__ & ~new_new_n8234__;
  assign new_new_n8238__ = ~new_new_n8235__ & new_new_n8237__;
  assign new_new_n8239__ = ~new_new_n8236__ & new_new_n8238__;
  assign new_new_n8240__ = pi23 & ~new_new_n8239__;
  assign new_new_n8241__ = ~pi23 & new_new_n8239__;
  assign new_new_n8242__ = ~new_new_n8240__ & ~new_new_n8241__;
  assign new_new_n8243__ = ~new_new_n8232__ & ~new_new_n8242__;
  assign new_new_n8244__ = ~new_new_n8231__ & ~new_new_n8243__;
  assign new_new_n8245__ = ~new_new_n8019__ & ~new_new_n8020__;
  assign new_new_n8246__ = new_new_n8024__ & new_new_n8245__;
  assign new_new_n8247__ = ~new_new_n8024__ & ~new_new_n8245__;
  assign new_new_n8248__ = ~new_new_n8246__ & ~new_new_n8247__;
  assign new_new_n8249__ = ~new_new_n8244__ & new_new_n8248__;
  assign new_new_n8250__ = new_new_n8244__ & ~new_new_n8248__;
  assign new_new_n8251__ = ~new_new_n1556__ & new_new_n6634__;
  assign new_new_n8252__ = ~new_new_n1466__ & new_new_n6629__;
  assign new_new_n8253__ = ~new_new_n1737__ & ~new_new_n6625__;
  assign new_new_n8254__ = ~new_new_n8251__ & ~new_new_n8252__;
  assign new_new_n8255__ = ~new_new_n8253__ & new_new_n8254__;
  assign new_new_n8256__ = ~new_new_n5671__ & new_new_n6631__;
  assign new_new_n8257__ = ~pi20 & ~new_new_n8256__;
  assign new_new_n8258__ = ~new_new_n5671__ & new_new_n7015__;
  assign new_new_n8259__ = ~new_new_n8257__ & ~new_new_n8258__;
  assign new_new_n8260__ = new_new_n8255__ & ~new_new_n8259__;
  assign new_new_n8261__ = pi20 & ~new_new_n8255__;
  assign new_new_n8262__ = ~new_new_n8260__ & ~new_new_n8261__;
  assign new_new_n8263__ = ~new_new_n8250__ & ~new_new_n8262__;
  assign new_new_n8264__ = ~new_new_n8249__ & ~new_new_n8263__;
  assign new_new_n8265__ = ~new_new_n8167__ & ~new_new_n8264__;
  assign new_new_n8266__ = ~new_new_n8166__ & ~new_new_n8265__;
  assign new_new_n8267__ = ~new_new_n8053__ & ~new_new_n8054__;
  assign new_new_n8268__ = ~new_new_n8058__ & new_new_n8267__;
  assign new_new_n8269__ = new_new_n8058__ & ~new_new_n8267__;
  assign new_new_n8270__ = ~new_new_n8268__ & ~new_new_n8269__;
  assign new_new_n8271__ = new_new_n8266__ & ~new_new_n8270__;
  assign new_new_n8272__ = ~new_new_n8266__ & new_new_n8270__;
  assign new_new_n8273__ = ~new_new_n4550__ & new_new_n6959__;
  assign new_new_n8274__ = ~new_new_n868__ & new_new_n7935__;
  assign new_new_n8275__ = ~new_new_n1061__ & new_new_n6964__;
  assign new_new_n8276__ = ~new_new_n1207__ & new_new_n6968__;
  assign new_new_n8277__ = ~new_new_n8274__ & ~new_new_n8275__;
  assign new_new_n8278__ = ~new_new_n8276__ & new_new_n8277__;
  assign new_new_n8279__ = ~new_new_n8273__ & new_new_n8278__;
  assign new_new_n8280__ = pi17 & ~new_new_n8279__;
  assign new_new_n8281__ = ~pi17 & new_new_n8279__;
  assign new_new_n8282__ = ~new_new_n8280__ & ~new_new_n8281__;
  assign new_new_n8283__ = ~new_new_n8272__ & new_new_n8282__;
  assign new_new_n8284__ = ~new_new_n8271__ & ~new_new_n8283__;
  assign new_new_n8285__ = new_new_n8148__ & new_new_n8284__;
  assign new_new_n8286__ = ~new_new_n7888__ & new_new_n8060__;
  assign new_new_n8287__ = new_new_n7888__ & ~new_new_n8060__;
  assign new_new_n8288__ = ~new_new_n8286__ & ~new_new_n8287__;
  assign new_new_n8289__ = new_new_n7947__ & new_new_n8288__;
  assign new_new_n8290__ = ~new_new_n7947__ & ~new_new_n8288__;
  assign new_new_n8291__ = ~new_new_n8289__ & ~new_new_n8290__;
  assign new_new_n8292__ = ~new_new_n7930__ & ~new_new_n8291__;
  assign new_new_n8293__ = ~new_new_n8148__ & ~new_new_n8284__;
  assign new_new_n8294__ = new_new_n7930__ & new_new_n8291__;
  assign new_new_n8295__ = ~new_new_n8292__ & ~new_new_n8293__;
  assign new_new_n8296__ = ~new_new_n8294__ & new_new_n8295__;
  assign new_new_n8297__ = ~new_new_n8285__ & ~new_new_n8296__;
  assign new_new_n8298__ = new_new_n8131__ & ~new_new_n8297__;
  assign new_new_n8299__ = ~pi10 & ~new_new_n466__;
  assign new_new_n8300__ = pi11 & ~new_new_n8299__;
  assign new_new_n8301__ = ~pi08 & ~pi09;
  assign new_new_n8302__ = ~pi10 & ~pi11;
  assign new_new_n8303__ = ~new_new_n8301__ & ~new_new_n8302__;
  assign new_new_n8304__ = ~new_new_n466__ & new_new_n8303__;
  assign new_new_n8305__ = ~new_new_n8300__ & ~new_new_n8304__;
  assign new_new_n8306__ = pi08 & pi09;
  assign new_new_n8307__ = ~new_new_n4168__ & ~new_new_n8299__;
  assign new_new_n8308__ = pi11 & new_new_n4168__;
  assign new_new_n8309__ = ~new_new_n8306__ & ~new_new_n8307__;
  assign new_new_n8310__ = ~new_new_n8308__ & new_new_n8309__;
  assign new_new_n8311__ = ~new_new_n8305__ & ~new_new_n8310__;
  assign new_new_n8312__ = ~new_new_n8131__ & new_new_n8297__;
  assign new_new_n8313__ = ~new_new_n8311__ & ~new_new_n8312__;
  assign new_new_n8314__ = ~new_new_n8298__ & ~new_new_n8313__;
  assign new_new_n8315__ = ~new_new_n8063__ & ~new_new_n8128__;
  assign new_new_n8316__ = ~new_new_n8064__ & ~new_new_n8315__;
  assign new_new_n8317__ = new_new_n8314__ & new_new_n8316__;
  assign new_new_n8318__ = ~new_new_n8314__ & ~new_new_n8316__;
  assign new_new_n8319__ = ~new_new_n3720__ & new_new_n6964__;
  assign new_new_n8320__ = ~new_new_n691__ & new_new_n7935__;
  assign new_new_n8321__ = ~new_new_n910__ & new_new_n6968__;
  assign new_new_n8322__ = ~new_new_n8319__ & ~new_new_n8320__;
  assign new_new_n8323__ = ~new_new_n8321__ & new_new_n8322__;
  assign new_new_n8324__ = new_new_n4042__ & new_new_n6958__;
  assign new_new_n8325__ = pi17 & ~new_new_n8324__;
  assign new_new_n8326__ = new_new_n4042__ & new_new_n7942__;
  assign new_new_n8327__ = ~new_new_n8325__ & ~new_new_n8326__;
  assign new_new_n8328__ = new_new_n8323__ & ~new_new_n8327__;
  assign new_new_n8329__ = ~pi17 & ~new_new_n8323__;
  assign new_new_n8330__ = ~new_new_n8328__ & ~new_new_n8329__;
  assign new_new_n8331__ = ~new_new_n1207__ & new_new_n6629__;
  assign new_new_n8332__ = ~new_new_n1061__ & ~new_new_n6625__;
  assign new_new_n8333__ = ~new_new_n868__ & new_new_n6634__;
  assign new_new_n8334__ = ~new_new_n4550__ & new_new_n6936__;
  assign new_new_n8335__ = ~new_new_n8331__ & ~new_new_n8332__;
  assign new_new_n8336__ = ~new_new_n8333__ & new_new_n8335__;
  assign new_new_n8337__ = ~new_new_n8334__ & new_new_n8336__;
  assign new_new_n8338__ = pi20 & ~new_new_n8337__;
  assign new_new_n8339__ = ~pi20 & new_new_n8337__;
  assign new_new_n8340__ = ~new_new_n8338__ & ~new_new_n8339__;
  assign new_new_n8341__ = new_new_n8092__ & ~new_new_n8117__;
  assign new_new_n8342__ = ~new_new_n8118__ & ~new_new_n8341__;
  assign new_new_n8343__ = ~new_new_n1325__ & new_new_n5183__;
  assign new_new_n8344__ = ~new_new_n4920__ & new_new_n5983__;
  assign new_new_n8345__ = new_new_n5212__ & new_new_n8344__;
  assign new_new_n8346__ = ~new_new_n3618__ & ~new_new_n5212__;
  assign new_new_n8347__ = ~new_new_n5981__ & ~new_new_n8346__;
  assign new_new_n8348__ = ~new_new_n8345__ & new_new_n8347__;
  assign new_new_n8349__ = new_new_n5195__ & ~new_new_n8348__;
  assign new_new_n8350__ = ~new_new_n8343__ & ~new_new_n8349__;
  assign new_new_n8351__ = ~new_new_n1556__ & new_new_n5185__;
  assign new_new_n8352__ = pi23 & ~new_new_n8351__;
  assign new_new_n8353__ = ~new_new_n1556__ & new_new_n5188__;
  assign new_new_n8354__ = ~pi23 & ~new_new_n8353__;
  assign new_new_n8355__ = pi20 & ~new_new_n8354__;
  assign new_new_n8356__ = ~new_new_n8352__ & ~new_new_n8355__;
  assign new_new_n8357__ = new_new_n8350__ & ~new_new_n8356__;
  assign new_new_n8358__ = ~pi23 & ~new_new_n8350__;
  assign new_new_n8359__ = ~new_new_n8357__ & ~new_new_n8358__;
  assign new_new_n8360__ = ~new_new_n8108__ & new_new_n8111__;
  assign new_new_n8361__ = ~new_new_n8107__ & ~new_new_n8360__;
  assign new_new_n8362__ = new_new_n8359__ & new_new_n8361__;
  assign new_new_n8363__ = ~new_new_n8359__ & ~new_new_n8361__;
  assign new_new_n8364__ = ~new_new_n8362__ & ~new_new_n8363__;
  assign new_new_n8365__ = ~new_new_n6903__ & ~new_new_n6904__;
  assign new_new_n8366__ = new_new_n6916__ & new_new_n8365__;
  assign new_new_n8367__ = ~new_new_n6916__ & ~new_new_n8365__;
  assign new_new_n8368__ = ~new_new_n8366__ & ~new_new_n8367__;
  assign new_new_n8369__ = new_new_n8364__ & ~new_new_n8368__;
  assign new_new_n8370__ = ~new_new_n8364__ & new_new_n8368__;
  assign new_new_n8371__ = ~new_new_n8369__ & ~new_new_n8370__;
  assign new_new_n8372__ = new_new_n8342__ & ~new_new_n8371__;
  assign new_new_n8373__ = ~new_new_n8342__ & new_new_n8371__;
  assign new_new_n8374__ = ~new_new_n8372__ & ~new_new_n8373__;
  assign new_new_n8375__ = new_new_n8340__ & ~new_new_n8374__;
  assign new_new_n8376__ = ~new_new_n8340__ & new_new_n8374__;
  assign new_new_n8377__ = ~new_new_n8375__ & ~new_new_n8376__;
  assign new_new_n8378__ = ~new_new_n8330__ & ~new_new_n8377__;
  assign new_new_n8379__ = ~new_new_n8081__ & ~new_new_n8124__;
  assign new_new_n8380__ = ~new_new_n8123__ & ~new_new_n8379__;
  assign new_new_n8381__ = new_new_n8330__ & new_new_n8377__;
  assign new_new_n8382__ = new_new_n8380__ & ~new_new_n8381__;
  assign new_new_n8383__ = ~new_new_n8378__ & ~new_new_n8382__;
  assign new_new_n8384__ = ~new_new_n3768__ & new_new_n6991__;
  assign new_new_n8385__ = ~new_new_n466__ & new_new_n6985__;
  assign new_new_n8386__ = ~new_new_n8384__ & ~new_new_n8385__;
  assign new_new_n8387__ = pi14 & ~new_new_n8386__;
  assign new_new_n8388__ = ~pi13 & new_new_n6994__;
  assign new_new_n8389__ = new_new_n6952__ & new_new_n8388__;
  assign new_new_n8390__ = new_new_n6952__ & new_new_n6994__;
  assign new_new_n8391__ = ~pi14 & new_new_n8386__;
  assign new_new_n8392__ = ~new_new_n8390__ & new_new_n8391__;
  assign new_new_n8393__ = ~new_new_n8387__ & ~new_new_n8389__;
  assign new_new_n8394__ = ~new_new_n8392__ & new_new_n8393__;
  assign new_new_n8395__ = new_new_n8383__ & ~new_new_n8394__;
  assign new_new_n8396__ = ~new_new_n8383__ & new_new_n8394__;
  assign new_new_n8397__ = ~new_new_n8395__ & ~new_new_n8396__;
  assign new_new_n8398__ = ~new_new_n910__ & new_new_n6964__;
  assign new_new_n8399__ = ~new_new_n691__ & new_new_n6968__;
  assign new_new_n8400__ = new_new_n3742__ & new_new_n6959__;
  assign new_new_n8401__ = ~new_new_n8398__ & ~new_new_n8399__;
  assign new_new_n8402__ = ~new_new_n8400__ & new_new_n8401__;
  assign new_new_n8403__ = ~new_new_n583__ & new_new_n6958__;
  assign new_new_n8404__ = ~pi17 & ~new_new_n8403__;
  assign new_new_n8405__ = ~new_new_n583__ & new_new_n7942__;
  assign new_new_n8406__ = ~new_new_n8404__ & ~new_new_n8405__;
  assign new_new_n8407__ = new_new_n8402__ & ~new_new_n8406__;
  assign new_new_n8408__ = pi17 & ~new_new_n8402__;
  assign new_new_n8409__ = ~new_new_n8407__ & ~new_new_n8408__;
  assign new_new_n8410__ = new_new_n8340__ & ~new_new_n8373__;
  assign new_new_n8411__ = ~new_new_n8372__ & ~new_new_n8410__;
  assign new_new_n8412__ = ~new_new_n8409__ & new_new_n8411__;
  assign new_new_n8413__ = new_new_n8409__ & ~new_new_n8411__;
  assign new_new_n8414__ = ~new_new_n8412__ & ~new_new_n8413__;
  assign new_new_n8415__ = ~new_new_n1207__ & ~new_new_n6625__;
  assign new_new_n8416__ = ~new_new_n3720__ & new_new_n6634__;
  assign new_new_n8417__ = ~new_new_n868__ & new_new_n6629__;
  assign new_new_n8418__ = ~new_new_n8415__ & ~new_new_n8416__;
  assign new_new_n8419__ = ~new_new_n8417__ & new_new_n8418__;
  assign new_new_n8420__ = ~new_new_n5927__ & new_new_n6631__;
  assign new_new_n8421__ = pi20 & ~new_new_n8420__;
  assign new_new_n8422__ = ~new_new_n5927__ & new_new_n6640__;
  assign new_new_n8423__ = ~new_new_n8421__ & ~new_new_n8422__;
  assign new_new_n8424__ = new_new_n8419__ & ~new_new_n8423__;
  assign new_new_n8425__ = ~pi20 & ~new_new_n8419__;
  assign new_new_n8426__ = ~new_new_n8424__ & ~new_new_n8425__;
  assign new_new_n8427__ = ~new_new_n6734__ & ~new_new_n6735__;
  assign new_new_n8428__ = ~new_new_n6918__ & new_new_n8427__;
  assign new_new_n8429__ = new_new_n6918__ & ~new_new_n8427__;
  assign new_new_n8430__ = ~new_new_n8428__ & ~new_new_n8429__;
  assign new_new_n8431__ = new_new_n8426__ & new_new_n8430__;
  assign new_new_n8432__ = ~new_new_n8426__ & ~new_new_n8430__;
  assign new_new_n8433__ = ~new_new_n8431__ & ~new_new_n8432__;
  assign new_new_n8434__ = ~new_new_n8363__ & ~new_new_n8368__;
  assign new_new_n8435__ = ~new_new_n8362__ & ~new_new_n8434__;
  assign new_new_n8436__ = new_new_n8433__ & ~new_new_n8435__;
  assign new_new_n8437__ = ~new_new_n8433__ & new_new_n8435__;
  assign new_new_n8438__ = ~new_new_n8436__ & ~new_new_n8437__;
  assign new_new_n8439__ = new_new_n8414__ & new_new_n8438__;
  assign new_new_n8440__ = ~new_new_n8414__ & ~new_new_n8438__;
  assign new_new_n8441__ = ~new_new_n8439__ & ~new_new_n8440__;
  assign new_new_n8442__ = new_new_n8397__ & ~new_new_n8441__;
  assign new_new_n8443__ = ~new_new_n8397__ & new_new_n8441__;
  assign new_new_n8444__ = ~new_new_n8442__ & ~new_new_n8443__;
  assign new_new_n8445__ = ~new_new_n8318__ & new_new_n8444__;
  assign new_new_n8446__ = ~new_new_n3768__ & new_new_n6985__;
  assign new_new_n8447__ = ~new_new_n583__ & new_new_n6991__;
  assign new_new_n8448__ = ~new_new_n8446__ & ~new_new_n8447__;
  assign new_new_n8449__ = new_new_n5194__ & new_new_n6994__;
  assign new_new_n8450__ = new_new_n8448__ & ~new_new_n8449__;
  assign new_new_n8451__ = pi14 & ~new_new_n8450__;
  assign new_new_n8452__ = ~new_new_n4170__ & new_new_n6994__;
  assign new_new_n8453__ = ~pi14 & new_new_n8448__;
  assign new_new_n8454__ = ~new_new_n8452__ & new_new_n8453__;
  assign new_new_n8455__ = pi13 & new_new_n4172__;
  assign new_new_n8456__ = ~pi13 & ~new_new_n466__;
  assign new_new_n8457__ = new_new_n8452__ & ~new_new_n8456__;
  assign new_new_n8458__ = ~new_new_n8455__ & new_new_n8457__;
  assign new_new_n8459__ = ~new_new_n8451__ & ~new_new_n8454__;
  assign new_new_n8460__ = ~new_new_n8458__ & new_new_n8459__;
  assign new_new_n8461__ = ~new_new_n8445__ & ~new_new_n8460__;
  assign new_new_n8462__ = ~new_new_n8378__ & ~new_new_n8381__;
  assign new_new_n8463__ = new_new_n8380__ & new_new_n8462__;
  assign new_new_n8464__ = ~new_new_n8380__ & ~new_new_n8462__;
  assign new_new_n8465__ = ~new_new_n8463__ & ~new_new_n8464__;
  assign new_new_n8466__ = ~pi10 & pi11;
  assign new_new_n8467__ = pi10 & ~pi11;
  assign new_new_n8468__ = ~new_new_n8466__ & ~new_new_n8467__;
  assign new_new_n8469__ = ~new_new_n8301__ & ~new_new_n8306__;
  assign new_new_n8470__ = ~new_new_n8468__ & new_new_n8469__;
  assign new_new_n8471__ = new_new_n6952__ & new_new_n8470__;
  assign new_new_n8472__ = pi10 & ~new_new_n8301__;
  assign new_new_n8473__ = ~pi10 & ~new_new_n8306__;
  assign new_new_n8474__ = ~new_new_n8472__ & ~new_new_n8473__;
  assign new_new_n8475__ = ~new_new_n466__ & new_new_n8474__;
  assign new_new_n8476__ = new_new_n8306__ & new_new_n8467__;
  assign new_new_n8477__ = ~pi10 & new_new_n8301__;
  assign new_new_n8478__ = pi11 & new_new_n8477__;
  assign new_new_n8479__ = ~new_new_n8476__ & ~new_new_n8478__;
  assign new_new_n8480__ = ~new_new_n3768__ & ~new_new_n8479__;
  assign new_new_n8481__ = ~new_new_n8475__ & ~new_new_n8480__;
  assign new_new_n8482__ = ~new_new_n8471__ & new_new_n8481__;
  assign new_new_n8483__ = pi11 & ~new_new_n8482__;
  assign new_new_n8484__ = ~pi11 & new_new_n8482__;
  assign new_new_n8485__ = ~new_new_n8483__ & ~new_new_n8484__;
  assign new_new_n8486__ = ~new_new_n910__ & new_new_n6985__;
  assign new_new_n8487__ = ~new_new_n3720__ & new_new_n6991__;
  assign new_new_n8488__ = ~new_new_n8486__ & ~new_new_n8487__;
  assign new_new_n8489__ = ~new_new_n691__ & new_new_n6994__;
  assign new_new_n8490__ = new_new_n4042__ & new_new_n8489__;
  assign new_new_n8491__ = new_new_n8488__ & ~new_new_n8490__;
  assign new_new_n8492__ = ~pi14 & ~new_new_n8491__;
  assign new_new_n8493__ = ~pi13 & new_new_n691__;
  assign new_new_n8494__ = pi13 & ~new_new_n691__;
  assign new_new_n8495__ = new_new_n6994__ & ~new_new_n8493__;
  assign new_new_n8496__ = ~new_new_n8494__ & new_new_n8495__;
  assign new_new_n8497__ = new_new_n4039__ & new_new_n8496__;
  assign new_new_n8498__ = ~new_new_n4040__ & new_new_n6994__;
  assign new_new_n8499__ = pi14 & new_new_n8488__;
  assign new_new_n8500__ = ~new_new_n8498__ & new_new_n8499__;
  assign new_new_n8501__ = ~new_new_n8497__ & ~new_new_n8500__;
  assign new_new_n8502__ = ~new_new_n8492__ & new_new_n8501__;
  assign new_new_n8503__ = ~new_new_n8271__ & ~new_new_n8272__;
  assign new_new_n8504__ = ~new_new_n8282__ & new_new_n8503__;
  assign new_new_n8505__ = new_new_n8282__ & ~new_new_n8503__;
  assign new_new_n8506__ = ~new_new_n8504__ & ~new_new_n8505__;
  assign new_new_n8507__ = ~new_new_n8502__ & ~new_new_n8506__;
  assign new_new_n8508__ = new_new_n8502__ & new_new_n8506__;
  assign new_new_n8509__ = new_new_n4926__ & new_new_n6959__;
  assign new_new_n8510__ = ~new_new_n1325__ & new_new_n6964__;
  assign new_new_n8511__ = ~new_new_n3618__ & new_new_n6968__;
  assign new_new_n8512__ = ~new_new_n8510__ & ~new_new_n8511__;
  assign new_new_n8513__ = ~new_new_n8509__ & new_new_n8512__;
  assign new_new_n8514__ = ~new_new_n1061__ & new_new_n6958__;
  assign new_new_n8515__ = ~pi17 & ~new_new_n8514__;
  assign new_new_n8516__ = ~new_new_n1061__ & new_new_n7942__;
  assign new_new_n8517__ = ~new_new_n8515__ & ~new_new_n8516__;
  assign new_new_n8518__ = new_new_n8513__ & ~new_new_n8517__;
  assign new_new_n8519__ = pi17 & ~new_new_n8513__;
  assign new_new_n8520__ = ~new_new_n8518__ & ~new_new_n8519__;
  assign new_new_n8521__ = ~new_new_n1737__ & new_new_n6634__;
  assign new_new_n8522__ = ~new_new_n1902__ & ~new_new_n6625__;
  assign new_new_n8523__ = ~new_new_n1660__ & new_new_n6629__;
  assign new_new_n8524__ = ~new_new_n8521__ & ~new_new_n8522__;
  assign new_new_n8525__ = ~new_new_n8523__ & new_new_n8524__;
  assign new_new_n8526__ = new_new_n5688__ & new_new_n6631__;
  assign new_new_n8527__ = ~pi20 & ~new_new_n8526__;
  assign new_new_n8528__ = new_new_n5688__ & new_new_n7015__;
  assign new_new_n8529__ = ~new_new_n8527__ & ~new_new_n8528__;
  assign new_new_n8530__ = new_new_n8525__ & ~new_new_n8529__;
  assign new_new_n8531__ = pi20 & ~new_new_n8525__;
  assign new_new_n8532__ = ~new_new_n8530__ & ~new_new_n8531__;
  assign new_new_n8533__ = ~new_new_n8209__ & ~new_new_n8210__;
  assign new_new_n8534__ = new_new_n5215__ & new_new_n6854__;
  assign new_new_n8535__ = ~new_new_n2130__ & new_new_n5183__;
  assign new_new_n8536__ = ~new_new_n8534__ & ~new_new_n8535__;
  assign new_new_n8537__ = ~new_new_n3535__ & new_new_n5213__;
  assign new_new_n8538__ = ~new_new_n2024__ & new_new_n5191__;
  assign new_new_n8539__ = ~new_new_n8537__ & ~new_new_n8538__;
  assign new_new_n8540__ = new_new_n8536__ & new_new_n8539__;
  assign new_new_n8541__ = pi23 & ~new_new_n8540__;
  assign new_new_n8542__ = new_new_n2024__ & ~new_new_n5213__;
  assign new_new_n8543__ = new_new_n5191__ & ~new_new_n8542__;
  assign new_new_n8544__ = ~pi23 & ~new_new_n8537__;
  assign new_new_n8545__ = ~new_new_n8543__ & new_new_n8544__;
  assign new_new_n8546__ = new_new_n8536__ & new_new_n8545__;
  assign new_new_n8547__ = ~new_new_n8541__ & ~new_new_n8546__;
  assign new_new_n8548__ = ~new_new_n333__ & ~new_new_n2572__;
  assign new_new_n8549__ = new_new_n873__ & ~new_new_n2313__;
  assign new_new_n8550__ = ~new_new_n8548__ & ~new_new_n8549__;
  assign new_new_n8551__ = new_new_n801__ & new_new_n6749__;
  assign new_new_n8552__ = new_new_n8550__ & ~new_new_n8551__;
  assign new_new_n8553__ = pi26 & ~new_new_n8552__;
  assign new_new_n8554__ = new_new_n512__ & ~new_new_n2420__;
  assign new_new_n8555__ = new_new_n6748__ & new_new_n8554__;
  assign new_new_n8556__ = ~new_new_n991__ & ~new_new_n8555__;
  assign new_new_n8557__ = new_new_n8550__ & ~new_new_n8556__;
  assign new_new_n8558__ = ~pi26 & new_new_n8550__;
  assign new_new_n8559__ = ~new_new_n6748__ & ~new_new_n8558__;
  assign new_new_n8560__ = ~new_new_n4899__ & new_new_n6748__;
  assign new_new_n8561__ = new_new_n2420__ & ~new_new_n8559__;
  assign new_new_n8562__ = ~new_new_n8560__ & new_new_n8561__;
  assign new_new_n8563__ = ~new_new_n8557__ & ~new_new_n8562__;
  assign new_new_n8564__ = ~new_new_n8553__ & new_new_n8563__;
  assign new_new_n8565__ = ~new_new_n7515__ & ~new_new_n7516__;
  assign new_new_n8566__ = ~new_new_n2848__ & new_new_n7065__;
  assign new_new_n8567__ = ~new_new_n2960__ & new_new_n7057__;
  assign new_new_n8568__ = new_new_n3460__ & ~new_new_n8567__;
  assign new_new_n8569__ = ~new_new_n8566__ & ~new_new_n8568__;
  assign new_new_n8570__ = ~new_new_n2886__ & new_new_n7065__;
  assign new_new_n8571__ = ~new_new_n7077__ & ~new_new_n8570__;
  assign new_new_n8572__ = new_new_n8569__ & new_new_n8571__;
  assign new_new_n8573__ = ~new_new_n8569__ & ~new_new_n8571__;
  assign new_new_n8574__ = ~new_new_n8572__ & ~new_new_n8573__;
  assign new_new_n8575__ = new_new_n4813__ & ~new_new_n8574__;
  assign new_new_n8576__ = ~new_new_n2886__ & new_new_n4815__;
  assign new_new_n8577__ = ~new_new_n2848__ & new_new_n4212__;
  assign new_new_n8578__ = ~new_new_n8576__ & ~new_new_n8577__;
  assign new_new_n8579__ = ~new_new_n8575__ & new_new_n8578__;
  assign new_new_n8580__ = new_new_n67__ & ~new_new_n3460__;
  assign new_new_n8581__ = pi29 & ~new_new_n8580__;
  assign new_new_n8582__ = new_new_n65__ & ~new_new_n3460__;
  assign new_new_n8583__ = ~pi29 & ~new_new_n8582__;
  assign new_new_n8584__ = pi26 & ~new_new_n8583__;
  assign new_new_n8585__ = ~new_new_n8581__ & ~new_new_n8584__;
  assign new_new_n8586__ = new_new_n8579__ & ~new_new_n8585__;
  assign new_new_n8587__ = ~pi29 & ~new_new_n8579__;
  assign new_new_n8588__ = ~new_new_n8586__ & ~new_new_n8587__;
  assign new_new_n8589__ = new_new_n8565__ & ~new_new_n8588__;
  assign new_new_n8590__ = ~new_new_n8565__ & new_new_n8588__;
  assign new_new_n8591__ = ~new_new_n8589__ & ~new_new_n8590__;
  assign new_new_n8592__ = new_new_n7697__ & new_new_n8591__;
  assign new_new_n8593__ = ~new_new_n7697__ & ~new_new_n8591__;
  assign new_new_n8594__ = ~new_new_n8592__ & ~new_new_n8593__;
  assign new_new_n8595__ = ~new_new_n7646__ & ~new_new_n7647__;
  assign new_new_n8596__ = ~new_new_n2960__ & new_new_n4815__;
  assign new_new_n8597__ = ~new_new_n3126__ & new_new_n4212__;
  assign new_new_n8598__ = ~new_new_n3164__ & ~new_new_n4818__;
  assign new_new_n8599__ = ~new_new_n8597__ & ~new_new_n8598__;
  assign new_new_n8600__ = ~new_new_n8596__ & new_new_n8599__;
  assign new_new_n8601__ = new_new_n4214__ & ~new_new_n7468__;
  assign new_new_n8602__ = pi29 & ~new_new_n8601__;
  assign new_new_n8603__ = new_new_n4825__ & ~new_new_n7468__;
  assign new_new_n8604__ = ~new_new_n8602__ & ~new_new_n8603__;
  assign new_new_n8605__ = new_new_n8600__ & ~new_new_n8604__;
  assign new_new_n8606__ = ~pi29 & ~new_new_n8600__;
  assign new_new_n8607__ = ~new_new_n8605__ & ~new_new_n8606__;
  assign new_new_n8608__ = new_new_n765__ & ~new_new_n3356__;
  assign new_new_n8609__ = ~new_new_n3254__ & new_new_n4815__;
  assign new_new_n8610__ = ~new_new_n3055__ & new_new_n3356__;
  assign new_new_n8611__ = new_new_n3254__ & ~new_new_n8610__;
  assign new_new_n8612__ = ~new_new_n3254__ & new_new_n8610__;
  assign new_new_n8613__ = new_new_n4813__ & ~new_new_n8611__;
  assign new_new_n8614__ = ~new_new_n8612__ & new_new_n8613__;
  assign new_new_n8615__ = ~new_new_n3055__ & new_new_n4212__;
  assign new_new_n8616__ = ~new_new_n3356__ & ~new_new_n4818__;
  assign new_new_n8617__ = ~new_new_n8609__ & ~new_new_n8615__;
  assign new_new_n8618__ = ~new_new_n8616__ & new_new_n8617__;
  assign new_new_n8619__ = ~new_new_n8614__ & new_new_n8618__;
  assign new_new_n8620__ = pi29 & new_new_n8619__;
  assign new_new_n8621__ = ~pi28 & ~new_new_n3356__;
  assign new_new_n8622__ = new_new_n3889__ & ~new_new_n8621__;
  assign new_new_n8623__ = ~new_new_n3055__ & ~new_new_n4209__;
  assign new_new_n8624__ = ~new_new_n68__ & ~new_new_n3356__;
  assign new_new_n8625__ = ~new_new_n8623__ & ~new_new_n8624__;
  assign new_new_n8626__ = ~new_new_n8622__ & ~new_new_n8625__;
  assign new_new_n8627__ = new_new_n8620__ & ~new_new_n8626__;
  assign new_new_n8628__ = ~new_new_n8608__ & ~new_new_n8627__;
  assign new_new_n8629__ = ~new_new_n3055__ & ~new_new_n4818__;
  assign new_new_n8630__ = ~new_new_n3164__ & new_new_n4815__;
  assign new_new_n8631__ = ~new_new_n3254__ & new_new_n4212__;
  assign new_new_n8632__ = ~new_new_n8629__ & ~new_new_n8630__;
  assign new_new_n8633__ = ~new_new_n8631__ & new_new_n8632__;
  assign new_new_n8634__ = ~new_new_n3357__ & ~new_new_n7560__;
  assign new_new_n8635__ = ~new_new_n8611__ & ~new_new_n8634__;
  assign new_new_n8636__ = new_new_n8611__ & new_new_n8634__;
  assign new_new_n8637__ = ~new_new_n8635__ & ~new_new_n8636__;
  assign new_new_n8638__ = new_new_n4214__ & ~new_new_n8637__;
  assign new_new_n8639__ = pi29 & ~new_new_n8638__;
  assign new_new_n8640__ = new_new_n4825__ & ~new_new_n8637__;
  assign new_new_n8641__ = ~new_new_n8639__ & ~new_new_n8640__;
  assign new_new_n8642__ = new_new_n8633__ & ~new_new_n8641__;
  assign new_new_n8643__ = ~pi29 & ~new_new_n8633__;
  assign new_new_n8644__ = ~new_new_n8642__ & ~new_new_n8643__;
  assign new_new_n8645__ = ~new_new_n8628__ & ~new_new_n8644__;
  assign new_new_n8646__ = ~new_new_n5052__ & ~new_new_n5059__;
  assign new_new_n8647__ = ~new_new_n3356__ & new_new_n8646__;
  assign new_new_n8648__ = new_new_n765__ & ~new_new_n3055__;
  assign new_new_n8649__ = ~new_new_n8647__ & new_new_n8648__;
  assign new_new_n8650__ = new_new_n8647__ & ~new_new_n8648__;
  assign new_new_n8651__ = ~new_new_n8649__ & ~new_new_n8650__;
  assign new_new_n8652__ = new_new_n8645__ & ~new_new_n8651__;
  assign new_new_n8653__ = ~new_new_n8645__ & new_new_n8651__;
  assign new_new_n8654__ = ~new_new_n3254__ & ~new_new_n4818__;
  assign new_new_n8655__ = ~new_new_n3164__ & new_new_n4212__;
  assign new_new_n8656__ = ~new_new_n3126__ & new_new_n4815__;
  assign new_new_n8657__ = new_new_n4813__ & ~new_new_n7570__;
  assign new_new_n8658__ = ~new_new_n8654__ & ~new_new_n8655__;
  assign new_new_n8659__ = ~new_new_n8656__ & new_new_n8658__;
  assign new_new_n8660__ = ~new_new_n8657__ & new_new_n8659__;
  assign new_new_n8661__ = ~pi29 & ~new_new_n8660__;
  assign new_new_n8662__ = pi29 & new_new_n8660__;
  assign new_new_n8663__ = ~new_new_n8661__ & ~new_new_n8662__;
  assign new_new_n8664__ = ~new_new_n8653__ & ~new_new_n8663__;
  assign new_new_n8665__ = ~new_new_n8652__ & ~new_new_n8664__;
  assign new_new_n8666__ = new_new_n8607__ & new_new_n8665__;
  assign new_new_n8667__ = ~new_new_n2960__ & new_new_n4212__;
  assign new_new_n8668__ = ~new_new_n3126__ & ~new_new_n4818__;
  assign new_new_n8669__ = ~new_new_n3460__ & new_new_n4815__;
  assign new_new_n8670__ = ~new_new_n8668__ & ~new_new_n8669__;
  assign new_new_n8671__ = ~new_new_n8667__ & new_new_n8670__;
  assign new_new_n8672__ = new_new_n4214__ & new_new_n7391__;
  assign new_new_n8673__ = pi29 & ~new_new_n8672__;
  assign new_new_n8674__ = new_new_n4825__ & new_new_n7391__;
  assign new_new_n8675__ = ~new_new_n8673__ & ~new_new_n8674__;
  assign new_new_n8676__ = new_new_n8671__ & ~new_new_n8675__;
  assign new_new_n8677__ = ~pi29 & ~new_new_n8671__;
  assign new_new_n8678__ = ~new_new_n8676__ & ~new_new_n8677__;
  assign new_new_n8679__ = ~new_new_n8666__ & ~new_new_n8678__;
  assign new_new_n8680__ = ~new_new_n7693__ & ~new_new_n8679__;
  assign new_new_n8681__ = ~new_new_n8607__ & ~new_new_n8665__;
  assign new_new_n8682__ = new_new_n7677__ & new_new_n7692__;
  assign new_new_n8683__ = ~new_new_n8678__ & ~new_new_n8682__;
  assign new_new_n8684__ = ~new_new_n8681__ & ~new_new_n8683__;
  assign new_new_n8685__ = ~new_new_n8680__ & ~new_new_n8684__;
  assign new_new_n8686__ = ~new_new_n8595__ & ~new_new_n8685__;
  assign new_new_n8687__ = ~new_new_n8666__ & ~new_new_n8682__;
  assign new_new_n8688__ = new_new_n8678__ & ~new_new_n8681__;
  assign new_new_n8689__ = ~new_new_n8687__ & new_new_n8688__;
  assign new_new_n8690__ = ~new_new_n8678__ & new_new_n8681__;
  assign new_new_n8691__ = new_new_n7693__ & new_new_n8595__;
  assign new_new_n8692__ = ~new_new_n8690__ & new_new_n8691__;
  assign new_new_n8693__ = ~new_new_n8689__ & ~new_new_n8692__;
  assign new_new_n8694__ = ~new_new_n8686__ & new_new_n8693__;
  assign new_new_n8695__ = ~new_new_n7580__ & ~new_new_n7581__;
  assign new_new_n8696__ = ~new_new_n7695__ & new_new_n8695__;
  assign new_new_n8697__ = new_new_n7695__ & ~new_new_n8695__;
  assign new_new_n8698__ = ~new_new_n8696__ & ~new_new_n8697__;
  assign new_new_n8699__ = ~new_new_n8694__ & ~new_new_n8698__;
  assign new_new_n8700__ = new_new_n8694__ & new_new_n8698__;
  assign new_new_n8701__ = ~new_new_n2960__ & ~new_new_n4818__;
  assign new_new_n8702__ = ~new_new_n2848__ & new_new_n4815__;
  assign new_new_n8703__ = ~new_new_n3460__ & new_new_n4212__;
  assign new_new_n8704__ = ~new_new_n8702__ & ~new_new_n8703__;
  assign new_new_n8705__ = ~new_new_n8701__ & new_new_n8704__;
  assign new_new_n8706__ = new_new_n4214__ & ~new_new_n7065__;
  assign new_new_n8707__ = pi29 & ~new_new_n8706__;
  assign new_new_n8708__ = new_new_n4825__ & ~new_new_n7065__;
  assign new_new_n8709__ = ~new_new_n8707__ & ~new_new_n8708__;
  assign new_new_n8710__ = new_new_n8705__ & ~new_new_n8709__;
  assign new_new_n8711__ = ~pi29 & ~new_new_n8705__;
  assign new_new_n8712__ = ~new_new_n8710__ & ~new_new_n8711__;
  assign new_new_n8713__ = ~new_new_n8700__ & new_new_n8712__;
  assign new_new_n8714__ = ~new_new_n8699__ & ~new_new_n8713__;
  assign new_new_n8715__ = ~new_new_n8594__ & ~new_new_n8714__;
  assign new_new_n8716__ = new_new_n8588__ & new_new_n8594__;
  assign new_new_n8717__ = ~new_new_n8715__ & ~new_new_n8716__;
  assign new_new_n8718__ = ~new_new_n7441__ & ~new_new_n7442__;
  assign new_new_n8719__ = ~new_new_n7699__ & new_new_n8718__;
  assign new_new_n8720__ = new_new_n7699__ & ~new_new_n8718__;
  assign new_new_n8721__ = ~new_new_n8719__ & ~new_new_n8720__;
  assign new_new_n8722__ = ~new_new_n8717__ & ~new_new_n8721__;
  assign new_new_n8723__ = new_new_n8717__ & new_new_n8721__;
  assign new_new_n8724__ = ~new_new_n2737__ & new_new_n4815__;
  assign new_new_n8725__ = ~new_new_n2886__ & new_new_n4212__;
  assign new_new_n8726__ = ~new_new_n2848__ & ~new_new_n4818__;
  assign new_new_n8727__ = new_new_n4813__ & ~new_new_n7378__;
  assign new_new_n8728__ = ~new_new_n8724__ & ~new_new_n8725__;
  assign new_new_n8729__ = ~new_new_n8726__ & new_new_n8728__;
  assign new_new_n8730__ = ~new_new_n8727__ & new_new_n8729__;
  assign new_new_n8731__ = ~pi29 & ~new_new_n8730__;
  assign new_new_n8732__ = pi29 & new_new_n8730__;
  assign new_new_n8733__ = ~new_new_n8731__ & ~new_new_n8732__;
  assign new_new_n8734__ = ~new_new_n8723__ & new_new_n8733__;
  assign new_new_n8735__ = ~new_new_n8722__ & ~new_new_n8734__;
  assign new_new_n8736__ = ~new_new_n7722__ & ~new_new_n7723__;
  assign new_new_n8737__ = new_new_n7764__ & ~new_new_n8736__;
  assign new_new_n8738__ = ~new_new_n7764__ & new_new_n8736__;
  assign new_new_n8739__ = ~new_new_n8737__ & ~new_new_n8738__;
  assign new_new_n8740__ = ~new_new_n8735__ & ~new_new_n8739__;
  assign new_new_n8741__ = new_new_n8735__ & new_new_n8739__;
  assign new_new_n8742__ = new_new_n4813__ & ~new_new_n7814__;
  assign new_new_n8743__ = ~new_new_n2886__ & ~new_new_n4818__;
  assign new_new_n8744__ = ~new_new_n2636__ & new_new_n4815__;
  assign new_new_n8745__ = ~new_new_n2737__ & new_new_n4212__;
  assign new_new_n8746__ = ~new_new_n8743__ & ~new_new_n8744__;
  assign new_new_n8747__ = ~new_new_n8745__ & new_new_n8746__;
  assign new_new_n8748__ = ~new_new_n8742__ & new_new_n8747__;
  assign new_new_n8749__ = pi29 & ~new_new_n8748__;
  assign new_new_n8750__ = new_new_n2636__ & new_new_n6793__;
  assign new_new_n8751__ = new_new_n4813__ & ~new_new_n6796__;
  assign new_new_n8752__ = new_new_n8747__ & ~new_new_n8751__;
  assign new_new_n8753__ = ~new_new_n2636__ & new_new_n8747__;
  assign new_new_n8754__ = new_new_n7811__ & new_new_n8753__;
  assign new_new_n8755__ = ~new_new_n8750__ & ~new_new_n8754__;
  assign new_new_n8756__ = ~new_new_n8752__ & new_new_n8755__;
  assign new_new_n8757__ = ~pi29 & ~new_new_n8756__;
  assign new_new_n8758__ = ~new_new_n8749__ & ~new_new_n8757__;
  assign new_new_n8759__ = ~new_new_n8741__ & ~new_new_n8758__;
  assign new_new_n8760__ = ~new_new_n8740__ & ~new_new_n8759__;
  assign new_new_n8761__ = ~new_new_n8564__ & ~new_new_n8760__;
  assign new_new_n8762__ = new_new_n8564__ & new_new_n8760__;
  assign new_new_n8763__ = ~new_new_n7782__ & ~new_new_n7783__;
  assign new_new_n8764__ = ~new_new_n7789__ & new_new_n8763__;
  assign new_new_n8765__ = new_new_n7789__ & ~new_new_n8763__;
  assign new_new_n8766__ = ~new_new_n8764__ & ~new_new_n8765__;
  assign new_new_n8767__ = ~new_new_n8762__ & ~new_new_n8766__;
  assign new_new_n8768__ = ~new_new_n8761__ & ~new_new_n8767__;
  assign new_new_n8769__ = ~new_new_n8547__ & ~new_new_n8768__;
  assign new_new_n8770__ = new_new_n8547__ & new_new_n8768__;
  assign new_new_n8771__ = ~new_new_n8769__ & ~new_new_n8770__;
  assign new_new_n8772__ = ~new_new_n8533__ & new_new_n8771__;
  assign new_new_n8773__ = ~new_new_n8222__ & new_new_n8772__;
  assign new_new_n8774__ = new_new_n8533__ & ~new_new_n8771__;
  assign new_new_n8775__ = ~new_new_n8772__ & ~new_new_n8774__;
  assign new_new_n8776__ = new_new_n8222__ & new_new_n8775__;
  assign new_new_n8777__ = new_new_n8533__ & new_new_n8776__;
  assign new_new_n8778__ = ~new_new_n8769__ & ~new_new_n8773__;
  assign new_new_n8779__ = ~new_new_n8777__ & new_new_n8778__;
  assign new_new_n8780__ = new_new_n8532__ & new_new_n8779__;
  assign new_new_n8781__ = ~new_new_n8532__ & ~new_new_n8779__;
  assign new_new_n8782__ = ~new_new_n8188__ & ~new_new_n8189__;
  assign new_new_n8783__ = ~new_new_n8224__ & new_new_n8782__;
  assign new_new_n8784__ = new_new_n8224__ & ~new_new_n8782__;
  assign new_new_n8785__ = ~new_new_n8783__ & ~new_new_n8784__;
  assign new_new_n8786__ = ~new_new_n8781__ & ~new_new_n8785__;
  assign new_new_n8787__ = ~new_new_n8780__ & ~new_new_n8786__;
  assign new_new_n8788__ = ~new_new_n8231__ & ~new_new_n8232__;
  assign new_new_n8789__ = new_new_n8242__ & new_new_n8788__;
  assign new_new_n8790__ = ~new_new_n8242__ & ~new_new_n8788__;
  assign new_new_n8791__ = ~new_new_n8789__ & ~new_new_n8790__;
  assign new_new_n8792__ = new_new_n8787__ & ~new_new_n8791__;
  assign new_new_n8793__ = ~new_new_n8787__ & new_new_n8791__;
  assign new_new_n8794__ = ~new_new_n1660__ & ~new_new_n6625__;
  assign new_new_n8795__ = ~new_new_n1466__ & new_new_n6634__;
  assign new_new_n8796__ = ~new_new_n1737__ & new_new_n6629__;
  assign new_new_n8797__ = ~new_new_n6410__ & new_new_n6936__;
  assign new_new_n8798__ = ~new_new_n8794__ & ~new_new_n8795__;
  assign new_new_n8799__ = ~new_new_n8796__ & new_new_n8798__;
  assign new_new_n8800__ = ~new_new_n8797__ & new_new_n8799__;
  assign new_new_n8801__ = pi20 & ~new_new_n8800__;
  assign new_new_n8802__ = ~pi20 & new_new_n8800__;
  assign new_new_n8803__ = ~new_new_n8801__ & ~new_new_n8802__;
  assign new_new_n8804__ = ~new_new_n8793__ & ~new_new_n8803__;
  assign new_new_n8805__ = ~new_new_n8792__ & ~new_new_n8804__;
  assign new_new_n8806__ = ~new_new_n8520__ & ~new_new_n8805__;
  assign new_new_n8807__ = new_new_n8520__ & new_new_n8805__;
  assign new_new_n8808__ = ~new_new_n8249__ & ~new_new_n8250__;
  assign new_new_n8809__ = new_new_n8262__ & ~new_new_n8808__;
  assign new_new_n8810__ = ~new_new_n8262__ & new_new_n8808__;
  assign new_new_n8811__ = ~new_new_n8809__ & ~new_new_n8810__;
  assign new_new_n8812__ = ~new_new_n8807__ & new_new_n8811__;
  assign new_new_n8813__ = ~new_new_n8806__ & ~new_new_n8812__;
  assign new_new_n8814__ = ~new_new_n8166__ & ~new_new_n8167__;
  assign new_new_n8815__ = ~new_new_n8264__ & new_new_n8814__;
  assign new_new_n8816__ = new_new_n8264__ & ~new_new_n8814__;
  assign new_new_n8817__ = ~new_new_n8815__ & ~new_new_n8816__;
  assign new_new_n8818__ = new_new_n8813__ & ~new_new_n8817__;
  assign new_new_n8819__ = ~new_new_n8813__ & new_new_n8817__;
  assign new_new_n8820__ = pi13 & new_new_n6994__;
  assign new_new_n8821__ = new_new_n5121__ & new_new_n8820__;
  assign new_new_n8822__ = ~new_new_n3720__ & new_new_n6985__;
  assign new_new_n8823__ = ~new_new_n868__ & new_new_n6991__;
  assign new_new_n8824__ = ~new_new_n8822__ & ~new_new_n8823__;
  assign new_new_n8825__ = ~new_new_n5129__ & new_new_n6994__;
  assign new_new_n8826__ = pi14 & ~new_new_n8825__;
  assign new_new_n8827__ = new_new_n5127__ & new_new_n8388__;
  assign new_new_n8828__ = ~new_new_n8826__ & ~new_new_n8827__;
  assign new_new_n8829__ = new_new_n8824__ & ~new_new_n8828__;
  assign new_new_n8830__ = new_new_n5116__ & new_new_n6994__;
  assign new_new_n8831__ = new_new_n8824__ & ~new_new_n8830__;
  assign new_new_n8832__ = ~pi14 & ~new_new_n8831__;
  assign new_new_n8833__ = ~new_new_n8821__ & ~new_new_n8832__;
  assign new_new_n8834__ = ~new_new_n8829__ & new_new_n8833__;
  assign new_new_n8835__ = ~new_new_n8819__ & ~new_new_n8834__;
  assign new_new_n8836__ = ~new_new_n8818__ & ~new_new_n8835__;
  assign new_new_n8837__ = ~new_new_n8508__ & ~new_new_n8836__;
  assign new_new_n8838__ = ~new_new_n8507__ & ~new_new_n8837__;
  assign new_new_n8839__ = new_new_n8485__ & ~new_new_n8838__;
  assign new_new_n8840__ = ~new_new_n8485__ & new_new_n8838__;
  assign new_new_n8841__ = ~new_new_n7948__ & ~new_new_n7949__;
  assign new_new_n8842__ = ~new_new_n8285__ & ~new_new_n8293__;
  assign new_new_n8843__ = new_new_n8841__ & ~new_new_n8842__;
  assign new_new_n8844__ = ~new_new_n8841__ & new_new_n8842__;
  assign new_new_n8845__ = ~new_new_n8843__ & ~new_new_n8844__;
  assign new_new_n8846__ = new_new_n8060__ & new_new_n8845__;
  assign new_new_n8847__ = ~new_new_n8060__ & ~new_new_n8845__;
  assign new_new_n8848__ = ~new_new_n8846__ & ~new_new_n8847__;
  assign new_new_n8849__ = ~new_new_n8840__ & new_new_n8848__;
  assign new_new_n8850__ = ~new_new_n8839__ & ~new_new_n8849__;
  assign new_new_n8851__ = ~pi10 & ~new_new_n910__;
  assign new_new_n8852__ = new_new_n8301__ & new_new_n8851__;
  assign new_new_n8853__ = pi11 & ~new_new_n8852__;
  assign new_new_n8854__ = pi09 & pi10;
  assign new_new_n8855__ = pi08 & new_new_n8854__;
  assign new_new_n8856__ = ~new_new_n910__ & new_new_n8855__;
  assign new_new_n8857__ = ~new_new_n8853__ & ~new_new_n8856__;
  assign new_new_n8858__ = new_new_n8468__ & new_new_n8469__;
  assign new_new_n8859__ = ~new_new_n583__ & new_new_n8858__;
  assign new_new_n8860__ = ~new_new_n691__ & new_new_n8474__;
  assign new_new_n8861__ = new_new_n3742__ & new_new_n8470__;
  assign new_new_n8862__ = ~new_new_n8859__ & ~new_new_n8860__;
  assign new_new_n8863__ = ~new_new_n8861__ & new_new_n8862__;
  assign new_new_n8864__ = ~new_new_n8857__ & new_new_n8863__;
  assign new_new_n8865__ = ~pi11 & ~new_new_n8863__;
  assign new_new_n8866__ = ~new_new_n8864__ & ~new_new_n8865__;
  assign new_new_n8867__ = ~new_new_n1061__ & new_new_n6991__;
  assign new_new_n8868__ = ~new_new_n1207__ & new_new_n6985__;
  assign new_new_n8869__ = ~new_new_n8867__ & ~new_new_n8868__;
  assign new_new_n8870__ = ~new_new_n868__ & new_new_n6994__;
  assign new_new_n8871__ = ~new_new_n4550__ & new_new_n8870__;
  assign new_new_n8872__ = new_new_n8869__ & ~new_new_n8871__;
  assign new_new_n8873__ = pi14 & ~new_new_n8872__;
  assign new_new_n8874__ = ~pi13 & ~new_new_n868__;
  assign new_new_n8875__ = pi13 & ~new_new_n4550__;
  assign new_new_n8876__ = new_new_n868__ & new_new_n4547__;
  assign new_new_n8877__ = new_new_n6994__ & ~new_new_n8876__;
  assign new_new_n8878__ = ~new_new_n8874__ & ~new_new_n8875__;
  assign new_new_n8879__ = new_new_n8877__ & new_new_n8878__;
  assign new_new_n8880__ = ~pi14 & new_new_n8869__;
  assign new_new_n8881__ = ~new_new_n8877__ & new_new_n8880__;
  assign new_new_n8882__ = ~new_new_n8873__ & ~new_new_n8881__;
  assign new_new_n8883__ = ~new_new_n8879__ & new_new_n8882__;
  assign new_new_n8884__ = ~new_new_n3618__ & new_new_n7935__;
  assign new_new_n8885__ = ~new_new_n5984__ & new_new_n6959__;
  assign new_new_n8886__ = ~new_new_n1556__ & new_new_n6964__;
  assign new_new_n8887__ = ~new_new_n1325__ & new_new_n6968__;
  assign new_new_n8888__ = ~new_new_n8884__ & ~new_new_n8886__;
  assign new_new_n8889__ = ~new_new_n8887__ & new_new_n8888__;
  assign new_new_n8890__ = ~new_new_n8885__ & new_new_n8889__;
  assign new_new_n8891__ = ~pi17 & ~new_new_n8890__;
  assign new_new_n8892__ = pi17 & new_new_n8890__;
  assign new_new_n8893__ = ~new_new_n8891__ & ~new_new_n8892__;
  assign new_new_n8894__ = ~new_new_n1325__ & new_new_n7935__;
  assign new_new_n8895__ = ~new_new_n1556__ & new_new_n6968__;
  assign new_new_n8896__ = ~new_new_n1466__ & new_new_n6964__;
  assign new_new_n8897__ = new_new_n5048__ & new_new_n6959__;
  assign new_new_n8898__ = ~new_new_n8894__ & ~new_new_n8895__;
  assign new_new_n8899__ = ~new_new_n8896__ & new_new_n8898__;
  assign new_new_n8900__ = ~new_new_n8897__ & new_new_n8899__;
  assign new_new_n8901__ = ~pi17 & ~new_new_n8900__;
  assign new_new_n8902__ = pi17 & new_new_n8900__;
  assign new_new_n8903__ = ~new_new_n8901__ & ~new_new_n8902__;
  assign new_new_n8904__ = new_new_n873__ & ~new_new_n2572__;
  assign new_new_n8905__ = ~new_new_n333__ & ~new_new_n2497__;
  assign new_new_n8906__ = ~new_new_n2313__ & new_new_n3311__;
  assign new_new_n8907__ = ~new_new_n8904__ & ~new_new_n8905__;
  assign new_new_n8908__ = ~new_new_n8906__ & new_new_n8907__;
  assign new_new_n8909__ = pi26 & ~new_new_n8908__;
  assign new_new_n8910__ = new_new_n4898__ & ~new_new_n7236__;
  assign new_new_n8911__ = new_new_n801__ & ~new_new_n7236__;
  assign new_new_n8912__ = ~pi26 & ~new_new_n8911__;
  assign new_new_n8913__ = ~new_new_n8910__ & ~new_new_n8912__;
  assign new_new_n8914__ = new_new_n8908__ & ~new_new_n8913__;
  assign new_new_n8915__ = ~new_new_n8909__ & ~new_new_n8914__;
  assign new_new_n8916__ = ~new_new_n8722__ & ~new_new_n8723__;
  assign new_new_n8917__ = new_new_n8733__ & new_new_n8916__;
  assign new_new_n8918__ = ~new_new_n8733__ & ~new_new_n8916__;
  assign new_new_n8919__ = ~new_new_n8917__ & ~new_new_n8918__;
  assign new_new_n8920__ = ~new_new_n4900__ & ~new_new_n6796__;
  assign new_new_n8921__ = ~new_new_n333__ & ~new_new_n2886__;
  assign new_new_n8922__ = ~new_new_n2636__ & new_new_n3311__;
  assign new_new_n8923__ = new_new_n873__ & ~new_new_n2737__;
  assign new_new_n8924__ = ~new_new_n8921__ & ~new_new_n8922__;
  assign new_new_n8925__ = ~new_new_n8923__ & new_new_n8924__;
  assign new_new_n8926__ = ~new_new_n8920__ & new_new_n8925__;
  assign new_new_n8927__ = ~new_new_n8750__ & ~new_new_n8926__;
  assign new_new_n8928__ = ~pi26 & ~new_new_n8927__;
  assign new_new_n8929__ = ~new_new_n4900__ & new_new_n7812__;
  assign new_new_n8930__ = new_new_n8925__ & ~new_new_n8929__;
  assign new_new_n8931__ = pi26 & ~new_new_n8930__;
  assign new_new_n8932__ = ~pi26 & new_new_n8925__;
  assign new_new_n8933__ = ~new_new_n2636__ & ~new_new_n8932__;
  assign new_new_n8934__ = new_new_n2636__ & ~new_new_n4899__;
  assign new_new_n8935__ = ~new_new_n8933__ & ~new_new_n8934__;
  assign new_new_n8936__ = new_new_n7811__ & new_new_n8935__;
  assign new_new_n8937__ = ~new_new_n8928__ & ~new_new_n8936__;
  assign new_new_n8938__ = ~new_new_n8931__ & new_new_n8937__;
  assign new_new_n8939__ = ~new_new_n7693__ & ~new_new_n8666__;
  assign new_new_n8940__ = ~new_new_n7692__ & ~new_new_n8681__;
  assign new_new_n8941__ = ~new_new_n8939__ & ~new_new_n8940__;
  assign new_new_n8942__ = ~new_new_n8595__ & new_new_n8678__;
  assign new_new_n8943__ = new_new_n8595__ & ~new_new_n8678__;
  assign new_new_n8944__ = ~new_new_n8942__ & ~new_new_n8943__;
  assign new_new_n8945__ = ~new_new_n7692__ & ~new_new_n8666__;
  assign new_new_n8946__ = new_new_n7677__ & ~new_new_n8681__;
  assign new_new_n8947__ = ~new_new_n8945__ & new_new_n8946__;
  assign new_new_n8948__ = ~new_new_n8941__ & ~new_new_n8944__;
  assign new_new_n8949__ = ~new_new_n8947__ & new_new_n8948__;
  assign new_new_n8950__ = new_new_n7693__ & new_new_n8665__;
  assign new_new_n8951__ = ~new_new_n8666__ & ~new_new_n8681__;
  assign new_new_n8952__ = ~new_new_n8682__ & new_new_n8951__;
  assign new_new_n8953__ = ~new_new_n7693__ & new_new_n8681__;
  assign new_new_n8954__ = ~new_new_n8950__ & ~new_new_n8953__;
  assign new_new_n8955__ = new_new_n8944__ & new_new_n8954__;
  assign new_new_n8956__ = ~new_new_n8952__ & new_new_n8955__;
  assign new_new_n8957__ = ~new_new_n8949__ & ~new_new_n8956__;
  assign new_new_n8958__ = new_new_n873__ & ~new_new_n2848__;
  assign new_new_n8959__ = ~new_new_n2886__ & new_new_n3311__;
  assign new_new_n8960__ = ~new_new_n333__ & ~new_new_n3460__;
  assign new_new_n8961__ = ~new_new_n4900__ & ~new_new_n8574__;
  assign new_new_n8962__ = ~new_new_n8958__ & ~new_new_n8959__;
  assign new_new_n8963__ = ~new_new_n8960__ & new_new_n8962__;
  assign new_new_n8964__ = ~new_new_n8961__ & new_new_n8963__;
  assign new_new_n8965__ = ~pi26 & ~new_new_n8964__;
  assign new_new_n8966__ = pi26 & new_new_n8964__;
  assign new_new_n8967__ = ~new_new_n8965__ & ~new_new_n8966__;
  assign new_new_n8968__ = ~new_new_n8652__ & ~new_new_n8653__;
  assign new_new_n8969__ = ~new_new_n8663__ & new_new_n8968__;
  assign new_new_n8970__ = new_new_n8663__ & ~new_new_n8968__;
  assign new_new_n8971__ = ~new_new_n8969__ & ~new_new_n8970__;
  assign new_new_n8972__ = ~new_new_n2960__ & new_new_n3311__;
  assign new_new_n8973__ = new_new_n873__ & ~new_new_n3126__;
  assign new_new_n8974__ = ~new_new_n333__ & ~new_new_n3164__;
  assign new_new_n8975__ = ~new_new_n8973__ & ~new_new_n8974__;
  assign new_new_n8976__ = ~new_new_n8972__ & new_new_n8975__;
  assign new_new_n8977__ = ~pi26 & ~new_new_n8976__;
  assign new_new_n8978__ = new_new_n512__ & ~new_new_n7468__;
  assign new_new_n8979__ = new_new_n801__ & ~new_new_n7468__;
  assign new_new_n8980__ = pi26 & ~new_new_n8979__;
  assign new_new_n8981__ = ~new_new_n8978__ & ~new_new_n8980__;
  assign new_new_n8982__ = new_new_n8976__ & ~new_new_n8981__;
  assign new_new_n8983__ = ~new_new_n8977__ & ~new_new_n8982__;
  assign new_new_n8984__ = new_new_n8626__ & ~new_new_n8983__;
  assign new_new_n8985__ = ~new_new_n333__ & ~new_new_n3254__;
  assign new_new_n8986__ = new_new_n873__ & ~new_new_n3164__;
  assign new_new_n8987__ = ~new_new_n4900__ & ~new_new_n7570__;
  assign new_new_n8988__ = ~new_new_n8985__ & ~new_new_n8986__;
  assign new_new_n8989__ = ~new_new_n8987__ & new_new_n8988__;
  assign new_new_n8990__ = ~pi26 & ~new_new_n8989__;
  assign new_new_n8991__ = ~new_new_n3126__ & new_new_n4898__;
  assign new_new_n8992__ = new_new_n801__ & ~new_new_n3126__;
  assign new_new_n8993__ = pi26 & ~new_new_n8992__;
  assign new_new_n8994__ = ~new_new_n8991__ & ~new_new_n8993__;
  assign new_new_n8995__ = new_new_n8989__ & ~new_new_n8994__;
  assign new_new_n8996__ = ~new_new_n8990__ & ~new_new_n8995__;
  assign new_new_n8997__ = ~new_new_n3356__ & new_new_n8623__;
  assign new_new_n8998__ = ~new_new_n3889__ & ~new_new_n8997__;
  assign new_new_n8999__ = pi28 & ~new_new_n8998__;
  assign new_new_n9000__ = ~new_new_n3356__ & ~new_new_n4211__;
  assign new_new_n9001__ = ~new_new_n3055__ & new_new_n4214__;
  assign new_new_n9002__ = ~new_new_n9000__ & ~new_new_n9001__;
  assign new_new_n9003__ = ~new_new_n8999__ & ~new_new_n9002__;
  assign new_new_n9004__ = ~new_new_n333__ & ~new_new_n3055__;
  assign new_new_n9005__ = ~new_new_n3164__ & new_new_n3311__;
  assign new_new_n9006__ = new_new_n873__ & ~new_new_n3254__;
  assign new_new_n9007__ = ~new_new_n9004__ & ~new_new_n9005__;
  assign new_new_n9008__ = ~new_new_n9006__ & new_new_n9007__;
  assign new_new_n9009__ = pi26 & ~new_new_n9008__;
  assign new_new_n9010__ = new_new_n4898__ & ~new_new_n8637__;
  assign new_new_n9011__ = new_new_n801__ & ~new_new_n8637__;
  assign new_new_n9012__ = ~pi26 & ~new_new_n9011__;
  assign new_new_n9013__ = ~new_new_n9010__ & ~new_new_n9012__;
  assign new_new_n9014__ = new_new_n9008__ & ~new_new_n9013__;
  assign new_new_n9015__ = ~new_new_n9009__ & ~new_new_n9014__;
  assign new_new_n9016__ = ~new_new_n3356__ & new_new_n4214__;
  assign new_new_n9017__ = new_new_n3055__ & new_new_n3356__;
  assign new_new_n9018__ = ~new_new_n110__ & ~new_new_n9017__;
  assign new_new_n9019__ = new_new_n873__ & ~new_new_n3356__;
  assign new_new_n9020__ = ~new_new_n9018__ & ~new_new_n9019__;
  assign new_new_n9021__ = ~new_new_n4900__ & new_new_n7682__;
  assign new_new_n9022__ = ~pi24 & ~new_new_n112__;
  assign new_new_n9023__ = ~new_new_n2502__ & ~new_new_n9022__;
  assign new_new_n9024__ = ~new_new_n9021__ & ~new_new_n9023__;
  assign new_new_n9025__ = ~new_new_n3055__ & ~new_new_n9024__;
  assign new_new_n9026__ = ~new_new_n3254__ & ~new_new_n4900__;
  assign new_new_n9027__ = new_new_n333__ & ~new_new_n9026__;
  assign new_new_n9028__ = ~new_new_n3356__ & ~new_new_n9027__;
  assign new_new_n9029__ = new_new_n550__ & ~new_new_n3055__;
  assign new_new_n9030__ = ~new_new_n110__ & ~new_new_n3254__;
  assign new_new_n9031__ = ~new_new_n9029__ & new_new_n9030__;
  assign new_new_n9032__ = ~new_new_n9028__ & ~new_new_n9031__;
  assign new_new_n9033__ = ~new_new_n9025__ & new_new_n9032__;
  assign new_new_n9034__ = pi26 & new_new_n9020__;
  assign new_new_n9035__ = new_new_n9033__ & new_new_n9034__;
  assign new_new_n9036__ = ~new_new_n9016__ & ~new_new_n9035__;
  assign new_new_n9037__ = new_new_n9015__ & ~new_new_n9036__;
  assign new_new_n9038__ = ~new_new_n9003__ & ~new_new_n9037__;
  assign new_new_n9039__ = ~new_new_n8996__ & ~new_new_n9038__;
  assign new_new_n9040__ = new_new_n9003__ & new_new_n9016__;
  assign new_new_n9041__ = new_new_n9015__ & new_new_n9040__;
  assign new_new_n9042__ = ~new_new_n9039__ & ~new_new_n9041__;
  assign new_new_n9043__ = ~new_new_n8984__ & new_new_n9042__;
  assign new_new_n9044__ = new_new_n8620__ & ~new_new_n9043__;
  assign new_new_n9045__ = ~pi29 & ~new_new_n8619__;
  assign new_new_n9046__ = new_new_n8983__ & ~new_new_n9045__;
  assign new_new_n9047__ = ~new_new_n8619__ & ~new_new_n8626__;
  assign new_new_n9048__ = ~new_new_n9045__ & ~new_new_n9047__;
  assign new_new_n9049__ = ~new_new_n8983__ & ~new_new_n9048__;
  assign new_new_n9050__ = new_new_n9042__ & ~new_new_n9049__;
  assign new_new_n9051__ = ~new_new_n9046__ & ~new_new_n9050__;
  assign new_new_n9052__ = ~new_new_n9044__ & ~new_new_n9051__;
  assign new_new_n9053__ = new_new_n8608__ & new_new_n8627__;
  assign new_new_n9054__ = new_new_n8628__ & new_new_n8644__;
  assign new_new_n9055__ = ~new_new_n8645__ & ~new_new_n9054__;
  assign new_new_n9056__ = ~new_new_n9053__ & ~new_new_n9055__;
  assign new_new_n9057__ = ~new_new_n9052__ & ~new_new_n9056__;
  assign new_new_n9058__ = new_new_n9052__ & new_new_n9056__;
  assign new_new_n9059__ = new_new_n873__ & ~new_new_n2960__;
  assign new_new_n9060__ = ~new_new_n333__ & ~new_new_n3126__;
  assign new_new_n9061__ = new_new_n3311__ & ~new_new_n3460__;
  assign new_new_n9062__ = ~new_new_n9060__ & ~new_new_n9061__;
  assign new_new_n9063__ = ~new_new_n9059__ & new_new_n9062__;
  assign new_new_n9064__ = pi26 & ~new_new_n9063__;
  assign new_new_n9065__ = new_new_n4898__ & new_new_n7391__;
  assign new_new_n9066__ = new_new_n801__ & new_new_n7391__;
  assign new_new_n9067__ = ~pi26 & ~new_new_n9066__;
  assign new_new_n9068__ = ~new_new_n9065__ & ~new_new_n9067__;
  assign new_new_n9069__ = new_new_n9063__ & ~new_new_n9068__;
  assign new_new_n9070__ = ~new_new_n9064__ & ~new_new_n9069__;
  assign new_new_n9071__ = ~new_new_n9058__ & new_new_n9070__;
  assign new_new_n9072__ = ~new_new_n9057__ & ~new_new_n9071__;
  assign new_new_n9073__ = new_new_n8971__ & ~new_new_n9072__;
  assign new_new_n9074__ = ~new_new_n8971__ & new_new_n9072__;
  assign new_new_n9075__ = ~new_new_n9073__ & ~new_new_n9074__;
  assign new_new_n9076__ = ~new_new_n333__ & ~new_new_n2960__;
  assign new_new_n9077__ = ~new_new_n2848__ & new_new_n3311__;
  assign new_new_n9078__ = new_new_n873__ & ~new_new_n3460__;
  assign new_new_n9079__ = ~new_new_n9077__ & ~new_new_n9078__;
  assign new_new_n9080__ = ~new_new_n9076__ & new_new_n9079__;
  assign new_new_n9081__ = pi26 & ~new_new_n9080__;
  assign new_new_n9082__ = new_new_n4898__ & ~new_new_n7065__;
  assign new_new_n9083__ = new_new_n801__ & ~new_new_n7065__;
  assign new_new_n9084__ = ~pi26 & ~new_new_n9083__;
  assign new_new_n9085__ = ~new_new_n9082__ & ~new_new_n9084__;
  assign new_new_n9086__ = new_new_n9080__ & ~new_new_n9085__;
  assign new_new_n9087__ = ~new_new_n9081__ & ~new_new_n9086__;
  assign new_new_n9088__ = new_new_n9075__ & new_new_n9087__;
  assign new_new_n9089__ = ~new_new_n9073__ & ~new_new_n9088__;
  assign new_new_n9090__ = new_new_n8967__ & new_new_n9089__;
  assign new_new_n9091__ = ~new_new_n8967__ & ~new_new_n9089__;
  assign new_new_n9092__ = ~new_new_n7693__ & ~new_new_n8682__;
  assign new_new_n9093__ = new_new_n8951__ & ~new_new_n9092__;
  assign new_new_n9094__ = ~new_new_n8951__ & new_new_n9092__;
  assign new_new_n9095__ = ~new_new_n9093__ & ~new_new_n9094__;
  assign new_new_n9096__ = ~new_new_n9091__ & new_new_n9095__;
  assign new_new_n9097__ = ~new_new_n9090__ & ~new_new_n9096__;
  assign new_new_n9098__ = ~new_new_n8957__ & new_new_n9097__;
  assign new_new_n9099__ = new_new_n8957__ & ~new_new_n9097__;
  assign new_new_n9100__ = ~new_new_n2737__ & new_new_n3311__;
  assign new_new_n9101__ = ~new_new_n333__ & ~new_new_n2848__;
  assign new_new_n9102__ = new_new_n873__ & ~new_new_n2886__;
  assign new_new_n9103__ = ~new_new_n4900__ & ~new_new_n7378__;
  assign new_new_n9104__ = ~new_new_n9100__ & ~new_new_n9101__;
  assign new_new_n9105__ = ~new_new_n9102__ & new_new_n9104__;
  assign new_new_n9106__ = ~new_new_n9103__ & new_new_n9105__;
  assign new_new_n9107__ = ~pi26 & ~new_new_n9106__;
  assign new_new_n9108__ = pi26 & new_new_n9106__;
  assign new_new_n9109__ = ~new_new_n9107__ & ~new_new_n9108__;
  assign new_new_n9110__ = ~new_new_n9099__ & ~new_new_n9109__;
  assign new_new_n9111__ = ~new_new_n9098__ & ~new_new_n9110__;
  assign new_new_n9112__ = new_new_n8938__ & ~new_new_n9111__;
  assign new_new_n9113__ = ~new_new_n8938__ & new_new_n9111__;
  assign new_new_n9114__ = ~new_new_n8699__ & ~new_new_n8700__;
  assign new_new_n9115__ = new_new_n8712__ & new_new_n9114__;
  assign new_new_n9116__ = ~new_new_n8712__ & ~new_new_n9114__;
  assign new_new_n9117__ = ~new_new_n9115__ & ~new_new_n9116__;
  assign new_new_n9118__ = ~new_new_n9113__ & ~new_new_n9117__;
  assign new_new_n9119__ = ~new_new_n9112__ & ~new_new_n9118__;
  assign new_new_n9120__ = ~new_new_n333__ & ~new_new_n2737__;
  assign new_new_n9121__ = new_new_n873__ & ~new_new_n2636__;
  assign new_new_n9122__ = ~new_new_n9120__ & ~new_new_n9121__;
  assign new_new_n9123__ = new_new_n801__ & new_new_n7772__;
  assign new_new_n9124__ = new_new_n9122__ & ~new_new_n9123__;
  assign new_new_n9125__ = pi26 & ~new_new_n9124__;
  assign new_new_n9126__ = new_new_n2497__ & new_new_n6797__;
  assign new_new_n9127__ = new_new_n801__ & ~new_new_n9126__;
  assign new_new_n9128__ = ~pi26 & ~new_new_n9127__;
  assign new_new_n9129__ = pi25 & new_new_n2497__;
  assign new_new_n9130__ = ~pi25 & ~new_new_n2497__;
  assign new_new_n9131__ = ~new_new_n110__ & ~new_new_n9129__;
  assign new_new_n9132__ = ~new_new_n9130__ & new_new_n9131__;
  assign new_new_n9133__ = ~new_new_n6797__ & new_new_n9132__;
  assign new_new_n9134__ = ~new_new_n9128__ & ~new_new_n9133__;
  assign new_new_n9135__ = new_new_n9122__ & ~new_new_n9134__;
  assign new_new_n9136__ = ~new_new_n9125__ & ~new_new_n9135__;
  assign new_new_n9137__ = new_new_n8594__ & new_new_n8714__;
  assign new_new_n9138__ = ~new_new_n8715__ & ~new_new_n9137__;
  assign new_new_n9139__ = ~new_new_n9136__ & new_new_n9138__;
  assign new_new_n9140__ = ~new_new_n9119__ & ~new_new_n9139__;
  assign new_new_n9141__ = new_new_n9136__ & ~new_new_n9138__;
  assign new_new_n9142__ = ~new_new_n9140__ & ~new_new_n9141__;
  assign new_new_n9143__ = ~new_new_n8919__ & ~new_new_n9142__;
  assign new_new_n9144__ = new_new_n8919__ & new_new_n9142__;
  assign new_new_n9145__ = ~new_new_n2572__ & new_new_n3311__;
  assign new_new_n9146__ = new_new_n873__ & ~new_new_n2497__;
  assign new_new_n9147__ = ~new_new_n333__ & ~new_new_n2636__;
  assign new_new_n9148__ = ~new_new_n4900__ & new_new_n6804__;
  assign new_new_n9149__ = ~new_new_n9145__ & ~new_new_n9146__;
  assign new_new_n9150__ = ~new_new_n9147__ & new_new_n9149__;
  assign new_new_n9151__ = ~new_new_n9148__ & new_new_n9150__;
  assign new_new_n9152__ = pi26 & ~new_new_n9151__;
  assign new_new_n9153__ = ~pi26 & new_new_n9151__;
  assign new_new_n9154__ = ~new_new_n9152__ & ~new_new_n9153__;
  assign new_new_n9155__ = ~new_new_n9144__ & new_new_n9154__;
  assign new_new_n9156__ = ~new_new_n9143__ & ~new_new_n9155__;
  assign new_new_n9157__ = ~new_new_n8915__ & new_new_n9156__;
  assign new_new_n9158__ = new_new_n8915__ & ~new_new_n9156__;
  assign new_new_n9159__ = ~new_new_n8740__ & ~new_new_n8741__;
  assign new_new_n9160__ = new_new_n8758__ & new_new_n9159__;
  assign new_new_n9161__ = ~new_new_n8758__ & ~new_new_n9159__;
  assign new_new_n9162__ = ~new_new_n9160__ & ~new_new_n9161__;
  assign new_new_n9163__ = ~new_new_n9158__ & ~new_new_n9162__;
  assign new_new_n9164__ = ~new_new_n9157__ & ~new_new_n9163__;
  assign new_new_n9165__ = ~new_new_n8761__ & ~new_new_n8762__;
  assign new_new_n9166__ = ~new_new_n8766__ & new_new_n9165__;
  assign new_new_n9167__ = new_new_n8766__ & ~new_new_n9165__;
  assign new_new_n9168__ = ~new_new_n9166__ & ~new_new_n9167__;
  assign new_new_n9169__ = ~new_new_n9164__ & new_new_n9168__;
  assign new_new_n9170__ = ~new_new_n2024__ & new_new_n5183__;
  assign new_new_n9171__ = ~new_new_n2224__ & new_new_n5191__;
  assign new_new_n9172__ = ~new_new_n9170__ & ~new_new_n9171__;
  assign new_new_n9173__ = ~new_new_n2130__ & ~new_new_n6036__;
  assign new_new_n9174__ = new_new_n5195__ & new_new_n9173__;
  assign new_new_n9175__ = new_new_n9172__ & ~new_new_n9174__;
  assign new_new_n9176__ = pi23 & ~new_new_n9175__;
  assign new_new_n9177__ = new_new_n2130__ & new_new_n6034__;
  assign new_new_n9178__ = new_new_n5195__ & ~new_new_n9177__;
  assign new_new_n9179__ = ~pi23 & ~new_new_n9178__;
  assign new_new_n9180__ = new_new_n2130__ & ~new_new_n6034__;
  assign new_new_n9181__ = ~pi22 & ~new_new_n9180__;
  assign new_new_n9182__ = ~new_new_n2130__ & new_new_n6036__;
  assign new_new_n9183__ = pi22 & ~new_new_n9182__;
  assign new_new_n9184__ = new_new_n5195__ & ~new_new_n9181__;
  assign new_new_n9185__ = ~new_new_n9183__ & new_new_n9184__;
  assign new_new_n9186__ = ~new_new_n9179__ & ~new_new_n9185__;
  assign new_new_n9187__ = new_new_n9172__ & ~new_new_n9186__;
  assign new_new_n9188__ = ~new_new_n9176__ & ~new_new_n9187__;
  assign new_new_n9189__ = new_new_n9164__ & ~new_new_n9168__;
  assign new_new_n9190__ = ~new_new_n9169__ & ~new_new_n9189__;
  assign new_new_n9191__ = ~new_new_n9188__ & new_new_n9190__;
  assign new_new_n9192__ = ~new_new_n9169__ & ~new_new_n9191__;
  assign new_new_n9193__ = ~new_new_n8222__ & ~new_new_n8775__;
  assign new_new_n9194__ = ~new_new_n8776__ & ~new_new_n9193__;
  assign new_new_n9195__ = ~new_new_n1823__ & ~new_new_n6625__;
  assign new_new_n9196__ = ~new_new_n1660__ & new_new_n6634__;
  assign new_new_n9197__ = ~new_new_n1902__ & new_new_n6629__;
  assign new_new_n9198__ = ~new_new_n5274__ & new_new_n6936__;
  assign new_new_n9199__ = ~new_new_n9195__ & ~new_new_n9196__;
  assign new_new_n9200__ = ~new_new_n9197__ & new_new_n9199__;
  assign new_new_n9201__ = ~new_new_n9198__ & new_new_n9200__;
  assign new_new_n9202__ = pi20 & ~new_new_n9201__;
  assign new_new_n9203__ = ~pi20 & new_new_n9201__;
  assign new_new_n9204__ = ~new_new_n9202__ & ~new_new_n9203__;
  assign new_new_n9205__ = new_new_n9194__ & ~new_new_n9204__;
  assign new_new_n9206__ = new_new_n9192__ & ~new_new_n9205__;
  assign new_new_n9207__ = ~new_new_n9194__ & new_new_n9204__;
  assign new_new_n9208__ = ~new_new_n9206__ & ~new_new_n9207__;
  assign new_new_n9209__ = new_new_n8903__ & new_new_n9208__;
  assign new_new_n9210__ = ~new_new_n8903__ & ~new_new_n9208__;
  assign new_new_n9211__ = new_new_n8532__ & ~new_new_n8779__;
  assign new_new_n9212__ = ~new_new_n8532__ & new_new_n8779__;
  assign new_new_n9213__ = ~new_new_n9211__ & ~new_new_n9212__;
  assign new_new_n9214__ = new_new_n8785__ & new_new_n9213__;
  assign new_new_n9215__ = ~new_new_n8785__ & ~new_new_n9213__;
  assign new_new_n9216__ = ~new_new_n9214__ & ~new_new_n9215__;
  assign new_new_n9217__ = ~new_new_n9210__ & ~new_new_n9216__;
  assign new_new_n9218__ = ~new_new_n9209__ & ~new_new_n9217__;
  assign new_new_n9219__ = ~new_new_n8792__ & ~new_new_n8793__;
  assign new_new_n9220__ = new_new_n8803__ & new_new_n9219__;
  assign new_new_n9221__ = ~new_new_n8803__ & ~new_new_n9219__;
  assign new_new_n9222__ = ~new_new_n9220__ & ~new_new_n9221__;
  assign new_new_n9223__ = new_new_n9218__ & new_new_n9222__;
  assign new_new_n9224__ = ~new_new_n9218__ & ~new_new_n9222__;
  assign new_new_n9225__ = ~new_new_n9223__ & ~new_new_n9224__;
  assign new_new_n9226__ = new_new_n8893__ & ~new_new_n9225__;
  assign new_new_n9227__ = ~new_new_n8893__ & new_new_n9225__;
  assign new_new_n9228__ = ~new_new_n9226__ & ~new_new_n9227__;
  assign new_new_n9229__ = new_new_n8883__ & new_new_n9228__;
  assign new_new_n9230__ = ~new_new_n8883__ & ~new_new_n9228__;
  assign new_new_n9231__ = ~new_new_n9192__ & new_new_n9204__;
  assign new_new_n9232__ = new_new_n9192__ & ~new_new_n9204__;
  assign new_new_n9233__ = ~new_new_n9231__ & ~new_new_n9232__;
  assign new_new_n9234__ = ~new_new_n8222__ & new_new_n8775__;
  assign new_new_n9235__ = new_new_n8222__ & ~new_new_n8775__;
  assign new_new_n9236__ = ~new_new_n9234__ & ~new_new_n9235__;
  assign new_new_n9237__ = new_new_n9233__ & new_new_n9236__;
  assign new_new_n9238__ = ~new_new_n9233__ & ~new_new_n9236__;
  assign new_new_n9239__ = ~new_new_n9237__ & ~new_new_n9238__;
  assign new_new_n9240__ = new_new_n9188__ & ~new_new_n9190__;
  assign new_new_n9241__ = ~new_new_n9191__ & ~new_new_n9240__;
  assign new_new_n9242__ = ~new_new_n3535__ & ~new_new_n6625__;
  assign new_new_n9243__ = ~new_new_n1902__ & new_new_n6634__;
  assign new_new_n9244__ = ~new_new_n1823__ & new_new_n6629__;
  assign new_new_n9245__ = ~new_new_n9242__ & ~new_new_n9243__;
  assign new_new_n9246__ = ~new_new_n9244__ & new_new_n9245__;
  assign new_new_n9247__ = ~new_new_n6487__ & new_new_n6631__;
  assign new_new_n9248__ = ~pi20 & ~new_new_n9247__;
  assign new_new_n9249__ = ~new_new_n6487__ & new_new_n7015__;
  assign new_new_n9250__ = ~new_new_n9248__ & ~new_new_n9249__;
  assign new_new_n9251__ = new_new_n9246__ & ~new_new_n9250__;
  assign new_new_n9252__ = pi20 & ~new_new_n9246__;
  assign new_new_n9253__ = ~new_new_n9251__ & ~new_new_n9252__;
  assign new_new_n9254__ = new_new_n9241__ & ~new_new_n9253__;
  assign new_new_n9255__ = ~new_new_n9241__ & new_new_n9253__;
  assign new_new_n9256__ = ~new_new_n9157__ & ~new_new_n9158__;
  assign new_new_n9257__ = ~new_new_n9162__ & new_new_n9256__;
  assign new_new_n9258__ = new_new_n9162__ & ~new_new_n9256__;
  assign new_new_n9259__ = ~new_new_n9257__ & ~new_new_n9258__;
  assign new_new_n9260__ = ~new_new_n9143__ & ~new_new_n9144__;
  assign new_new_n9261__ = new_new_n9154__ & new_new_n9260__;
  assign new_new_n9262__ = ~new_new_n9154__ & ~new_new_n9260__;
  assign new_new_n9263__ = ~new_new_n9261__ & ~new_new_n9262__;
  assign new_new_n9264__ = ~new_new_n2572__ & new_new_n5191__;
  assign new_new_n9265__ = ~new_new_n2313__ & new_new_n5183__;
  assign new_new_n9266__ = ~new_new_n9264__ & ~new_new_n9265__;
  assign new_new_n9267__ = new_new_n2420__ & ~new_new_n6748__;
  assign new_new_n9268__ = new_new_n5195__ & ~new_new_n9267__;
  assign new_new_n9269__ = pi23 & ~new_new_n9268__;
  assign new_new_n9270__ = ~pi22 & new_new_n2420__;
  assign new_new_n9271__ = pi22 & ~new_new_n2420__;
  assign new_new_n9272__ = new_new_n5195__ & ~new_new_n9270__;
  assign new_new_n9273__ = ~new_new_n9271__ & new_new_n9272__;
  assign new_new_n9274__ = new_new_n6748__ & new_new_n9273__;
  assign new_new_n9275__ = ~new_new_n9269__ & ~new_new_n9274__;
  assign new_new_n9276__ = new_new_n9266__ & ~new_new_n9275__;
  assign new_new_n9277__ = new_new_n5195__ & new_new_n6749__;
  assign new_new_n9278__ = new_new_n9266__ & ~new_new_n9277__;
  assign new_new_n9279__ = ~pi23 & ~new_new_n9278__;
  assign new_new_n9280__ = ~new_new_n9276__ & ~new_new_n9279__;
  assign new_new_n9281__ = ~new_new_n9119__ & new_new_n9136__;
  assign new_new_n9282__ = new_new_n9119__ & ~new_new_n9136__;
  assign new_new_n9283__ = ~new_new_n9281__ & ~new_new_n9282__;
  assign new_new_n9284__ = new_new_n8594__ & ~new_new_n8714__;
  assign new_new_n9285__ = ~new_new_n8594__ & new_new_n8714__;
  assign new_new_n9286__ = ~new_new_n9284__ & ~new_new_n9285__;
  assign new_new_n9287__ = new_new_n9283__ & new_new_n9286__;
  assign new_new_n9288__ = ~new_new_n9283__ & ~new_new_n9286__;
  assign new_new_n9289__ = ~new_new_n9287__ & ~new_new_n9288__;
  assign new_new_n9290__ = new_new_n9280__ & ~new_new_n9289__;
  assign new_new_n9291__ = ~new_new_n9280__ & new_new_n9289__;
  assign new_new_n9292__ = ~new_new_n2572__ & new_new_n5213__;
  assign new_new_n9293__ = ~new_new_n2497__ & new_new_n5183__;
  assign new_new_n9294__ = new_new_n5215__ & new_new_n6804__;
  assign new_new_n9295__ = ~new_new_n9292__ & ~new_new_n9293__;
  assign new_new_n9296__ = ~new_new_n9294__ & new_new_n9295__;
  assign new_new_n9297__ = ~new_new_n2636__ & new_new_n5185__;
  assign new_new_n9298__ = pi23 & ~new_new_n9297__;
  assign new_new_n9299__ = ~new_new_n2636__ & new_new_n5188__;
  assign new_new_n9300__ = ~pi23 & ~new_new_n9299__;
  assign new_new_n9301__ = pi20 & ~new_new_n9300__;
  assign new_new_n9302__ = ~new_new_n9298__ & ~new_new_n9301__;
  assign new_new_n9303__ = new_new_n9296__ & ~new_new_n9302__;
  assign new_new_n9304__ = ~pi23 & ~new_new_n9296__;
  assign new_new_n9305__ = ~new_new_n9303__ & ~new_new_n9304__;
  assign new_new_n9306__ = ~new_new_n9098__ & ~new_new_n9099__;
  assign new_new_n9307__ = ~new_new_n9109__ & new_new_n9306__;
  assign new_new_n9308__ = new_new_n9109__ & ~new_new_n9306__;
  assign new_new_n9309__ = ~new_new_n9307__ & ~new_new_n9308__;
  assign new_new_n9310__ = ~new_new_n9305__ & new_new_n9309__;
  assign new_new_n9311__ = new_new_n9305__ & ~new_new_n9309__;
  assign new_new_n9312__ = ~new_new_n9090__ & ~new_new_n9091__;
  assign new_new_n9313__ = ~new_new_n9095__ & new_new_n9312__;
  assign new_new_n9314__ = new_new_n9095__ & ~new_new_n9312__;
  assign new_new_n9315__ = ~new_new_n9313__ & ~new_new_n9314__;
  assign new_new_n9316__ = ~new_new_n9057__ & ~new_new_n9058__;
  assign new_new_n9317__ = ~new_new_n9070__ & new_new_n9316__;
  assign new_new_n9318__ = new_new_n9070__ & ~new_new_n9316__;
  assign new_new_n9319__ = ~new_new_n9317__ & ~new_new_n9318__;
  assign new_new_n9320__ = ~new_new_n8620__ & new_new_n9042__;
  assign new_new_n9321__ = new_new_n9052__ & ~new_new_n9320__;
  assign new_new_n9322__ = new_new_n8620__ & ~new_new_n8983__;
  assign new_new_n9323__ = ~new_new_n9042__ & new_new_n9322__;
  assign new_new_n9324__ = ~new_new_n9321__ & ~new_new_n9323__;
  assign new_new_n9325__ = new_new_n8626__ & ~new_new_n9324__;
  assign new_new_n9326__ = ~new_new_n8983__ & new_new_n9042__;
  assign new_new_n9327__ = ~new_new_n9048__ & ~new_new_n9326__;
  assign new_new_n9328__ = ~new_new_n9052__ & ~new_new_n9327__;
  assign new_new_n9329__ = ~pi29 & ~new_new_n9042__;
  assign new_new_n9330__ = ~new_new_n9048__ & ~new_new_n9329__;
  assign new_new_n9331__ = new_new_n8983__ & ~new_new_n9330__;
  assign new_new_n9332__ = ~new_new_n9328__ & ~new_new_n9331__;
  assign new_new_n9333__ = ~new_new_n9325__ & ~new_new_n9332__;
  assign new_new_n9334__ = ~new_new_n8996__ & ~new_new_n9003__;
  assign new_new_n9335__ = new_new_n8996__ & new_new_n9003__;
  assign new_new_n9336__ = ~new_new_n9334__ & ~new_new_n9335__;
  assign new_new_n9337__ = new_new_n9016__ & ~new_new_n9336__;
  assign new_new_n9338__ = new_new_n9035__ & new_new_n9334__;
  assign new_new_n9339__ = ~new_new_n9337__ & ~new_new_n9338__;
  assign new_new_n9340__ = new_new_n9015__ & ~new_new_n9339__;
  assign new_new_n9341__ = ~new_new_n9037__ & new_new_n9336__;
  assign new_new_n9342__ = ~new_new_n9340__ & ~new_new_n9341__;
  assign new_new_n9343__ = ~new_new_n2960__ & new_new_n5183__;
  assign new_new_n9344__ = ~new_new_n3460__ & new_new_n5213__;
  assign new_new_n9345__ = ~new_new_n5212__ & ~new_new_n7388__;
  assign new_new_n9346__ = new_new_n5195__ & ~new_new_n9345__;
  assign new_new_n9347__ = new_new_n7391__ & new_new_n9346__;
  assign new_new_n9348__ = ~new_new_n9343__ & ~new_new_n9344__;
  assign new_new_n9349__ = ~new_new_n9347__ & new_new_n9348__;
  assign new_new_n9350__ = ~pi23 & ~new_new_n9349__;
  assign new_new_n9351__ = ~new_new_n3126__ & new_new_n5186__;
  assign new_new_n9352__ = pi23 & ~new_new_n9351__;
  assign new_new_n9353__ = ~new_new_n3126__ & new_new_n5189__;
  assign new_new_n9354__ = ~new_new_n9352__ & ~new_new_n9353__;
  assign new_new_n9355__ = new_new_n9349__ & ~new_new_n9354__;
  assign new_new_n9356__ = ~new_new_n9350__ & ~new_new_n9355__;
  assign new_new_n9357__ = pi26 & ~new_new_n349__;
  assign new_new_n9358__ = ~new_new_n146__ & new_new_n9357__;
  assign new_new_n9359__ = ~new_new_n9017__ & new_new_n9358__;
  assign new_new_n9360__ = new_new_n9033__ & ~new_new_n9359__;
  assign new_new_n9361__ = pi26 & ~new_new_n9020__;
  assign new_new_n9362__ = ~new_new_n9033__ & new_new_n9361__;
  assign new_new_n9363__ = ~new_new_n9360__ & ~new_new_n9362__;
  assign new_new_n9364__ = ~new_new_n104__ & ~new_new_n3055__;
  assign new_new_n9365__ = ~new_new_n3356__ & new_new_n9364__;
  assign new_new_n9366__ = ~new_new_n99__ & ~new_new_n9365__;
  assign new_new_n9367__ = pi25 & ~new_new_n9366__;
  assign new_new_n9368__ = ~new_new_n389__ & ~new_new_n3356__;
  assign new_new_n9369__ = new_new_n801__ & ~new_new_n3055__;
  assign new_new_n9370__ = ~new_new_n9368__ & ~new_new_n9369__;
  assign new_new_n9371__ = ~new_new_n9367__ & ~new_new_n9370__;
  assign new_new_n9372__ = pi22 & new_new_n5179__;
  assign new_new_n9373__ = ~pi22 & new_new_n5181__;
  assign new_new_n9374__ = ~new_new_n9372__ & ~new_new_n9373__;
  assign new_new_n9375__ = new_new_n5215__ & new_new_n7682__;
  assign new_new_n9376__ = new_new_n9374__ & ~new_new_n9375__;
  assign new_new_n9377__ = ~new_new_n3055__ & ~new_new_n9376__;
  assign new_new_n9378__ = ~new_new_n3254__ & new_new_n5195__;
  assign new_new_n9379__ = ~new_new_n3356__ & new_new_n5191__;
  assign new_new_n9380__ = ~new_new_n9378__ & ~new_new_n9379__;
  assign new_new_n9381__ = ~new_new_n3055__ & new_new_n5212__;
  assign new_new_n9382__ = new_new_n3356__ & new_new_n9381__;
  assign new_new_n9383__ = ~new_new_n9380__ & ~new_new_n9382__;
  assign new_new_n9384__ = ~new_new_n9377__ & ~new_new_n9383__;
  assign new_new_n9385__ = ~pi22 & ~new_new_n3356__;
  assign new_new_n9386__ = new_new_n5181__ & ~new_new_n9385__;
  assign new_new_n9387__ = ~new_new_n3055__ & ~new_new_n5179__;
  assign new_new_n9388__ = new_new_n3356__ & ~new_new_n9387__;
  assign new_new_n9389__ = ~new_new_n5186__ & ~new_new_n9386__;
  assign new_new_n9390__ = ~new_new_n9388__ & new_new_n9389__;
  assign new_new_n9391__ = pi23 & ~new_new_n9390__;
  assign new_new_n9392__ = new_new_n9384__ & new_new_n9391__;
  assign new_new_n9393__ = ~new_new_n110__ & ~new_new_n3356__;
  assign new_new_n9394__ = ~new_new_n9392__ & ~new_new_n9393__;
  assign new_new_n9395__ = ~new_new_n3164__ & new_new_n5213__;
  assign new_new_n9396__ = ~new_new_n3055__ & new_new_n5191__;
  assign new_new_n9397__ = ~new_new_n3254__ & new_new_n5183__;
  assign new_new_n9398__ = ~new_new_n9395__ & ~new_new_n9396__;
  assign new_new_n9399__ = ~new_new_n9397__ & new_new_n9398__;
  assign new_new_n9400__ = new_new_n5195__ & ~new_new_n8637__;
  assign new_new_n9401__ = ~pi23 & ~new_new_n9400__;
  assign new_new_n9402__ = new_new_n5974__ & ~new_new_n8637__;
  assign new_new_n9403__ = ~new_new_n9401__ & ~new_new_n9402__;
  assign new_new_n9404__ = new_new_n9399__ & ~new_new_n9403__;
  assign new_new_n9405__ = pi23 & ~new_new_n9399__;
  assign new_new_n9406__ = ~new_new_n9404__ & ~new_new_n9405__;
  assign new_new_n9407__ = ~new_new_n9394__ & new_new_n9406__;
  assign new_new_n9408__ = ~new_new_n9371__ & ~new_new_n9407__;
  assign new_new_n9409__ = new_new_n9371__ & new_new_n9407__;
  assign new_new_n9410__ = ~new_new_n3254__ & new_new_n5191__;
  assign new_new_n9411__ = ~new_new_n3126__ & new_new_n5213__;
  assign new_new_n9412__ = ~new_new_n3164__ & new_new_n5183__;
  assign new_new_n9413__ = new_new_n5215__ & ~new_new_n7570__;
  assign new_new_n9414__ = ~new_new_n9410__ & ~new_new_n9411__;
  assign new_new_n9415__ = ~new_new_n9412__ & new_new_n9414__;
  assign new_new_n9416__ = ~new_new_n9413__ & new_new_n9415__;
  assign new_new_n9417__ = pi23 & ~new_new_n9416__;
  assign new_new_n9418__ = ~pi23 & new_new_n9416__;
  assign new_new_n9419__ = ~new_new_n9417__ & ~new_new_n9418__;
  assign new_new_n9420__ = ~new_new_n9409__ & ~new_new_n9419__;
  assign new_new_n9421__ = ~new_new_n9408__ & ~new_new_n9420__;
  assign new_new_n9422__ = ~new_new_n9363__ & ~new_new_n9421__;
  assign new_new_n9423__ = new_new_n9363__ & new_new_n9421__;
  assign new_new_n9424__ = ~new_new_n2960__ & new_new_n5213__;
  assign new_new_n9425__ = ~new_new_n3126__ & new_new_n5183__;
  assign new_new_n9426__ = ~new_new_n3164__ & new_new_n5191__;
  assign new_new_n9427__ = new_new_n5215__ & ~new_new_n7468__;
  assign new_new_n9428__ = ~new_new_n9425__ & ~new_new_n9426__;
  assign new_new_n9429__ = ~new_new_n9424__ & new_new_n9428__;
  assign new_new_n9430__ = ~new_new_n9427__ & new_new_n9429__;
  assign new_new_n9431__ = ~pi23 & ~new_new_n9430__;
  assign new_new_n9432__ = pi23 & new_new_n9430__;
  assign new_new_n9433__ = ~new_new_n9431__ & ~new_new_n9432__;
  assign new_new_n9434__ = ~new_new_n9423__ & new_new_n9433__;
  assign new_new_n9435__ = ~new_new_n9422__ & ~new_new_n9434__;
  assign new_new_n9436__ = ~new_new_n9035__ & ~new_new_n9435__;
  assign new_new_n9437__ = ~new_new_n9356__ & ~new_new_n9436__;
  assign new_new_n9438__ = new_new_n9015__ & ~new_new_n9016__;
  assign new_new_n9439__ = ~new_new_n9015__ & new_new_n9016__;
  assign new_new_n9440__ = ~new_new_n9438__ & ~new_new_n9439__;
  assign new_new_n9441__ = ~new_new_n9437__ & new_new_n9440__;
  assign new_new_n9442__ = new_new_n9035__ & new_new_n9438__;
  assign new_new_n9443__ = ~new_new_n9356__ & ~new_new_n9442__;
  assign new_new_n9444__ = ~new_new_n9435__ & ~new_new_n9443__;
  assign new_new_n9445__ = ~new_new_n9441__ & ~new_new_n9444__;
  assign new_new_n9446__ = new_new_n9342__ & new_new_n9445__;
  assign new_new_n9447__ = ~new_new_n9342__ & ~new_new_n9445__;
  assign new_new_n9448__ = new_new_n5215__ & ~new_new_n7065__;
  assign new_new_n9449__ = ~new_new_n2960__ & new_new_n5191__;
  assign new_new_n9450__ = ~new_new_n3460__ & new_new_n5183__;
  assign new_new_n9451__ = ~new_new_n9449__ & ~new_new_n9450__;
  assign new_new_n9452__ = ~new_new_n9448__ & new_new_n9451__;
  assign new_new_n9453__ = ~new_new_n2848__ & new_new_n5213__;
  assign new_new_n9454__ = new_new_n9452__ & ~new_new_n9453__;
  assign new_new_n9455__ = ~pi23 & ~new_new_n9454__;
  assign new_new_n9456__ = pi23 & new_new_n9454__;
  assign new_new_n9457__ = ~new_new_n9455__ & ~new_new_n9456__;
  assign new_new_n9458__ = ~new_new_n9447__ & ~new_new_n9457__;
  assign new_new_n9459__ = ~new_new_n9446__ & ~new_new_n9458__;
  assign new_new_n9460__ = new_new_n9333__ & new_new_n9459__;
  assign new_new_n9461__ = ~new_new_n9333__ & ~new_new_n9459__;
  assign new_new_n9462__ = ~new_new_n3460__ & new_new_n5191__;
  assign new_new_n9463__ = ~new_new_n2886__ & new_new_n5213__;
  assign new_new_n9464__ = ~new_new_n2848__ & new_new_n5183__;
  assign new_new_n9465__ = new_new_n5215__ & ~new_new_n8574__;
  assign new_new_n9466__ = ~new_new_n9462__ & ~new_new_n9463__;
  assign new_new_n9467__ = ~new_new_n9464__ & new_new_n9466__;
  assign new_new_n9468__ = ~new_new_n9465__ & new_new_n9467__;
  assign new_new_n9469__ = pi23 & ~new_new_n9468__;
  assign new_new_n9470__ = ~pi23 & new_new_n9468__;
  assign new_new_n9471__ = ~new_new_n9469__ & ~new_new_n9470__;
  assign new_new_n9472__ = ~new_new_n9461__ & ~new_new_n9471__;
  assign new_new_n9473__ = ~new_new_n9460__ & ~new_new_n9472__;
  assign new_new_n9474__ = new_new_n9319__ & ~new_new_n9473__;
  assign new_new_n9475__ = ~new_new_n9319__ & new_new_n9473__;
  assign new_new_n9476__ = new_new_n5215__ & ~new_new_n7378__;
  assign new_new_n9477__ = ~new_new_n2737__ & new_new_n5213__;
  assign new_new_n9478__ = ~new_new_n2886__ & new_new_n5183__;
  assign new_new_n9479__ = ~new_new_n9477__ & ~new_new_n9478__;
  assign new_new_n9480__ = ~new_new_n9476__ & new_new_n9479__;
  assign new_new_n9481__ = ~pi23 & ~new_new_n9480__;
  assign new_new_n9482__ = ~new_new_n2848__ & new_new_n5186__;
  assign new_new_n9483__ = pi23 & ~new_new_n9482__;
  assign new_new_n9484__ = ~new_new_n2848__ & new_new_n5189__;
  assign new_new_n9485__ = ~new_new_n9483__ & ~new_new_n9484__;
  assign new_new_n9486__ = new_new_n9480__ & ~new_new_n9485__;
  assign new_new_n9487__ = ~new_new_n9481__ & ~new_new_n9486__;
  assign new_new_n9488__ = ~new_new_n9475__ & new_new_n9487__;
  assign new_new_n9489__ = ~new_new_n9474__ & ~new_new_n9488__;
  assign new_new_n9490__ = ~new_new_n9075__ & ~new_new_n9087__;
  assign new_new_n9491__ = ~new_new_n9088__ & ~new_new_n9490__;
  assign new_new_n9492__ = ~new_new_n2737__ & new_new_n5183__;
  assign new_new_n9493__ = ~new_new_n2886__ & new_new_n5191__;
  assign new_new_n9494__ = ~new_new_n2636__ & new_new_n5213__;
  assign new_new_n9495__ = ~new_new_n9492__ & ~new_new_n9493__;
  assign new_new_n9496__ = ~new_new_n9494__ & new_new_n9495__;
  assign new_new_n9497__ = pi23 & ~new_new_n9496__;
  assign new_new_n9498__ = pi23 & new_new_n5974__;
  assign new_new_n9499__ = ~new_new_n2636__ & ~new_new_n9498__;
  assign new_new_n9500__ = ~pi23 & new_new_n9496__;
  assign new_new_n9501__ = new_new_n2636__ & ~new_new_n9500__;
  assign new_new_n9502__ = ~new_new_n9499__ & ~new_new_n9501__;
  assign new_new_n9503__ = ~new_new_n7811__ & new_new_n9502__;
  assign new_new_n9504__ = ~new_new_n7878__ & new_new_n9500__;
  assign new_new_n9505__ = new_new_n2636__ & ~new_new_n9498__;
  assign new_new_n9506__ = ~new_new_n2636__ & ~new_new_n9500__;
  assign new_new_n9507__ = ~new_new_n9505__ & ~new_new_n9506__;
  assign new_new_n9508__ = new_new_n7811__ & new_new_n9507__;
  assign new_new_n9509__ = ~new_new_n9497__ & ~new_new_n9504__;
  assign new_new_n9510__ = ~new_new_n9503__ & new_new_n9509__;
  assign new_new_n9511__ = ~new_new_n9508__ & new_new_n9510__;
  assign new_new_n9512__ = new_new_n9491__ & new_new_n9511__;
  assign new_new_n9513__ = ~new_new_n9489__ & ~new_new_n9512__;
  assign new_new_n9514__ = ~new_new_n9491__ & ~new_new_n9511__;
  assign new_new_n9515__ = ~new_new_n9513__ & ~new_new_n9514__;
  assign new_new_n9516__ = ~new_new_n9315__ & ~new_new_n9515__;
  assign new_new_n9517__ = new_new_n9315__ & new_new_n9515__;
  assign new_new_n9518__ = ~new_new_n2636__ & new_new_n5183__;
  assign new_new_n9519__ = ~new_new_n2737__ & new_new_n5191__;
  assign new_new_n9520__ = ~new_new_n9518__ & ~new_new_n9519__;
  assign new_new_n9521__ = new_new_n5195__ & ~new_new_n9126__;
  assign new_new_n9522__ = pi23 & ~new_new_n9521__;
  assign new_new_n9523__ = ~pi22 & new_new_n2497__;
  assign new_new_n9524__ = pi22 & ~new_new_n2497__;
  assign new_new_n9525__ = new_new_n5195__ & ~new_new_n9523__;
  assign new_new_n9526__ = ~new_new_n9524__ & new_new_n9525__;
  assign new_new_n9527__ = ~new_new_n6797__ & new_new_n9526__;
  assign new_new_n9528__ = ~new_new_n9522__ & ~new_new_n9527__;
  assign new_new_n9529__ = new_new_n9520__ & ~new_new_n9528__;
  assign new_new_n9530__ = new_new_n5195__ & new_new_n7772__;
  assign new_new_n9531__ = new_new_n9520__ & ~new_new_n9530__;
  assign new_new_n9532__ = ~pi23 & ~new_new_n9531__;
  assign new_new_n9533__ = ~new_new_n9529__ & ~new_new_n9532__;
  assign new_new_n9534__ = ~new_new_n9517__ & new_new_n9533__;
  assign new_new_n9535__ = ~new_new_n9516__ & ~new_new_n9534__;
  assign new_new_n9536__ = ~new_new_n9311__ & new_new_n9535__;
  assign new_new_n9537__ = ~new_new_n9310__ & ~new_new_n9536__;
  assign new_new_n9538__ = ~new_new_n9112__ & ~new_new_n9113__;
  assign new_new_n9539__ = ~new_new_n9117__ & new_new_n9538__;
  assign new_new_n9540__ = new_new_n9117__ & ~new_new_n9538__;
  assign new_new_n9541__ = ~new_new_n9539__ & ~new_new_n9540__;
  assign new_new_n9542__ = new_new_n9537__ & ~new_new_n9541__;
  assign new_new_n9543__ = ~new_new_n9537__ & new_new_n9541__;
  assign new_new_n9544__ = new_new_n5215__ & ~new_new_n7236__;
  assign new_new_n9545__ = ~new_new_n2497__ & new_new_n5191__;
  assign new_new_n9546__ = ~new_new_n2572__ & new_new_n5183__;
  assign new_new_n9547__ = ~new_new_n2313__ & new_new_n5213__;
  assign new_new_n9548__ = ~new_new_n9545__ & ~new_new_n9546__;
  assign new_new_n9549__ = ~new_new_n9547__ & new_new_n9548__;
  assign new_new_n9550__ = ~new_new_n9544__ & new_new_n9549__;
  assign new_new_n9551__ = pi23 & new_new_n9550__;
  assign new_new_n9552__ = ~pi23 & ~new_new_n9550__;
  assign new_new_n9553__ = ~new_new_n9551__ & ~new_new_n9552__;
  assign new_new_n9554__ = ~new_new_n9543__ & new_new_n9553__;
  assign new_new_n9555__ = ~new_new_n9542__ & ~new_new_n9554__;
  assign new_new_n9556__ = ~new_new_n9291__ & ~new_new_n9555__;
  assign new_new_n9557__ = ~new_new_n9290__ & ~new_new_n9556__;
  assign new_new_n9558__ = ~new_new_n9263__ & ~new_new_n9557__;
  assign new_new_n9559__ = new_new_n9263__ & new_new_n9557__;
  assign new_new_n9560__ = ~new_new_n2420__ & new_new_n5183__;
  assign new_new_n9561__ = ~new_new_n2224__ & new_new_n5213__;
  assign new_new_n9562__ = ~new_new_n2313__ & new_new_n5191__;
  assign new_new_n9563__ = ~new_new_n9560__ & ~new_new_n9561__;
  assign new_new_n9564__ = ~new_new_n9562__ & new_new_n9563__;
  assign new_new_n9565__ = new_new_n5195__ & new_new_n6521__;
  assign new_new_n9566__ = ~pi23 & ~new_new_n9565__;
  assign new_new_n9567__ = new_new_n5974__ & new_new_n6521__;
  assign new_new_n9568__ = ~new_new_n9566__ & ~new_new_n9567__;
  assign new_new_n9569__ = new_new_n9564__ & ~new_new_n9568__;
  assign new_new_n9570__ = pi23 & ~new_new_n9564__;
  assign new_new_n9571__ = ~new_new_n9569__ & ~new_new_n9570__;
  assign new_new_n9572__ = ~new_new_n9559__ & ~new_new_n9571__;
  assign new_new_n9573__ = ~new_new_n9558__ & ~new_new_n9572__;
  assign new_new_n9574__ = new_new_n9259__ & ~new_new_n9573__;
  assign new_new_n9575__ = ~new_new_n9259__ & new_new_n9573__;
  assign new_new_n9576__ = ~new_new_n2224__ & new_new_n5183__;
  assign new_new_n9577__ = ~new_new_n2024__ & new_new_n5213__;
  assign new_new_n9578__ = ~new_new_n2420__ & new_new_n5191__;
  assign new_new_n9579__ = new_new_n5215__ & new_new_n7313__;
  assign new_new_n9580__ = ~new_new_n9576__ & ~new_new_n9577__;
  assign new_new_n9581__ = ~new_new_n9578__ & new_new_n9580__;
  assign new_new_n9582__ = ~new_new_n9579__ & new_new_n9581__;
  assign new_new_n9583__ = ~pi23 & ~new_new_n9582__;
  assign new_new_n9584__ = pi23 & new_new_n9582__;
  assign new_new_n9585__ = ~new_new_n9583__ & ~new_new_n9584__;
  assign new_new_n9586__ = ~new_new_n9575__ & new_new_n9585__;
  assign new_new_n9587__ = ~new_new_n9574__ & ~new_new_n9586__;
  assign new_new_n9588__ = ~new_new_n9255__ & ~new_new_n9587__;
  assign new_new_n9589__ = ~new_new_n9254__ & ~new_new_n9588__;
  assign new_new_n9590__ = new_new_n9239__ & ~new_new_n9589__;
  assign new_new_n9591__ = ~new_new_n9239__ & new_new_n9589__;
  assign new_new_n9592__ = ~new_new_n5671__ & new_new_n6959__;
  assign new_new_n9593__ = ~new_new_n1737__ & new_new_n6964__;
  assign new_new_n9594__ = ~new_new_n1466__ & new_new_n6968__;
  assign new_new_n9595__ = ~new_new_n9593__ & ~new_new_n9594__;
  assign new_new_n9596__ = ~new_new_n9592__ & new_new_n9595__;
  assign new_new_n9597__ = ~new_new_n1556__ & new_new_n6958__;
  assign new_new_n9598__ = pi17 & ~new_new_n9597__;
  assign new_new_n9599__ = ~new_new_n1556__ & new_new_n8160__;
  assign new_new_n9600__ = ~new_new_n9598__ & ~new_new_n9599__;
  assign new_new_n9601__ = new_new_n9596__ & ~new_new_n9600__;
  assign new_new_n9602__ = ~pi17 & ~new_new_n9596__;
  assign new_new_n9603__ = ~new_new_n9601__ & ~new_new_n9602__;
  assign new_new_n9604__ = ~new_new_n9591__ & new_new_n9603__;
  assign new_new_n9605__ = ~new_new_n9590__ & ~new_new_n9604__;
  assign new_new_n9606__ = ~new_new_n9209__ & ~new_new_n9210__;
  assign new_new_n9607__ = ~new_new_n9216__ & new_new_n9606__;
  assign new_new_n9608__ = new_new_n9216__ & ~new_new_n9606__;
  assign new_new_n9609__ = ~new_new_n9607__ & ~new_new_n9608__;
  assign new_new_n9610__ = new_new_n9605__ & ~new_new_n9609__;
  assign new_new_n9611__ = ~new_new_n9605__ & new_new_n9609__;
  assign new_new_n9612__ = ~new_new_n3618__ & new_new_n6991__;
  assign new_new_n9613__ = ~new_new_n1061__ & new_new_n6985__;
  assign new_new_n9614__ = ~new_new_n9612__ & ~new_new_n9613__;
  assign new_new_n9615__ = ~new_new_n1207__ & new_new_n6994__;
  assign new_new_n9616__ = ~new_new_n5235__ & new_new_n9615__;
  assign new_new_n9617__ = new_new_n9614__ & ~new_new_n9616__;
  assign new_new_n9618__ = pi14 & ~new_new_n9617__;
  assign new_new_n9619__ = ~pi13 & ~new_new_n1207__;
  assign new_new_n9620__ = new_new_n1207__ & new_new_n5235__;
  assign new_new_n9621__ = new_new_n6994__ & ~new_new_n9620__;
  assign new_new_n9622__ = pi13 & ~new_new_n5235__;
  assign new_new_n9623__ = ~new_new_n9619__ & ~new_new_n9622__;
  assign new_new_n9624__ = new_new_n9621__ & new_new_n9623__;
  assign new_new_n9625__ = ~pi14 & new_new_n9614__;
  assign new_new_n9626__ = ~new_new_n9621__ & new_new_n9625__;
  assign new_new_n9627__ = ~new_new_n9618__ & ~new_new_n9624__;
  assign new_new_n9628__ = ~new_new_n9626__ & new_new_n9627__;
  assign new_new_n9629__ = ~new_new_n9611__ & new_new_n9628__;
  assign new_new_n9630__ = ~new_new_n9610__ & ~new_new_n9629__;
  assign new_new_n9631__ = ~new_new_n9230__ & ~new_new_n9630__;
  assign new_new_n9632__ = ~new_new_n9229__ & ~new_new_n9631__;
  assign new_new_n9633__ = ~new_new_n8866__ & ~new_new_n9632__;
  assign new_new_n9634__ = new_new_n8866__ & new_new_n9632__;
  assign new_new_n9635__ = ~pi13 & new_new_n3720__;
  assign new_new_n9636__ = pi13 & ~new_new_n3720__;
  assign new_new_n9637__ = new_new_n6994__ & ~new_new_n9635__;
  assign new_new_n9638__ = ~new_new_n9636__ & new_new_n9637__;
  assign new_new_n9639__ = ~new_new_n4032__ & new_new_n9638__;
  assign new_new_n9640__ = ~new_new_n868__ & new_new_n6985__;
  assign new_new_n9641__ = ~new_new_n1207__ & new_new_n6991__;
  assign new_new_n9642__ = ~new_new_n9640__ & ~new_new_n9641__;
  assign new_new_n9643__ = ~new_new_n3720__ & new_new_n6994__;
  assign new_new_n9644__ = new_new_n4032__ & new_new_n9643__;
  assign new_new_n9645__ = new_new_n9642__ & ~new_new_n9644__;
  assign new_new_n9646__ = ~pi14 & ~new_new_n9645__;
  assign new_new_n9647__ = new_new_n3720__ & new_new_n4032__;
  assign new_new_n9648__ = new_new_n6994__ & ~new_new_n9647__;
  assign new_new_n9649__ = pi14 & new_new_n9642__;
  assign new_new_n9650__ = ~new_new_n9648__ & new_new_n9649__;
  assign new_new_n9651__ = ~new_new_n9639__ & ~new_new_n9646__;
  assign new_new_n9652__ = ~new_new_n9650__ & new_new_n9651__;
  assign new_new_n9653__ = new_new_n8893__ & ~new_new_n9223__;
  assign new_new_n9654__ = ~new_new_n9224__ & ~new_new_n9653__;
  assign new_new_n9655__ = ~new_new_n8806__ & ~new_new_n8807__;
  assign new_new_n9656__ = new_new_n8811__ & new_new_n9655__;
  assign new_new_n9657__ = ~new_new_n8811__ & ~new_new_n9655__;
  assign new_new_n9658__ = ~new_new_n9656__ & ~new_new_n9657__;
  assign new_new_n9659__ = new_new_n9654__ & ~new_new_n9658__;
  assign new_new_n9660__ = ~new_new_n9654__ & new_new_n9658__;
  assign new_new_n9661__ = ~new_new_n9659__ & ~new_new_n9660__;
  assign new_new_n9662__ = new_new_n9652__ & new_new_n9661__;
  assign new_new_n9663__ = ~new_new_n9652__ & ~new_new_n9661__;
  assign new_new_n9664__ = ~new_new_n9662__ & ~new_new_n9663__;
  assign new_new_n9665__ = ~new_new_n9634__ & ~new_new_n9664__;
  assign new_new_n9666__ = ~new_new_n9633__ & ~new_new_n9665__;
  assign new_new_n9667__ = ~new_new_n583__ & new_new_n8474__;
  assign new_new_n9668__ = ~new_new_n691__ & ~new_new_n8479__;
  assign new_new_n9669__ = new_new_n3768__ & new_new_n8468__;
  assign new_new_n9670__ = new_new_n4144__ & ~new_new_n8468__;
  assign new_new_n9671__ = new_new_n8469__ & ~new_new_n9669__;
  assign new_new_n9672__ = ~new_new_n9670__ & new_new_n9671__;
  assign new_new_n9673__ = ~new_new_n9668__ & ~new_new_n9672__;
  assign new_new_n9674__ = ~new_new_n9667__ & new_new_n9673__;
  assign new_new_n9675__ = pi11 & ~new_new_n9674__;
  assign new_new_n9676__ = new_new_n583__ & new_new_n8479__;
  assign new_new_n9677__ = new_new_n8474__ & ~new_new_n9676__;
  assign new_new_n9678__ = ~pi11 & ~new_new_n9677__;
  assign new_new_n9679__ = new_new_n9673__ & new_new_n9678__;
  assign new_new_n9680__ = ~new_new_n9675__ & ~new_new_n9679__;
  assign new_new_n9681__ = ~new_new_n8818__ & ~new_new_n8819__;
  assign new_new_n9682__ = new_new_n8834__ & ~new_new_n9681__;
  assign new_new_n9683__ = ~new_new_n8834__ & new_new_n9681__;
  assign new_new_n9684__ = ~new_new_n9682__ & ~new_new_n9683__;
  assign new_new_n9685__ = new_new_n9680__ & new_new_n9684__;
  assign new_new_n9686__ = ~new_new_n9680__ & ~new_new_n9684__;
  assign new_new_n9687__ = ~new_new_n9685__ & ~new_new_n9686__;
  assign new_new_n9688__ = ~new_new_n9652__ & ~new_new_n9660__;
  assign new_new_n9689__ = ~new_new_n9659__ & ~new_new_n9688__;
  assign new_new_n9690__ = new_new_n9687__ & new_new_n9689__;
  assign new_new_n9691__ = ~new_new_n9687__ & ~new_new_n9689__;
  assign new_new_n9692__ = ~new_new_n9690__ & ~new_new_n9691__;
  assign new_new_n9693__ = new_new_n9666__ & new_new_n9692__;
  assign new_new_n9694__ = ~pi07 & ~new_new_n466__;
  assign new_new_n9695__ = pi08 & ~new_new_n9694__;
  assign new_new_n9696__ = ~pi07 & ~pi08;
  assign new_new_n9697__ = ~pi05 & ~pi06;
  assign new_new_n9698__ = ~new_new_n9696__ & ~new_new_n9697__;
  assign new_new_n9699__ = ~new_new_n466__ & new_new_n9698__;
  assign new_new_n9700__ = ~new_new_n9695__ & ~new_new_n9699__;
  assign new_new_n9701__ = pi05 & pi06;
  assign new_new_n9702__ = ~new_new_n4168__ & ~new_new_n9694__;
  assign new_new_n9703__ = pi08 & new_new_n4168__;
  assign new_new_n9704__ = ~new_new_n9701__ & ~new_new_n9702__;
  assign new_new_n9705__ = ~new_new_n9703__ & new_new_n9704__;
  assign new_new_n9706__ = ~new_new_n9700__ & ~new_new_n9705__;
  assign new_new_n9707__ = ~new_new_n9666__ & ~new_new_n9692__;
  assign new_new_n9708__ = ~new_new_n9706__ & ~new_new_n9707__;
  assign new_new_n9709__ = ~new_new_n9693__ & ~new_new_n9708__;
  assign new_new_n9710__ = ~new_new_n3720__ & new_new_n8474__;
  assign new_new_n9711__ = ~new_new_n868__ & ~new_new_n8479__;
  assign new_new_n9712__ = ~new_new_n9710__ & ~new_new_n9711__;
  assign new_new_n9713__ = ~new_new_n5129__ & new_new_n8469__;
  assign new_new_n9714__ = pi11 & ~new_new_n9713__;
  assign new_new_n9715__ = pi10 & new_new_n910__;
  assign new_new_n9716__ = ~new_new_n8851__ & ~new_new_n9715__;
  assign new_new_n9717__ = new_new_n8469__ & ~new_new_n9716__;
  assign new_new_n9718__ = new_new_n4036__ & new_new_n9717__;
  assign new_new_n9719__ = ~new_new_n9714__ & ~new_new_n9718__;
  assign new_new_n9720__ = new_new_n9712__ & ~new_new_n9719__;
  assign new_new_n9721__ = new_new_n5116__ & new_new_n8469__;
  assign new_new_n9722__ = new_new_n9712__ & ~new_new_n9721__;
  assign new_new_n9723__ = ~pi11 & ~new_new_n9722__;
  assign new_new_n9724__ = ~new_new_n9720__ & ~new_new_n9723__;
  assign new_new_n9725__ = ~new_new_n3618__ & new_new_n6985__;
  assign new_new_n9726__ = ~new_new_n1325__ & new_new_n6991__;
  assign new_new_n9727__ = ~new_new_n9725__ & ~new_new_n9726__;
  assign new_new_n9728__ = ~new_new_n1061__ & new_new_n6994__;
  assign new_new_n9729__ = new_new_n4926__ & new_new_n9728__;
  assign new_new_n9730__ = new_new_n9727__ & ~new_new_n9729__;
  assign new_new_n9731__ = pi14 & ~new_new_n9730__;
  assign new_new_n9732__ = pi13 & new_new_n4926__;
  assign new_new_n9733__ = ~new_new_n4927__ & new_new_n6994__;
  assign new_new_n9734__ = ~pi13 & ~new_new_n1061__;
  assign new_new_n9735__ = ~new_new_n9732__ & ~new_new_n9734__;
  assign new_new_n9736__ = new_new_n9733__ & new_new_n9735__;
  assign new_new_n9737__ = ~pi14 & new_new_n9727__;
  assign new_new_n9738__ = ~new_new_n9733__ & new_new_n9737__;
  assign new_new_n9739__ = ~new_new_n9731__ & ~new_new_n9736__;
  assign new_new_n9740__ = ~new_new_n9738__ & new_new_n9739__;
  assign new_new_n9741__ = ~new_new_n1466__ & new_new_n7935__;
  assign new_new_n9742__ = ~new_new_n1660__ & new_new_n6964__;
  assign new_new_n9743__ = ~new_new_n1737__ & new_new_n6968__;
  assign new_new_n9744__ = ~new_new_n9741__ & ~new_new_n9742__;
  assign new_new_n9745__ = ~new_new_n9743__ & new_new_n9744__;
  assign new_new_n9746__ = ~new_new_n6410__ & new_new_n6958__;
  assign new_new_n9747__ = pi17 & ~new_new_n9746__;
  assign new_new_n9748__ = ~new_new_n6410__ & new_new_n7942__;
  assign new_new_n9749__ = ~new_new_n9747__ & ~new_new_n9748__;
  assign new_new_n9750__ = new_new_n9745__ & ~new_new_n9749__;
  assign new_new_n9751__ = ~pi17 & ~new_new_n9745__;
  assign new_new_n9752__ = ~new_new_n9750__ & ~new_new_n9751__;
  assign new_new_n9753__ = ~new_new_n9574__ & ~new_new_n9575__;
  assign new_new_n9754__ = pi23 & ~new_new_n9582__;
  assign new_new_n9755__ = ~pi23 & new_new_n9582__;
  assign new_new_n9756__ = ~new_new_n9754__ & ~new_new_n9755__;
  assign new_new_n9757__ = new_new_n9753__ & new_new_n9756__;
  assign new_new_n9758__ = ~new_new_n9753__ & ~new_new_n9756__;
  assign new_new_n9759__ = ~new_new_n9757__ & ~new_new_n9758__;
  assign new_new_n9760__ = ~new_new_n3535__ & new_new_n6634__;
  assign new_new_n9761__ = ~new_new_n2024__ & ~new_new_n6625__;
  assign new_new_n9762__ = ~new_new_n2130__ & new_new_n6629__;
  assign new_new_n9763__ = ~new_new_n9760__ & ~new_new_n9761__;
  assign new_new_n9764__ = ~new_new_n9762__ & new_new_n9763__;
  assign new_new_n9765__ = new_new_n6631__ & new_new_n6854__;
  assign new_new_n9766__ = pi20 & ~new_new_n9765__;
  assign new_new_n9767__ = new_new_n6640__ & new_new_n6854__;
  assign new_new_n9768__ = ~new_new_n9766__ & ~new_new_n9767__;
  assign new_new_n9769__ = new_new_n9764__ & ~new_new_n9768__;
  assign new_new_n9770__ = ~pi20 & ~new_new_n9764__;
  assign new_new_n9771__ = ~new_new_n9769__ & ~new_new_n9770__;
  assign new_new_n9772__ = ~new_new_n9290__ & ~new_new_n9291__;
  assign new_new_n9773__ = new_new_n9555__ & ~new_new_n9772__;
  assign new_new_n9774__ = ~new_new_n9555__ & new_new_n9772__;
  assign new_new_n9775__ = ~new_new_n9773__ & ~new_new_n9774__;
  assign new_new_n9776__ = ~new_new_n2420__ & ~new_new_n6625__;
  assign new_new_n9777__ = ~new_new_n2024__ & new_new_n6634__;
  assign new_new_n9778__ = ~new_new_n2224__ & new_new_n6629__;
  assign new_new_n9779__ = ~new_new_n9776__ & ~new_new_n9777__;
  assign new_new_n9780__ = ~new_new_n9778__ & new_new_n9779__;
  assign new_new_n9781__ = new_new_n6631__ & new_new_n7313__;
  assign new_new_n9782__ = pi20 & ~new_new_n9781__;
  assign new_new_n9783__ = new_new_n6640__ & new_new_n7313__;
  assign new_new_n9784__ = ~new_new_n9782__ & ~new_new_n9783__;
  assign new_new_n9785__ = new_new_n9780__ & ~new_new_n9784__;
  assign new_new_n9786__ = ~pi20 & ~new_new_n9780__;
  assign new_new_n9787__ = ~new_new_n9785__ & ~new_new_n9786__;
  assign new_new_n9788__ = ~new_new_n9310__ & ~new_new_n9311__;
  assign new_new_n9789__ = new_new_n9535__ & new_new_n9788__;
  assign new_new_n9790__ = ~new_new_n9535__ & ~new_new_n9788__;
  assign new_new_n9791__ = ~new_new_n9789__ & ~new_new_n9790__;
  assign new_new_n9792__ = ~new_new_n2313__ & new_new_n6629__;
  assign new_new_n9793__ = ~new_new_n2420__ & new_new_n6634__;
  assign new_new_n9794__ = ~new_new_n6751__ & new_new_n6936__;
  assign new_new_n9795__ = ~new_new_n9792__ & ~new_new_n9793__;
  assign new_new_n9796__ = ~new_new_n9794__ & new_new_n9795__;
  assign new_new_n9797__ = ~pi18 & ~pi19;
  assign new_new_n9798__ = ~new_new_n2572__ & new_new_n9797__;
  assign new_new_n9799__ = pi20 & ~new_new_n9798__;
  assign new_new_n9800__ = pi18 & pi19;
  assign new_new_n9801__ = ~new_new_n2572__ & new_new_n9800__;
  assign new_new_n9802__ = ~pi20 & ~new_new_n9801__;
  assign new_new_n9803__ = pi17 & ~new_new_n9802__;
  assign new_new_n9804__ = ~new_new_n9799__ & ~new_new_n9803__;
  assign new_new_n9805__ = new_new_n9796__ & ~new_new_n9804__;
  assign new_new_n9806__ = ~pi20 & ~new_new_n9796__;
  assign new_new_n9807__ = ~new_new_n9805__ & ~new_new_n9806__;
  assign new_new_n9808__ = ~new_new_n2497__ & new_new_n6629__;
  assign new_new_n9809__ = ~new_new_n2636__ & ~new_new_n6625__;
  assign new_new_n9810__ = ~new_new_n2572__ & new_new_n6634__;
  assign new_new_n9811__ = ~new_new_n9808__ & ~new_new_n9809__;
  assign new_new_n9812__ = ~new_new_n9810__ & new_new_n9811__;
  assign new_new_n9813__ = new_new_n6631__ & new_new_n6804__;
  assign new_new_n9814__ = ~pi20 & ~new_new_n9813__;
  assign new_new_n9815__ = new_new_n6804__ & new_new_n7015__;
  assign new_new_n9816__ = ~new_new_n9814__ & ~new_new_n9815__;
  assign new_new_n9817__ = new_new_n9812__ & ~new_new_n9816__;
  assign new_new_n9818__ = pi20 & ~new_new_n9812__;
  assign new_new_n9819__ = ~new_new_n9817__ & ~new_new_n9818__;
  assign new_new_n9820__ = ~new_new_n2636__ & new_new_n6629__;
  assign new_new_n9821__ = ~new_new_n2737__ & ~new_new_n6625__;
  assign new_new_n9822__ = ~new_new_n9820__ & ~new_new_n9821__;
  assign new_new_n9823__ = new_new_n6631__ & ~new_new_n9126__;
  assign new_new_n9824__ = pi20 & ~new_new_n9823__;
  assign new_new_n9825__ = ~pi19 & new_new_n2497__;
  assign new_new_n9826__ = pi19 & ~new_new_n2497__;
  assign new_new_n9827__ = new_new_n6631__ & ~new_new_n9825__;
  assign new_new_n9828__ = ~new_new_n9826__ & new_new_n9827__;
  assign new_new_n9829__ = ~new_new_n6797__ & new_new_n9828__;
  assign new_new_n9830__ = ~new_new_n9824__ & ~new_new_n9829__;
  assign new_new_n9831__ = new_new_n9822__ & ~new_new_n9830__;
  assign new_new_n9832__ = new_new_n6631__ & new_new_n7772__;
  assign new_new_n9833__ = new_new_n9822__ & ~new_new_n9832__;
  assign new_new_n9834__ = ~pi20 & ~new_new_n9833__;
  assign new_new_n9835__ = ~new_new_n9831__ & ~new_new_n9834__;
  assign new_new_n9836__ = ~new_new_n9460__ & ~new_new_n9461__;
  assign new_new_n9837__ = ~new_new_n9471__ & new_new_n9836__;
  assign new_new_n9838__ = new_new_n9471__ & ~new_new_n9836__;
  assign new_new_n9839__ = ~new_new_n9837__ & ~new_new_n9838__;
  assign new_new_n9840__ = ~new_new_n9835__ & ~new_new_n9839__;
  assign new_new_n9841__ = new_new_n9835__ & new_new_n9839__;
  assign new_new_n9842__ = ~pi20 & new_new_n6936__;
  assign new_new_n9843__ = ~new_new_n2636__ & new_new_n9842__;
  assign new_new_n9844__ = ~new_new_n2886__ & ~new_new_n6625__;
  assign new_new_n9845__ = ~new_new_n2636__ & new_new_n6634__;
  assign new_new_n9846__ = ~new_new_n2737__ & new_new_n6629__;
  assign new_new_n9847__ = ~new_new_n9844__ & ~new_new_n9845__;
  assign new_new_n9848__ = ~new_new_n9846__ & new_new_n9847__;
  assign new_new_n9849__ = pi20 & new_new_n2636__;
  assign new_new_n9850__ = new_new_n9848__ & new_new_n9849__;
  assign new_new_n9851__ = ~new_new_n9843__ & ~new_new_n9850__;
  assign new_new_n9852__ = ~new_new_n7811__ & ~new_new_n9851__;
  assign new_new_n9853__ = new_new_n2636__ & new_new_n9842__;
  assign new_new_n9854__ = pi20 & ~new_new_n2636__;
  assign new_new_n9855__ = new_new_n9848__ & new_new_n9854__;
  assign new_new_n9856__ = ~new_new_n9853__ & ~new_new_n9855__;
  assign new_new_n9857__ = new_new_n7811__ & ~new_new_n9856__;
  assign new_new_n9858__ = ~pi20 & ~new_new_n9848__;
  assign new_new_n9859__ = pi20 & ~new_new_n7015__;
  assign new_new_n9860__ = new_new_n9848__ & new_new_n9859__;
  assign new_new_n9861__ = ~new_new_n9858__ & ~new_new_n9860__;
  assign new_new_n9862__ = ~new_new_n9852__ & new_new_n9861__;
  assign new_new_n9863__ = ~new_new_n9857__ & new_new_n9862__;
  assign new_new_n9864__ = new_new_n6936__ & ~new_new_n7378__;
  assign new_new_n9865__ = ~new_new_n2886__ & new_new_n6629__;
  assign new_new_n9866__ = ~new_new_n2737__ & new_new_n6634__;
  assign new_new_n9867__ = ~new_new_n9865__ & ~new_new_n9866__;
  assign new_new_n9868__ = ~new_new_n9864__ & new_new_n9867__;
  assign new_new_n9869__ = ~new_new_n2848__ & new_new_n9797__;
  assign new_new_n9870__ = pi20 & ~new_new_n9869__;
  assign new_new_n9871__ = ~new_new_n2848__ & new_new_n9800__;
  assign new_new_n9872__ = ~pi20 & ~new_new_n9871__;
  assign new_new_n9873__ = pi17 & ~new_new_n9872__;
  assign new_new_n9874__ = ~new_new_n9870__ & ~new_new_n9873__;
  assign new_new_n9875__ = new_new_n9868__ & ~new_new_n9874__;
  assign new_new_n9876__ = ~pi20 & ~new_new_n9868__;
  assign new_new_n9877__ = ~new_new_n9875__ & ~new_new_n9876__;
  assign new_new_n9878__ = ~new_new_n2848__ & new_new_n6629__;
  assign new_new_n9879__ = ~new_new_n2886__ & new_new_n6634__;
  assign new_new_n9880__ = ~new_new_n3460__ & ~new_new_n6625__;
  assign new_new_n9881__ = new_new_n6936__ & ~new_new_n8574__;
  assign new_new_n9882__ = ~new_new_n9878__ & ~new_new_n9879__;
  assign new_new_n9883__ = ~new_new_n9880__ & new_new_n9882__;
  assign new_new_n9884__ = ~new_new_n9881__ & new_new_n9883__;
  assign new_new_n9885__ = pi20 & ~new_new_n9884__;
  assign new_new_n9886__ = ~pi20 & new_new_n9884__;
  assign new_new_n9887__ = ~new_new_n9885__ & ~new_new_n9886__;
  assign new_new_n9888__ = ~new_new_n9408__ & ~new_new_n9409__;
  assign new_new_n9889__ = new_new_n9419__ & ~new_new_n9888__;
  assign new_new_n9890__ = ~new_new_n9419__ & new_new_n9888__;
  assign new_new_n9891__ = ~new_new_n9889__ & ~new_new_n9890__;
  assign new_new_n9892__ = new_new_n6936__ & ~new_new_n7468__;
  assign new_new_n9893__ = ~new_new_n3126__ & new_new_n6629__;
  assign new_new_n9894__ = ~new_new_n3164__ & ~new_new_n6625__;
  assign new_new_n9895__ = ~new_new_n2960__ & new_new_n6634__;
  assign new_new_n9896__ = ~new_new_n9893__ & ~new_new_n9894__;
  assign new_new_n9897__ = ~new_new_n9895__ & new_new_n9896__;
  assign new_new_n9898__ = ~new_new_n9892__ & new_new_n9897__;
  assign new_new_n9899__ = ~pi20 & ~new_new_n9898__;
  assign new_new_n9900__ = pi20 & new_new_n9898__;
  assign new_new_n9901__ = ~new_new_n9899__ & ~new_new_n9900__;
  assign new_new_n9902__ = ~new_new_n3356__ & new_new_n9387__;
  assign new_new_n9903__ = ~new_new_n5181__ & ~new_new_n9902__;
  assign new_new_n9904__ = pi22 & ~new_new_n9903__;
  assign new_new_n9905__ = ~new_new_n3356__ & ~new_new_n5182__;
  assign new_new_n9906__ = ~new_new_n3055__ & new_new_n5195__;
  assign new_new_n9907__ = ~new_new_n9905__ & ~new_new_n9906__;
  assign new_new_n9908__ = ~new_new_n9904__ & ~new_new_n9907__;
  assign new_new_n9909__ = ~new_new_n3254__ & new_new_n6629__;
  assign new_new_n9910__ = ~new_new_n3164__ & new_new_n6634__;
  assign new_new_n9911__ = ~new_new_n3055__ & ~new_new_n6625__;
  assign new_new_n9912__ = new_new_n6936__ & ~new_new_n8637__;
  assign new_new_n9913__ = ~new_new_n9909__ & ~new_new_n9910__;
  assign new_new_n9914__ = ~new_new_n9911__ & new_new_n9913__;
  assign new_new_n9915__ = ~new_new_n9912__ & new_new_n9914__;
  assign new_new_n9916__ = pi20 & ~new_new_n9915__;
  assign new_new_n9917__ = ~pi20 & new_new_n9915__;
  assign new_new_n9918__ = ~new_new_n9916__ & ~new_new_n9917__;
  assign new_new_n9919__ = ~new_new_n3356__ & new_new_n5195__;
  assign new_new_n9920__ = pi19 & new_new_n6619__;
  assign new_new_n9921__ = ~new_new_n6623__ & ~new_new_n9920__;
  assign new_new_n9922__ = ~new_new_n9017__ & new_new_n9921__;
  assign new_new_n9923__ = ~new_new_n3254__ & new_new_n6631__;
  assign new_new_n9924__ = new_new_n6625__ & ~new_new_n9923__;
  assign new_new_n9925__ = ~new_new_n3055__ & ~new_new_n6633__;
  assign new_new_n9926__ = new_new_n9923__ & ~new_new_n9925__;
  assign new_new_n9927__ = new_new_n3356__ & ~new_new_n9926__;
  assign new_new_n9928__ = ~new_new_n9924__ & ~new_new_n9927__;
  assign new_new_n9929__ = pi20 & ~new_new_n9922__;
  assign new_new_n9930__ = ~new_new_n9928__ & new_new_n9929__;
  assign new_new_n9931__ = ~new_new_n9919__ & ~new_new_n9930__;
  assign new_new_n9932__ = new_new_n9918__ & ~new_new_n9931__;
  assign new_new_n9933__ = new_new_n9908__ & new_new_n9932__;
  assign new_new_n9934__ = ~new_new_n9908__ & ~new_new_n9932__;
  assign new_new_n9935__ = new_new_n6936__ & ~new_new_n7570__;
  assign new_new_n9936__ = ~new_new_n3126__ & new_new_n6634__;
  assign new_new_n9937__ = ~new_new_n3164__ & new_new_n6629__;
  assign new_new_n9938__ = ~new_new_n3254__ & ~new_new_n6625__;
  assign new_new_n9939__ = ~new_new_n9936__ & ~new_new_n9937__;
  assign new_new_n9940__ = ~new_new_n9938__ & new_new_n9939__;
  assign new_new_n9941__ = ~new_new_n9935__ & new_new_n9940__;
  assign new_new_n9942__ = pi20 & ~new_new_n9941__;
  assign new_new_n9943__ = ~pi20 & new_new_n9941__;
  assign new_new_n9944__ = ~new_new_n9942__ & ~new_new_n9943__;
  assign new_new_n9945__ = ~new_new_n9934__ & new_new_n9944__;
  assign new_new_n9946__ = ~new_new_n9933__ & ~new_new_n9945__;
  assign new_new_n9947__ = new_new_n9901__ & new_new_n9946__;
  assign new_new_n9948__ = pi23 & new_new_n9390__;
  assign new_new_n9949__ = new_new_n9384__ & new_new_n9948__;
  assign new_new_n9950__ = ~new_new_n9384__ & new_new_n9391__;
  assign new_new_n9951__ = new_new_n9946__ & ~new_new_n9950__;
  assign new_new_n9952__ = ~new_new_n9901__ & ~new_new_n9951__;
  assign new_new_n9953__ = ~pi23 & ~new_new_n9384__;
  assign new_new_n9954__ = ~new_new_n9949__ & ~new_new_n9953__;
  assign new_new_n9955__ = ~new_new_n9952__ & new_new_n9954__;
  assign new_new_n9956__ = ~new_new_n9947__ & ~new_new_n9955__;
  assign new_new_n9957__ = ~new_new_n3460__ & new_new_n6634__;
  assign new_new_n9958__ = ~new_new_n3126__ & ~new_new_n6625__;
  assign new_new_n9959__ = ~new_new_n2960__ & new_new_n6629__;
  assign new_new_n9960__ = ~new_new_n9957__ & ~new_new_n9958__;
  assign new_new_n9961__ = ~new_new_n9959__ & new_new_n9960__;
  assign new_new_n9962__ = new_new_n6631__ & new_new_n7391__;
  assign new_new_n9963__ = pi20 & ~new_new_n9962__;
  assign new_new_n9964__ = new_new_n6640__ & new_new_n7391__;
  assign new_new_n9965__ = ~new_new_n9963__ & ~new_new_n9964__;
  assign new_new_n9966__ = new_new_n9961__ & ~new_new_n9965__;
  assign new_new_n9967__ = ~pi20 & ~new_new_n9961__;
  assign new_new_n9968__ = ~new_new_n9966__ & ~new_new_n9967__;
  assign new_new_n9969__ = ~new_new_n9956__ & new_new_n9968__;
  assign new_new_n9970__ = new_new_n9956__ & ~new_new_n9968__;
  assign new_new_n9971__ = new_new_n9392__ & new_new_n9393__;
  assign new_new_n9972__ = new_new_n9394__ & ~new_new_n9406__;
  assign new_new_n9973__ = ~new_new_n9407__ & ~new_new_n9972__;
  assign new_new_n9974__ = ~new_new_n9971__ & ~new_new_n9973__;
  assign new_new_n9975__ = ~new_new_n9970__ & new_new_n9974__;
  assign new_new_n9976__ = ~new_new_n9969__ & ~new_new_n9975__;
  assign new_new_n9977__ = new_new_n9891__ & ~new_new_n9976__;
  assign new_new_n9978__ = ~new_new_n9891__ & new_new_n9976__;
  assign new_new_n9979__ = ~new_new_n3460__ & new_new_n6629__;
  assign new_new_n9980__ = ~new_new_n2848__ & new_new_n6634__;
  assign new_new_n9981__ = ~new_new_n2960__ & ~new_new_n6625__;
  assign new_new_n9982__ = new_new_n6936__ & ~new_new_n7065__;
  assign new_new_n9983__ = ~new_new_n9979__ & ~new_new_n9980__;
  assign new_new_n9984__ = ~new_new_n9981__ & new_new_n9983__;
  assign new_new_n9985__ = ~new_new_n9982__ & new_new_n9984__;
  assign new_new_n9986__ = pi20 & ~new_new_n9985__;
  assign new_new_n9987__ = ~pi20 & new_new_n9985__;
  assign new_new_n9988__ = ~new_new_n9986__ & ~new_new_n9987__;
  assign new_new_n9989__ = ~new_new_n9978__ & ~new_new_n9988__;
  assign new_new_n9990__ = ~new_new_n9977__ & ~new_new_n9989__;
  assign new_new_n9991__ = ~new_new_n9887__ & ~new_new_n9990__;
  assign new_new_n9992__ = new_new_n9887__ & new_new_n9990__;
  assign new_new_n9993__ = ~new_new_n9422__ & ~new_new_n9423__;
  assign new_new_n9994__ = ~new_new_n9433__ & new_new_n9993__;
  assign new_new_n9995__ = new_new_n9433__ & ~new_new_n9993__;
  assign new_new_n9996__ = ~new_new_n9994__ & ~new_new_n9995__;
  assign new_new_n9997__ = ~new_new_n9992__ & ~new_new_n9996__;
  assign new_new_n9998__ = ~new_new_n9991__ & ~new_new_n9997__;
  assign new_new_n9999__ = new_new_n9877__ & ~new_new_n9998__;
  assign new_new_n10000__ = ~new_new_n9877__ & new_new_n9998__;
  assign new_new_n10001__ = new_new_n9035__ & new_new_n9435__;
  assign new_new_n10002__ = ~new_new_n9436__ & ~new_new_n10001__;
  assign new_new_n10003__ = ~new_new_n9035__ & new_new_n9439__;
  assign new_new_n10004__ = ~new_new_n9438__ & ~new_new_n10003__;
  assign new_new_n10005__ = new_new_n10002__ & ~new_new_n10004__;
  assign new_new_n10006__ = ~new_new_n10002__ & new_new_n10004__;
  assign new_new_n10007__ = ~new_new_n10005__ & ~new_new_n10006__;
  assign new_new_n10008__ = new_new_n9356__ & new_new_n10007__;
  assign new_new_n10009__ = ~new_new_n9356__ & ~new_new_n10007__;
  assign new_new_n10010__ = ~new_new_n10008__ & ~new_new_n10009__;
  assign new_new_n10011__ = ~new_new_n10000__ & new_new_n10010__;
  assign new_new_n10012__ = ~new_new_n9999__ & ~new_new_n10011__;
  assign new_new_n10013__ = ~new_new_n9863__ & new_new_n10012__;
  assign new_new_n10014__ = new_new_n9863__ & ~new_new_n10012__;
  assign new_new_n10015__ = ~new_new_n2848__ & new_new_n5195__;
  assign new_new_n10016__ = pi22 & ~new_new_n9342__;
  assign new_new_n10017__ = ~pi22 & new_new_n9342__;
  assign new_new_n10018__ = ~new_new_n10016__ & ~new_new_n10017__;
  assign new_new_n10019__ = new_new_n10015__ & ~new_new_n10018__;
  assign new_new_n10020__ = pi23 & ~new_new_n9342__;
  assign new_new_n10021__ = ~pi23 & new_new_n9342__;
  assign new_new_n10022__ = ~new_new_n10020__ & ~new_new_n10021__;
  assign new_new_n10023__ = ~new_new_n10015__ & new_new_n10022__;
  assign new_new_n10024__ = ~new_new_n10019__ & ~new_new_n10023__;
  assign new_new_n10025__ = new_new_n9452__ & ~new_new_n10024__;
  assign new_new_n10026__ = ~new_new_n9452__ & ~new_new_n10022__;
  assign new_new_n10027__ = ~new_new_n10025__ & ~new_new_n10026__;
  assign new_new_n10028__ = ~new_new_n9445__ & ~new_new_n10027__;
  assign new_new_n10029__ = new_new_n9445__ & new_new_n10027__;
  assign new_new_n10030__ = ~new_new_n10028__ & ~new_new_n10029__;
  assign new_new_n10031__ = ~new_new_n10014__ & new_new_n10030__;
  assign new_new_n10032__ = ~new_new_n10013__ & ~new_new_n10031__;
  assign new_new_n10033__ = ~new_new_n9841__ & ~new_new_n10032__;
  assign new_new_n10034__ = ~new_new_n9840__ & ~new_new_n10033__;
  assign new_new_n10035__ = new_new_n9819__ & ~new_new_n10034__;
  assign new_new_n10036__ = ~new_new_n9819__ & new_new_n10034__;
  assign new_new_n10037__ = ~new_new_n9474__ & ~new_new_n9475__;
  assign new_new_n10038__ = ~new_new_n9487__ & ~new_new_n10037__;
  assign new_new_n10039__ = new_new_n9487__ & new_new_n10037__;
  assign new_new_n10040__ = ~new_new_n10038__ & ~new_new_n10039__;
  assign new_new_n10041__ = ~new_new_n10036__ & ~new_new_n10040__;
  assign new_new_n10042__ = ~new_new_n10035__ & ~new_new_n10041__;
  assign new_new_n10043__ = new_new_n9491__ & ~new_new_n9511__;
  assign new_new_n10044__ = ~new_new_n9491__ & new_new_n9511__;
  assign new_new_n10045__ = ~new_new_n10043__ & ~new_new_n10044__;
  assign new_new_n10046__ = new_new_n9489__ & new_new_n10045__;
  assign new_new_n10047__ = ~new_new_n9489__ & ~new_new_n10045__;
  assign new_new_n10048__ = ~new_new_n10046__ & ~new_new_n10047__;
  assign new_new_n10049__ = new_new_n10042__ & new_new_n10048__;
  assign new_new_n10050__ = ~new_new_n10042__ & ~new_new_n10048__;
  assign new_new_n10051__ = new_new_n6936__ & ~new_new_n7236__;
  assign new_new_n10052__ = ~new_new_n2497__ & ~new_new_n6625__;
  assign new_new_n10053__ = ~new_new_n2313__ & new_new_n6634__;
  assign new_new_n10054__ = ~new_new_n2572__ & new_new_n6629__;
  assign new_new_n10055__ = ~new_new_n10052__ & ~new_new_n10053__;
  assign new_new_n10056__ = ~new_new_n10054__ & new_new_n10055__;
  assign new_new_n10057__ = ~new_new_n10051__ & new_new_n10056__;
  assign new_new_n10058__ = pi20 & ~new_new_n10057__;
  assign new_new_n10059__ = ~pi20 & new_new_n10057__;
  assign new_new_n10060__ = ~new_new_n10058__ & ~new_new_n10059__;
  assign new_new_n10061__ = ~new_new_n10050__ & ~new_new_n10060__;
  assign new_new_n10062__ = ~new_new_n10049__ & ~new_new_n10061__;
  assign new_new_n10063__ = new_new_n9807__ & ~new_new_n10062__;
  assign new_new_n10064__ = ~new_new_n9807__ & new_new_n10062__;
  assign new_new_n10065__ = ~new_new_n9516__ & ~new_new_n9517__;
  assign new_new_n10066__ = new_new_n9533__ & ~new_new_n10065__;
  assign new_new_n10067__ = ~new_new_n9533__ & new_new_n10065__;
  assign new_new_n10068__ = ~new_new_n10066__ & ~new_new_n10067__;
  assign new_new_n10069__ = ~new_new_n10064__ & ~new_new_n10068__;
  assign new_new_n10070__ = ~new_new_n10063__ & ~new_new_n10069__;
  assign new_new_n10071__ = ~new_new_n9791__ & ~new_new_n10070__;
  assign new_new_n10072__ = new_new_n9791__ & new_new_n10070__;
  assign new_new_n10073__ = ~new_new_n2313__ & ~new_new_n6625__;
  assign new_new_n10074__ = ~new_new_n2420__ & new_new_n6629__;
  assign new_new_n10075__ = ~new_new_n2224__ & new_new_n6634__;
  assign new_new_n10076__ = new_new_n6521__ & new_new_n6936__;
  assign new_new_n10077__ = ~new_new_n10073__ & ~new_new_n10074__;
  assign new_new_n10078__ = ~new_new_n10075__ & new_new_n10077__;
  assign new_new_n10079__ = ~new_new_n10076__ & new_new_n10078__;
  assign new_new_n10080__ = pi20 & ~new_new_n10079__;
  assign new_new_n10081__ = ~pi20 & new_new_n10079__;
  assign new_new_n10082__ = ~new_new_n10080__ & ~new_new_n10081__;
  assign new_new_n10083__ = ~new_new_n10072__ & ~new_new_n10082__;
  assign new_new_n10084__ = ~new_new_n10071__ & ~new_new_n10083__;
  assign new_new_n10085__ = new_new_n9787__ & ~new_new_n10084__;
  assign new_new_n10086__ = ~new_new_n9787__ & new_new_n10084__;
  assign new_new_n10087__ = ~new_new_n9542__ & ~new_new_n9543__;
  assign new_new_n10088__ = new_new_n9553__ & ~new_new_n10087__;
  assign new_new_n10089__ = ~new_new_n9553__ & new_new_n10087__;
  assign new_new_n10090__ = ~new_new_n10088__ & ~new_new_n10089__;
  assign new_new_n10091__ = ~new_new_n10086__ & ~new_new_n10090__;
  assign new_new_n10092__ = ~new_new_n10085__ & ~new_new_n10091__;
  assign new_new_n10093__ = new_new_n9775__ & ~new_new_n10092__;
  assign new_new_n10094__ = ~new_new_n9775__ & new_new_n10092__;
  assign new_new_n10095__ = ~new_new_n2224__ & ~new_new_n6625__;
  assign new_new_n10096__ = ~new_new_n2024__ & new_new_n6629__;
  assign new_new_n10097__ = ~new_new_n2130__ & new_new_n6634__;
  assign new_new_n10098__ = ~new_new_n6036__ & new_new_n6936__;
  assign new_new_n10099__ = ~new_new_n10095__ & ~new_new_n10096__;
  assign new_new_n10100__ = ~new_new_n10097__ & new_new_n10099__;
  assign new_new_n10101__ = ~new_new_n10098__ & new_new_n10100__;
  assign new_new_n10102__ = pi20 & ~new_new_n10101__;
  assign new_new_n10103__ = ~pi20 & new_new_n10101__;
  assign new_new_n10104__ = ~new_new_n10102__ & ~new_new_n10103__;
  assign new_new_n10105__ = ~new_new_n10094__ & ~new_new_n10104__;
  assign new_new_n10106__ = ~new_new_n10093__ & ~new_new_n10105__;
  assign new_new_n10107__ = new_new_n9771__ & ~new_new_n10106__;
  assign new_new_n10108__ = ~new_new_n9771__ & new_new_n10106__;
  assign new_new_n10109__ = ~new_new_n9558__ & ~new_new_n9559__;
  assign new_new_n10110__ = new_new_n9571__ & ~new_new_n10109__;
  assign new_new_n10111__ = ~new_new_n9571__ & new_new_n10109__;
  assign new_new_n10112__ = ~new_new_n10110__ & ~new_new_n10111__;
  assign new_new_n10113__ = ~new_new_n10108__ & new_new_n10112__;
  assign new_new_n10114__ = ~new_new_n10107__ & ~new_new_n10113__;
  assign new_new_n10115__ = ~new_new_n9759__ & ~new_new_n10114__;
  assign new_new_n10116__ = new_new_n9759__ & new_new_n10114__;
  assign new_new_n10117__ = ~new_new_n3535__ & new_new_n6629__;
  assign new_new_n10118__ = ~new_new_n2130__ & ~new_new_n6625__;
  assign new_new_n10119__ = new_new_n5501__ & ~new_new_n6633__;
  assign new_new_n10120__ = new_new_n1823__ & ~new_new_n10119__;
  assign new_new_n10121__ = ~new_new_n6633__ & new_new_n7273__;
  assign new_new_n10122__ = new_new_n6631__ & ~new_new_n10120__;
  assign new_new_n10123__ = ~new_new_n10121__ & new_new_n10122__;
  assign new_new_n10124__ = ~new_new_n10117__ & ~new_new_n10118__;
  assign new_new_n10125__ = ~new_new_n10123__ & new_new_n10124__;
  assign new_new_n10126__ = ~pi20 & new_new_n10125__;
  assign new_new_n10127__ = pi20 & ~new_new_n10125__;
  assign new_new_n10128__ = ~new_new_n10126__ & ~new_new_n10127__;
  assign new_new_n10129__ = ~new_new_n10116__ & ~new_new_n10128__;
  assign new_new_n10130__ = ~new_new_n10115__ & ~new_new_n10129__;
  assign new_new_n10131__ = ~new_new_n9752__ & new_new_n10130__;
  assign new_new_n10132__ = new_new_n9752__ & ~new_new_n10130__;
  assign new_new_n10133__ = ~new_new_n9241__ & ~new_new_n9587__;
  assign new_new_n10134__ = new_new_n9241__ & new_new_n9587__;
  assign new_new_n10135__ = ~new_new_n10133__ & ~new_new_n10134__;
  assign new_new_n10136__ = new_new_n9253__ & new_new_n10135__;
  assign new_new_n10137__ = ~new_new_n9253__ & ~new_new_n10135__;
  assign new_new_n10138__ = ~new_new_n10136__ & ~new_new_n10137__;
  assign new_new_n10139__ = ~new_new_n10132__ & ~new_new_n10138__;
  assign new_new_n10140__ = ~new_new_n10131__ & ~new_new_n10139__;
  assign new_new_n10141__ = new_new_n9740__ & ~new_new_n10140__;
  assign new_new_n10142__ = ~new_new_n9740__ & new_new_n10140__;
  assign new_new_n10143__ = ~new_new_n9590__ & ~new_new_n9591__;
  assign new_new_n10144__ = new_new_n9603__ & new_new_n10143__;
  assign new_new_n10145__ = ~new_new_n9603__ & ~new_new_n10143__;
  assign new_new_n10146__ = ~new_new_n10144__ & ~new_new_n10145__;
  assign new_new_n10147__ = ~new_new_n10142__ & ~new_new_n10146__;
  assign new_new_n10148__ = ~new_new_n10141__ & ~new_new_n10147__;
  assign new_new_n10149__ = new_new_n9724__ & new_new_n10148__;
  assign new_new_n10150__ = ~new_new_n9724__ & ~new_new_n10148__;
  assign new_new_n10151__ = ~new_new_n10149__ & ~new_new_n10150__;
  assign new_new_n10152__ = ~new_new_n9610__ & ~new_new_n9611__;
  assign new_new_n10153__ = new_new_n9628__ & new_new_n10152__;
  assign new_new_n10154__ = ~new_new_n9628__ & ~new_new_n10152__;
  assign new_new_n10155__ = ~new_new_n10153__ & ~new_new_n10154__;
  assign new_new_n10156__ = new_new_n10151__ & ~new_new_n10155__;
  assign new_new_n10157__ = ~new_new_n10151__ & new_new_n10155__;
  assign new_new_n10158__ = ~new_new_n10156__ & ~new_new_n10157__;
  assign new_new_n10159__ = ~new_new_n10141__ & ~new_new_n10142__;
  assign new_new_n10160__ = ~new_new_n10146__ & new_new_n10159__;
  assign new_new_n10161__ = new_new_n10146__ & ~new_new_n10159__;
  assign new_new_n10162__ = ~new_new_n10160__ & ~new_new_n10161__;
  assign new_new_n10163__ = new_new_n8344__ & new_new_n8388__;
  assign new_new_n10164__ = ~new_new_n1556__ & new_new_n6991__;
  assign new_new_n10165__ = ~new_new_n1325__ & new_new_n6985__;
  assign new_new_n10166__ = ~new_new_n10164__ & ~new_new_n10165__;
  assign new_new_n10167__ = ~new_new_n5746__ & new_new_n6994__;
  assign new_new_n10168__ = ~pi14 & ~new_new_n10167__;
  assign new_new_n10169__ = new_new_n5061__ & new_new_n8820__;
  assign new_new_n10170__ = ~new_new_n10168__ & ~new_new_n10169__;
  assign new_new_n10171__ = new_new_n10166__ & ~new_new_n10170__;
  assign new_new_n10172__ = new_new_n5756__ & new_new_n6994__;
  assign new_new_n10173__ = new_new_n10166__ & ~new_new_n10172__;
  assign new_new_n10174__ = pi14 & ~new_new_n10173__;
  assign new_new_n10175__ = ~new_new_n10163__ & ~new_new_n10174__;
  assign new_new_n10176__ = ~new_new_n10171__ & new_new_n10175__;
  assign new_new_n10177__ = ~new_new_n10131__ & ~new_new_n10132__;
  assign new_new_n10178__ = ~new_new_n9254__ & ~new_new_n9255__;
  assign new_new_n10179__ = ~new_new_n9587__ & new_new_n10178__;
  assign new_new_n10180__ = new_new_n9587__ & ~new_new_n10178__;
  assign new_new_n10181__ = ~new_new_n10179__ & ~new_new_n10180__;
  assign new_new_n10182__ = new_new_n10177__ & ~new_new_n10181__;
  assign new_new_n10183__ = ~new_new_n10177__ & new_new_n10181__;
  assign new_new_n10184__ = ~new_new_n10182__ & ~new_new_n10183__;
  assign new_new_n10185__ = ~new_new_n10176__ & ~new_new_n10184__;
  assign new_new_n10186__ = new_new_n10176__ & new_new_n10184__;
  assign new_new_n10187__ = ~new_new_n10115__ & ~new_new_n10116__;
  assign new_new_n10188__ = new_new_n10128__ & ~new_new_n10187__;
  assign new_new_n10189__ = ~new_new_n10128__ & new_new_n10187__;
  assign new_new_n10190__ = ~new_new_n10188__ & ~new_new_n10189__;
  assign new_new_n10191__ = ~new_new_n1823__ & new_new_n6968__;
  assign new_new_n10192__ = ~new_new_n1902__ & new_new_n7935__;
  assign new_new_n10193__ = ~new_new_n3535__ & new_new_n6964__;
  assign new_new_n10194__ = ~new_new_n6487__ & new_new_n6959__;
  assign new_new_n10195__ = ~new_new_n10191__ & ~new_new_n10192__;
  assign new_new_n10196__ = ~new_new_n10193__ & new_new_n10195__;
  assign new_new_n10197__ = ~new_new_n10194__ & new_new_n10196__;
  assign new_new_n10198__ = ~pi17 & ~new_new_n10197__;
  assign new_new_n10199__ = pi17 & new_new_n10197__;
  assign new_new_n10200__ = ~new_new_n10198__ & ~new_new_n10199__;
  assign new_new_n10201__ = ~new_new_n10093__ & ~new_new_n10094__;
  assign new_new_n10202__ = ~new_new_n10104__ & new_new_n10201__;
  assign new_new_n10203__ = new_new_n10104__ & ~new_new_n10201__;
  assign new_new_n10204__ = ~new_new_n10202__ & ~new_new_n10203__;
  assign new_new_n10205__ = ~new_new_n10200__ & ~new_new_n10204__;
  assign new_new_n10206__ = ~new_new_n2024__ & new_new_n6964__;
  assign new_new_n10207__ = ~new_new_n2130__ & new_new_n6968__;
  assign new_new_n10208__ = ~new_new_n10206__ & ~new_new_n10207__;
  assign new_new_n10209__ = ~new_new_n3535__ & ~new_new_n6853__;
  assign new_new_n10210__ = new_new_n6958__ & new_new_n10209__;
  assign new_new_n10211__ = new_new_n10208__ & ~new_new_n10210__;
  assign new_new_n10212__ = ~pi17 & ~new_new_n10211__;
  assign new_new_n10213__ = ~new_new_n6850__ & new_new_n6958__;
  assign new_new_n10214__ = pi17 & ~new_new_n10213__;
  assign new_new_n10215__ = new_new_n3535__ & new_new_n5500__;
  assign new_new_n10216__ = pi16 & ~new_new_n10215__;
  assign new_new_n10217__ = ~pi16 & ~new_new_n6853__;
  assign new_new_n10218__ = new_new_n6958__ & ~new_new_n10216__;
  assign new_new_n10219__ = ~new_new_n10217__ & new_new_n10218__;
  assign new_new_n10220__ = ~new_new_n10214__ & ~new_new_n10219__;
  assign new_new_n10221__ = new_new_n10208__ & ~new_new_n10220__;
  assign new_new_n10222__ = ~new_new_n10212__ & ~new_new_n10221__;
  assign new_new_n10223__ = ~new_new_n10071__ & ~new_new_n10072__;
  assign new_new_n10224__ = ~new_new_n10082__ & new_new_n10223__;
  assign new_new_n10225__ = new_new_n10082__ & ~new_new_n10223__;
  assign new_new_n10226__ = ~new_new_n10224__ & ~new_new_n10225__;
  assign new_new_n10227__ = new_new_n10222__ & new_new_n10226__;
  assign new_new_n10228__ = ~new_new_n10222__ & ~new_new_n10226__;
  assign new_new_n10229__ = ~new_new_n10035__ & ~new_new_n10036__;
  assign new_new_n10230__ = new_new_n10040__ & ~new_new_n10229__;
  assign new_new_n10231__ = ~new_new_n10040__ & new_new_n10229__;
  assign new_new_n10232__ = ~new_new_n10230__ & ~new_new_n10231__;
  assign new_new_n10233__ = ~new_new_n10049__ & ~new_new_n10050__;
  assign new_new_n10234__ = ~new_new_n10060__ & new_new_n10233__;
  assign new_new_n10235__ = new_new_n10060__ & ~new_new_n10233__;
  assign new_new_n10236__ = ~new_new_n10234__ & ~new_new_n10235__;
  assign new_new_n10237__ = ~new_new_n2313__ & new_new_n6964__;
  assign new_new_n10238__ = ~new_new_n2224__ & new_new_n7935__;
  assign new_new_n10239__ = ~new_new_n2420__ & new_new_n6968__;
  assign new_new_n10240__ = new_new_n6521__ & new_new_n6959__;
  assign new_new_n10241__ = ~new_new_n10237__ & ~new_new_n10238__;
  assign new_new_n10242__ = ~new_new_n10239__ & new_new_n10241__;
  assign new_new_n10243__ = ~new_new_n10240__ & new_new_n10242__;
  assign new_new_n10244__ = new_new_n10236__ & new_new_n10243__;
  assign new_new_n10245__ = pi17 & ~new_new_n10243__;
  assign new_new_n10246__ = ~new_new_n10244__ & ~new_new_n10245__;
  assign new_new_n10247__ = ~new_new_n2024__ & new_new_n7935__;
  assign new_new_n10248__ = ~new_new_n2224__ & new_new_n6968__;
  assign new_new_n10249__ = ~new_new_n2420__ & new_new_n6964__;
  assign new_new_n10250__ = new_new_n6959__ & new_new_n7313__;
  assign new_new_n10251__ = ~new_new_n10247__ & ~new_new_n10248__;
  assign new_new_n10252__ = ~new_new_n10249__ & new_new_n10251__;
  assign new_new_n10253__ = ~new_new_n10250__ & new_new_n10252__;
  assign new_new_n10254__ = new_new_n10246__ & ~new_new_n10253__;
  assign new_new_n10255__ = ~new_new_n10236__ & ~new_new_n10243__;
  assign new_new_n10256__ = ~new_new_n2572__ & new_new_n6964__;
  assign new_new_n10257__ = ~new_new_n2313__ & new_new_n6968__;
  assign new_new_n10258__ = ~new_new_n10256__ & ~new_new_n10257__;
  assign new_new_n10259__ = new_new_n6958__ & ~new_new_n9267__;
  assign new_new_n10260__ = pi17 & ~new_new_n10259__;
  assign new_new_n10261__ = ~pi16 & new_new_n2420__;
  assign new_new_n10262__ = pi16 & ~new_new_n2420__;
  assign new_new_n10263__ = new_new_n6958__ & ~new_new_n10261__;
  assign new_new_n10264__ = ~new_new_n10262__ & new_new_n10263__;
  assign new_new_n10265__ = new_new_n6748__ & new_new_n10264__;
  assign new_new_n10266__ = ~new_new_n10260__ & ~new_new_n10265__;
  assign new_new_n10267__ = new_new_n10258__ & ~new_new_n10266__;
  assign new_new_n10268__ = new_new_n6749__ & new_new_n6958__;
  assign new_new_n10269__ = new_new_n10258__ & ~new_new_n10268__;
  assign new_new_n10270__ = ~pi17 & ~new_new_n10269__;
  assign new_new_n10271__ = ~new_new_n10267__ & ~new_new_n10270__;
  assign new_new_n10272__ = ~new_new_n9840__ & ~new_new_n9841__;
  assign new_new_n10273__ = ~new_new_n10032__ & new_new_n10272__;
  assign new_new_n10274__ = new_new_n10032__ & ~new_new_n10272__;
  assign new_new_n10275__ = ~new_new_n10273__ & ~new_new_n10274__;
  assign new_new_n10276__ = ~new_new_n10271__ & new_new_n10275__;
  assign new_new_n10277__ = new_new_n10271__ & ~new_new_n10275__;
  assign new_new_n10278__ = ~new_new_n2636__ & new_new_n6964__;
  assign new_new_n10279__ = ~new_new_n2497__ & new_new_n6968__;
  assign new_new_n10280__ = ~new_new_n2572__ & new_new_n7935__;
  assign new_new_n10281__ = ~new_new_n10278__ & ~new_new_n10279__;
  assign new_new_n10282__ = ~new_new_n10280__ & new_new_n10281__;
  assign new_new_n10283__ = new_new_n6804__ & new_new_n6958__;
  assign new_new_n10284__ = pi17 & ~new_new_n10283__;
  assign new_new_n10285__ = new_new_n6804__ & new_new_n7942__;
  assign new_new_n10286__ = ~new_new_n10284__ & ~new_new_n10285__;
  assign new_new_n10287__ = new_new_n10282__ & ~new_new_n10286__;
  assign new_new_n10288__ = ~pi17 & ~new_new_n10282__;
  assign new_new_n10289__ = ~new_new_n10287__ & ~new_new_n10288__;
  assign new_new_n10290__ = ~new_new_n9999__ & ~new_new_n10000__;
  assign new_new_n10291__ = new_new_n10010__ & new_new_n10290__;
  assign new_new_n10292__ = ~new_new_n10010__ & ~new_new_n10290__;
  assign new_new_n10293__ = ~new_new_n10291__ & ~new_new_n10292__;
  assign new_new_n10294__ = new_new_n10289__ & new_new_n10293__;
  assign new_new_n10295__ = ~new_new_n10289__ & ~new_new_n10293__;
  assign new_new_n10296__ = ~new_new_n2636__ & new_new_n6968__;
  assign new_new_n10297__ = ~new_new_n2737__ & new_new_n6964__;
  assign new_new_n10298__ = ~new_new_n10296__ & ~new_new_n10297__;
  assign new_new_n10299__ = new_new_n6958__ & ~new_new_n9126__;
  assign new_new_n10300__ = pi17 & ~new_new_n10299__;
  assign new_new_n10301__ = ~pi16 & new_new_n2497__;
  assign new_new_n10302__ = pi16 & ~new_new_n2497__;
  assign new_new_n10303__ = new_new_n6958__ & ~new_new_n10301__;
  assign new_new_n10304__ = ~new_new_n10302__ & new_new_n10303__;
  assign new_new_n10305__ = ~new_new_n6797__ & new_new_n10304__;
  assign new_new_n10306__ = ~new_new_n10300__ & ~new_new_n10305__;
  assign new_new_n10307__ = new_new_n10298__ & ~new_new_n10306__;
  assign new_new_n10308__ = new_new_n6958__ & new_new_n7772__;
  assign new_new_n10309__ = new_new_n10298__ & ~new_new_n10308__;
  assign new_new_n10310__ = ~pi17 & ~new_new_n10309__;
  assign new_new_n10311__ = ~new_new_n10307__ & ~new_new_n10310__;
  assign new_new_n10312__ = ~new_new_n2737__ & new_new_n7935__;
  assign new_new_n10313__ = ~new_new_n2848__ & new_new_n6964__;
  assign new_new_n10314__ = ~new_new_n2886__ & new_new_n6968__;
  assign new_new_n10315__ = ~new_new_n10312__ & ~new_new_n10313__;
  assign new_new_n10316__ = ~new_new_n10314__ & new_new_n10315__;
  assign new_new_n10317__ = new_new_n6958__ & ~new_new_n7378__;
  assign new_new_n10318__ = pi17 & ~new_new_n10317__;
  assign new_new_n10319__ = ~new_new_n7378__ & new_new_n7942__;
  assign new_new_n10320__ = ~new_new_n10318__ & ~new_new_n10319__;
  assign new_new_n10321__ = new_new_n10316__ & ~new_new_n10320__;
  assign new_new_n10322__ = ~pi17 & ~new_new_n10316__;
  assign new_new_n10323__ = ~new_new_n10321__ & ~new_new_n10322__;
  assign new_new_n10324__ = ~new_new_n9947__ & new_new_n9955__;
  assign new_new_n10325__ = ~new_new_n9901__ & ~new_new_n9946__;
  assign new_new_n10326__ = ~new_new_n9947__ & ~new_new_n10325__;
  assign new_new_n10327__ = ~new_new_n9384__ & ~new_new_n9948__;
  assign new_new_n10328__ = ~new_new_n9949__ & ~new_new_n10327__;
  assign new_new_n10329__ = ~new_new_n10326__ & ~new_new_n10328__;
  assign new_new_n10330__ = ~new_new_n10324__ & ~new_new_n10329__;
  assign new_new_n10331__ = new_new_n6959__ & new_new_n7391__;
  assign new_new_n10332__ = ~new_new_n3460__ & new_new_n7935__;
  assign new_new_n10333__ = ~new_new_n2960__ & new_new_n6968__;
  assign new_new_n10334__ = ~new_new_n10332__ & ~new_new_n10333__;
  assign new_new_n10335__ = ~new_new_n10331__ & new_new_n10334__;
  assign new_new_n10336__ = ~pi17 & ~new_new_n10335__;
  assign new_new_n10337__ = ~pi15 & ~pi16;
  assign new_new_n10338__ = ~new_new_n3126__ & new_new_n10337__;
  assign new_new_n10339__ = pi17 & ~new_new_n10338__;
  assign new_new_n10340__ = pi15 & pi16;
  assign new_new_n10341__ = ~new_new_n3126__ & new_new_n10340__;
  assign new_new_n10342__ = ~pi17 & ~new_new_n10341__;
  assign new_new_n10343__ = pi14 & ~new_new_n10342__;
  assign new_new_n10344__ = ~new_new_n10339__ & ~new_new_n10343__;
  assign new_new_n10345__ = new_new_n10335__ & ~new_new_n10344__;
  assign new_new_n10346__ = ~new_new_n10336__ & ~new_new_n10345__;
  assign new_new_n10347__ = new_new_n9918__ & ~new_new_n9919__;
  assign new_new_n10348__ = ~new_new_n9918__ & new_new_n9919__;
  assign new_new_n10349__ = ~new_new_n9930__ & ~new_new_n10348__;
  assign new_new_n10350__ = ~new_new_n10347__ & ~new_new_n10349__;
  assign new_new_n10351__ = new_new_n6936__ & new_new_n7682__;
  assign new_new_n10352__ = ~new_new_n6629__ & ~new_new_n10351__;
  assign new_new_n10353__ = ~new_new_n3055__ & ~new_new_n10352__;
  assign new_new_n10354__ = ~new_new_n9928__ & ~new_new_n10353__;
  assign new_new_n10355__ = ~new_new_n3055__ & ~new_new_n6622__;
  assign new_new_n10356__ = ~new_new_n6619__ & new_new_n10355__;
  assign new_new_n10357__ = new_new_n3356__ & ~new_new_n10356__;
  assign new_new_n10358__ = pi20 & new_new_n9921__;
  assign new_new_n10359__ = ~new_new_n10357__ & new_new_n10358__;
  assign new_new_n10360__ = ~new_new_n10354__ & new_new_n10359__;
  assign new_new_n10361__ = new_new_n10354__ & ~new_new_n10359__;
  assign new_new_n10362__ = ~new_new_n10360__ & ~new_new_n10361__;
  assign new_new_n10363__ = new_new_n6628__ & ~new_new_n10356__;
  assign new_new_n10364__ = ~new_new_n3356__ & new_new_n10355__;
  assign new_new_n10365__ = ~new_new_n6619__ & ~new_new_n10364__;
  assign new_new_n10366__ = pi19 & ~new_new_n10365__;
  assign new_new_n10367__ = ~new_new_n10357__ & ~new_new_n10363__;
  assign new_new_n10368__ = ~new_new_n10366__ & new_new_n10367__;
  assign new_new_n10369__ = ~new_new_n3055__ & new_new_n6964__;
  assign new_new_n10370__ = ~new_new_n3164__ & new_new_n7935__;
  assign new_new_n10371__ = ~new_new_n3254__ & new_new_n6968__;
  assign new_new_n10372__ = ~new_new_n10369__ & ~new_new_n10370__;
  assign new_new_n10373__ = ~new_new_n10371__ & new_new_n10372__;
  assign new_new_n10374__ = ~pi17 & ~new_new_n10373__;
  assign new_new_n10375__ = new_new_n8160__ & ~new_new_n8637__;
  assign new_new_n10376__ = new_new_n6958__ & ~new_new_n8637__;
  assign new_new_n10377__ = ~pi17 & ~new_new_n10376__;
  assign new_new_n10378__ = new_new_n10373__ & ~new_new_n10375__;
  assign new_new_n10379__ = ~new_new_n10377__ & new_new_n10378__;
  assign new_new_n10380__ = ~new_new_n10374__ & ~new_new_n10379__;
  assign new_new_n10381__ = ~new_new_n3356__ & new_new_n6631__;
  assign new_new_n10382__ = ~new_new_n10380__ & new_new_n10381__;
  assign new_new_n10383__ = ~new_new_n3254__ & new_new_n6964__;
  assign new_new_n10384__ = ~new_new_n3164__ & new_new_n6968__;
  assign new_new_n10385__ = new_new_n6959__ & ~new_new_n7570__;
  assign new_new_n10386__ = ~new_new_n10383__ & ~new_new_n10384__;
  assign new_new_n10387__ = ~new_new_n10385__ & new_new_n10386__;
  assign new_new_n10388__ = ~new_new_n3126__ & new_new_n6958__;
  assign new_new_n10389__ = ~pi17 & ~new_new_n10388__;
  assign new_new_n10390__ = ~new_new_n3126__ & new_new_n7942__;
  assign new_new_n10391__ = ~new_new_n10389__ & ~new_new_n10390__;
  assign new_new_n10392__ = new_new_n10387__ & ~new_new_n10391__;
  assign new_new_n10393__ = pi17 & ~new_new_n10387__;
  assign new_new_n10394__ = ~new_new_n10392__ & ~new_new_n10393__;
  assign new_new_n10395__ = ~new_new_n10382__ & ~new_new_n10394__;
  assign new_new_n10396__ = new_new_n10368__ & ~new_new_n10395__;
  assign new_new_n10397__ = new_new_n6959__ & new_new_n7682__;
  assign new_new_n10398__ = ~new_new_n6968__ & ~new_new_n10397__;
  assign new_new_n10399__ = ~new_new_n3055__ & ~new_new_n10398__;
  assign new_new_n10400__ = ~new_new_n3254__ & new_new_n6958__;
  assign new_new_n10401__ = ~new_new_n6964__ & ~new_new_n10400__;
  assign new_new_n10402__ = ~new_new_n3055__ & new_new_n6955__;
  assign new_new_n10403__ = new_new_n10400__ & ~new_new_n10402__;
  assign new_new_n10404__ = new_new_n3356__ & ~new_new_n10403__;
  assign new_new_n10405__ = ~new_new_n10401__ & ~new_new_n10404__;
  assign new_new_n10406__ = ~new_new_n10399__ & ~new_new_n10405__;
  assign new_new_n10407__ = ~pi16 & ~new_new_n3356__;
  assign new_new_n10408__ = new_new_n6957__ & ~new_new_n10407__;
  assign new_new_n10409__ = ~new_new_n3055__ & ~new_new_n6956__;
  assign new_new_n10410__ = new_new_n3356__ & ~new_new_n10409__;
  assign new_new_n10411__ = pi17 & ~new_new_n6961__;
  assign new_new_n10412__ = ~new_new_n10408__ & new_new_n10411__;
  assign new_new_n10413__ = ~new_new_n10410__ & new_new_n10412__;
  assign new_new_n10414__ = new_new_n10406__ & ~new_new_n10413__;
  assign new_new_n10415__ = pi17 & new_new_n10414__;
  assign new_new_n10416__ = new_new_n10379__ & new_new_n10415__;
  assign new_new_n10417__ = ~new_new_n10382__ & ~new_new_n10416__;
  assign new_new_n10418__ = new_new_n10394__ & ~new_new_n10417__;
  assign new_new_n10419__ = ~new_new_n10396__ & ~new_new_n10418__;
  assign new_new_n10420__ = new_new_n10362__ & ~new_new_n10419__;
  assign new_new_n10421__ = ~new_new_n10362__ & new_new_n10419__;
  assign new_new_n10422__ = ~new_new_n2960__ & new_new_n7935__;
  assign new_new_n10423__ = ~new_new_n3126__ & new_new_n6968__;
  assign new_new_n10424__ = ~new_new_n3164__ & new_new_n6964__;
  assign new_new_n10425__ = new_new_n6959__ & ~new_new_n7468__;
  assign new_new_n10426__ = ~new_new_n10423__ & ~new_new_n10424__;
  assign new_new_n10427__ = ~new_new_n10422__ & new_new_n10426__;
  assign new_new_n10428__ = ~new_new_n10425__ & new_new_n10427__;
  assign new_new_n10429__ = pi17 & ~new_new_n10428__;
  assign new_new_n10430__ = ~pi17 & new_new_n10428__;
  assign new_new_n10431__ = ~new_new_n10429__ & ~new_new_n10430__;
  assign new_new_n10432__ = ~new_new_n10421__ & new_new_n10431__;
  assign new_new_n10433__ = ~new_new_n10420__ & ~new_new_n10432__;
  assign new_new_n10434__ = ~new_new_n10350__ & new_new_n10433__;
  assign new_new_n10435__ = ~new_new_n10346__ & ~new_new_n10434__;
  assign new_new_n10436__ = ~new_new_n10346__ & new_new_n10347__;
  assign new_new_n10437__ = new_new_n10433__ & ~new_new_n10436__;
  assign new_new_n10438__ = ~new_new_n10347__ & ~new_new_n10348__;
  assign new_new_n10439__ = ~new_new_n9930__ & ~new_new_n10438__;
  assign new_new_n10440__ = ~new_new_n10437__ & new_new_n10439__;
  assign new_new_n10441__ = ~new_new_n10435__ & ~new_new_n10440__;
  assign new_new_n10442__ = ~new_new_n9933__ & ~new_new_n9934__;
  assign new_new_n10443__ = new_new_n9944__ & new_new_n10442__;
  assign new_new_n10444__ = ~new_new_n9944__ & ~new_new_n10442__;
  assign new_new_n10445__ = ~new_new_n10443__ & ~new_new_n10444__;
  assign new_new_n10446__ = new_new_n10441__ & ~new_new_n10445__;
  assign new_new_n10447__ = ~new_new_n10441__ & new_new_n10445__;
  assign new_new_n10448__ = ~new_new_n2960__ & new_new_n6964__;
  assign new_new_n10449__ = ~new_new_n2848__ & new_new_n7935__;
  assign new_new_n10450__ = ~new_new_n3460__ & new_new_n6968__;
  assign new_new_n10451__ = ~new_new_n10449__ & ~new_new_n10450__;
  assign new_new_n10452__ = ~new_new_n10448__ & new_new_n10451__;
  assign new_new_n10453__ = new_new_n6959__ & ~new_new_n7065__;
  assign new_new_n10454__ = new_new_n10452__ & ~new_new_n10453__;
  assign new_new_n10455__ = pi17 & ~new_new_n10454__;
  assign new_new_n10456__ = ~pi17 & new_new_n10454__;
  assign new_new_n10457__ = ~new_new_n10455__ & ~new_new_n10456__;
  assign new_new_n10458__ = ~new_new_n10447__ & ~new_new_n10457__;
  assign new_new_n10459__ = ~new_new_n10446__ & ~new_new_n10458__;
  assign new_new_n10460__ = new_new_n10330__ & ~new_new_n10459__;
  assign new_new_n10461__ = ~new_new_n10330__ & new_new_n10459__;
  assign new_new_n10462__ = ~new_new_n3460__ & new_new_n6964__;
  assign new_new_n10463__ = ~new_new_n2848__ & new_new_n6968__;
  assign new_new_n10464__ = ~new_new_n2886__ & new_new_n7935__;
  assign new_new_n10465__ = new_new_n6959__ & ~new_new_n8574__;
  assign new_new_n10466__ = ~new_new_n10462__ & ~new_new_n10463__;
  assign new_new_n10467__ = ~new_new_n10464__ & new_new_n10466__;
  assign new_new_n10468__ = ~new_new_n10465__ & new_new_n10467__;
  assign new_new_n10469__ = pi17 & ~new_new_n10468__;
  assign new_new_n10470__ = ~pi17 & new_new_n10468__;
  assign new_new_n10471__ = ~new_new_n10469__ & ~new_new_n10470__;
  assign new_new_n10472__ = ~new_new_n10461__ & ~new_new_n10471__;
  assign new_new_n10473__ = ~new_new_n10460__ & ~new_new_n10472__;
  assign new_new_n10474__ = ~new_new_n10323__ & new_new_n10473__;
  assign new_new_n10475__ = new_new_n10323__ & ~new_new_n10473__;
  assign new_new_n10476__ = ~new_new_n9969__ & ~new_new_n9970__;
  assign new_new_n10477__ = new_new_n9974__ & new_new_n10476__;
  assign new_new_n10478__ = ~new_new_n9974__ & ~new_new_n10476__;
  assign new_new_n10479__ = ~new_new_n10477__ & ~new_new_n10478__;
  assign new_new_n10480__ = ~new_new_n10475__ & ~new_new_n10479__;
  assign new_new_n10481__ = ~new_new_n10474__ & ~new_new_n10480__;
  assign new_new_n10482__ = ~new_new_n9977__ & ~new_new_n9978__;
  assign new_new_n10483__ = new_new_n9988__ & new_new_n10482__;
  assign new_new_n10484__ = ~new_new_n9988__ & ~new_new_n10482__;
  assign new_new_n10485__ = ~new_new_n10483__ & ~new_new_n10484__;
  assign new_new_n10486__ = new_new_n10481__ & ~new_new_n10485__;
  assign new_new_n10487__ = ~new_new_n10481__ & new_new_n10485__;
  assign new_new_n10488__ = ~new_new_n2886__ & new_new_n6964__;
  assign new_new_n10489__ = ~new_new_n2636__ & new_new_n7935__;
  assign new_new_n10490__ = ~new_new_n2737__ & new_new_n6968__;
  assign new_new_n10491__ = ~new_new_n10488__ & ~new_new_n10489__;
  assign new_new_n10492__ = ~new_new_n10490__ & new_new_n10491__;
  assign new_new_n10493__ = ~pi17 & new_new_n10492__;
  assign new_new_n10494__ = ~new_new_n7942__ & new_new_n10493__;
  assign new_new_n10495__ = ~new_new_n2636__ & new_new_n6959__;
  assign new_new_n10496__ = ~new_new_n10493__ & ~new_new_n10495__;
  assign new_new_n10497__ = ~pi17 & ~new_new_n2636__;
  assign new_new_n10498__ = ~new_new_n10496__ & ~new_new_n10497__;
  assign new_new_n10499__ = ~new_new_n7811__ & new_new_n10498__;
  assign new_new_n10500__ = pi17 & new_new_n6959__;
  assign new_new_n10501__ = new_new_n2636__ & new_new_n10500__;
  assign new_new_n10502__ = new_new_n10492__ & new_new_n10497__;
  assign new_new_n10503__ = ~new_new_n10501__ & ~new_new_n10502__;
  assign new_new_n10504__ = new_new_n7811__ & ~new_new_n10503__;
  assign new_new_n10505__ = pi17 & ~new_new_n10492__;
  assign new_new_n10506__ = ~new_new_n10494__ & ~new_new_n10505__;
  assign new_new_n10507__ = ~new_new_n10499__ & new_new_n10506__;
  assign new_new_n10508__ = ~new_new_n10504__ & new_new_n10507__;
  assign new_new_n10509__ = ~new_new_n10487__ & ~new_new_n10508__;
  assign new_new_n10510__ = ~new_new_n10486__ & ~new_new_n10509__;
  assign new_new_n10511__ = ~new_new_n10311__ & new_new_n10510__;
  assign new_new_n10512__ = new_new_n10311__ & ~new_new_n10510__;
  assign new_new_n10513__ = ~new_new_n9991__ & ~new_new_n9992__;
  assign new_new_n10514__ = ~new_new_n9996__ & new_new_n10513__;
  assign new_new_n10515__ = new_new_n9996__ & ~new_new_n10513__;
  assign new_new_n10516__ = ~new_new_n10514__ & ~new_new_n10515__;
  assign new_new_n10517__ = ~new_new_n10512__ & ~new_new_n10516__;
  assign new_new_n10518__ = ~new_new_n10511__ & ~new_new_n10517__;
  assign new_new_n10519__ = ~new_new_n10295__ & new_new_n10518__;
  assign new_new_n10520__ = ~new_new_n10294__ & ~new_new_n10519__;
  assign new_new_n10521__ = ~new_new_n10013__ & ~new_new_n10014__;
  assign new_new_n10522__ = new_new_n9445__ & ~new_new_n10027__;
  assign new_new_n10523__ = ~new_new_n9445__ & new_new_n10027__;
  assign new_new_n10524__ = ~new_new_n10522__ & ~new_new_n10523__;
  assign new_new_n10525__ = new_new_n10521__ & new_new_n10524__;
  assign new_new_n10526__ = ~new_new_n10521__ & ~new_new_n10524__;
  assign new_new_n10527__ = ~new_new_n10525__ & ~new_new_n10526__;
  assign new_new_n10528__ = new_new_n10520__ & ~new_new_n10527__;
  assign new_new_n10529__ = ~new_new_n10520__ & new_new_n10527__;
  assign new_new_n10530__ = ~new_new_n2313__ & new_new_n7935__;
  assign new_new_n10531__ = ~new_new_n2497__ & new_new_n6964__;
  assign new_new_n10532__ = ~new_new_n2572__ & new_new_n6968__;
  assign new_new_n10533__ = ~new_new_n10530__ & ~new_new_n10531__;
  assign new_new_n10534__ = ~new_new_n10532__ & new_new_n10533__;
  assign new_new_n10535__ = new_new_n6958__ & ~new_new_n7236__;
  assign new_new_n10536__ = ~pi17 & ~new_new_n10535__;
  assign new_new_n10537__ = ~new_new_n7236__ & new_new_n8160__;
  assign new_new_n10538__ = ~new_new_n10536__ & ~new_new_n10537__;
  assign new_new_n10539__ = new_new_n10534__ & ~new_new_n10538__;
  assign new_new_n10540__ = pi17 & ~new_new_n10534__;
  assign new_new_n10541__ = ~new_new_n10539__ & ~new_new_n10540__;
  assign new_new_n10542__ = ~new_new_n10529__ & new_new_n10541__;
  assign new_new_n10543__ = ~new_new_n10528__ & ~new_new_n10542__;
  assign new_new_n10544__ = ~new_new_n10277__ & ~new_new_n10543__;
  assign new_new_n10545__ = ~new_new_n10276__ & ~new_new_n10544__;
  assign new_new_n10546__ = ~new_new_n10243__ & new_new_n10545__;
  assign new_new_n10547__ = pi17 & ~new_new_n10546__;
  assign new_new_n10548__ = ~new_new_n10255__ & ~new_new_n10547__;
  assign new_new_n10549__ = new_new_n10253__ & ~new_new_n10548__;
  assign new_new_n10550__ = ~pi17 & ~new_new_n10253__;
  assign new_new_n10551__ = new_new_n10236__ & ~new_new_n10550__;
  assign new_new_n10552__ = ~new_new_n10545__ & ~new_new_n10551__;
  assign new_new_n10553__ = ~new_new_n10254__ & ~new_new_n10552__;
  assign new_new_n10554__ = ~new_new_n10549__ & new_new_n10553__;
  assign new_new_n10555__ = new_new_n10232__ & ~new_new_n10554__;
  assign new_new_n10556__ = pi17 & ~new_new_n10236__;
  assign new_new_n10557__ = ~pi17 & new_new_n10243__;
  assign new_new_n10558__ = new_new_n10236__ & ~new_new_n10243__;
  assign new_new_n10559__ = ~new_new_n10545__ & ~new_new_n10557__;
  assign new_new_n10560__ = ~new_new_n10558__ & new_new_n10559__;
  assign new_new_n10561__ = ~new_new_n10556__ & ~new_new_n10560__;
  assign new_new_n10562__ = new_new_n10253__ & ~new_new_n10561__;
  assign new_new_n10563__ = ~pi17 & ~new_new_n10236__;
  assign new_new_n10564__ = new_new_n10246__ & ~new_new_n10545__;
  assign new_new_n10565__ = ~new_new_n10563__ & ~new_new_n10564__;
  assign new_new_n10566__ = ~new_new_n10253__ & ~new_new_n10565__;
  assign new_new_n10567__ = ~new_new_n10562__ & ~new_new_n10566__;
  assign new_new_n10568__ = ~new_new_n10555__ & new_new_n10567__;
  assign new_new_n10569__ = ~new_new_n2024__ & new_new_n6968__;
  assign new_new_n10570__ = ~new_new_n2224__ & new_new_n6964__;
  assign new_new_n10571__ = ~new_new_n10569__ & ~new_new_n10570__;
  assign new_new_n10572__ = new_new_n6958__ & new_new_n9173__;
  assign new_new_n10573__ = new_new_n10571__ & ~new_new_n10572__;
  assign new_new_n10574__ = pi17 & ~new_new_n10573__;
  assign new_new_n10575__ = new_new_n6958__ & ~new_new_n9177__;
  assign new_new_n10576__ = ~pi17 & ~new_new_n10575__;
  assign new_new_n10577__ = ~pi16 & ~new_new_n9180__;
  assign new_new_n10578__ = pi16 & ~new_new_n9182__;
  assign new_new_n10579__ = new_new_n6958__ & ~new_new_n10577__;
  assign new_new_n10580__ = ~new_new_n10578__ & new_new_n10579__;
  assign new_new_n10581__ = ~new_new_n10576__ & ~new_new_n10580__;
  assign new_new_n10582__ = new_new_n10571__ & ~new_new_n10581__;
  assign new_new_n10583__ = ~new_new_n10574__ & ~new_new_n10582__;
  assign new_new_n10584__ = new_new_n10568__ & ~new_new_n10583__;
  assign new_new_n10585__ = ~new_new_n10568__ & new_new_n10583__;
  assign new_new_n10586__ = ~new_new_n10063__ & ~new_new_n10064__;
  assign new_new_n10587__ = ~new_new_n8967__ & ~new_new_n9533__;
  assign new_new_n10588__ = new_new_n8967__ & new_new_n9533__;
  assign new_new_n10589__ = ~new_new_n10587__ & ~new_new_n10588__;
  assign new_new_n10590__ = new_new_n9089__ & ~new_new_n9515__;
  assign new_new_n10591__ = ~new_new_n9089__ & new_new_n9515__;
  assign new_new_n10592__ = ~new_new_n10590__ & ~new_new_n10591__;
  assign new_new_n10593__ = new_new_n9095__ & ~new_new_n10592__;
  assign new_new_n10594__ = ~new_new_n9095__ & new_new_n10592__;
  assign new_new_n10595__ = ~new_new_n10593__ & ~new_new_n10594__;
  assign new_new_n10596__ = new_new_n10589__ & ~new_new_n10595__;
  assign new_new_n10597__ = ~new_new_n10589__ & new_new_n10595__;
  assign new_new_n10598__ = ~new_new_n10596__ & ~new_new_n10597__;
  assign new_new_n10599__ = ~new_new_n10586__ & new_new_n10598__;
  assign new_new_n10600__ = new_new_n10586__ & ~new_new_n10598__;
  assign new_new_n10601__ = ~new_new_n10599__ & ~new_new_n10600__;
  assign new_new_n10602__ = ~new_new_n10585__ & ~new_new_n10601__;
  assign new_new_n10603__ = ~new_new_n10584__ & ~new_new_n10602__;
  assign new_new_n10604__ = ~new_new_n10228__ & ~new_new_n10603__;
  assign new_new_n10605__ = ~new_new_n10227__ & ~new_new_n10604__;
  assign new_new_n10606__ = ~new_new_n9553__ & new_new_n9787__;
  assign new_new_n10607__ = new_new_n9553__ & ~new_new_n9787__;
  assign new_new_n10608__ = ~new_new_n10606__ & ~new_new_n10607__;
  assign new_new_n10609__ = new_new_n10087__ & ~new_new_n10608__;
  assign new_new_n10610__ = ~new_new_n10087__ & new_new_n10608__;
  assign new_new_n10611__ = ~new_new_n10609__ & ~new_new_n10610__;
  assign new_new_n10612__ = new_new_n10084__ & new_new_n10611__;
  assign new_new_n10613__ = ~new_new_n10084__ & ~new_new_n10611__;
  assign new_new_n10614__ = ~new_new_n10612__ & ~new_new_n10613__;
  assign new_new_n10615__ = new_new_n10605__ & new_new_n10614__;
  assign new_new_n10616__ = ~new_new_n3535__ & new_new_n6968__;
  assign new_new_n10617__ = ~new_new_n2130__ & new_new_n6964__;
  assign new_new_n10618__ = ~new_new_n10616__ & ~new_new_n10617__;
  assign new_new_n10619__ = ~new_new_n5520__ & new_new_n6958__;
  assign new_new_n10620__ = pi17 & ~new_new_n10619__;
  assign new_new_n10621__ = ~pi16 & new_new_n1823__;
  assign new_new_n10622__ = pi16 & ~new_new_n1823__;
  assign new_new_n10623__ = new_new_n6958__ & ~new_new_n10621__;
  assign new_new_n10624__ = ~new_new_n10622__ & new_new_n10623__;
  assign new_new_n10625__ = new_new_n5501__ & new_new_n10624__;
  assign new_new_n10626__ = ~new_new_n10620__ & ~new_new_n10625__;
  assign new_new_n10627__ = new_new_n10618__ & ~new_new_n10626__;
  assign new_new_n10628__ = new_new_n6553__ & new_new_n6958__;
  assign new_new_n10629__ = new_new_n10618__ & ~new_new_n10628__;
  assign new_new_n10630__ = ~pi17 & ~new_new_n10629__;
  assign new_new_n10631__ = ~new_new_n10627__ & ~new_new_n10630__;
  assign new_new_n10632__ = ~new_new_n10615__ & new_new_n10631__;
  assign new_new_n10633__ = new_new_n10200__ & new_new_n10204__;
  assign new_new_n10634__ = ~new_new_n10605__ & ~new_new_n10614__;
  assign new_new_n10635__ = ~new_new_n10633__ & ~new_new_n10634__;
  assign new_new_n10636__ = ~new_new_n10632__ & new_new_n10635__;
  assign new_new_n10637__ = ~new_new_n10205__ & ~new_new_n10636__;
  assign new_new_n10638__ = ~new_new_n10107__ & ~new_new_n10108__;
  assign new_new_n10639__ = new_new_n10112__ & new_new_n10638__;
  assign new_new_n10640__ = ~new_new_n10112__ & ~new_new_n10638__;
  assign new_new_n10641__ = ~new_new_n10639__ & ~new_new_n10640__;
  assign new_new_n10642__ = ~new_new_n10637__ & ~new_new_n10641__;
  assign new_new_n10643__ = new_new_n10637__ & new_new_n10641__;
  assign new_new_n10644__ = ~new_new_n1823__ & new_new_n6964__;
  assign new_new_n10645__ = ~new_new_n1902__ & new_new_n6968__;
  assign new_new_n10646__ = ~new_new_n1660__ & new_new_n7935__;
  assign new_new_n10647__ = ~new_new_n5274__ & new_new_n6959__;
  assign new_new_n10648__ = ~new_new_n10644__ & ~new_new_n10645__;
  assign new_new_n10649__ = ~new_new_n10646__ & new_new_n10648__;
  assign new_new_n10650__ = ~new_new_n10647__ & new_new_n10649__;
  assign new_new_n10651__ = pi17 & ~new_new_n10650__;
  assign new_new_n10652__ = ~pi17 & new_new_n10650__;
  assign new_new_n10653__ = ~new_new_n10651__ & ~new_new_n10652__;
  assign new_new_n10654__ = ~new_new_n10643__ & new_new_n10653__;
  assign new_new_n10655__ = ~new_new_n10642__ & ~new_new_n10654__;
  assign new_new_n10656__ = ~new_new_n10190__ & ~new_new_n10655__;
  assign new_new_n10657__ = ~new_new_n1660__ & new_new_n6968__;
  assign new_new_n10658__ = ~new_new_n1902__ & new_new_n6964__;
  assign new_new_n10659__ = ~new_new_n10657__ & ~new_new_n10658__;
  assign new_new_n10660__ = ~new_new_n1737__ & new_new_n6958__;
  assign new_new_n10661__ = new_new_n5688__ & new_new_n10660__;
  assign new_new_n10662__ = new_new_n10659__ & ~new_new_n10661__;
  assign new_new_n10663__ = pi17 & ~new_new_n10662__;
  assign new_new_n10664__ = new_new_n1737__ & ~new_new_n5688__;
  assign new_new_n10665__ = new_new_n6958__ & ~new_new_n10664__;
  assign new_new_n10666__ = pi17 & ~new_new_n10665__;
  assign new_new_n10667__ = ~pi16 & new_new_n1737__;
  assign new_new_n10668__ = pi16 & ~new_new_n5688__;
  assign new_new_n10669__ = new_new_n6958__ & ~new_new_n10667__;
  assign new_new_n10670__ = ~new_new_n10668__ & new_new_n10669__;
  assign new_new_n10671__ = new_new_n10659__ & ~new_new_n10670__;
  assign new_new_n10672__ = ~new_new_n10666__ & new_new_n10671__;
  assign new_new_n10673__ = ~new_new_n10663__ & ~new_new_n10672__;
  assign new_new_n10674__ = new_new_n10190__ & new_new_n10655__;
  assign new_new_n10675__ = new_new_n10673__ & ~new_new_n10674__;
  assign new_new_n10676__ = ~new_new_n10656__ & ~new_new_n10675__;
  assign new_new_n10677__ = ~new_new_n10186__ & new_new_n10676__;
  assign new_new_n10678__ = ~new_new_n10185__ & ~new_new_n10677__;
  assign new_new_n10679__ = new_new_n10162__ & new_new_n10678__;
  assign new_new_n10680__ = ~new_new_n10162__ & ~new_new_n10678__;
  assign new_new_n10681__ = ~new_new_n1207__ & ~new_new_n8479__;
  assign new_new_n10682__ = ~new_new_n3720__ & new_new_n8858__;
  assign new_new_n10683__ = ~new_new_n868__ & new_new_n8474__;
  assign new_new_n10684__ = ~new_new_n5927__ & new_new_n8470__;
  assign new_new_n10685__ = ~new_new_n10681__ & ~new_new_n10682__;
  assign new_new_n10686__ = ~new_new_n10683__ & new_new_n10685__;
  assign new_new_n10687__ = ~new_new_n10684__ & new_new_n10686__;
  assign new_new_n10688__ = ~pi11 & new_new_n10687__;
  assign new_new_n10689__ = pi11 & ~new_new_n10687__;
  assign new_new_n10690__ = ~new_new_n10688__ & ~new_new_n10689__;
  assign new_new_n10691__ = ~new_new_n10680__ & new_new_n10690__;
  assign new_new_n10692__ = ~new_new_n10679__ & ~new_new_n10691__;
  assign new_new_n10693__ = ~new_new_n10158__ & ~new_new_n10692__;
  assign new_new_n10694__ = ~new_new_n9697__ & ~new_new_n9701__;
  assign new_new_n10695__ = pi07 & ~pi08;
  assign new_new_n10696__ = ~pi07 & pi08;
  assign new_new_n10697__ = ~new_new_n10695__ & ~new_new_n10696__;
  assign new_new_n10698__ = new_new_n10694__ & new_new_n10697__;
  assign new_new_n10699__ = ~new_new_n3768__ & new_new_n10698__;
  assign new_new_n10700__ = pi07 & ~new_new_n9697__;
  assign new_new_n10701__ = ~pi07 & ~new_new_n9701__;
  assign new_new_n10702__ = ~new_new_n10700__ & ~new_new_n10701__;
  assign new_new_n10703__ = ~new_new_n583__ & new_new_n10702__;
  assign new_new_n10704__ = new_new_n4141__ & new_new_n10697__;
  assign new_new_n10705__ = new_new_n10694__ & ~new_new_n10704__;
  assign new_new_n10706__ = ~new_new_n4144__ & new_new_n10705__;
  assign new_new_n10707__ = ~new_new_n10699__ & ~new_new_n10703__;
  assign new_new_n10708__ = ~new_new_n10706__ & new_new_n10707__;
  assign new_new_n10709__ = ~pi06 & ~pi07;
  assign new_new_n10710__ = ~new_new_n691__ & new_new_n10709__;
  assign new_new_n10711__ = pi08 & ~new_new_n10710__;
  assign new_new_n10712__ = pi06 & pi07;
  assign new_new_n10713__ = ~new_new_n691__ & new_new_n10712__;
  assign new_new_n10714__ = ~pi08 & ~new_new_n10713__;
  assign new_new_n10715__ = pi05 & ~new_new_n10714__;
  assign new_new_n10716__ = ~new_new_n10711__ & ~new_new_n10715__;
  assign new_new_n10717__ = new_new_n10708__ & ~new_new_n10716__;
  assign new_new_n10718__ = ~pi08 & ~new_new_n10708__;
  assign new_new_n10719__ = ~new_new_n10717__ & ~new_new_n10718__;
  assign new_new_n10720__ = new_new_n10158__ & new_new_n10692__;
  assign new_new_n10721__ = ~new_new_n10693__ & ~new_new_n10720__;
  assign new_new_n10722__ = ~new_new_n10719__ & new_new_n10721__;
  assign new_new_n10723__ = ~new_new_n10693__ & ~new_new_n10722__;
  assign new_new_n10724__ = ~pi04 & ~new_new_n466__;
  assign new_new_n10725__ = pi05 & ~new_new_n10724__;
  assign new_new_n10726__ = ~pi02 & ~pi03;
  assign new_new_n10727__ = ~pi04 & ~pi05;
  assign new_new_n10728__ = ~new_new_n10726__ & ~new_new_n10727__;
  assign new_new_n10729__ = ~new_new_n466__ & new_new_n10728__;
  assign new_new_n10730__ = ~new_new_n10725__ & ~new_new_n10729__;
  assign new_new_n10731__ = pi02 & pi03;
  assign new_new_n10732__ = ~new_new_n4168__ & ~new_new_n10724__;
  assign new_new_n10733__ = pi05 & new_new_n4168__;
  assign new_new_n10734__ = ~new_new_n10731__ & ~new_new_n10732__;
  assign new_new_n10735__ = ~new_new_n10733__ & new_new_n10734__;
  assign new_new_n10736__ = ~new_new_n10730__ & ~new_new_n10735__;
  assign new_new_n10737__ = ~new_new_n10185__ & ~new_new_n10186__;
  assign new_new_n10738__ = new_new_n10676__ & new_new_n10737__;
  assign new_new_n10739__ = ~new_new_n10676__ & ~new_new_n10737__;
  assign new_new_n10740__ = ~new_new_n10738__ & ~new_new_n10739__;
  assign new_new_n10741__ = ~new_new_n1737__ & new_new_n6991__;
  assign new_new_n10742__ = ~new_new_n1466__ & new_new_n6985__;
  assign new_new_n10743__ = ~new_new_n10741__ & ~new_new_n10742__;
  assign new_new_n10744__ = ~new_new_n1556__ & new_new_n6994__;
  assign new_new_n10745__ = ~new_new_n5671__ & new_new_n10744__;
  assign new_new_n10746__ = new_new_n10743__ & ~new_new_n10745__;
  assign new_new_n10747__ = ~pi14 & ~new_new_n10746__;
  assign new_new_n10748__ = pi13 & ~new_new_n1556__;
  assign new_new_n10749__ = new_new_n1556__ & new_new_n5671__;
  assign new_new_n10750__ = new_new_n6994__ & ~new_new_n10749__;
  assign new_new_n10751__ = ~pi13 & ~new_new_n5671__;
  assign new_new_n10752__ = ~new_new_n10748__ & ~new_new_n10751__;
  assign new_new_n10753__ = new_new_n10750__ & new_new_n10752__;
  assign new_new_n10754__ = pi14 & new_new_n10743__;
  assign new_new_n10755__ = ~new_new_n10750__ & new_new_n10754__;
  assign new_new_n10756__ = ~new_new_n10747__ & ~new_new_n10753__;
  assign new_new_n10757__ = ~new_new_n10755__ & new_new_n10756__;
  assign new_new_n10758__ = ~new_new_n10642__ & ~new_new_n10643__;
  assign new_new_n10759__ = new_new_n10653__ & ~new_new_n10758__;
  assign new_new_n10760__ = ~new_new_n10653__ & new_new_n10758__;
  assign new_new_n10761__ = ~new_new_n10759__ & ~new_new_n10760__;
  assign new_new_n10762__ = new_new_n10757__ & new_new_n10761__;
  assign new_new_n10763__ = ~new_new_n10757__ & ~new_new_n10761__;
  assign new_new_n10764__ = ~new_new_n10227__ & ~new_new_n10228__;
  assign new_new_n10765__ = new_new_n10603__ & ~new_new_n10764__;
  assign new_new_n10766__ = ~new_new_n10603__ & new_new_n10764__;
  assign new_new_n10767__ = ~new_new_n10765__ & ~new_new_n10766__;
  assign new_new_n10768__ = ~new_new_n3535__ & new_new_n6991__;
  assign new_new_n10769__ = ~new_new_n1823__ & new_new_n6985__;
  assign new_new_n10770__ = ~pi13 & ~pi14;
  assign new_new_n10771__ = pi13 & pi14;
  assign new_new_n10772__ = ~new_new_n10770__ & ~new_new_n10771__;
  assign new_new_n10773__ = new_new_n6487__ & new_new_n10772__;
  assign new_new_n10774__ = new_new_n1902__ & ~new_new_n10772__;
  assign new_new_n10775__ = new_new_n6994__ & ~new_new_n10774__;
  assign new_new_n10776__ = ~new_new_n10773__ & new_new_n10775__;
  assign new_new_n10777__ = ~new_new_n10768__ & ~new_new_n10769__;
  assign new_new_n10778__ = ~new_new_n10776__ & new_new_n10777__;
  assign new_new_n10779__ = pi14 & ~new_new_n10778__;
  assign new_new_n10780__ = ~pi14 & new_new_n10778__;
  assign new_new_n10781__ = ~new_new_n10779__ & ~new_new_n10780__;
  assign new_new_n10782__ = new_new_n10232__ & ~new_new_n10545__;
  assign new_new_n10783__ = new_new_n10236__ & ~new_new_n10782__;
  assign new_new_n10784__ = ~new_new_n10232__ & new_new_n10545__;
  assign new_new_n10785__ = ~new_new_n10236__ & ~new_new_n10784__;
  assign new_new_n10786__ = pi17 & new_new_n10253__;
  assign new_new_n10787__ = ~new_new_n10550__ & ~new_new_n10786__;
  assign new_new_n10788__ = ~new_new_n10783__ & ~new_new_n10787__;
  assign new_new_n10789__ = ~new_new_n10785__ & new_new_n10788__;
  assign new_new_n10790__ = ~new_new_n10782__ & ~new_new_n10784__;
  assign new_new_n10791__ = ~new_new_n10244__ & ~new_new_n10255__;
  assign new_new_n10792__ = ~new_new_n10253__ & ~new_new_n10791__;
  assign new_new_n10793__ = new_new_n10253__ & new_new_n10791__;
  assign new_new_n10794__ = new_new_n10790__ & ~new_new_n10792__;
  assign new_new_n10795__ = ~new_new_n10793__ & new_new_n10794__;
  assign new_new_n10796__ = ~new_new_n10236__ & ~new_new_n10782__;
  assign new_new_n10797__ = new_new_n10236__ & ~new_new_n10784__;
  assign new_new_n10798__ = new_new_n10787__ & ~new_new_n10796__;
  assign new_new_n10799__ = ~new_new_n10797__ & new_new_n10798__;
  assign new_new_n10800__ = ~new_new_n10789__ & ~new_new_n10799__;
  assign new_new_n10801__ = ~new_new_n10795__ & new_new_n10800__;
  assign new_new_n10802__ = ~new_new_n2024__ & new_new_n6991__;
  assign new_new_n10803__ = ~new_new_n2130__ & new_new_n6985__;
  assign new_new_n10804__ = ~new_new_n10802__ & ~new_new_n10803__;
  assign new_new_n10805__ = new_new_n6994__ & new_new_n10209__;
  assign new_new_n10806__ = new_new_n10804__ & ~new_new_n10805__;
  assign new_new_n10807__ = pi14 & ~new_new_n10806__;
  assign new_new_n10808__ = ~pi13 & ~new_new_n10215__;
  assign new_new_n10809__ = pi13 & ~new_new_n6853__;
  assign new_new_n10810__ = new_new_n6994__ & ~new_new_n10808__;
  assign new_new_n10811__ = ~new_new_n10809__ & new_new_n10810__;
  assign new_new_n10812__ = ~new_new_n6850__ & new_new_n6994__;
  assign new_new_n10813__ = ~pi14 & new_new_n10804__;
  assign new_new_n10814__ = ~new_new_n10812__ & new_new_n10813__;
  assign new_new_n10815__ = ~new_new_n10811__ & ~new_new_n10814__;
  assign new_new_n10816__ = ~new_new_n10807__ & new_new_n10815__;
  assign new_new_n10817__ = ~new_new_n2420__ & new_new_n6991__;
  assign new_new_n10818__ = ~new_new_n2224__ & new_new_n6985__;
  assign new_new_n10819__ = ~new_new_n10817__ & ~new_new_n10818__;
  assign new_new_n10820__ = ~new_new_n2024__ & new_new_n6994__;
  assign new_new_n10821__ = new_new_n7313__ & new_new_n10820__;
  assign new_new_n10822__ = new_new_n10819__ & ~new_new_n10821__;
  assign new_new_n10823__ = pi14 & ~new_new_n10822__;
  assign new_new_n10824__ = pi13 & new_new_n7313__;
  assign new_new_n10825__ = new_new_n2024__ & ~new_new_n7313__;
  assign new_new_n10826__ = new_new_n6994__ & ~new_new_n10825__;
  assign new_new_n10827__ = ~pi13 & ~new_new_n2024__;
  assign new_new_n10828__ = ~new_new_n10824__ & ~new_new_n10827__;
  assign new_new_n10829__ = new_new_n10826__ & new_new_n10828__;
  assign new_new_n10830__ = ~pi14 & new_new_n10819__;
  assign new_new_n10831__ = ~new_new_n10826__ & new_new_n10830__;
  assign new_new_n10832__ = ~new_new_n10823__ & ~new_new_n10829__;
  assign new_new_n10833__ = ~new_new_n10831__ & new_new_n10832__;
  assign new_new_n10834__ = new_new_n6750__ & new_new_n8820__;
  assign new_new_n10835__ = ~new_new_n2572__ & new_new_n6991__;
  assign new_new_n10836__ = ~new_new_n2313__ & new_new_n6985__;
  assign new_new_n10837__ = ~new_new_n10835__ & ~new_new_n10836__;
  assign new_new_n10838__ = new_new_n6994__ & ~new_new_n9267__;
  assign new_new_n10839__ = pi14 & ~new_new_n10838__;
  assign new_new_n10840__ = ~new_new_n2420__ & new_new_n8388__;
  assign new_new_n10841__ = new_new_n6748__ & new_new_n10840__;
  assign new_new_n10842__ = ~new_new_n10839__ & ~new_new_n10841__;
  assign new_new_n10843__ = new_new_n10837__ & ~new_new_n10842__;
  assign new_new_n10844__ = new_new_n6749__ & new_new_n6994__;
  assign new_new_n10845__ = new_new_n10837__ & ~new_new_n10844__;
  assign new_new_n10846__ = ~pi14 & ~new_new_n10845__;
  assign new_new_n10847__ = ~new_new_n10834__ & ~new_new_n10846__;
  assign new_new_n10848__ = ~new_new_n10843__ & new_new_n10847__;
  assign new_new_n10849__ = ~new_new_n10511__ & ~new_new_n10512__;
  assign new_new_n10850__ = ~new_new_n10516__ & new_new_n10849__;
  assign new_new_n10851__ = new_new_n10516__ & ~new_new_n10849__;
  assign new_new_n10852__ = ~new_new_n10850__ & ~new_new_n10851__;
  assign new_new_n10853__ = ~new_new_n10848__ & new_new_n10852__;
  assign new_new_n10854__ = ~new_new_n2572__ & new_new_n6985__;
  assign new_new_n10855__ = ~new_new_n2497__ & new_new_n6991__;
  assign new_new_n10856__ = ~new_new_n10854__ & ~new_new_n10855__;
  assign new_new_n10857__ = ~new_new_n2313__ & new_new_n6994__;
  assign new_new_n10858__ = ~new_new_n7236__ & new_new_n10857__;
  assign new_new_n10859__ = new_new_n10856__ & ~new_new_n10858__;
  assign new_new_n10860__ = ~pi14 & ~new_new_n10859__;
  assign new_new_n10861__ = pi13 & ~new_new_n2313__;
  assign new_new_n10862__ = new_new_n2313__ & new_new_n7236__;
  assign new_new_n10863__ = new_new_n6994__ & ~new_new_n10862__;
  assign new_new_n10864__ = ~pi13 & ~new_new_n7236__;
  assign new_new_n10865__ = ~new_new_n10861__ & ~new_new_n10864__;
  assign new_new_n10866__ = new_new_n10863__ & new_new_n10865__;
  assign new_new_n10867__ = pi14 & new_new_n10856__;
  assign new_new_n10868__ = ~new_new_n10863__ & new_new_n10867__;
  assign new_new_n10869__ = ~new_new_n10860__ & ~new_new_n10866__;
  assign new_new_n10870__ = ~new_new_n10868__ & new_new_n10869__;
  assign new_new_n10871__ = ~new_new_n2636__ & new_new_n6991__;
  assign new_new_n10872__ = ~new_new_n2497__ & new_new_n6985__;
  assign new_new_n10873__ = ~new_new_n10871__ & ~new_new_n10872__;
  assign new_new_n10874__ = ~new_new_n2572__ & ~new_new_n6801__;
  assign new_new_n10875__ = new_new_n6994__ & new_new_n10874__;
  assign new_new_n10876__ = new_new_n10873__ & ~new_new_n10875__;
  assign new_new_n10877__ = pi14 & ~new_new_n10876__;
  assign new_new_n10878__ = pi13 & new_new_n2572__;
  assign new_new_n10879__ = ~pi13 & ~new_new_n2572__;
  assign new_new_n10880__ = new_new_n6994__ & ~new_new_n10878__;
  assign new_new_n10881__ = ~new_new_n10879__ & new_new_n10880__;
  assign new_new_n10882__ = new_new_n6801__ & new_new_n10881__;
  assign new_new_n10883__ = ~new_new_n6802__ & new_new_n6994__;
  assign new_new_n10884__ = ~pi14 & new_new_n10873__;
  assign new_new_n10885__ = ~new_new_n10883__ & new_new_n10884__;
  assign new_new_n10886__ = ~new_new_n10882__ & ~new_new_n10885__;
  assign new_new_n10887__ = ~new_new_n10877__ & new_new_n10886__;
  assign new_new_n10888__ = ~new_new_n10474__ & ~new_new_n10475__;
  assign new_new_n10889__ = ~new_new_n10479__ & new_new_n10888__;
  assign new_new_n10890__ = new_new_n10479__ & ~new_new_n10888__;
  assign new_new_n10891__ = ~new_new_n10889__ & ~new_new_n10890__;
  assign new_new_n10892__ = new_new_n10887__ & new_new_n10891__;
  assign new_new_n10893__ = ~new_new_n10887__ & ~new_new_n10891__;
  assign new_new_n10894__ = ~new_new_n10460__ & ~new_new_n10461__;
  assign new_new_n10895__ = new_new_n10471__ & new_new_n10894__;
  assign new_new_n10896__ = ~new_new_n10471__ & ~new_new_n10894__;
  assign new_new_n10897__ = ~new_new_n10895__ & ~new_new_n10896__;
  assign new_new_n10898__ = new_new_n6958__ & ~new_new_n7065__;
  assign new_new_n10899__ = pi17 & new_new_n10445__;
  assign new_new_n10900__ = ~pi17 & ~new_new_n10445__;
  assign new_new_n10901__ = ~new_new_n10899__ & ~new_new_n10900__;
  assign new_new_n10902__ = ~new_new_n10898__ & ~new_new_n10901__;
  assign new_new_n10903__ = pi16 & new_new_n10445__;
  assign new_new_n10904__ = ~pi16 & ~new_new_n10445__;
  assign new_new_n10905__ = ~new_new_n10903__ & ~new_new_n10904__;
  assign new_new_n10906__ = new_new_n10898__ & ~new_new_n10905__;
  assign new_new_n10907__ = ~new_new_n10902__ & ~new_new_n10906__;
  assign new_new_n10908__ = new_new_n10452__ & ~new_new_n10907__;
  assign new_new_n10909__ = ~new_new_n10452__ & new_new_n10901__;
  assign new_new_n10910__ = ~new_new_n10908__ & ~new_new_n10909__;
  assign new_new_n10911__ = ~new_new_n10441__ & new_new_n10910__;
  assign new_new_n10912__ = new_new_n10441__ & ~new_new_n10910__;
  assign new_new_n10913__ = ~new_new_n10911__ & ~new_new_n10912__;
  assign new_new_n10914__ = ~new_new_n2886__ & new_new_n6985__;
  assign new_new_n10915__ = ~new_new_n2848__ & new_new_n6991__;
  assign new_new_n10916__ = ~new_new_n10914__ & ~new_new_n10915__;
  assign new_new_n10917__ = ~new_new_n2737__ & new_new_n6994__;
  assign new_new_n10918__ = ~new_new_n7378__ & new_new_n10917__;
  assign new_new_n10919__ = new_new_n10916__ & ~new_new_n10918__;
  assign new_new_n10920__ = pi14 & ~new_new_n10919__;
  assign new_new_n10921__ = ~pi13 & ~new_new_n2737__;
  assign new_new_n10922__ = new_new_n2737__ & new_new_n7378__;
  assign new_new_n10923__ = new_new_n6994__ & ~new_new_n10922__;
  assign new_new_n10924__ = pi13 & ~new_new_n7378__;
  assign new_new_n10925__ = ~new_new_n10921__ & ~new_new_n10924__;
  assign new_new_n10926__ = new_new_n10923__ & new_new_n10925__;
  assign new_new_n10927__ = ~pi14 & new_new_n10916__;
  assign new_new_n10928__ = ~new_new_n10923__ & new_new_n10927__;
  assign new_new_n10929__ = ~new_new_n10920__ & ~new_new_n10926__;
  assign new_new_n10930__ = ~new_new_n10928__ & new_new_n10929__;
  assign new_new_n10931__ = ~new_new_n10346__ & new_new_n10433__;
  assign new_new_n10932__ = new_new_n9930__ & ~new_new_n10347__;
  assign new_new_n10933__ = new_new_n10931__ & new_new_n10932__;
  assign new_new_n10934__ = new_new_n10346__ & ~new_new_n10433__;
  assign new_new_n10935__ = ~new_new_n10931__ & ~new_new_n10934__;
  assign new_new_n10936__ = ~new_new_n10439__ & ~new_new_n10932__;
  assign new_new_n10937__ = new_new_n10935__ & new_new_n10936__;
  assign new_new_n10938__ = ~new_new_n9919__ & new_new_n9930__;
  assign new_new_n10939__ = ~new_new_n10438__ & ~new_new_n10938__;
  assign new_new_n10940__ = ~new_new_n10935__ & new_new_n10939__;
  assign new_new_n10941__ = ~new_new_n10933__ & ~new_new_n10937__;
  assign new_new_n10942__ = ~new_new_n10940__ & new_new_n10941__;
  assign new_new_n10943__ = ~new_new_n10930__ & ~new_new_n10942__;
  assign new_new_n10944__ = new_new_n10930__ & new_new_n10942__;
  assign new_new_n10945__ = ~new_new_n2960__ & new_new_n6991__;
  assign new_new_n10946__ = ~new_new_n3460__ & new_new_n6985__;
  assign new_new_n10947__ = ~new_new_n10945__ & ~new_new_n10946__;
  assign new_new_n10948__ = ~new_new_n2848__ & new_new_n6994__;
  assign new_new_n10949__ = ~new_new_n7065__ & new_new_n10948__;
  assign new_new_n10950__ = new_new_n10947__ & ~new_new_n10949__;
  assign new_new_n10951__ = ~pi14 & ~new_new_n10950__;
  assign new_new_n10952__ = new_new_n2848__ & new_new_n7065__;
  assign new_new_n10953__ = new_new_n6994__ & ~new_new_n10952__;
  assign new_new_n10954__ = pi14 & new_new_n10947__;
  assign new_new_n10955__ = ~new_new_n10953__ & new_new_n10954__;
  assign new_new_n10956__ = ~pi13 & ~new_new_n8566__;
  assign new_new_n10957__ = pi13 & ~new_new_n7067__;
  assign new_new_n10958__ = new_new_n6994__ & ~new_new_n10956__;
  assign new_new_n10959__ = ~new_new_n10957__ & new_new_n10958__;
  assign new_new_n10960__ = ~new_new_n10951__ & ~new_new_n10955__;
  assign new_new_n10961__ = ~new_new_n10959__ & new_new_n10960__;
  assign new_new_n10962__ = ~new_new_n10368__ & new_new_n10394__;
  assign new_new_n10963__ = new_new_n10368__ & ~new_new_n10394__;
  assign new_new_n10964__ = ~new_new_n10962__ & ~new_new_n10963__;
  assign new_new_n10965__ = ~new_new_n10417__ & new_new_n10964__;
  assign new_new_n10966__ = ~new_new_n10415__ & ~new_new_n10417__;
  assign new_new_n10967__ = ~new_new_n10418__ & ~new_new_n10964__;
  assign new_new_n10968__ = ~new_new_n10966__ & new_new_n10967__;
  assign new_new_n10969__ = ~new_new_n10965__ & ~new_new_n10968__;
  assign new_new_n10970__ = ~new_new_n10961__ & ~new_new_n10969__;
  assign new_new_n10971__ = new_new_n10961__ & new_new_n10969__;
  assign new_new_n10972__ = new_new_n10380__ & ~new_new_n10415__;
  assign new_new_n10973__ = ~new_new_n10416__ & ~new_new_n10972__;
  assign new_new_n10974__ = ~new_new_n10381__ & ~new_new_n10973__;
  assign new_new_n10975__ = new_new_n10382__ & ~new_new_n10415__;
  assign new_new_n10976__ = ~new_new_n10974__ & ~new_new_n10975__;
  assign new_new_n10977__ = ~new_new_n10406__ & new_new_n10413__;
  assign new_new_n10978__ = ~new_new_n10414__ & ~new_new_n10977__;
  assign new_new_n10979__ = ~new_new_n3126__ & new_new_n6985__;
  assign new_new_n10980__ = ~new_new_n3164__ & new_new_n6991__;
  assign new_new_n10981__ = ~new_new_n10979__ & ~new_new_n10980__;
  assign new_new_n10982__ = ~new_new_n2960__ & new_new_n6994__;
  assign new_new_n10983__ = ~new_new_n7468__ & new_new_n10982__;
  assign new_new_n10984__ = new_new_n10981__ & ~new_new_n10983__;
  assign new_new_n10985__ = pi14 & ~new_new_n10984__;
  assign new_new_n10986__ = ~pi13 & ~new_new_n2960__;
  assign new_new_n10987__ = new_new_n2960__ & new_new_n7468__;
  assign new_new_n10988__ = new_new_n6994__ & ~new_new_n10987__;
  assign new_new_n10989__ = pi13 & ~new_new_n7468__;
  assign new_new_n10990__ = ~new_new_n10986__ & ~new_new_n10989__;
  assign new_new_n10991__ = new_new_n10988__ & new_new_n10990__;
  assign new_new_n10992__ = ~pi14 & new_new_n10981__;
  assign new_new_n10993__ = ~new_new_n10988__ & new_new_n10992__;
  assign new_new_n10994__ = ~new_new_n10985__ & ~new_new_n10991__;
  assign new_new_n10995__ = ~new_new_n10993__ & new_new_n10994__;
  assign new_new_n10996__ = new_new_n10978__ & new_new_n10995__;
  assign new_new_n10997__ = ~new_new_n10978__ & ~new_new_n10995__;
  assign new_new_n10998__ = ~new_new_n6987__ & ~new_new_n6989__;
  assign new_new_n10999__ = ~new_new_n3055__ & ~new_new_n6981__;
  assign new_new_n11000__ = ~new_new_n6983__ & new_new_n10999__;
  assign new_new_n11001__ = new_new_n3356__ & ~new_new_n11000__;
  assign new_new_n11002__ = new_new_n10998__ & ~new_new_n11001__;
  assign new_new_n11003__ = pi14 & ~new_new_n11002__;
  assign new_new_n11004__ = ~new_new_n3356__ & new_new_n6991__;
  assign new_new_n11005__ = ~new_new_n3055__ & new_new_n6985__;
  assign new_new_n11006__ = new_new_n8610__ & new_new_n10772__;
  assign new_new_n11007__ = new_new_n3254__ & ~new_new_n11006__;
  assign new_new_n11008__ = ~new_new_n3254__ & new_new_n11006__;
  assign new_new_n11009__ = new_new_n6994__ & ~new_new_n11007__;
  assign new_new_n11010__ = ~new_new_n11008__ & new_new_n11009__;
  assign new_new_n11011__ = ~new_new_n11004__ & ~new_new_n11005__;
  assign new_new_n11012__ = ~new_new_n11010__ & new_new_n11011__;
  assign new_new_n11013__ = new_new_n11003__ & new_new_n11012__;
  assign new_new_n11014__ = ~new_new_n3356__ & new_new_n6958__;
  assign new_new_n11015__ = ~new_new_n11013__ & ~new_new_n11014__;
  assign new_new_n11016__ = ~new_new_n3254__ & new_new_n6985__;
  assign new_new_n11017__ = ~new_new_n3055__ & new_new_n6991__;
  assign new_new_n11018__ = ~new_new_n11016__ & ~new_new_n11017__;
  assign new_new_n11019__ = ~new_new_n3164__ & new_new_n6994__;
  assign new_new_n11020__ = ~new_new_n8637__ & new_new_n11019__;
  assign new_new_n11021__ = new_new_n11018__ & ~new_new_n11020__;
  assign new_new_n11022__ = ~pi14 & ~new_new_n11021__;
  assign new_new_n11023__ = pi13 & ~new_new_n3164__;
  assign new_new_n11024__ = new_new_n3164__ & new_new_n8637__;
  assign new_new_n11025__ = new_new_n6994__ & ~new_new_n11024__;
  assign new_new_n11026__ = ~pi13 & ~new_new_n8637__;
  assign new_new_n11027__ = ~new_new_n11023__ & ~new_new_n11026__;
  assign new_new_n11028__ = new_new_n11025__ & new_new_n11027__;
  assign new_new_n11029__ = pi14 & new_new_n11018__;
  assign new_new_n11030__ = ~new_new_n11025__ & new_new_n11029__;
  assign new_new_n11031__ = ~new_new_n11022__ & ~new_new_n11028__;
  assign new_new_n11032__ = ~new_new_n11030__ & new_new_n11031__;
  assign new_new_n11033__ = ~new_new_n11015__ & ~new_new_n11032__;
  assign new_new_n11034__ = ~new_new_n3254__ & new_new_n6991__;
  assign new_new_n11035__ = ~new_new_n3164__ & new_new_n6985__;
  assign new_new_n11036__ = ~new_new_n11034__ & ~new_new_n11035__;
  assign new_new_n11037__ = ~new_new_n3126__ & new_new_n6994__;
  assign new_new_n11038__ = ~new_new_n7570__ & new_new_n11037__;
  assign new_new_n11039__ = new_new_n11036__ & ~new_new_n11038__;
  assign new_new_n11040__ = ~pi14 & ~new_new_n11039__;
  assign new_new_n11041__ = pi13 & ~new_new_n3126__;
  assign new_new_n11042__ = new_new_n3126__ & new_new_n7570__;
  assign new_new_n11043__ = new_new_n6994__ & ~new_new_n11042__;
  assign new_new_n11044__ = ~pi13 & ~new_new_n7570__;
  assign new_new_n11045__ = ~new_new_n11041__ & ~new_new_n11044__;
  assign new_new_n11046__ = new_new_n11043__ & new_new_n11045__;
  assign new_new_n11047__ = pi14 & new_new_n11036__;
  assign new_new_n11048__ = ~new_new_n11043__ & new_new_n11047__;
  assign new_new_n11049__ = ~new_new_n11040__ & ~new_new_n11046__;
  assign new_new_n11050__ = ~new_new_n11048__ & new_new_n11049__;
  assign new_new_n11051__ = new_new_n11033__ & ~new_new_n11050__;
  assign new_new_n11052__ = ~new_new_n11033__ & new_new_n11050__;
  assign new_new_n11053__ = ~new_new_n3356__ & new_new_n10409__;
  assign new_new_n11054__ = ~new_new_n6957__ & ~new_new_n11053__;
  assign new_new_n11055__ = pi16 & ~new_new_n11054__;
  assign new_new_n11056__ = ~new_new_n3356__ & ~new_new_n6967__;
  assign new_new_n11057__ = ~new_new_n3055__ & new_new_n6958__;
  assign new_new_n11058__ = ~new_new_n11056__ & ~new_new_n11057__;
  assign new_new_n11059__ = ~new_new_n11055__ & ~new_new_n11058__;
  assign new_new_n11060__ = ~new_new_n11052__ & new_new_n11059__;
  assign new_new_n11061__ = ~new_new_n11051__ & ~new_new_n11060__;
  assign new_new_n11062__ = ~new_new_n10997__ & ~new_new_n11061__;
  assign new_new_n11063__ = ~new_new_n10996__ & ~new_new_n11062__;
  assign new_new_n11064__ = new_new_n10976__ & ~new_new_n11063__;
  assign new_new_n11065__ = ~new_new_n10976__ & new_new_n11063__;
  assign new_new_n11066__ = ~new_new_n2960__ & new_new_n6985__;
  assign new_new_n11067__ = ~new_new_n3126__ & new_new_n6991__;
  assign new_new_n11068__ = ~new_new_n11066__ & ~new_new_n11067__;
  assign new_new_n11069__ = ~new_new_n3460__ & new_new_n6994__;
  assign new_new_n11070__ = new_new_n7388__ & new_new_n11069__;
  assign new_new_n11071__ = new_new_n11068__ & ~new_new_n11070__;
  assign new_new_n11072__ = pi14 & ~new_new_n11071__;
  assign new_new_n11073__ = new_new_n6994__ & ~new_new_n7389__;
  assign new_new_n11074__ = ~pi14 & new_new_n11068__;
  assign new_new_n11075__ = ~new_new_n11073__ & new_new_n11074__;
  assign new_new_n11076__ = new_new_n3460__ & ~new_new_n7388__;
  assign new_new_n11077__ = ~pi13 & ~new_new_n11076__;
  assign new_new_n11078__ = pi13 & ~new_new_n7390__;
  assign new_new_n11079__ = new_new_n6994__ & ~new_new_n11077__;
  assign new_new_n11080__ = ~new_new_n11078__ & new_new_n11079__;
  assign new_new_n11081__ = ~new_new_n11072__ & ~new_new_n11075__;
  assign new_new_n11082__ = ~new_new_n11080__ & new_new_n11081__;
  assign new_new_n11083__ = ~new_new_n11065__ & new_new_n11082__;
  assign new_new_n11084__ = ~new_new_n11064__ & ~new_new_n11083__;
  assign new_new_n11085__ = ~new_new_n10971__ & ~new_new_n11084__;
  assign new_new_n11086__ = ~new_new_n10970__ & ~new_new_n11085__;
  assign new_new_n11087__ = ~new_new_n10420__ & ~new_new_n10421__;
  assign new_new_n11088__ = ~new_new_n10431__ & ~new_new_n11087__;
  assign new_new_n11089__ = new_new_n10431__ & new_new_n11087__;
  assign new_new_n11090__ = ~new_new_n11088__ & ~new_new_n11089__;
  assign new_new_n11091__ = new_new_n11086__ & ~new_new_n11090__;
  assign new_new_n11092__ = ~new_new_n11086__ & new_new_n11090__;
  assign new_new_n11093__ = ~new_new_n3460__ & new_new_n6991__;
  assign new_new_n11094__ = ~new_new_n2848__ & new_new_n6985__;
  assign new_new_n11095__ = ~new_new_n11093__ & ~new_new_n11094__;
  assign new_new_n11096__ = ~new_new_n2886__ & new_new_n6994__;
  assign new_new_n11097__ = ~new_new_n8574__ & new_new_n11096__;
  assign new_new_n11098__ = new_new_n11095__ & ~new_new_n11097__;
  assign new_new_n11099__ = ~pi14 & ~new_new_n11098__;
  assign new_new_n11100__ = pi13 & ~new_new_n2886__;
  assign new_new_n11101__ = new_new_n2886__ & new_new_n8574__;
  assign new_new_n11102__ = new_new_n6994__ & ~new_new_n11101__;
  assign new_new_n11103__ = ~pi13 & ~new_new_n8574__;
  assign new_new_n11104__ = ~new_new_n11100__ & ~new_new_n11103__;
  assign new_new_n11105__ = new_new_n11102__ & new_new_n11104__;
  assign new_new_n11106__ = pi14 & new_new_n11095__;
  assign new_new_n11107__ = ~new_new_n11102__ & new_new_n11106__;
  assign new_new_n11108__ = ~new_new_n11099__ & ~new_new_n11105__;
  assign new_new_n11109__ = ~new_new_n11107__ & new_new_n11108__;
  assign new_new_n11110__ = ~new_new_n11092__ & new_new_n11109__;
  assign new_new_n11111__ = ~new_new_n11091__ & ~new_new_n11110__;
  assign new_new_n11112__ = ~new_new_n10944__ & ~new_new_n11111__;
  assign new_new_n11113__ = ~new_new_n10943__ & ~new_new_n11112__;
  assign new_new_n11114__ = new_new_n10913__ & new_new_n11113__;
  assign new_new_n11115__ = ~new_new_n10913__ & ~new_new_n11113__;
  assign new_new_n11116__ = ~new_new_n2737__ & new_new_n6985__;
  assign new_new_n11117__ = new_new_n7814__ & new_new_n10772__;
  assign new_new_n11118__ = new_new_n2636__ & ~new_new_n10772__;
  assign new_new_n11119__ = new_new_n6994__ & ~new_new_n11118__;
  assign new_new_n11120__ = ~new_new_n11117__ & new_new_n11119__;
  assign new_new_n11121__ = ~new_new_n11116__ & ~new_new_n11120__;
  assign new_new_n11122__ = new_new_n2886__ & ~new_new_n6985__;
  assign new_new_n11123__ = new_new_n6991__ & ~new_new_n11122__;
  assign new_new_n11124__ = new_new_n11121__ & ~new_new_n11123__;
  assign new_new_n11125__ = ~pi14 & ~new_new_n11124__;
  assign new_new_n11126__ = ~new_new_n2886__ & new_new_n6991__;
  assign new_new_n11127__ = new_new_n11121__ & ~new_new_n11126__;
  assign new_new_n11128__ = pi14 & new_new_n11127__;
  assign new_new_n11129__ = ~new_new_n11125__ & ~new_new_n11128__;
  assign new_new_n11130__ = ~new_new_n11115__ & ~new_new_n11129__;
  assign new_new_n11131__ = ~new_new_n11114__ & ~new_new_n11130__;
  assign new_new_n11132__ = new_new_n10897__ & ~new_new_n11131__;
  assign new_new_n11133__ = ~new_new_n10897__ & new_new_n11131__;
  assign new_new_n11134__ = new_new_n7773__ & new_new_n8388__;
  assign new_new_n11135__ = ~new_new_n2636__ & new_new_n6985__;
  assign new_new_n11136__ = ~new_new_n2737__ & new_new_n6991__;
  assign new_new_n11137__ = ~new_new_n11135__ & ~new_new_n11136__;
  assign new_new_n11138__ = new_new_n6994__ & ~new_new_n9126__;
  assign new_new_n11139__ = ~pi14 & ~new_new_n11138__;
  assign new_new_n11140__ = ~new_new_n2497__ & new_new_n8820__;
  assign new_new_n11141__ = ~new_new_n6797__ & new_new_n11140__;
  assign new_new_n11142__ = ~new_new_n11139__ & ~new_new_n11141__;
  assign new_new_n11143__ = new_new_n11137__ & ~new_new_n11142__;
  assign new_new_n11144__ = new_new_n6994__ & new_new_n7772__;
  assign new_new_n11145__ = new_new_n11137__ & ~new_new_n11144__;
  assign new_new_n11146__ = pi14 & ~new_new_n11145__;
  assign new_new_n11147__ = ~new_new_n11134__ & ~new_new_n11146__;
  assign new_new_n11148__ = ~new_new_n11143__ & new_new_n11147__;
  assign new_new_n11149__ = ~new_new_n11133__ & new_new_n11148__;
  assign new_new_n11150__ = ~new_new_n11132__ & ~new_new_n11149__;
  assign new_new_n11151__ = ~new_new_n10893__ & ~new_new_n11150__;
  assign new_new_n11152__ = ~new_new_n10892__ & ~new_new_n11151__;
  assign new_new_n11153__ = new_new_n10870__ & new_new_n11152__;
  assign new_new_n11154__ = ~new_new_n10870__ & ~new_new_n11152__;
  assign new_new_n11155__ = ~new_new_n10486__ & ~new_new_n10487__;
  assign new_new_n11156__ = new_new_n10508__ & ~new_new_n11155__;
  assign new_new_n11157__ = ~new_new_n10508__ & new_new_n11155__;
  assign new_new_n11158__ = ~new_new_n11156__ & ~new_new_n11157__;
  assign new_new_n11159__ = ~new_new_n11154__ & new_new_n11158__;
  assign new_new_n11160__ = ~new_new_n11153__ & ~new_new_n11159__;
  assign new_new_n11161__ = new_new_n10848__ & ~new_new_n10852__;
  assign new_new_n11162__ = ~new_new_n10853__ & ~new_new_n11161__;
  assign new_new_n11163__ = new_new_n11160__ & new_new_n11162__;
  assign new_new_n11164__ = ~new_new_n10853__ & ~new_new_n11163__;
  assign new_new_n11165__ = ~new_new_n10294__ & ~new_new_n10295__;
  assign new_new_n11166__ = new_new_n10518__ & ~new_new_n11165__;
  assign new_new_n11167__ = ~new_new_n10518__ & new_new_n11165__;
  assign new_new_n11168__ = ~new_new_n11166__ & ~new_new_n11167__;
  assign new_new_n11169__ = new_new_n11164__ & ~new_new_n11168__;
  assign new_new_n11170__ = ~new_new_n11164__ & new_new_n11168__;
  assign new_new_n11171__ = new_new_n2224__ & ~new_new_n10772__;
  assign new_new_n11172__ = ~new_new_n6521__ & new_new_n10772__;
  assign new_new_n11173__ = new_new_n6994__ & ~new_new_n11171__;
  assign new_new_n11174__ = ~new_new_n11172__ & new_new_n11173__;
  assign new_new_n11175__ = ~new_new_n2420__ & new_new_n6985__;
  assign new_new_n11176__ = ~new_new_n2313__ & new_new_n6991__;
  assign new_new_n11177__ = ~new_new_n11175__ & ~new_new_n11176__;
  assign new_new_n11178__ = ~new_new_n11174__ & new_new_n11177__;
  assign new_new_n11179__ = pi14 & ~new_new_n11178__;
  assign new_new_n11180__ = ~new_new_n6991__ & ~new_new_n11175__;
  assign new_new_n11181__ = pi13 & new_new_n6981__;
  assign new_new_n11182__ = ~pi13 & new_new_n6983__;
  assign new_new_n11183__ = ~new_new_n11181__ & ~new_new_n11182__;
  assign new_new_n11184__ = new_new_n2313__ & new_new_n11183__;
  assign new_new_n11185__ = ~new_new_n11180__ & ~new_new_n11184__;
  assign new_new_n11186__ = ~pi14 & ~new_new_n11185__;
  assign new_new_n11187__ = ~new_new_n11174__ & new_new_n11186__;
  assign new_new_n11188__ = ~new_new_n11179__ & ~new_new_n11187__;
  assign new_new_n11189__ = ~new_new_n11170__ & ~new_new_n11188__;
  assign new_new_n11190__ = ~new_new_n11169__ & ~new_new_n11189__;
  assign new_new_n11191__ = ~new_new_n10833__ & ~new_new_n11190__;
  assign new_new_n11192__ = new_new_n10833__ & new_new_n11190__;
  assign new_new_n11193__ = ~new_new_n10528__ & ~new_new_n10529__;
  assign new_new_n11194__ = ~new_new_n10541__ & new_new_n11193__;
  assign new_new_n11195__ = new_new_n10541__ & ~new_new_n11193__;
  assign new_new_n11196__ = ~new_new_n11194__ & ~new_new_n11195__;
  assign new_new_n11197__ = ~new_new_n11192__ & new_new_n11196__;
  assign new_new_n11198__ = ~new_new_n11191__ & ~new_new_n11197__;
  assign new_new_n11199__ = ~new_new_n10276__ & ~new_new_n10277__;
  assign new_new_n11200__ = ~new_new_n10543__ & new_new_n11199__;
  assign new_new_n11201__ = new_new_n10543__ & ~new_new_n11199__;
  assign new_new_n11202__ = ~new_new_n11200__ & ~new_new_n11201__;
  assign new_new_n11203__ = new_new_n11198__ & new_new_n11202__;
  assign new_new_n11204__ = ~new_new_n11198__ & ~new_new_n11202__;
  assign new_new_n11205__ = ~new_new_n2024__ & new_new_n6985__;
  assign new_new_n11206__ = ~new_new_n2224__ & new_new_n6991__;
  assign new_new_n11207__ = ~new_new_n11205__ & ~new_new_n11206__;
  assign new_new_n11208__ = new_new_n6994__ & new_new_n9173__;
  assign new_new_n11209__ = new_new_n11207__ & ~new_new_n11208__;
  assign new_new_n11210__ = pi14 & ~new_new_n11209__;
  assign new_new_n11211__ = ~pi13 & ~new_new_n9180__;
  assign new_new_n11212__ = pi13 & ~new_new_n9182__;
  assign new_new_n11213__ = new_new_n6994__ & ~new_new_n11211__;
  assign new_new_n11214__ = ~new_new_n11212__ & new_new_n11213__;
  assign new_new_n11215__ = new_new_n6994__ & ~new_new_n9177__;
  assign new_new_n11216__ = ~pi14 & new_new_n11207__;
  assign new_new_n11217__ = ~new_new_n11215__ & new_new_n11216__;
  assign new_new_n11218__ = ~new_new_n11214__ & ~new_new_n11217__;
  assign new_new_n11219__ = ~new_new_n11210__ & new_new_n11218__;
  assign new_new_n11220__ = ~new_new_n11204__ & new_new_n11219__;
  assign new_new_n11221__ = ~new_new_n11203__ & ~new_new_n11220__;
  assign new_new_n11222__ = ~new_new_n10816__ & new_new_n11221__;
  assign new_new_n11223__ = new_new_n10816__ & ~new_new_n11221__;
  assign new_new_n11224__ = ~new_new_n10245__ & ~new_new_n10557__;
  assign new_new_n11225__ = new_new_n10790__ & ~new_new_n11224__;
  assign new_new_n11226__ = ~new_new_n10790__ & new_new_n11224__;
  assign new_new_n11227__ = ~new_new_n11225__ & ~new_new_n11226__;
  assign new_new_n11228__ = ~new_new_n11223__ & new_new_n11227__;
  assign new_new_n11229__ = ~new_new_n11222__ & ~new_new_n11228__;
  assign new_new_n11230__ = ~new_new_n10801__ & ~new_new_n11229__;
  assign new_new_n11231__ = new_new_n10801__ & new_new_n11229__;
  assign new_new_n11232__ = ~new_new_n3535__ & new_new_n6985__;
  assign new_new_n11233__ = ~new_new_n2130__ & new_new_n6991__;
  assign new_new_n11234__ = ~new_new_n11232__ & ~new_new_n11233__;
  assign new_new_n11235__ = ~new_new_n5520__ & new_new_n6994__;
  assign new_new_n11236__ = pi14 & ~new_new_n11235__;
  assign new_new_n11237__ = new_new_n7273__ & new_new_n8388__;
  assign new_new_n11238__ = ~new_new_n11236__ & ~new_new_n11237__;
  assign new_new_n11239__ = new_new_n11234__ & ~new_new_n11238__;
  assign new_new_n11240__ = new_new_n6553__ & new_new_n6994__;
  assign new_new_n11241__ = new_new_n11234__ & ~new_new_n11240__;
  assign new_new_n11242__ = ~pi14 & ~new_new_n11241__;
  assign new_new_n11243__ = new_new_n1823__ & new_new_n8820__;
  assign new_new_n11244__ = new_new_n5501__ & new_new_n11243__;
  assign new_new_n11245__ = ~new_new_n11242__ & ~new_new_n11244__;
  assign new_new_n11246__ = ~new_new_n11239__ & new_new_n11245__;
  assign new_new_n11247__ = ~new_new_n11231__ & new_new_n11246__;
  assign new_new_n11248__ = ~new_new_n11230__ & ~new_new_n11247__;
  assign new_new_n11249__ = ~new_new_n10781__ & ~new_new_n11248__;
  assign new_new_n11250__ = new_new_n10781__ & new_new_n11248__;
  assign new_new_n11251__ = ~new_new_n10584__ & ~new_new_n10585__;
  assign new_new_n11252__ = new_new_n10601__ & new_new_n11251__;
  assign new_new_n11253__ = ~new_new_n10601__ & ~new_new_n11251__;
  assign new_new_n11254__ = ~new_new_n11252__ & ~new_new_n11253__;
  assign new_new_n11255__ = ~new_new_n11250__ & ~new_new_n11254__;
  assign new_new_n11256__ = ~new_new_n11249__ & ~new_new_n11255__;
  assign new_new_n11257__ = new_new_n10767__ & ~new_new_n11256__;
  assign new_new_n11258__ = ~new_new_n10767__ & new_new_n11256__;
  assign new_new_n11259__ = ~new_new_n1902__ & new_new_n6985__;
  assign new_new_n11260__ = ~new_new_n1823__ & new_new_n6991__;
  assign new_new_n11261__ = ~new_new_n11259__ & ~new_new_n11260__;
  assign new_new_n11262__ = ~new_new_n1660__ & new_new_n6994__;
  assign new_new_n11263__ = ~new_new_n5274__ & new_new_n11262__;
  assign new_new_n11264__ = new_new_n11261__ & ~new_new_n11263__;
  assign new_new_n11265__ = ~pi14 & ~new_new_n11264__;
  assign new_new_n11266__ = pi13 & ~new_new_n1660__;
  assign new_new_n11267__ = ~pi13 & ~new_new_n5274__;
  assign new_new_n11268__ = new_new_n1660__ & new_new_n5273__;
  assign new_new_n11269__ = new_new_n6994__ & ~new_new_n11268__;
  assign new_new_n11270__ = ~new_new_n11266__ & ~new_new_n11267__;
  assign new_new_n11271__ = new_new_n11269__ & new_new_n11270__;
  assign new_new_n11272__ = pi14 & new_new_n11261__;
  assign new_new_n11273__ = ~new_new_n11269__ & new_new_n11272__;
  assign new_new_n11274__ = ~new_new_n11265__ & ~new_new_n11273__;
  assign new_new_n11275__ = ~new_new_n11271__ & new_new_n11274__;
  assign new_new_n11276__ = ~new_new_n11258__ & new_new_n11275__;
  assign new_new_n11277__ = ~new_new_n11257__ & ~new_new_n11276__;
  assign new_new_n11278__ = new_new_n1737__ & ~new_new_n10772__;
  assign new_new_n11279__ = ~new_new_n5688__ & new_new_n10772__;
  assign new_new_n11280__ = new_new_n6994__ & ~new_new_n11278__;
  assign new_new_n11281__ = ~new_new_n11279__ & new_new_n11280__;
  assign new_new_n11282__ = ~new_new_n1660__ & new_new_n6985__;
  assign new_new_n11283__ = ~new_new_n1902__ & new_new_n6991__;
  assign new_new_n11284__ = ~new_new_n11282__ & ~new_new_n11283__;
  assign new_new_n11285__ = ~new_new_n11281__ & new_new_n11284__;
  assign new_new_n11286__ = pi14 & ~new_new_n11285__;
  assign new_new_n11287__ = ~new_new_n6991__ & ~new_new_n11282__;
  assign new_new_n11288__ = new_new_n1902__ & new_new_n11183__;
  assign new_new_n11289__ = ~new_new_n11287__ & ~new_new_n11288__;
  assign new_new_n11290__ = ~pi14 & ~new_new_n11289__;
  assign new_new_n11291__ = ~new_new_n11281__ & new_new_n11290__;
  assign new_new_n11292__ = ~new_new_n11286__ & ~new_new_n11291__;
  assign new_new_n11293__ = ~new_new_n11277__ & ~new_new_n11292__;
  assign new_new_n11294__ = new_new_n11277__ & new_new_n11292__;
  assign new_new_n11295__ = ~new_new_n11293__ & ~new_new_n11294__;
  assign new_new_n11296__ = ~new_new_n10615__ & ~new_new_n10634__;
  assign new_new_n11297__ = ~new_new_n10631__ & new_new_n11296__;
  assign new_new_n11298__ = new_new_n10631__ & ~new_new_n11296__;
  assign new_new_n11299__ = ~new_new_n11297__ & ~new_new_n11298__;
  assign new_new_n11300__ = new_new_n11295__ & ~new_new_n11299__;
  assign new_new_n11301__ = ~new_new_n11293__ & ~new_new_n11300__;
  assign new_new_n11302__ = ~new_new_n10205__ & new_new_n10636__;
  assign new_new_n11303__ = new_new_n10205__ & ~new_new_n10605__;
  assign new_new_n11304__ = new_new_n10631__ & new_new_n10633__;
  assign new_new_n11305__ = ~new_new_n11303__ & ~new_new_n11304__;
  assign new_new_n11306__ = ~new_new_n10614__ & ~new_new_n11305__;
  assign new_new_n11307__ = ~new_new_n10605__ & new_new_n10633__;
  assign new_new_n11308__ = new_new_n10205__ & new_new_n10631__;
  assign new_new_n11309__ = ~new_new_n11307__ & ~new_new_n11308__;
  assign new_new_n11310__ = new_new_n11299__ & ~new_new_n11309__;
  assign new_new_n11311__ = ~new_new_n11302__ & ~new_new_n11306__;
  assign new_new_n11312__ = ~new_new_n11310__ & new_new_n11311__;
  assign new_new_n11313__ = ~new_new_n11301__ & ~new_new_n11312__;
  assign new_new_n11314__ = new_new_n11301__ & new_new_n11312__;
  assign new_new_n11315__ = ~new_new_n1660__ & new_new_n6991__;
  assign new_new_n11316__ = ~new_new_n1737__ & new_new_n6985__;
  assign new_new_n11317__ = ~new_new_n11315__ & ~new_new_n11316__;
  assign new_new_n11318__ = new_new_n5881__ & new_new_n6994__;
  assign new_new_n11319__ = new_new_n11317__ & ~new_new_n11318__;
  assign new_new_n11320__ = pi14 & ~new_new_n11319__;
  assign new_new_n11321__ = ~pi13 & ~new_new_n5665__;
  assign new_new_n11322__ = pi13 & ~new_new_n5875__;
  assign new_new_n11323__ = new_new_n6994__ & ~new_new_n11321__;
  assign new_new_n11324__ = ~new_new_n11322__ & new_new_n11323__;
  assign new_new_n11325__ = ~new_new_n5874__ & new_new_n6994__;
  assign new_new_n11326__ = ~pi14 & new_new_n11317__;
  assign new_new_n11327__ = ~new_new_n11325__ & new_new_n11326__;
  assign new_new_n11328__ = ~new_new_n11320__ & ~new_new_n11327__;
  assign new_new_n11329__ = ~new_new_n11324__ & new_new_n11328__;
  assign new_new_n11330__ = ~new_new_n11314__ & ~new_new_n11329__;
  assign new_new_n11331__ = ~new_new_n11313__ & ~new_new_n11330__;
  assign new_new_n11332__ = ~new_new_n10763__ & ~new_new_n11331__;
  assign new_new_n11333__ = ~new_new_n10762__ & ~new_new_n11332__;
  assign new_new_n11334__ = ~new_new_n1556__ & new_new_n6985__;
  assign new_new_n11335__ = ~new_new_n1466__ & new_new_n6991__;
  assign new_new_n11336__ = ~new_new_n11334__ & ~new_new_n11335__;
  assign new_new_n11337__ = ~new_new_n1325__ & new_new_n6994__;
  assign new_new_n11338__ = new_new_n5048__ & new_new_n11337__;
  assign new_new_n11339__ = new_new_n11336__ & ~new_new_n11338__;
  assign new_new_n11340__ = pi14 & ~new_new_n11339__;
  assign new_new_n11341__ = pi13 & new_new_n5048__;
  assign new_new_n11342__ = new_new_n1325__ & ~new_new_n5048__;
  assign new_new_n11343__ = new_new_n6994__ & ~new_new_n11342__;
  assign new_new_n11344__ = ~pi13 & ~new_new_n1325__;
  assign new_new_n11345__ = ~new_new_n11341__ & ~new_new_n11344__;
  assign new_new_n11346__ = new_new_n11343__ & new_new_n11345__;
  assign new_new_n11347__ = ~pi14 & new_new_n11336__;
  assign new_new_n11348__ = ~new_new_n11343__ & new_new_n11347__;
  assign new_new_n11349__ = ~new_new_n11340__ & ~new_new_n11346__;
  assign new_new_n11350__ = ~new_new_n11348__ & new_new_n11349__;
  assign new_new_n11351__ = ~new_new_n11333__ & ~new_new_n11350__;
  assign new_new_n11352__ = new_new_n11333__ & new_new_n11350__;
  assign new_new_n11353__ = ~new_new_n10656__ & ~new_new_n10674__;
  assign new_new_n11354__ = ~new_new_n10673__ & new_new_n11353__;
  assign new_new_n11355__ = new_new_n10673__ & ~new_new_n11353__;
  assign new_new_n11356__ = ~new_new_n11354__ & ~new_new_n11355__;
  assign new_new_n11357__ = ~new_new_n11352__ & new_new_n11356__;
  assign new_new_n11358__ = ~new_new_n11351__ & ~new_new_n11357__;
  assign new_new_n11359__ = new_new_n10740__ & ~new_new_n11358__;
  assign new_new_n11360__ = ~new_new_n10740__ & new_new_n11358__;
  assign new_new_n11361__ = ~new_new_n1207__ & new_new_n8474__;
  assign new_new_n11362__ = ~new_new_n1061__ & ~new_new_n8479__;
  assign new_new_n11363__ = ~new_new_n4550__ & new_new_n8470__;
  assign new_new_n11364__ = ~new_new_n11361__ & ~new_new_n11362__;
  assign new_new_n11365__ = ~new_new_n11363__ & new_new_n11364__;
  assign new_new_n11366__ = ~new_new_n868__ & new_new_n8469__;
  assign new_new_n11367__ = pi11 & ~new_new_n11366__;
  assign new_new_n11368__ = ~pi10 & new_new_n8469__;
  assign new_new_n11369__ = ~new_new_n868__ & new_new_n11368__;
  assign new_new_n11370__ = ~new_new_n11367__ & ~new_new_n11369__;
  assign new_new_n11371__ = new_new_n11365__ & ~new_new_n11370__;
  assign new_new_n11372__ = ~pi11 & ~new_new_n11365__;
  assign new_new_n11373__ = ~new_new_n11371__ & ~new_new_n11372__;
  assign new_new_n11374__ = ~new_new_n11360__ & new_new_n11373__;
  assign new_new_n11375__ = ~new_new_n11359__ & ~new_new_n11374__;
  assign new_new_n11376__ = ~new_new_n583__ & new_new_n10698__;
  assign new_new_n11377__ = ~new_new_n691__ & new_new_n10702__;
  assign new_new_n11378__ = new_new_n10694__ & ~new_new_n10697__;
  assign new_new_n11379__ = new_new_n3742__ & new_new_n11378__;
  assign new_new_n11380__ = ~new_new_n11376__ & ~new_new_n11377__;
  assign new_new_n11381__ = ~new_new_n11379__ & new_new_n11380__;
  assign new_new_n11382__ = ~new_new_n910__ & new_new_n10709__;
  assign new_new_n11383__ = pi08 & ~new_new_n11382__;
  assign new_new_n11384__ = ~new_new_n910__ & new_new_n10712__;
  assign new_new_n11385__ = ~pi08 & ~new_new_n11384__;
  assign new_new_n11386__ = pi05 & ~new_new_n11385__;
  assign new_new_n11387__ = ~new_new_n11383__ & ~new_new_n11386__;
  assign new_new_n11388__ = new_new_n11381__ & ~new_new_n11387__;
  assign new_new_n11389__ = ~pi08 & ~new_new_n11381__;
  assign new_new_n11390__ = ~new_new_n11388__ & ~new_new_n11389__;
  assign new_new_n11391__ = ~new_new_n11375__ & new_new_n11390__;
  assign new_new_n11392__ = new_new_n11375__ & ~new_new_n11390__;
  assign new_new_n11393__ = ~new_new_n10679__ & ~new_new_n10680__;
  assign new_new_n11394__ = ~new_new_n10690__ & ~new_new_n11393__;
  assign new_new_n11395__ = new_new_n10690__ & new_new_n11393__;
  assign new_new_n11396__ = ~new_new_n11394__ & ~new_new_n11395__;
  assign new_new_n11397__ = ~new_new_n11392__ & ~new_new_n11396__;
  assign new_new_n11398__ = ~new_new_n11391__ & ~new_new_n11397__;
  assign new_new_n11399__ = ~new_new_n10736__ & ~new_new_n11398__;
  assign new_new_n11400__ = new_new_n10719__ & ~new_new_n10721__;
  assign new_new_n11401__ = ~new_new_n10722__ & ~new_new_n11400__;
  assign new_new_n11402__ = new_new_n10736__ & new_new_n11398__;
  assign new_new_n11403__ = ~new_new_n11401__ & ~new_new_n11402__;
  assign new_new_n11404__ = ~new_new_n11399__ & ~new_new_n11403__;
  assign new_new_n11405__ = ~new_new_n10723__ & new_new_n11404__;
  assign new_new_n11406__ = new_new_n6952__ & new_new_n11378__;
  assign new_new_n11407__ = new_new_n9701__ & new_new_n10695__;
  assign new_new_n11408__ = new_new_n9697__ & new_new_n10696__;
  assign new_new_n11409__ = ~new_new_n11407__ & ~new_new_n11408__;
  assign new_new_n11410__ = ~new_new_n3768__ & ~new_new_n11409__;
  assign new_new_n11411__ = ~new_new_n466__ & new_new_n10702__;
  assign new_new_n11412__ = ~new_new_n11410__ & ~new_new_n11411__;
  assign new_new_n11413__ = ~new_new_n11406__ & new_new_n11412__;
  assign new_new_n11414__ = pi08 & ~new_new_n11413__;
  assign new_new_n11415__ = ~pi08 & new_new_n11413__;
  assign new_new_n11416__ = ~new_new_n11414__ & ~new_new_n11415__;
  assign new_new_n11417__ = ~new_new_n9229__ & ~new_new_n9230__;
  assign new_new_n11418__ = ~new_new_n9630__ & new_new_n11417__;
  assign new_new_n11419__ = new_new_n9630__ & ~new_new_n11417__;
  assign new_new_n11420__ = ~new_new_n11418__ & ~new_new_n11419__;
  assign new_new_n11421__ = ~new_new_n10149__ & new_new_n10155__;
  assign new_new_n11422__ = ~new_new_n10150__ & ~new_new_n11421__;
  assign new_new_n11423__ = new_new_n11420__ & ~new_new_n11422__;
  assign new_new_n11424__ = ~new_new_n11420__ & new_new_n11422__;
  assign new_new_n11425__ = ~new_new_n910__ & new_new_n8474__;
  assign new_new_n11426__ = ~new_new_n3720__ & ~new_new_n8479__;
  assign new_new_n11427__ = new_new_n4042__ & new_new_n8470__;
  assign new_new_n11428__ = ~new_new_n11425__ & ~new_new_n11426__;
  assign new_new_n11429__ = ~new_new_n11427__ & new_new_n11428__;
  assign new_new_n11430__ = ~new_new_n691__ & new_new_n8469__;
  assign new_new_n11431__ = pi11 & ~new_new_n11430__;
  assign new_new_n11432__ = ~new_new_n691__ & new_new_n11368__;
  assign new_new_n11433__ = ~new_new_n11431__ & ~new_new_n11432__;
  assign new_new_n11434__ = new_new_n11429__ & ~new_new_n11433__;
  assign new_new_n11435__ = ~pi11 & ~new_new_n11429__;
  assign new_new_n11436__ = ~new_new_n11434__ & ~new_new_n11435__;
  assign new_new_n11437__ = ~new_new_n11424__ & ~new_new_n11436__;
  assign new_new_n11438__ = ~new_new_n11423__ & ~new_new_n11437__;
  assign new_new_n11439__ = ~new_new_n9633__ & ~new_new_n9634__;
  assign new_new_n11440__ = ~new_new_n9664__ & new_new_n11439__;
  assign new_new_n11441__ = new_new_n9664__ & ~new_new_n11439__;
  assign new_new_n11442__ = ~new_new_n11440__ & ~new_new_n11441__;
  assign new_new_n11443__ = ~new_new_n11438__ & new_new_n11442__;
  assign new_new_n11444__ = new_new_n11438__ & ~new_new_n11442__;
  assign new_new_n11445__ = ~new_new_n11443__ & ~new_new_n11444__;
  assign new_new_n11446__ = new_new_n11416__ & new_new_n11445__;
  assign new_new_n11447__ = ~new_new_n11416__ & ~new_new_n11445__;
  assign new_new_n11448__ = ~new_new_n11446__ & ~new_new_n11447__;
  assign new_new_n11449__ = new_new_n11405__ & new_new_n11448__;
  assign new_new_n11450__ = new_new_n10723__ & ~new_new_n11404__;
  assign new_new_n11451__ = ~new_new_n3768__ & new_new_n10702__;
  assign new_new_n11452__ = new_new_n466__ & new_new_n10697__;
  assign new_new_n11453__ = ~new_new_n4172__ & ~new_new_n10697__;
  assign new_new_n11454__ = new_new_n10694__ & ~new_new_n11452__;
  assign new_new_n11455__ = ~new_new_n11453__ & new_new_n11454__;
  assign new_new_n11456__ = ~new_new_n11451__ & ~new_new_n11455__;
  assign new_new_n11457__ = ~new_new_n583__ & new_new_n10709__;
  assign new_new_n11458__ = pi08 & ~new_new_n11457__;
  assign new_new_n11459__ = ~new_new_n583__ & new_new_n10712__;
  assign new_new_n11460__ = ~pi08 & ~new_new_n11459__;
  assign new_new_n11461__ = pi05 & ~new_new_n11460__;
  assign new_new_n11462__ = ~new_new_n11458__ & ~new_new_n11461__;
  assign new_new_n11463__ = new_new_n11456__ & ~new_new_n11462__;
  assign new_new_n11464__ = ~pi08 & ~new_new_n11456__;
  assign new_new_n11465__ = ~new_new_n11463__ & ~new_new_n11464__;
  assign new_new_n11466__ = ~pi03 & ~pi04;
  assign new_new_n11467__ = pi03 & pi04;
  assign new_new_n11468__ = ~new_new_n11466__ & ~new_new_n11467__;
  assign new_new_n11469__ = ~new_new_n10726__ & ~new_new_n10731__;
  assign new_new_n11470__ = ~new_new_n11468__ & ~new_new_n11469__;
  assign new_new_n11471__ = new_new_n7191__ & new_new_n11470__;
  assign new_new_n11472__ = ~new_new_n583__ & new_new_n11471__;
  assign new_new_n11473__ = ~pi04 & ~new_new_n10731__;
  assign new_new_n11474__ = pi04 & ~new_new_n10726__;
  assign new_new_n11475__ = ~new_new_n11473__ & ~new_new_n11474__;
  assign new_new_n11476__ = ~new_new_n3768__ & new_new_n11475__;
  assign new_new_n11477__ = pi04 & pi05;
  assign new_new_n11478__ = ~new_new_n10727__ & ~new_new_n11477__;
  assign new_new_n11479__ = new_new_n466__ & ~new_new_n11478__;
  assign new_new_n11480__ = ~pi02 & pi03;
  assign new_new_n11481__ = pi02 & ~pi03;
  assign new_new_n11482__ = ~new_new_n11480__ & ~new_new_n11481__;
  assign new_new_n11483__ = ~new_new_n4172__ & new_new_n11478__;
  assign new_new_n11484__ = ~new_new_n11479__ & ~new_new_n11482__;
  assign new_new_n11485__ = ~new_new_n11483__ & new_new_n11484__;
  assign new_new_n11486__ = ~new_new_n11472__ & ~new_new_n11476__;
  assign new_new_n11487__ = ~new_new_n11485__ & new_new_n11486__;
  assign new_new_n11488__ = pi05 & ~new_new_n11487__;
  assign new_new_n11489__ = ~pi05 & new_new_n11487__;
  assign new_new_n11490__ = ~new_new_n11488__ & ~new_new_n11489__;
  assign new_new_n11491__ = ~new_new_n3720__ & ~new_new_n11409__;
  assign new_new_n11492__ = ~new_new_n691__ & new_new_n10698__;
  assign new_new_n11493__ = ~new_new_n910__ & new_new_n10702__;
  assign new_new_n11494__ = ~new_new_n11491__ & ~new_new_n11492__;
  assign new_new_n11495__ = ~new_new_n11493__ & new_new_n11494__;
  assign new_new_n11496__ = new_new_n4042__ & new_new_n10694__;
  assign new_new_n11497__ = pi08 & ~new_new_n11496__;
  assign new_new_n11498__ = pi07 & new_new_n10694__;
  assign new_new_n11499__ = new_new_n4042__ & new_new_n11498__;
  assign new_new_n11500__ = ~new_new_n11497__ & ~new_new_n11499__;
  assign new_new_n11501__ = new_new_n11495__ & ~new_new_n11500__;
  assign new_new_n11502__ = ~pi08 & ~new_new_n11495__;
  assign new_new_n11503__ = ~new_new_n11501__ & ~new_new_n11502__;
  assign new_new_n11504__ = ~new_new_n11351__ & ~new_new_n11352__;
  assign new_new_n11505__ = ~new_new_n11356__ & new_new_n11504__;
  assign new_new_n11506__ = new_new_n11356__ & ~new_new_n11504__;
  assign new_new_n11507__ = ~new_new_n11505__ & ~new_new_n11506__;
  assign new_new_n11508__ = ~new_new_n1325__ & new_new_n8474__;
  assign new_new_n11509__ = ~new_new_n5981__ & ~new_new_n8344__;
  assign new_new_n11510__ = new_new_n8470__ & ~new_new_n11509__;
  assign new_new_n11511__ = ~new_new_n11508__ & ~new_new_n11510__;
  assign new_new_n11512__ = ~new_new_n3618__ & new_new_n8858__;
  assign new_new_n11513__ = ~new_new_n1556__ & ~new_new_n8479__;
  assign new_new_n11514__ = ~new_new_n11512__ & ~new_new_n11513__;
  assign new_new_n11515__ = new_new_n11511__ & new_new_n11514__;
  assign new_new_n11516__ = ~pi11 & ~new_new_n11515__;
  assign new_new_n11517__ = ~new_new_n8858__ & ~new_new_n11513__;
  assign new_new_n11518__ = new_new_n3618__ & new_new_n8479__;
  assign new_new_n11519__ = ~new_new_n11517__ & ~new_new_n11518__;
  assign new_new_n11520__ = pi11 & ~new_new_n11519__;
  assign new_new_n11521__ = new_new_n11511__ & new_new_n11520__;
  assign new_new_n11522__ = ~new_new_n11516__ & ~new_new_n11521__;
  assign new_new_n11523__ = ~new_new_n1466__ & ~new_new_n8479__;
  assign new_new_n11524__ = ~new_new_n1325__ & new_new_n8858__;
  assign new_new_n11525__ = ~new_new_n1556__ & new_new_n8474__;
  assign new_new_n11526__ = ~new_new_n11523__ & ~new_new_n11524__;
  assign new_new_n11527__ = ~new_new_n11525__ & new_new_n11526__;
  assign new_new_n11528__ = new_new_n5048__ & new_new_n8469__;
  assign new_new_n11529__ = pi11 & ~new_new_n11528__;
  assign new_new_n11530__ = pi10 & new_new_n8469__;
  assign new_new_n11531__ = new_new_n5048__ & new_new_n11530__;
  assign new_new_n11532__ = ~new_new_n11529__ & ~new_new_n11531__;
  assign new_new_n11533__ = new_new_n11527__ & ~new_new_n11532__;
  assign new_new_n11534__ = ~pi11 & ~new_new_n11527__;
  assign new_new_n11535__ = ~new_new_n11533__ & ~new_new_n11534__;
  assign new_new_n11536__ = ~new_new_n1660__ & ~new_new_n8479__;
  assign new_new_n11537__ = ~new_new_n1466__ & new_new_n8858__;
  assign new_new_n11538__ = ~new_new_n1737__ & new_new_n8474__;
  assign new_new_n11539__ = ~new_new_n11536__ & ~new_new_n11537__;
  assign new_new_n11540__ = ~new_new_n11538__ & new_new_n11539__;
  assign new_new_n11541__ = ~new_new_n6410__ & new_new_n8469__;
  assign new_new_n11542__ = pi11 & ~new_new_n11541__;
  assign new_new_n11543__ = ~new_new_n6410__ & new_new_n11530__;
  assign new_new_n11544__ = ~new_new_n11542__ & ~new_new_n11543__;
  assign new_new_n11545__ = new_new_n11540__ & ~new_new_n11544__;
  assign new_new_n11546__ = ~pi11 & ~new_new_n11540__;
  assign new_new_n11547__ = ~new_new_n11545__ & ~new_new_n11546__;
  assign new_new_n11548__ = ~new_new_n3535__ & new_new_n8474__;
  assign new_new_n11549__ = ~new_new_n2130__ & ~new_new_n8479__;
  assign new_new_n11550__ = ~new_new_n11548__ & ~new_new_n11549__;
  assign new_new_n11551__ = ~new_new_n5520__ & new_new_n8469__;
  assign new_new_n11552__ = pi11 & ~new_new_n11551__;
  assign new_new_n11553__ = ~pi10 & new_new_n1823__;
  assign new_new_n11554__ = pi10 & ~new_new_n1823__;
  assign new_new_n11555__ = new_new_n8469__ & ~new_new_n11553__;
  assign new_new_n11556__ = ~new_new_n11554__ & new_new_n11555__;
  assign new_new_n11557__ = new_new_n5501__ & new_new_n11556__;
  assign new_new_n11558__ = ~new_new_n11552__ & ~new_new_n11557__;
  assign new_new_n11559__ = new_new_n11550__ & ~new_new_n11558__;
  assign new_new_n11560__ = new_new_n6553__ & new_new_n8469__;
  assign new_new_n11561__ = new_new_n11550__ & ~new_new_n11560__;
  assign new_new_n11562__ = ~pi11 & ~new_new_n11561__;
  assign new_new_n11563__ = ~new_new_n11559__ & ~new_new_n11562__;
  assign new_new_n11564__ = ~new_new_n11191__ & ~new_new_n11192__;
  assign new_new_n11565__ = new_new_n11196__ & new_new_n11564__;
  assign new_new_n11566__ = ~new_new_n11196__ & ~new_new_n11564__;
  assign new_new_n11567__ = ~new_new_n11565__ & ~new_new_n11566__;
  assign new_new_n11568__ = new_new_n11563__ & new_new_n11567__;
  assign new_new_n11569__ = ~new_new_n11169__ & ~new_new_n11170__;
  assign new_new_n11570__ = new_new_n11188__ & ~new_new_n11569__;
  assign new_new_n11571__ = ~new_new_n11188__ & new_new_n11569__;
  assign new_new_n11572__ = ~new_new_n11570__ & ~new_new_n11571__;
  assign new_new_n11573__ = ~new_new_n11160__ & ~new_new_n11162__;
  assign new_new_n11574__ = ~new_new_n11163__ & ~new_new_n11573__;
  assign new_new_n11575__ = ~new_new_n6036__ & new_new_n8470__;
  assign new_new_n11576__ = ~new_new_n2024__ & new_new_n8474__;
  assign new_new_n11577__ = ~new_new_n2224__ & ~new_new_n8479__;
  assign new_new_n11578__ = ~new_new_n11576__ & ~new_new_n11577__;
  assign new_new_n11579__ = ~new_new_n11575__ & new_new_n11578__;
  assign new_new_n11580__ = ~new_new_n2130__ & new_new_n8469__;
  assign new_new_n11581__ = pi11 & ~new_new_n11580__;
  assign new_new_n11582__ = ~new_new_n2130__ & new_new_n11368__;
  assign new_new_n11583__ = ~new_new_n11581__ & ~new_new_n11582__;
  assign new_new_n11584__ = new_new_n11579__ & ~new_new_n11583__;
  assign new_new_n11585__ = ~pi11 & ~new_new_n11579__;
  assign new_new_n11586__ = ~new_new_n11584__ & ~new_new_n11585__;
  assign new_new_n11587__ = ~new_new_n11574__ & new_new_n11586__;
  assign new_new_n11588__ = new_new_n11574__ & ~new_new_n11586__;
  assign new_new_n11589__ = ~new_new_n10892__ & ~new_new_n10893__;
  assign new_new_n11590__ = ~new_new_n11150__ & new_new_n11589__;
  assign new_new_n11591__ = new_new_n11150__ & ~new_new_n11589__;
  assign new_new_n11592__ = ~new_new_n11590__ & ~new_new_n11591__;
  assign new_new_n11593__ = ~new_new_n2313__ & ~new_new_n8479__;
  assign new_new_n11594__ = ~new_new_n2224__ & new_new_n8858__;
  assign new_new_n11595__ = ~new_new_n2420__ & new_new_n8474__;
  assign new_new_n11596__ = new_new_n6521__ & new_new_n8470__;
  assign new_new_n11597__ = ~new_new_n11593__ & ~new_new_n11594__;
  assign new_new_n11598__ = ~new_new_n11595__ & new_new_n11597__;
  assign new_new_n11599__ = ~new_new_n11596__ & new_new_n11598__;
  assign new_new_n11600__ = ~pi11 & new_new_n11599__;
  assign new_new_n11601__ = ~new_new_n11153__ & ~new_new_n11154__;
  assign new_new_n11602__ = new_new_n11158__ & new_new_n11601__;
  assign new_new_n11603__ = ~new_new_n11158__ & ~new_new_n11601__;
  assign new_new_n11604__ = ~new_new_n11602__ & ~new_new_n11603__;
  assign new_new_n11605__ = ~new_new_n11599__ & new_new_n11604__;
  assign new_new_n11606__ = ~new_new_n11600__ & ~new_new_n11605__;
  assign new_new_n11607__ = ~new_new_n2224__ & new_new_n8474__;
  assign new_new_n11608__ = ~new_new_n2024__ & new_new_n8858__;
  assign new_new_n11609__ = ~new_new_n2420__ & ~new_new_n8479__;
  assign new_new_n11610__ = new_new_n7313__ & new_new_n8470__;
  assign new_new_n11611__ = ~new_new_n11607__ & ~new_new_n11608__;
  assign new_new_n11612__ = ~new_new_n11609__ & new_new_n11611__;
  assign new_new_n11613__ = ~new_new_n11610__ & new_new_n11612__;
  assign new_new_n11614__ = ~new_new_n11606__ & new_new_n11613__;
  assign new_new_n11615__ = new_new_n11599__ & new_new_n11604__;
  assign new_new_n11616__ = ~new_new_n2313__ & new_new_n8474__;
  assign new_new_n11617__ = ~new_new_n2572__ & ~new_new_n8479__;
  assign new_new_n11618__ = ~new_new_n11616__ & ~new_new_n11617__;
  assign new_new_n11619__ = new_new_n6749__ & new_new_n8469__;
  assign new_new_n11620__ = new_new_n11618__ & ~new_new_n11619__;
  assign new_new_n11621__ = pi11 & ~new_new_n11620__;
  assign new_new_n11622__ = new_new_n8469__ & ~new_new_n9267__;
  assign new_new_n11623__ = ~pi11 & ~new_new_n11622__;
  assign new_new_n11624__ = pi10 & new_new_n2420__;
  assign new_new_n11625__ = ~pi10 & ~new_new_n2420__;
  assign new_new_n11626__ = new_new_n8469__ & ~new_new_n11624__;
  assign new_new_n11627__ = ~new_new_n11625__ & new_new_n11626__;
  assign new_new_n11628__ = new_new_n6748__ & new_new_n11627__;
  assign new_new_n11629__ = ~new_new_n11623__ & ~new_new_n11628__;
  assign new_new_n11630__ = new_new_n11618__ & ~new_new_n11629__;
  assign new_new_n11631__ = ~new_new_n11621__ & ~new_new_n11630__;
  assign new_new_n11632__ = ~new_new_n10943__ & ~new_new_n10944__;
  assign new_new_n11633__ = ~new_new_n11111__ & new_new_n11632__;
  assign new_new_n11634__ = new_new_n11111__ & ~new_new_n11632__;
  assign new_new_n11635__ = ~new_new_n11633__ & ~new_new_n11634__;
  assign new_new_n11636__ = ~new_new_n2737__ & ~new_new_n8479__;
  assign new_new_n11637__ = ~new_new_n2636__ & new_new_n8474__;
  assign new_new_n11638__ = new_new_n7774__ & ~new_new_n8468__;
  assign new_new_n11639__ = new_new_n2497__ & new_new_n8468__;
  assign new_new_n11640__ = new_new_n8469__ & ~new_new_n11639__;
  assign new_new_n11641__ = ~new_new_n11638__ & new_new_n11640__;
  assign new_new_n11642__ = ~new_new_n11636__ & ~new_new_n11637__;
  assign new_new_n11643__ = ~new_new_n11641__ & new_new_n11642__;
  assign new_new_n11644__ = pi11 & ~new_new_n11643__;
  assign new_new_n11645__ = ~pi11 & new_new_n11643__;
  assign new_new_n11646__ = ~new_new_n11644__ & ~new_new_n11645__;
  assign new_new_n11647__ = ~new_new_n11064__ & ~new_new_n11065__;
  assign new_new_n11648__ = new_new_n11082__ & new_new_n11647__;
  assign new_new_n11649__ = ~new_new_n11082__ & ~new_new_n11647__;
  assign new_new_n11650__ = ~new_new_n11648__ & ~new_new_n11649__;
  assign new_new_n11651__ = ~new_new_n2737__ & new_new_n8474__;
  assign new_new_n11652__ = ~new_new_n2886__ & ~new_new_n8479__;
  assign new_new_n11653__ = new_new_n2636__ & new_new_n8468__;
  assign new_new_n11654__ = new_new_n7814__ & ~new_new_n8468__;
  assign new_new_n11655__ = new_new_n8469__ & ~new_new_n11653__;
  assign new_new_n11656__ = ~new_new_n11654__ & new_new_n11655__;
  assign new_new_n11657__ = ~new_new_n11651__ & ~new_new_n11652__;
  assign new_new_n11658__ = ~new_new_n11656__ & new_new_n11657__;
  assign new_new_n11659__ = ~new_new_n10970__ & ~new_new_n10971__;
  assign new_new_n11660__ = ~new_new_n11084__ & new_new_n11659__;
  assign new_new_n11661__ = new_new_n11084__ & ~new_new_n11659__;
  assign new_new_n11662__ = ~new_new_n11660__ & ~new_new_n11661__;
  assign new_new_n11663__ = ~new_new_n2848__ & ~new_new_n8479__;
  assign new_new_n11664__ = ~new_new_n2737__ & new_new_n8858__;
  assign new_new_n11665__ = ~new_new_n2886__ & new_new_n8474__;
  assign new_new_n11666__ = ~new_new_n7378__ & new_new_n8470__;
  assign new_new_n11667__ = ~new_new_n11663__ & ~new_new_n11664__;
  assign new_new_n11668__ = ~new_new_n11665__ & new_new_n11667__;
  assign new_new_n11669__ = ~new_new_n11666__ & new_new_n11668__;
  assign new_new_n11670__ = ~new_new_n11662__ & new_new_n11669__;
  assign new_new_n11671__ = pi11 & ~new_new_n11669__;
  assign new_new_n11672__ = ~new_new_n11670__ & ~new_new_n11671__;
  assign new_new_n11673__ = ~new_new_n11658__ & new_new_n11672__;
  assign new_new_n11674__ = new_new_n11662__ & ~new_new_n11669__;
  assign new_new_n11675__ = ~new_new_n2848__ & new_new_n8474__;
  assign new_new_n11676__ = ~new_new_n3460__ & ~new_new_n8479__;
  assign new_new_n11677__ = ~new_new_n2886__ & new_new_n8858__;
  assign new_new_n11678__ = new_new_n8470__ & ~new_new_n8574__;
  assign new_new_n11679__ = ~new_new_n11675__ & ~new_new_n11676__;
  assign new_new_n11680__ = ~new_new_n11677__ & new_new_n11679__;
  assign new_new_n11681__ = ~new_new_n11678__ & new_new_n11680__;
  assign new_new_n11682__ = pi11 & ~new_new_n11681__;
  assign new_new_n11683__ = ~pi11 & new_new_n11681__;
  assign new_new_n11684__ = ~new_new_n11682__ & ~new_new_n11683__;
  assign new_new_n11685__ = ~new_new_n10996__ & ~new_new_n10997__;
  assign new_new_n11686__ = ~new_new_n11061__ & new_new_n11685__;
  assign new_new_n11687__ = new_new_n11061__ & ~new_new_n11685__;
  assign new_new_n11688__ = ~new_new_n11686__ & ~new_new_n11687__;
  assign new_new_n11689__ = ~new_new_n11684__ & ~new_new_n11688__;
  assign new_new_n11690__ = new_new_n11684__ & new_new_n11688__;
  assign new_new_n11691__ = ~new_new_n2960__ & ~new_new_n8479__;
  assign new_new_n11692__ = ~new_new_n3460__ & new_new_n8474__;
  assign new_new_n11693__ = ~new_new_n2848__ & new_new_n8858__;
  assign new_new_n11694__ = ~new_new_n11692__ & ~new_new_n11693__;
  assign new_new_n11695__ = ~new_new_n11691__ & new_new_n11694__;
  assign new_new_n11696__ = ~new_new_n7065__ & new_new_n8469__;
  assign new_new_n11697__ = pi11 & ~new_new_n11696__;
  assign new_new_n11698__ = ~new_new_n7065__ & new_new_n11530__;
  assign new_new_n11699__ = ~new_new_n11697__ & ~new_new_n11698__;
  assign new_new_n11700__ = new_new_n11695__ & ~new_new_n11699__;
  assign new_new_n11701__ = ~pi11 & ~new_new_n11695__;
  assign new_new_n11702__ = ~new_new_n11700__ & ~new_new_n11701__;
  assign new_new_n11703__ = ~new_new_n2960__ & new_new_n8474__;
  assign new_new_n11704__ = ~new_new_n7388__ & new_new_n8468__;
  assign new_new_n11705__ = new_new_n8469__ & ~new_new_n11704__;
  assign new_new_n11706__ = new_new_n7391__ & new_new_n11705__;
  assign new_new_n11707__ = ~new_new_n3126__ & ~new_new_n8479__;
  assign new_new_n11708__ = ~new_new_n3460__ & new_new_n8858__;
  assign new_new_n11709__ = ~new_new_n11707__ & ~new_new_n11708__;
  assign new_new_n11710__ = ~new_new_n11703__ & new_new_n11709__;
  assign new_new_n11711__ = ~new_new_n11706__ & new_new_n11710__;
  assign new_new_n11712__ = pi11 & ~new_new_n11711__;
  assign new_new_n11713__ = ~pi11 & new_new_n11711__;
  assign new_new_n11714__ = ~new_new_n11712__ & ~new_new_n11713__;
  assign new_new_n11715__ = new_new_n11013__ & new_new_n11014__;
  assign new_new_n11716__ = ~new_new_n11032__ & ~new_new_n11715__;
  assign new_new_n11717__ = new_new_n11015__ & ~new_new_n11716__;
  assign new_new_n11718__ = ~new_new_n11015__ & new_new_n11716__;
  assign new_new_n11719__ = ~new_new_n11717__ & ~new_new_n11718__;
  assign new_new_n11720__ = new_new_n11714__ & new_new_n11719__;
  assign new_new_n11721__ = ~new_new_n11714__ & ~new_new_n11719__;
  assign new_new_n11722__ = ~new_new_n2960__ & new_new_n8858__;
  assign new_new_n11723__ = ~new_new_n3164__ & ~new_new_n8479__;
  assign new_new_n11724__ = ~new_new_n3126__ & new_new_n8474__;
  assign new_new_n11725__ = ~new_new_n11723__ & ~new_new_n11724__;
  assign new_new_n11726__ = ~new_new_n11722__ & new_new_n11725__;
  assign new_new_n11727__ = ~new_new_n7468__ & new_new_n8469__;
  assign new_new_n11728__ = pi11 & ~new_new_n11727__;
  assign new_new_n11729__ = ~new_new_n7468__ & new_new_n11530__;
  assign new_new_n11730__ = ~new_new_n11728__ & ~new_new_n11729__;
  assign new_new_n11731__ = new_new_n11726__ & ~new_new_n11730__;
  assign new_new_n11732__ = ~pi11 & ~new_new_n11726__;
  assign new_new_n11733__ = ~new_new_n11731__ & ~new_new_n11732__;
  assign new_new_n11734__ = new_new_n7682__ & new_new_n8470__;
  assign new_new_n11735__ = ~new_new_n8474__ & ~new_new_n11734__;
  assign new_new_n11736__ = ~new_new_n3055__ & ~new_new_n11735__;
  assign new_new_n11737__ = ~new_new_n3254__ & new_new_n8469__;
  assign new_new_n11738__ = ~new_new_n3356__ & ~new_new_n8479__;
  assign new_new_n11739__ = ~new_new_n11737__ & ~new_new_n11738__;
  assign new_new_n11740__ = ~new_new_n3055__ & ~new_new_n8468__;
  assign new_new_n11741__ = new_new_n3356__ & new_new_n11740__;
  assign new_new_n11742__ = ~new_new_n11739__ & ~new_new_n11741__;
  assign new_new_n11743__ = ~new_new_n11736__ & ~new_new_n11742__;
  assign new_new_n11744__ = ~new_new_n3356__ & ~new_new_n8306__;
  assign new_new_n11745__ = ~pi10 & ~new_new_n3356__;
  assign new_new_n11746__ = ~new_new_n3055__ & ~new_new_n8301__;
  assign new_new_n11747__ = ~new_new_n8306__ & new_new_n11746__;
  assign new_new_n11748__ = ~new_new_n11744__ & ~new_new_n11745__;
  assign new_new_n11749__ = ~new_new_n11747__ & new_new_n11748__;
  assign new_new_n11750__ = ~new_new_n8477__ & ~new_new_n11749__;
  assign new_new_n11751__ = pi11 & ~new_new_n11750__;
  assign new_new_n11752__ = new_new_n11743__ & new_new_n11751__;
  assign new_new_n11753__ = ~new_new_n3254__ & new_new_n8474__;
  assign new_new_n11754__ = ~new_new_n3164__ & new_new_n8858__;
  assign new_new_n11755__ = ~new_new_n3055__ & ~new_new_n8479__;
  assign new_new_n11756__ = new_new_n8470__ & ~new_new_n8637__;
  assign new_new_n11757__ = ~new_new_n11753__ & ~new_new_n11754__;
  assign new_new_n11758__ = ~new_new_n11755__ & new_new_n11757__;
  assign new_new_n11759__ = ~new_new_n11756__ & new_new_n11758__;
  assign new_new_n11760__ = new_new_n11752__ & new_new_n11759__;
  assign new_new_n11761__ = pi11 & ~new_new_n11759__;
  assign new_new_n11762__ = pi12 & new_new_n11759__;
  assign new_new_n11763__ = ~new_new_n3356__ & ~new_new_n6981__;
  assign new_new_n11764__ = ~new_new_n11761__ & new_new_n11763__;
  assign new_new_n11765__ = ~new_new_n11762__ & new_new_n11764__;
  assign new_new_n11766__ = ~new_new_n11760__ & ~new_new_n11765__;
  assign new_new_n11767__ = ~new_new_n6983__ & ~new_new_n10999__;
  assign new_new_n11768__ = pi13 & ~new_new_n3356__;
  assign new_new_n11769__ = ~new_new_n11767__ & new_new_n11768__;
  assign new_new_n11770__ = new_new_n11767__ & ~new_new_n11768__;
  assign new_new_n11771__ = new_new_n3356__ & new_new_n6983__;
  assign new_new_n11772__ = ~new_new_n11769__ & ~new_new_n11771__;
  assign new_new_n11773__ = ~new_new_n11770__ & new_new_n11772__;
  assign new_new_n11774__ = ~new_new_n11766__ & new_new_n11773__;
  assign new_new_n11775__ = new_new_n11766__ & ~new_new_n11773__;
  assign new_new_n11776__ = ~new_new_n3254__ & ~new_new_n8479__;
  assign new_new_n11777__ = ~new_new_n3126__ & new_new_n8858__;
  assign new_new_n11778__ = ~new_new_n3164__ & new_new_n8474__;
  assign new_new_n11779__ = ~new_new_n7570__ & new_new_n8470__;
  assign new_new_n11780__ = ~new_new_n11776__ & ~new_new_n11777__;
  assign new_new_n11781__ = ~new_new_n11778__ & new_new_n11780__;
  assign new_new_n11782__ = ~new_new_n11779__ & new_new_n11781__;
  assign new_new_n11783__ = pi11 & ~new_new_n11782__;
  assign new_new_n11784__ = ~pi11 & new_new_n11782__;
  assign new_new_n11785__ = ~new_new_n11783__ & ~new_new_n11784__;
  assign new_new_n11786__ = ~new_new_n11775__ & new_new_n11785__;
  assign new_new_n11787__ = ~new_new_n11774__ & ~new_new_n11786__;
  assign new_new_n11788__ = new_new_n11003__ & ~new_new_n11012__;
  assign new_new_n11789__ = new_new_n11787__ & ~new_new_n11788__;
  assign new_new_n11790__ = ~new_new_n11733__ & ~new_new_n11789__;
  assign new_new_n11791__ = pi14 & new_new_n11002__;
  assign new_new_n11792__ = new_new_n11012__ & ~new_new_n11791__;
  assign new_new_n11793__ = new_new_n11733__ & new_new_n11787__;
  assign new_new_n11794__ = pi14 & ~new_new_n11012__;
  assign new_new_n11795__ = ~new_new_n11792__ & ~new_new_n11794__;
  assign new_new_n11796__ = ~new_new_n11793__ & new_new_n11795__;
  assign new_new_n11797__ = ~new_new_n11790__ & ~new_new_n11796__;
  assign new_new_n11798__ = ~new_new_n11721__ & ~new_new_n11797__;
  assign new_new_n11799__ = ~new_new_n11720__ & ~new_new_n11798__;
  assign new_new_n11800__ = new_new_n11702__ & new_new_n11799__;
  assign new_new_n11801__ = ~new_new_n11702__ & ~new_new_n11799__;
  assign new_new_n11802__ = ~new_new_n11051__ & ~new_new_n11052__;
  assign new_new_n11803__ = ~new_new_n11059__ & ~new_new_n11802__;
  assign new_new_n11804__ = new_new_n11059__ & new_new_n11802__;
  assign new_new_n11805__ = ~new_new_n11803__ & ~new_new_n11804__;
  assign new_new_n11806__ = ~new_new_n11801__ & ~new_new_n11805__;
  assign new_new_n11807__ = ~new_new_n11800__ & ~new_new_n11806__;
  assign new_new_n11808__ = ~new_new_n11690__ & ~new_new_n11807__;
  assign new_new_n11809__ = ~new_new_n11689__ & ~new_new_n11808__;
  assign new_new_n11810__ = ~new_new_n11669__ & ~new_new_n11809__;
  assign new_new_n11811__ = pi11 & ~new_new_n11810__;
  assign new_new_n11812__ = ~new_new_n11674__ & ~new_new_n11811__;
  assign new_new_n11813__ = new_new_n11658__ & ~new_new_n11812__;
  assign new_new_n11814__ = ~pi11 & ~new_new_n11658__;
  assign new_new_n11815__ = ~new_new_n11662__ & ~new_new_n11814__;
  assign new_new_n11816__ = new_new_n11809__ & ~new_new_n11815__;
  assign new_new_n11817__ = ~new_new_n11673__ & ~new_new_n11816__;
  assign new_new_n11818__ = ~new_new_n11813__ & new_new_n11817__;
  assign new_new_n11819__ = new_new_n11650__ & ~new_new_n11818__;
  assign new_new_n11820__ = pi11 & new_new_n11662__;
  assign new_new_n11821__ = pi11 & new_new_n11669__;
  assign new_new_n11822__ = ~new_new_n11674__ & ~new_new_n11821__;
  assign new_new_n11823__ = new_new_n11809__ & ~new_new_n11822__;
  assign new_new_n11824__ = ~new_new_n11820__ & ~new_new_n11823__;
  assign new_new_n11825__ = new_new_n11658__ & ~new_new_n11824__;
  assign new_new_n11826__ = ~pi11 & new_new_n11662__;
  assign new_new_n11827__ = new_new_n11672__ & new_new_n11809__;
  assign new_new_n11828__ = ~new_new_n11826__ & ~new_new_n11827__;
  assign new_new_n11829__ = ~new_new_n11658__ & ~new_new_n11828__;
  assign new_new_n11830__ = ~new_new_n11825__ & ~new_new_n11829__;
  assign new_new_n11831__ = ~new_new_n11819__ & new_new_n11830__;
  assign new_new_n11832__ = new_new_n11646__ & ~new_new_n11831__;
  assign new_new_n11833__ = ~new_new_n11646__ & new_new_n11831__;
  assign new_new_n11834__ = ~new_new_n11091__ & ~new_new_n11092__;
  assign new_new_n11835__ = new_new_n11109__ & new_new_n11834__;
  assign new_new_n11836__ = ~new_new_n11109__ & ~new_new_n11834__;
  assign new_new_n11837__ = ~new_new_n11835__ & ~new_new_n11836__;
  assign new_new_n11838__ = ~new_new_n11833__ & ~new_new_n11837__;
  assign new_new_n11839__ = ~new_new_n11832__ & ~new_new_n11838__;
  assign new_new_n11840__ = ~new_new_n11635__ & ~new_new_n11839__;
  assign new_new_n11841__ = new_new_n11635__ & new_new_n11839__;
  assign new_new_n11842__ = ~new_new_n2572__ & new_new_n8858__;
  assign new_new_n11843__ = ~new_new_n2636__ & ~new_new_n8479__;
  assign new_new_n11844__ = ~new_new_n2497__ & new_new_n8474__;
  assign new_new_n11845__ = new_new_n6804__ & new_new_n8470__;
  assign new_new_n11846__ = ~new_new_n11842__ & ~new_new_n11843__;
  assign new_new_n11847__ = ~new_new_n11844__ & new_new_n11846__;
  assign new_new_n11848__ = ~new_new_n11845__ & new_new_n11847__;
  assign new_new_n11849__ = pi11 & ~new_new_n11848__;
  assign new_new_n11850__ = ~pi11 & new_new_n11848__;
  assign new_new_n11851__ = ~new_new_n11849__ & ~new_new_n11850__;
  assign new_new_n11852__ = ~new_new_n11841__ & new_new_n11851__;
  assign new_new_n11853__ = ~new_new_n11840__ & ~new_new_n11852__;
  assign new_new_n11854__ = ~new_new_n2572__ & new_new_n8474__;
  assign new_new_n11855__ = ~new_new_n2497__ & ~new_new_n8479__;
  assign new_new_n11856__ = ~new_new_n2313__ & new_new_n8858__;
  assign new_new_n11857__ = ~new_new_n11854__ & ~new_new_n11855__;
  assign new_new_n11858__ = ~new_new_n11856__ & new_new_n11857__;
  assign new_new_n11859__ = ~new_new_n7236__ & new_new_n8469__;
  assign new_new_n11860__ = ~pi11 & ~new_new_n11859__;
  assign new_new_n11861__ = ~new_new_n7236__ & new_new_n11368__;
  assign new_new_n11862__ = ~new_new_n11860__ & ~new_new_n11861__;
  assign new_new_n11863__ = new_new_n11858__ & ~new_new_n11862__;
  assign new_new_n11864__ = pi11 & ~new_new_n11858__;
  assign new_new_n11865__ = ~new_new_n11863__ & ~new_new_n11864__;
  assign new_new_n11866__ = new_new_n11853__ & ~new_new_n11865__;
  assign new_new_n11867__ = ~new_new_n11853__ & new_new_n11865__;
  assign new_new_n11868__ = ~new_new_n10441__ & new_new_n11129__;
  assign new_new_n11869__ = new_new_n10441__ & ~new_new_n11129__;
  assign new_new_n11870__ = ~new_new_n11868__ & ~new_new_n11869__;
  assign new_new_n11871__ = new_new_n10910__ & ~new_new_n11870__;
  assign new_new_n11872__ = ~new_new_n10910__ & new_new_n11870__;
  assign new_new_n11873__ = ~new_new_n11871__ & ~new_new_n11872__;
  assign new_new_n11874__ = new_new_n11113__ & new_new_n11873__;
  assign new_new_n11875__ = ~new_new_n11113__ & ~new_new_n11873__;
  assign new_new_n11876__ = ~new_new_n11874__ & ~new_new_n11875__;
  assign new_new_n11877__ = ~new_new_n11867__ & ~new_new_n11876__;
  assign new_new_n11878__ = ~new_new_n11866__ & ~new_new_n11877__;
  assign new_new_n11879__ = new_new_n11631__ & new_new_n11878__;
  assign new_new_n11880__ = ~new_new_n11631__ & ~new_new_n11878__;
  assign new_new_n11881__ = ~new_new_n11132__ & ~new_new_n11133__;
  assign new_new_n11882__ = new_new_n11148__ & new_new_n11881__;
  assign new_new_n11883__ = ~new_new_n11148__ & ~new_new_n11881__;
  assign new_new_n11884__ = ~new_new_n11882__ & ~new_new_n11883__;
  assign new_new_n11885__ = ~new_new_n11880__ & new_new_n11884__;
  assign new_new_n11886__ = ~new_new_n11879__ & ~new_new_n11885__;
  assign new_new_n11887__ = new_new_n11599__ & ~new_new_n11886__;
  assign new_new_n11888__ = pi11 & ~new_new_n11887__;
  assign new_new_n11889__ = ~new_new_n11615__ & ~new_new_n11888__;
  assign new_new_n11890__ = ~new_new_n11613__ & ~new_new_n11889__;
  assign new_new_n11891__ = ~pi11 & new_new_n11613__;
  assign new_new_n11892__ = ~new_new_n11604__ & ~new_new_n11891__;
  assign new_new_n11893__ = new_new_n11886__ & ~new_new_n11892__;
  assign new_new_n11894__ = ~new_new_n11614__ & ~new_new_n11893__;
  assign new_new_n11895__ = ~new_new_n11890__ & new_new_n11894__;
  assign new_new_n11896__ = ~new_new_n11592__ & ~new_new_n11895__;
  assign new_new_n11897__ = pi11 & new_new_n11604__;
  assign new_new_n11898__ = pi11 & ~new_new_n11599__;
  assign new_new_n11899__ = ~new_new_n11615__ & ~new_new_n11898__;
  assign new_new_n11900__ = new_new_n11886__ & ~new_new_n11899__;
  assign new_new_n11901__ = ~new_new_n11897__ & ~new_new_n11900__;
  assign new_new_n11902__ = ~new_new_n11613__ & ~new_new_n11901__;
  assign new_new_n11903__ = ~pi11 & new_new_n11604__;
  assign new_new_n11904__ = ~new_new_n11606__ & new_new_n11886__;
  assign new_new_n11905__ = ~new_new_n11903__ & ~new_new_n11904__;
  assign new_new_n11906__ = new_new_n11613__ & ~new_new_n11905__;
  assign new_new_n11907__ = ~new_new_n11902__ & ~new_new_n11906__;
  assign new_new_n11908__ = ~new_new_n11896__ & new_new_n11907__;
  assign new_new_n11909__ = ~new_new_n11588__ & ~new_new_n11908__;
  assign new_new_n11910__ = ~new_new_n11587__ & ~new_new_n11909__;
  assign new_new_n11911__ = new_new_n11572__ & ~new_new_n11910__;
  assign new_new_n11912__ = new_new_n6854__ & new_new_n8470__;
  assign new_new_n11913__ = ~new_new_n2130__ & new_new_n8474__;
  assign new_new_n11914__ = ~new_new_n2024__ & ~new_new_n8479__;
  assign new_new_n11915__ = ~new_new_n11913__ & ~new_new_n11914__;
  assign new_new_n11916__ = ~new_new_n11912__ & new_new_n11915__;
  assign new_new_n11917__ = ~new_new_n3535__ & new_new_n8469__;
  assign new_new_n11918__ = ~pi11 & ~new_new_n11917__;
  assign new_new_n11919__ = ~new_new_n3535__ & new_new_n11530__;
  assign new_new_n11920__ = ~new_new_n11918__ & ~new_new_n11919__;
  assign new_new_n11921__ = new_new_n11916__ & ~new_new_n11920__;
  assign new_new_n11922__ = pi11 & ~new_new_n11916__;
  assign new_new_n11923__ = ~new_new_n11921__ & ~new_new_n11922__;
  assign new_new_n11924__ = ~new_new_n11911__ & new_new_n11923__;
  assign new_new_n11925__ = ~new_new_n11563__ & ~new_new_n11567__;
  assign new_new_n11926__ = ~new_new_n11572__ & new_new_n11910__;
  assign new_new_n11927__ = ~new_new_n11925__ & ~new_new_n11926__;
  assign new_new_n11928__ = ~new_new_n11924__ & new_new_n11927__;
  assign new_new_n11929__ = ~new_new_n11568__ & ~new_new_n11928__;
  assign new_new_n11930__ = ~new_new_n3535__ & ~new_new_n8479__;
  assign new_new_n11931__ = ~new_new_n1902__ & new_new_n8858__;
  assign new_new_n11932__ = ~new_new_n1823__ & new_new_n8474__;
  assign new_new_n11933__ = ~new_new_n11930__ & ~new_new_n11931__;
  assign new_new_n11934__ = ~new_new_n11932__ & new_new_n11933__;
  assign new_new_n11935__ = ~new_new_n6487__ & new_new_n8469__;
  assign new_new_n11936__ = pi11 & ~new_new_n11935__;
  assign new_new_n11937__ = ~new_new_n6487__ & new_new_n11530__;
  assign new_new_n11938__ = ~new_new_n11936__ & ~new_new_n11937__;
  assign new_new_n11939__ = new_new_n11934__ & ~new_new_n11938__;
  assign new_new_n11940__ = ~pi11 & ~new_new_n11934__;
  assign new_new_n11941__ = ~new_new_n11939__ & ~new_new_n11940__;
  assign new_new_n11942__ = new_new_n11929__ & ~new_new_n11941__;
  assign new_new_n11943__ = ~new_new_n11929__ & new_new_n11941__;
  assign new_new_n11944__ = ~new_new_n11203__ & ~new_new_n11204__;
  assign new_new_n11945__ = ~new_new_n11219__ & new_new_n11944__;
  assign new_new_n11946__ = new_new_n11219__ & ~new_new_n11944__;
  assign new_new_n11947__ = ~new_new_n11945__ & ~new_new_n11946__;
  assign new_new_n11948__ = ~new_new_n11943__ & ~new_new_n11947__;
  assign new_new_n11949__ = ~new_new_n11942__ & ~new_new_n11948__;
  assign new_new_n11950__ = ~new_new_n11222__ & ~new_new_n11223__;
  assign new_new_n11951__ = new_new_n11227__ & new_new_n11950__;
  assign new_new_n11952__ = ~new_new_n11227__ & ~new_new_n11950__;
  assign new_new_n11953__ = ~new_new_n11951__ & ~new_new_n11952__;
  assign new_new_n11954__ = ~new_new_n11949__ & ~new_new_n11953__;
  assign new_new_n11955__ = new_new_n11949__ & new_new_n11953__;
  assign new_new_n11956__ = ~new_new_n1823__ & ~new_new_n8479__;
  assign new_new_n11957__ = ~new_new_n1902__ & new_new_n8474__;
  assign new_new_n11958__ = ~new_new_n1660__ & new_new_n8858__;
  assign new_new_n11959__ = ~new_new_n11956__ & ~new_new_n11957__;
  assign new_new_n11960__ = ~new_new_n11958__ & new_new_n11959__;
  assign new_new_n11961__ = ~new_new_n5274__ & new_new_n8469__;
  assign new_new_n11962__ = pi11 & ~new_new_n11961__;
  assign new_new_n11963__ = ~new_new_n5274__ & new_new_n11530__;
  assign new_new_n11964__ = ~new_new_n11962__ & ~new_new_n11963__;
  assign new_new_n11965__ = new_new_n11960__ & ~new_new_n11964__;
  assign new_new_n11966__ = ~pi11 & ~new_new_n11960__;
  assign new_new_n11967__ = ~new_new_n11965__ & ~new_new_n11966__;
  assign new_new_n11968__ = ~new_new_n11955__ & ~new_new_n11967__;
  assign new_new_n11969__ = ~new_new_n11954__ & ~new_new_n11968__;
  assign new_new_n11970__ = ~new_new_n1902__ & ~new_new_n8479__;
  assign new_new_n11971__ = ~new_new_n1660__ & new_new_n8474__;
  assign new_new_n11972__ = ~new_new_n1737__ & new_new_n8858__;
  assign new_new_n11973__ = ~new_new_n11970__ & ~new_new_n11971__;
  assign new_new_n11974__ = ~new_new_n11972__ & new_new_n11973__;
  assign new_new_n11975__ = new_new_n5688__ & new_new_n8469__;
  assign new_new_n11976__ = pi11 & ~new_new_n11975__;
  assign new_new_n11977__ = new_new_n5688__ & new_new_n11530__;
  assign new_new_n11978__ = ~new_new_n11976__ & ~new_new_n11977__;
  assign new_new_n11979__ = new_new_n11974__ & ~new_new_n11978__;
  assign new_new_n11980__ = ~pi11 & ~new_new_n11974__;
  assign new_new_n11981__ = ~new_new_n11979__ & ~new_new_n11980__;
  assign new_new_n11982__ = new_new_n11969__ & new_new_n11981__;
  assign new_new_n11983__ = ~new_new_n11969__ & ~new_new_n11981__;
  assign new_new_n11984__ = ~new_new_n11230__ & ~new_new_n11231__;
  assign new_new_n11985__ = ~new_new_n11246__ & new_new_n11984__;
  assign new_new_n11986__ = new_new_n11246__ & ~new_new_n11984__;
  assign new_new_n11987__ = ~new_new_n11985__ & ~new_new_n11986__;
  assign new_new_n11988__ = ~new_new_n11983__ & ~new_new_n11987__;
  assign new_new_n11989__ = ~new_new_n11982__ & ~new_new_n11988__;
  assign new_new_n11990__ = new_new_n11547__ & ~new_new_n11989__;
  assign new_new_n11991__ = ~new_new_n11547__ & new_new_n11989__;
  assign new_new_n11992__ = pi14 & ~new_new_n10601__;
  assign new_new_n11993__ = ~pi14 & new_new_n10601__;
  assign new_new_n11994__ = ~new_new_n11992__ & ~new_new_n11993__;
  assign new_new_n11995__ = new_new_n11248__ & new_new_n11994__;
  assign new_new_n11996__ = ~new_new_n11248__ & ~new_new_n11994__;
  assign new_new_n11997__ = ~new_new_n11995__ & ~new_new_n11996__;
  assign new_new_n11998__ = new_new_n11251__ & ~new_new_n11997__;
  assign new_new_n11999__ = ~new_new_n11251__ & new_new_n11997__;
  assign new_new_n12000__ = ~new_new_n11998__ & ~new_new_n11999__;
  assign new_new_n12001__ = new_new_n10778__ & new_new_n12000__;
  assign new_new_n12002__ = ~new_new_n10778__ & ~new_new_n12000__;
  assign new_new_n12003__ = ~new_new_n12001__ & ~new_new_n12002__;
  assign new_new_n12004__ = ~new_new_n11991__ & new_new_n12003__;
  assign new_new_n12005__ = ~new_new_n11990__ & ~new_new_n12004__;
  assign new_new_n12006__ = ~new_new_n11257__ & ~new_new_n11258__;
  assign new_new_n12007__ = new_new_n11275__ & new_new_n12006__;
  assign new_new_n12008__ = ~new_new_n11275__ & ~new_new_n12006__;
  assign new_new_n12009__ = ~new_new_n12007__ & ~new_new_n12008__;
  assign new_new_n12010__ = new_new_n12005__ & ~new_new_n12009__;
  assign new_new_n12011__ = ~new_new_n12005__ & new_new_n12009__;
  assign new_new_n12012__ = ~new_new_n1737__ & ~new_new_n8479__;
  assign new_new_n12013__ = ~new_new_n1466__ & new_new_n8474__;
  assign new_new_n12014__ = ~new_new_n1556__ & new_new_n8858__;
  assign new_new_n12015__ = ~new_new_n12012__ & ~new_new_n12013__;
  assign new_new_n12016__ = ~new_new_n12014__ & new_new_n12015__;
  assign new_new_n12017__ = ~new_new_n5671__ & new_new_n8469__;
  assign new_new_n12018__ = pi11 & ~new_new_n12017__;
  assign new_new_n12019__ = ~new_new_n5671__ & new_new_n11530__;
  assign new_new_n12020__ = ~new_new_n12018__ & ~new_new_n12019__;
  assign new_new_n12021__ = new_new_n12016__ & ~new_new_n12020__;
  assign new_new_n12022__ = ~pi11 & ~new_new_n12016__;
  assign new_new_n12023__ = ~new_new_n12021__ & ~new_new_n12022__;
  assign new_new_n12024__ = ~new_new_n12011__ & ~new_new_n12023__;
  assign new_new_n12025__ = ~new_new_n12010__ & ~new_new_n12024__;
  assign new_new_n12026__ = ~new_new_n11535__ & ~new_new_n12025__;
  assign new_new_n12027__ = new_new_n11535__ & new_new_n12025__;
  assign new_new_n12028__ = ~new_new_n11295__ & new_new_n11299__;
  assign new_new_n12029__ = ~new_new_n11300__ & ~new_new_n12028__;
  assign new_new_n12030__ = ~new_new_n12027__ & ~new_new_n12029__;
  assign new_new_n12031__ = ~new_new_n12026__ & ~new_new_n12030__;
  assign new_new_n12032__ = ~new_new_n11522__ & ~new_new_n12031__;
  assign new_new_n12033__ = new_new_n11522__ & new_new_n12031__;
  assign new_new_n12034__ = ~new_new_n11313__ & ~new_new_n11314__;
  assign new_new_n12035__ = new_new_n11329__ & ~new_new_n12034__;
  assign new_new_n12036__ = ~new_new_n11329__ & new_new_n12034__;
  assign new_new_n12037__ = ~new_new_n12035__ & ~new_new_n12036__;
  assign new_new_n12038__ = ~new_new_n12033__ & ~new_new_n12037__;
  assign new_new_n12039__ = ~new_new_n12032__ & ~new_new_n12038__;
  assign new_new_n12040__ = ~new_new_n10762__ & ~new_new_n10763__;
  assign new_new_n12041__ = ~new_new_n11331__ & new_new_n12040__;
  assign new_new_n12042__ = new_new_n11331__ & ~new_new_n12040__;
  assign new_new_n12043__ = ~new_new_n12041__ & ~new_new_n12042__;
  assign new_new_n12044__ = new_new_n12039__ & new_new_n12043__;
  assign new_new_n12045__ = ~new_new_n12039__ & ~new_new_n12043__;
  assign new_new_n12046__ = ~new_new_n3618__ & new_new_n8474__;
  assign new_new_n12047__ = ~new_new_n1061__ & new_new_n8858__;
  assign new_new_n12048__ = ~new_new_n1325__ & ~new_new_n8479__;
  assign new_new_n12049__ = new_new_n4926__ & new_new_n8470__;
  assign new_new_n12050__ = ~new_new_n12046__ & ~new_new_n12047__;
  assign new_new_n12051__ = ~new_new_n12048__ & new_new_n12050__;
  assign new_new_n12052__ = ~new_new_n12049__ & new_new_n12051__;
  assign new_new_n12053__ = pi11 & ~new_new_n12052__;
  assign new_new_n12054__ = ~pi11 & new_new_n12052__;
  assign new_new_n12055__ = ~new_new_n12053__ & ~new_new_n12054__;
  assign new_new_n12056__ = ~new_new_n12045__ & ~new_new_n12055__;
  assign new_new_n12057__ = ~new_new_n12044__ & ~new_new_n12056__;
  assign new_new_n12058__ = ~new_new_n11507__ & ~new_new_n12057__;
  assign new_new_n12059__ = new_new_n11507__ & new_new_n12057__;
  assign new_new_n12060__ = ~new_new_n1207__ & new_new_n8858__;
  assign new_new_n12061__ = ~new_new_n1061__ & new_new_n8474__;
  assign new_new_n12062__ = ~new_new_n3618__ & ~new_new_n8479__;
  assign new_new_n12063__ = ~new_new_n5235__ & new_new_n8470__;
  assign new_new_n12064__ = ~new_new_n12060__ & ~new_new_n12061__;
  assign new_new_n12065__ = ~new_new_n12062__ & new_new_n12064__;
  assign new_new_n12066__ = ~new_new_n12063__ & new_new_n12065__;
  assign new_new_n12067__ = pi11 & ~new_new_n12066__;
  assign new_new_n12068__ = ~pi11 & new_new_n12066__;
  assign new_new_n12069__ = ~new_new_n12067__ & ~new_new_n12068__;
  assign new_new_n12070__ = ~new_new_n12059__ & ~new_new_n12069__;
  assign new_new_n12071__ = ~new_new_n12058__ & ~new_new_n12070__;
  assign new_new_n12072__ = ~new_new_n11503__ & new_new_n12071__;
  assign new_new_n12073__ = new_new_n11503__ & ~new_new_n12071__;
  assign new_new_n12074__ = ~new_new_n12072__ & ~new_new_n12073__;
  assign new_new_n12075__ = ~new_new_n11359__ & ~new_new_n11360__;
  assign new_new_n12076__ = new_new_n11373__ & new_new_n12075__;
  assign new_new_n12077__ = ~new_new_n11373__ & ~new_new_n12075__;
  assign new_new_n12078__ = ~new_new_n12076__ & ~new_new_n12077__;
  assign new_new_n12079__ = new_new_n12074__ & new_new_n12078__;
  assign new_new_n12080__ = ~new_new_n12074__ & ~new_new_n12078__;
  assign new_new_n12081__ = ~new_new_n12079__ & ~new_new_n12080__;
  assign new_new_n12082__ = ~new_new_n11490__ & new_new_n12081__;
  assign new_new_n12083__ = new_new_n11490__ & ~new_new_n12081__;
  assign new_new_n12084__ = ~new_new_n12032__ & ~new_new_n12033__;
  assign new_new_n12085__ = new_new_n12037__ & ~new_new_n12084__;
  assign new_new_n12086__ = ~new_new_n12037__ & new_new_n12084__;
  assign new_new_n12087__ = ~new_new_n12085__ & ~new_new_n12086__;
  assign new_new_n12088__ = ~new_new_n12026__ & ~new_new_n12027__;
  assign new_new_n12089__ = new_new_n12029__ & new_new_n12088__;
  assign new_new_n12090__ = ~new_new_n12029__ & ~new_new_n12088__;
  assign new_new_n12091__ = ~new_new_n12089__ & ~new_new_n12090__;
  assign new_new_n12092__ = ~new_new_n1325__ & new_new_n10702__;
  assign new_new_n12093__ = new_new_n8344__ & ~new_new_n10697__;
  assign new_new_n12094__ = ~new_new_n3618__ & new_new_n10697__;
  assign new_new_n12095__ = ~new_new_n5981__ & ~new_new_n12094__;
  assign new_new_n12096__ = ~new_new_n12093__ & new_new_n12095__;
  assign new_new_n12097__ = new_new_n10694__ & ~new_new_n12096__;
  assign new_new_n12098__ = ~new_new_n12092__ & ~new_new_n12097__;
  assign new_new_n12099__ = ~new_new_n1556__ & new_new_n10709__;
  assign new_new_n12100__ = pi08 & ~new_new_n12099__;
  assign new_new_n12101__ = ~new_new_n1556__ & new_new_n10712__;
  assign new_new_n12102__ = ~pi08 & ~new_new_n12101__;
  assign new_new_n12103__ = pi05 & ~new_new_n12102__;
  assign new_new_n12104__ = ~new_new_n12100__ & ~new_new_n12103__;
  assign new_new_n12105__ = new_new_n12098__ & ~new_new_n12104__;
  assign new_new_n12106__ = ~pi08 & ~new_new_n12098__;
  assign new_new_n12107__ = ~new_new_n12105__ & ~new_new_n12106__;
  assign new_new_n12108__ = ~new_new_n11990__ & ~new_new_n11991__;
  assign new_new_n12109__ = new_new_n12003__ & new_new_n12108__;
  assign new_new_n12110__ = ~new_new_n12003__ & ~new_new_n12108__;
  assign new_new_n12111__ = ~new_new_n12109__ & ~new_new_n12110__;
  assign new_new_n12112__ = ~new_new_n12107__ & ~new_new_n12111__;
  assign new_new_n12113__ = new_new_n12107__ & new_new_n12111__;
  assign new_new_n12114__ = ~new_new_n1466__ & new_new_n10698__;
  assign new_new_n12115__ = ~new_new_n1660__ & ~new_new_n11409__;
  assign new_new_n12116__ = ~new_new_n1737__ & new_new_n10702__;
  assign new_new_n12117__ = ~new_new_n12114__ & ~new_new_n12115__;
  assign new_new_n12118__ = ~new_new_n12116__ & new_new_n12117__;
  assign new_new_n12119__ = ~new_new_n6410__ & new_new_n10694__;
  assign new_new_n12120__ = ~pi08 & ~new_new_n12119__;
  assign new_new_n12121__ = ~pi07 & new_new_n10694__;
  assign new_new_n12122__ = ~new_new_n6410__ & new_new_n12121__;
  assign new_new_n12123__ = ~new_new_n12120__ & ~new_new_n12122__;
  assign new_new_n12124__ = new_new_n12118__ & ~new_new_n12123__;
  assign new_new_n12125__ = pi08 & ~new_new_n12118__;
  assign new_new_n12126__ = ~new_new_n12124__ & ~new_new_n12125__;
  assign new_new_n12127__ = ~new_new_n11942__ & ~new_new_n11943__;
  assign new_new_n12128__ = new_new_n11947__ & ~new_new_n12127__;
  assign new_new_n12129__ = ~new_new_n11947__ & new_new_n12127__;
  assign new_new_n12130__ = ~new_new_n12128__ & ~new_new_n12129__;
  assign new_new_n12131__ = ~new_new_n12126__ & ~new_new_n12130__;
  assign new_new_n12132__ = ~new_new_n11568__ & new_new_n11928__;
  assign new_new_n12133__ = ~new_new_n11572__ & new_new_n11925__;
  assign new_new_n12134__ = new_new_n11568__ & new_new_n11923__;
  assign new_new_n12135__ = ~new_new_n12133__ & ~new_new_n12134__;
  assign new_new_n12136__ = new_new_n11910__ & ~new_new_n12135__;
  assign new_new_n12137__ = ~new_new_n11911__ & ~new_new_n11926__;
  assign new_new_n12138__ = ~new_new_n11923__ & new_new_n12137__;
  assign new_new_n12139__ = new_new_n11923__ & ~new_new_n12137__;
  assign new_new_n12140__ = ~new_new_n12138__ & ~new_new_n12139__;
  assign new_new_n12141__ = new_new_n11568__ & ~new_new_n11572__;
  assign new_new_n12142__ = new_new_n11923__ & new_new_n11925__;
  assign new_new_n12143__ = ~new_new_n12141__ & ~new_new_n12142__;
  assign new_new_n12144__ = new_new_n12140__ & ~new_new_n12143__;
  assign new_new_n12145__ = ~new_new_n12132__ & ~new_new_n12136__;
  assign new_new_n12146__ = ~new_new_n12144__ & new_new_n12145__;
  assign new_new_n12147__ = ~new_new_n6487__ & new_new_n11378__;
  assign new_new_n12148__ = ~new_new_n3535__ & ~new_new_n11409__;
  assign new_new_n12149__ = ~new_new_n1823__ & new_new_n10702__;
  assign new_new_n12150__ = ~new_new_n12148__ & ~new_new_n12149__;
  assign new_new_n12151__ = ~new_new_n12147__ & new_new_n12150__;
  assign new_new_n12152__ = ~new_new_n1902__ & new_new_n10694__;
  assign new_new_n12153__ = ~pi08 & ~new_new_n12152__;
  assign new_new_n12154__ = ~new_new_n1902__ & new_new_n11498__;
  assign new_new_n12155__ = ~new_new_n12153__ & ~new_new_n12154__;
  assign new_new_n12156__ = new_new_n12151__ & ~new_new_n12155__;
  assign new_new_n12157__ = pi08 & ~new_new_n12151__;
  assign new_new_n12158__ = ~new_new_n12156__ & ~new_new_n12157__;
  assign new_new_n12159__ = new_new_n11592__ & ~new_new_n11886__;
  assign new_new_n12160__ = new_new_n11604__ & ~new_new_n12159__;
  assign new_new_n12161__ = ~new_new_n11592__ & new_new_n11886__;
  assign new_new_n12162__ = ~new_new_n11604__ & ~new_new_n12161__;
  assign new_new_n12163__ = pi11 & ~new_new_n11613__;
  assign new_new_n12164__ = ~new_new_n11891__ & ~new_new_n12163__;
  assign new_new_n12165__ = ~new_new_n12160__ & ~new_new_n12164__;
  assign new_new_n12166__ = ~new_new_n12162__ & new_new_n12165__;
  assign new_new_n12167__ = ~new_new_n11604__ & ~new_new_n12159__;
  assign new_new_n12168__ = new_new_n11604__ & ~new_new_n12161__;
  assign new_new_n12169__ = new_new_n12164__ & ~new_new_n12167__;
  assign new_new_n12170__ = ~new_new_n12168__ & new_new_n12169__;
  assign new_new_n12171__ = ~new_new_n12159__ & ~new_new_n12161__;
  assign new_new_n12172__ = new_new_n11599__ & ~new_new_n11604__;
  assign new_new_n12173__ = ~new_new_n11605__ & ~new_new_n12172__;
  assign new_new_n12174__ = new_new_n11613__ & new_new_n12173__;
  assign new_new_n12175__ = ~new_new_n11613__ & ~new_new_n12173__;
  assign new_new_n12176__ = ~new_new_n12174__ & ~new_new_n12175__;
  assign new_new_n12177__ = new_new_n12171__ & new_new_n12176__;
  assign new_new_n12178__ = ~new_new_n12166__ & ~new_new_n12177__;
  assign new_new_n12179__ = ~new_new_n12170__ & new_new_n12178__;
  assign new_new_n12180__ = ~new_new_n11600__ & ~new_new_n11898__;
  assign new_new_n12181__ = new_new_n12171__ & new_new_n12180__;
  assign new_new_n12182__ = ~new_new_n12171__ & ~new_new_n12180__;
  assign new_new_n12183__ = ~new_new_n12181__ & ~new_new_n12182__;
  assign new_new_n12184__ = ~new_new_n11879__ & ~new_new_n11880__;
  assign new_new_n12185__ = new_new_n11884__ & new_new_n12184__;
  assign new_new_n12186__ = ~new_new_n11884__ & ~new_new_n12184__;
  assign new_new_n12187__ = ~new_new_n12185__ & ~new_new_n12186__;
  assign new_new_n12188__ = ~pi14 & new_new_n11865__;
  assign new_new_n12189__ = pi14 & ~new_new_n11865__;
  assign new_new_n12190__ = ~new_new_n12188__ & ~new_new_n12189__;
  assign new_new_n12191__ = new_new_n11853__ & ~new_new_n12190__;
  assign new_new_n12192__ = ~new_new_n11853__ & new_new_n12190__;
  assign new_new_n12193__ = ~new_new_n12191__ & ~new_new_n12192__;
  assign new_new_n12194__ = new_new_n11113__ & ~new_new_n11124__;
  assign new_new_n12195__ = ~new_new_n11113__ & new_new_n11127__;
  assign new_new_n12196__ = ~new_new_n12194__ & ~new_new_n12195__;
  assign new_new_n12197__ = new_new_n10913__ & ~new_new_n12196__;
  assign new_new_n12198__ = ~new_new_n10913__ & new_new_n12196__;
  assign new_new_n12199__ = ~new_new_n12197__ & ~new_new_n12198__;
  assign new_new_n12200__ = new_new_n12193__ & new_new_n12199__;
  assign new_new_n12201__ = ~new_new_n12193__ & ~new_new_n12199__;
  assign new_new_n12202__ = ~new_new_n12200__ & ~new_new_n12201__;
  assign new_new_n12203__ = ~new_new_n11840__ & ~new_new_n11841__;
  assign new_new_n12204__ = new_new_n11851__ & new_new_n12203__;
  assign new_new_n12205__ = ~new_new_n11851__ & ~new_new_n12203__;
  assign new_new_n12206__ = ~new_new_n12204__ & ~new_new_n12205__;
  assign new_new_n12207__ = ~new_new_n11650__ & ~new_new_n11809__;
  assign new_new_n12208__ = new_new_n11650__ & new_new_n11809__;
  assign new_new_n12209__ = ~new_new_n12207__ & ~new_new_n12208__;
  assign new_new_n12210__ = ~new_new_n11670__ & ~new_new_n11674__;
  assign new_new_n12211__ = ~new_new_n11658__ & new_new_n12210__;
  assign new_new_n12212__ = new_new_n11658__ & ~new_new_n12210__;
  assign new_new_n12213__ = ~new_new_n12211__ & ~new_new_n12212__;
  assign new_new_n12214__ = new_new_n12209__ & new_new_n12213__;
  assign new_new_n12215__ = pi11 & new_new_n11658__;
  assign new_new_n12216__ = ~new_new_n11814__ & ~new_new_n12215__;
  assign new_new_n12217__ = ~new_new_n11662__ & ~new_new_n12208__;
  assign new_new_n12218__ = new_new_n11662__ & ~new_new_n12207__;
  assign new_new_n12219__ = new_new_n12216__ & ~new_new_n12217__;
  assign new_new_n12220__ = ~new_new_n12218__ & new_new_n12219__;
  assign new_new_n12221__ = new_new_n11662__ & ~new_new_n12208__;
  assign new_new_n12222__ = ~new_new_n11662__ & ~new_new_n12207__;
  assign new_new_n12223__ = ~new_new_n12216__ & ~new_new_n12221__;
  assign new_new_n12224__ = ~new_new_n12222__ & new_new_n12223__;
  assign new_new_n12225__ = ~new_new_n12214__ & ~new_new_n12220__;
  assign new_new_n12226__ = ~new_new_n12224__ & new_new_n12225__;
  assign new_new_n12227__ = ~new_new_n7236__ & new_new_n11378__;
  assign new_new_n12228__ = ~new_new_n2497__ & ~new_new_n11409__;
  assign new_new_n12229__ = ~new_new_n2572__ & new_new_n10702__;
  assign new_new_n12230__ = ~new_new_n12228__ & ~new_new_n12229__;
  assign new_new_n12231__ = ~new_new_n12227__ & new_new_n12230__;
  assign new_new_n12232__ = ~new_new_n2313__ & new_new_n10694__;
  assign new_new_n12233__ = ~pi08 & ~new_new_n12232__;
  assign new_new_n12234__ = ~new_new_n2313__ & new_new_n11498__;
  assign new_new_n12235__ = ~new_new_n12233__ & ~new_new_n12234__;
  assign new_new_n12236__ = new_new_n12231__ & ~new_new_n12235__;
  assign new_new_n12237__ = pi08 & ~new_new_n12231__;
  assign new_new_n12238__ = ~new_new_n12236__ & ~new_new_n12237__;
  assign new_new_n12239__ = new_new_n12226__ & ~new_new_n12238__;
  assign new_new_n12240__ = ~new_new_n12226__ & new_new_n12238__;
  assign new_new_n12241__ = ~new_new_n11793__ & new_new_n11797__;
  assign new_new_n12242__ = ~new_new_n11003__ & new_new_n11733__;
  assign new_new_n12243__ = ~new_new_n11787__ & ~new_new_n12242__;
  assign new_new_n12244__ = ~new_new_n11797__ & ~new_new_n12243__;
  assign new_new_n12245__ = ~new_new_n11012__ & new_new_n11791__;
  assign new_new_n12246__ = ~new_new_n11792__ & ~new_new_n12245__;
  assign new_new_n12247__ = ~new_new_n12244__ & new_new_n12246__;
  assign new_new_n12248__ = ~new_new_n12241__ & ~new_new_n12247__;
  assign new_new_n12249__ = ~new_new_n11774__ & ~new_new_n11775__;
  assign new_new_n12250__ = ~new_new_n11785__ & ~new_new_n12249__;
  assign new_new_n12251__ = new_new_n11785__ & new_new_n12249__;
  assign new_new_n12252__ = ~new_new_n12250__ & ~new_new_n12251__;
  assign new_new_n12253__ = ~new_new_n2960__ & new_new_n10698__;
  assign new_new_n12254__ = ~new_new_n3164__ & ~new_new_n11409__;
  assign new_new_n12255__ = ~new_new_n3126__ & new_new_n10702__;
  assign new_new_n12256__ = ~new_new_n12254__ & ~new_new_n12255__;
  assign new_new_n12257__ = ~new_new_n12253__ & new_new_n12256__;
  assign new_new_n12258__ = ~new_new_n7468__ & new_new_n10694__;
  assign new_new_n12259__ = ~pi08 & ~new_new_n12258__;
  assign new_new_n12260__ = ~new_new_n7468__ & new_new_n12121__;
  assign new_new_n12261__ = ~new_new_n12259__ & ~new_new_n12260__;
  assign new_new_n12262__ = new_new_n12257__ & ~new_new_n12261__;
  assign new_new_n12263__ = pi08 & ~new_new_n12257__;
  assign new_new_n12264__ = ~new_new_n12262__ & ~new_new_n12263__;
  assign new_new_n12265__ = ~new_new_n3356__ & new_new_n11746__;
  assign new_new_n12266__ = ~new_new_n8306__ & ~new_new_n12265__;
  assign new_new_n12267__ = pi10 & ~new_new_n12266__;
  assign new_new_n12268__ = ~new_new_n3356__ & ~new_new_n8473__;
  assign new_new_n12269__ = ~new_new_n11747__ & ~new_new_n12268__;
  assign new_new_n12270__ = ~new_new_n12267__ & ~new_new_n12269__;
  assign new_new_n12271__ = ~pi06 & pi07;
  assign new_new_n12272__ = ~pi05 & new_new_n12271__;
  assign new_new_n12273__ = pi06 & ~pi07;
  assign new_new_n12274__ = pi05 & new_new_n12273__;
  assign new_new_n12275__ = ~new_new_n12272__ & ~new_new_n12274__;
  assign new_new_n12276__ = ~new_new_n10694__ & new_new_n12275__;
  assign new_new_n12277__ = ~new_new_n3055__ & new_new_n10694__;
  assign new_new_n12278__ = new_new_n3356__ & ~new_new_n12277__;
  assign new_new_n12279__ = ~new_new_n12276__ & ~new_new_n12278__;
  assign new_new_n12280__ = new_new_n7682__ & new_new_n11378__;
  assign new_new_n12281__ = new_new_n12275__ & ~new_new_n12280__;
  assign new_new_n12282__ = ~new_new_n3055__ & ~new_new_n12281__;
  assign new_new_n12283__ = ~new_new_n3254__ & new_new_n10694__;
  assign new_new_n12284__ = ~new_new_n3356__ & ~new_new_n11409__;
  assign new_new_n12285__ = ~new_new_n12283__ & ~new_new_n12284__;
  assign new_new_n12286__ = ~new_new_n3055__ & ~new_new_n10697__;
  assign new_new_n12287__ = new_new_n3356__ & new_new_n12286__;
  assign new_new_n12288__ = ~new_new_n12285__ & ~new_new_n12287__;
  assign new_new_n12289__ = ~new_new_n12282__ & ~new_new_n12288__;
  assign new_new_n12290__ = pi08 & ~new_new_n12279__;
  assign new_new_n12291__ = new_new_n12289__ & new_new_n12290__;
  assign new_new_n12292__ = ~new_new_n8637__ & new_new_n11378__;
  assign new_new_n12293__ = ~new_new_n3164__ & new_new_n10698__;
  assign new_new_n12294__ = ~new_new_n3055__ & ~new_new_n11409__;
  assign new_new_n12295__ = ~new_new_n3254__ & new_new_n10702__;
  assign new_new_n12296__ = ~new_new_n12293__ & ~new_new_n12294__;
  assign new_new_n12297__ = ~new_new_n12295__ & new_new_n12296__;
  assign new_new_n12298__ = ~new_new_n12292__ & new_new_n12297__;
  assign new_new_n12299__ = new_new_n12291__ & new_new_n12298__;
  assign new_new_n12300__ = pi09 & ~new_new_n12298__;
  assign new_new_n12301__ = pi08 & new_new_n12298__;
  assign new_new_n12302__ = ~new_new_n12300__ & ~new_new_n12301__;
  assign new_new_n12303__ = new_new_n11744__ & ~new_new_n12302__;
  assign new_new_n12304__ = ~new_new_n12299__ & ~new_new_n12303__;
  assign new_new_n12305__ = ~new_new_n12270__ & new_new_n12304__;
  assign new_new_n12306__ = new_new_n12270__ & ~new_new_n12304__;
  assign new_new_n12307__ = ~new_new_n3254__ & ~new_new_n11409__;
  assign new_new_n12308__ = ~new_new_n3164__ & new_new_n10702__;
  assign new_new_n12309__ = ~new_new_n3126__ & new_new_n10698__;
  assign new_new_n12310__ = ~new_new_n7570__ & new_new_n11378__;
  assign new_new_n12311__ = ~new_new_n12307__ & ~new_new_n12308__;
  assign new_new_n12312__ = ~new_new_n12309__ & new_new_n12311__;
  assign new_new_n12313__ = ~new_new_n12310__ & new_new_n12312__;
  assign new_new_n12314__ = pi08 & ~new_new_n12313__;
  assign new_new_n12315__ = ~pi08 & new_new_n12313__;
  assign new_new_n12316__ = ~new_new_n12314__ & ~new_new_n12315__;
  assign new_new_n12317__ = ~new_new_n12306__ & ~new_new_n12316__;
  assign new_new_n12318__ = ~new_new_n12305__ & ~new_new_n12317__;
  assign new_new_n12319__ = ~new_new_n12264__ & ~new_new_n12318__;
  assign new_new_n12320__ = ~pi11 & ~new_new_n11743__;
  assign new_new_n12321__ = pi11 & new_new_n11743__;
  assign new_new_n12322__ = ~new_new_n12320__ & ~new_new_n12321__;
  assign new_new_n12323__ = ~new_new_n11751__ & ~new_new_n12322__;
  assign new_new_n12324__ = ~new_new_n12319__ & new_new_n12323__;
  assign new_new_n12325__ = ~new_new_n11743__ & ~new_new_n11750__;
  assign new_new_n12326__ = ~new_new_n12318__ & ~new_new_n12325__;
  assign new_new_n12327__ = new_new_n12264__ & ~new_new_n12326__;
  assign new_new_n12328__ = ~new_new_n12324__ & ~new_new_n12327__;
  assign new_new_n12329__ = ~pi12 & ~new_new_n3356__;
  assign new_new_n12330__ = new_new_n11752__ & new_new_n12329__;
  assign new_new_n12331__ = ~pi11 & new_new_n3356__;
  assign new_new_n12332__ = ~new_new_n12329__ & ~new_new_n12331__;
  assign new_new_n12333__ = ~new_new_n11752__ & new_new_n12332__;
  assign new_new_n12334__ = new_new_n11759__ & new_new_n12333__;
  assign new_new_n12335__ = ~new_new_n11759__ & ~new_new_n12333__;
  assign new_new_n12336__ = ~new_new_n12330__ & ~new_new_n12334__;
  assign new_new_n12337__ = ~new_new_n12335__ & new_new_n12336__;
  assign new_new_n12338__ = ~new_new_n12328__ & ~new_new_n12337__;
  assign new_new_n12339__ = new_new_n12328__ & new_new_n12337__;
  assign new_new_n12340__ = ~new_new_n3460__ & new_new_n10698__;
  assign new_new_n12341__ = ~new_new_n7388__ & new_new_n10697__;
  assign new_new_n12342__ = new_new_n10694__ & ~new_new_n12341__;
  assign new_new_n12343__ = new_new_n7391__ & new_new_n12342__;
  assign new_new_n12344__ = ~new_new_n3126__ & ~new_new_n11409__;
  assign new_new_n12345__ = ~new_new_n2960__ & new_new_n10702__;
  assign new_new_n12346__ = ~new_new_n12340__ & ~new_new_n12344__;
  assign new_new_n12347__ = ~new_new_n12345__ & new_new_n12346__;
  assign new_new_n12348__ = ~new_new_n12343__ & new_new_n12347__;
  assign new_new_n12349__ = ~pi08 & ~new_new_n12348__;
  assign new_new_n12350__ = pi08 & new_new_n12348__;
  assign new_new_n12351__ = ~new_new_n12349__ & ~new_new_n12350__;
  assign new_new_n12352__ = ~new_new_n12339__ & ~new_new_n12351__;
  assign new_new_n12353__ = ~new_new_n12338__ & ~new_new_n12352__;
  assign new_new_n12354__ = ~new_new_n12252__ & new_new_n12353__;
  assign new_new_n12355__ = new_new_n12252__ & ~new_new_n12353__;
  assign new_new_n12356__ = ~new_new_n2960__ & ~new_new_n11409__;
  assign new_new_n12357__ = ~new_new_n2848__ & new_new_n10698__;
  assign new_new_n12358__ = ~new_new_n3460__ & new_new_n10702__;
  assign new_new_n12359__ = ~new_new_n12357__ & ~new_new_n12358__;
  assign new_new_n12360__ = ~new_new_n12356__ & new_new_n12359__;
  assign new_new_n12361__ = ~new_new_n7065__ & new_new_n11378__;
  assign new_new_n12362__ = new_new_n12360__ & ~new_new_n12361__;
  assign new_new_n12363__ = pi08 & ~new_new_n12362__;
  assign new_new_n12364__ = ~pi08 & new_new_n12362__;
  assign new_new_n12365__ = ~new_new_n12363__ & ~new_new_n12364__;
  assign new_new_n12366__ = ~new_new_n12355__ & ~new_new_n12365__;
  assign new_new_n12367__ = ~new_new_n12354__ & ~new_new_n12366__;
  assign new_new_n12368__ = new_new_n12248__ & ~new_new_n12367__;
  assign new_new_n12369__ = ~new_new_n12248__ & new_new_n12367__;
  assign new_new_n12370__ = ~new_new_n3460__ & ~new_new_n11409__;
  assign new_new_n12371__ = ~new_new_n2848__ & new_new_n10702__;
  assign new_new_n12372__ = ~new_new_n2886__ & new_new_n10698__;
  assign new_new_n12373__ = ~new_new_n8574__ & new_new_n11378__;
  assign new_new_n12374__ = ~new_new_n12370__ & ~new_new_n12371__;
  assign new_new_n12375__ = ~new_new_n12372__ & new_new_n12374__;
  assign new_new_n12376__ = ~new_new_n12373__ & new_new_n12375__;
  assign new_new_n12377__ = pi08 & ~new_new_n12376__;
  assign new_new_n12378__ = ~pi08 & new_new_n12376__;
  assign new_new_n12379__ = ~new_new_n12377__ & ~new_new_n12378__;
  assign new_new_n12380__ = ~new_new_n12369__ & ~new_new_n12379__;
  assign new_new_n12381__ = ~new_new_n12368__ & ~new_new_n12380__;
  assign new_new_n12382__ = new_new_n11013__ & ~new_new_n11714__;
  assign new_new_n12383__ = ~new_new_n11013__ & new_new_n11714__;
  assign new_new_n12384__ = ~new_new_n12382__ & ~new_new_n12383__;
  assign new_new_n12385__ = new_new_n11032__ & new_new_n12384__;
  assign new_new_n12386__ = ~new_new_n11032__ & ~new_new_n12384__;
  assign new_new_n12387__ = ~new_new_n12385__ & ~new_new_n12386__;
  assign new_new_n12388__ = new_new_n11014__ & ~new_new_n12387__;
  assign new_new_n12389__ = ~new_new_n11014__ & new_new_n12387__;
  assign new_new_n12390__ = ~new_new_n12388__ & ~new_new_n12389__;
  assign new_new_n12391__ = new_new_n11797__ & new_new_n12390__;
  assign new_new_n12392__ = ~new_new_n11797__ & ~new_new_n12390__;
  assign new_new_n12393__ = ~new_new_n12391__ & ~new_new_n12392__;
  assign new_new_n12394__ = ~new_new_n12381__ & ~new_new_n12393__;
  assign new_new_n12395__ = ~new_new_n2886__ & new_new_n10702__;
  assign new_new_n12396__ = ~new_new_n2848__ & ~new_new_n11409__;
  assign new_new_n12397__ = ~new_new_n2737__ & new_new_n10698__;
  assign new_new_n12398__ = ~new_new_n7378__ & new_new_n11378__;
  assign new_new_n12399__ = ~new_new_n12395__ & ~new_new_n12396__;
  assign new_new_n12400__ = ~new_new_n12397__ & new_new_n12399__;
  assign new_new_n12401__ = ~new_new_n12398__ & new_new_n12400__;
  assign new_new_n12402__ = pi08 & ~new_new_n12401__;
  assign new_new_n12403__ = ~pi08 & new_new_n12401__;
  assign new_new_n12404__ = ~new_new_n12402__ & ~new_new_n12403__;
  assign new_new_n12405__ = new_new_n12381__ & new_new_n12393__;
  assign new_new_n12406__ = ~new_new_n12404__ & ~new_new_n12405__;
  assign new_new_n12407__ = ~new_new_n12394__ & ~new_new_n12406__;
  assign new_new_n12408__ = pi08 & ~new_new_n12121__;
  assign new_new_n12409__ = ~new_new_n2886__ & ~new_new_n11409__;
  assign new_new_n12410__ = ~new_new_n2636__ & new_new_n10698__;
  assign new_new_n12411__ = ~new_new_n2737__ & new_new_n10702__;
  assign new_new_n12412__ = ~new_new_n12409__ & ~new_new_n12410__;
  assign new_new_n12413__ = ~new_new_n12411__ & new_new_n12412__;
  assign new_new_n12414__ = new_new_n12408__ & new_new_n12413__;
  assign new_new_n12415__ = ~pi08 & new_new_n11498__;
  assign new_new_n12416__ = new_new_n2636__ & new_new_n12415__;
  assign new_new_n12417__ = pi08 & ~new_new_n2636__;
  assign new_new_n12418__ = new_new_n12413__ & new_new_n12417__;
  assign new_new_n12419__ = ~new_new_n12416__ & ~new_new_n12418__;
  assign new_new_n12420__ = new_new_n7811__ & ~new_new_n12419__;
  assign new_new_n12421__ = ~new_new_n2636__ & new_new_n12415__;
  assign new_new_n12422__ = pi08 & new_new_n2636__;
  assign new_new_n12423__ = new_new_n12413__ & new_new_n12422__;
  assign new_new_n12424__ = ~new_new_n12421__ & ~new_new_n12423__;
  assign new_new_n12425__ = ~new_new_n7811__ & ~new_new_n12424__;
  assign new_new_n12426__ = ~pi08 & ~new_new_n12413__;
  assign new_new_n12427__ = ~new_new_n12414__ & ~new_new_n12426__;
  assign new_new_n12428__ = ~new_new_n12420__ & new_new_n12427__;
  assign new_new_n12429__ = ~new_new_n12425__ & new_new_n12428__;
  assign new_new_n12430__ = new_new_n12407__ & ~new_new_n12429__;
  assign new_new_n12431__ = ~new_new_n12407__ & new_new_n12429__;
  assign new_new_n12432__ = new_new_n11702__ & ~new_new_n11799__;
  assign new_new_n12433__ = ~new_new_n11702__ & new_new_n11799__;
  assign new_new_n12434__ = ~new_new_n12432__ & ~new_new_n12433__;
  assign new_new_n12435__ = new_new_n11805__ & new_new_n12434__;
  assign new_new_n12436__ = ~new_new_n11805__ & ~new_new_n12434__;
  assign new_new_n12437__ = ~new_new_n12435__ & ~new_new_n12436__;
  assign new_new_n12438__ = ~new_new_n12431__ & ~new_new_n12437__;
  assign new_new_n12439__ = ~new_new_n12430__ & ~new_new_n12438__;
  assign new_new_n12440__ = new_new_n11061__ & new_new_n11801__;
  assign new_new_n12441__ = new_new_n11052__ & ~new_new_n11059__;
  assign new_new_n12442__ = new_new_n11051__ & new_new_n11059__;
  assign new_new_n12443__ = ~new_new_n12441__ & ~new_new_n12442__;
  assign new_new_n12444__ = ~new_new_n12434__ & new_new_n12443__;
  assign new_new_n12445__ = ~new_new_n11061__ & new_new_n11800__;
  assign new_new_n12446__ = ~new_new_n12440__ & ~new_new_n12445__;
  assign new_new_n12447__ = ~new_new_n12444__ & new_new_n12446__;
  assign new_new_n12448__ = ~new_new_n11684__ & ~new_new_n12447__;
  assign new_new_n12449__ = new_new_n11051__ & new_new_n11801__;
  assign new_new_n12450__ = new_new_n11033__ & new_new_n11801__;
  assign new_new_n12451__ = ~new_new_n11033__ & ~new_new_n11801__;
  assign new_new_n12452__ = ~new_new_n11050__ & ~new_new_n11800__;
  assign new_new_n12453__ = ~new_new_n12451__ & new_new_n12452__;
  assign new_new_n12454__ = ~new_new_n12450__ & ~new_new_n12453__;
  assign new_new_n12455__ = new_new_n11059__ & ~new_new_n12454__;
  assign new_new_n12456__ = ~new_new_n11051__ & new_new_n11800__;
  assign new_new_n12457__ = new_new_n11050__ & new_new_n12451__;
  assign new_new_n12458__ = ~new_new_n12456__ & ~new_new_n12457__;
  assign new_new_n12459__ = ~new_new_n11059__ & ~new_new_n12458__;
  assign new_new_n12460__ = new_new_n11052__ & new_new_n11800__;
  assign new_new_n12461__ = ~new_new_n12449__ & ~new_new_n12460__;
  assign new_new_n12462__ = ~new_new_n12455__ & new_new_n12461__;
  assign new_new_n12463__ = ~new_new_n12459__ & new_new_n12462__;
  assign new_new_n12464__ = new_new_n11684__ & ~new_new_n12463__;
  assign new_new_n12465__ = ~new_new_n12448__ & ~new_new_n12464__;
  assign new_new_n12466__ = new_new_n11685__ & new_new_n12465__;
  assign new_new_n12467__ = ~new_new_n11685__ & ~new_new_n12465__;
  assign new_new_n12468__ = ~new_new_n12466__ & ~new_new_n12467__;
  assign new_new_n12469__ = ~new_new_n12439__ & ~new_new_n12468__;
  assign new_new_n12470__ = new_new_n12439__ & new_new_n12468__;
  assign new_new_n12471__ = ~new_new_n2636__ & new_new_n10702__;
  assign new_new_n12472__ = ~new_new_n2737__ & ~new_new_n11409__;
  assign new_new_n12473__ = ~new_new_n12471__ & ~new_new_n12472__;
  assign new_new_n12474__ = ~new_new_n9126__ & new_new_n10694__;
  assign new_new_n12475__ = pi08 & ~new_new_n12474__;
  assign new_new_n12476__ = ~pi07 & new_new_n2497__;
  assign new_new_n12477__ = pi07 & ~new_new_n2497__;
  assign new_new_n12478__ = new_new_n10694__ & ~new_new_n12476__;
  assign new_new_n12479__ = ~new_new_n12477__ & new_new_n12478__;
  assign new_new_n12480__ = ~new_new_n6797__ & new_new_n12479__;
  assign new_new_n12481__ = ~new_new_n12475__ & ~new_new_n12480__;
  assign new_new_n12482__ = new_new_n12473__ & ~new_new_n12481__;
  assign new_new_n12483__ = new_new_n7772__ & new_new_n10694__;
  assign new_new_n12484__ = new_new_n12473__ & ~new_new_n12483__;
  assign new_new_n12485__ = ~pi08 & ~new_new_n12484__;
  assign new_new_n12486__ = ~new_new_n12482__ & ~new_new_n12485__;
  assign new_new_n12487__ = ~new_new_n12470__ & ~new_new_n12486__;
  assign new_new_n12488__ = ~new_new_n12469__ & ~new_new_n12487__;
  assign new_new_n12489__ = ~pi11 & new_new_n11669__;
  assign new_new_n12490__ = ~new_new_n11671__ & ~new_new_n12489__;
  assign new_new_n12491__ = new_new_n12209__ & new_new_n12490__;
  assign new_new_n12492__ = ~new_new_n12209__ & ~new_new_n12490__;
  assign new_new_n12493__ = ~new_new_n12491__ & ~new_new_n12492__;
  assign new_new_n12494__ = ~new_new_n12488__ & new_new_n12493__;
  assign new_new_n12495__ = new_new_n12488__ & ~new_new_n12493__;
  assign new_new_n12496__ = ~new_new_n2572__ & new_new_n10698__;
  assign new_new_n12497__ = ~new_new_n2497__ & new_new_n10702__;
  assign new_new_n12498__ = new_new_n6804__ & new_new_n11378__;
  assign new_new_n12499__ = ~new_new_n12496__ & ~new_new_n12497__;
  assign new_new_n12500__ = ~new_new_n12498__ & new_new_n12499__;
  assign new_new_n12501__ = ~new_new_n2636__ & new_new_n10709__;
  assign new_new_n12502__ = pi08 & ~new_new_n12501__;
  assign new_new_n12503__ = ~new_new_n2636__ & new_new_n10712__;
  assign new_new_n12504__ = ~pi08 & ~new_new_n12503__;
  assign new_new_n12505__ = pi05 & ~new_new_n12504__;
  assign new_new_n12506__ = ~new_new_n12502__ & ~new_new_n12505__;
  assign new_new_n12507__ = new_new_n12500__ & ~new_new_n12506__;
  assign new_new_n12508__ = ~pi08 & ~new_new_n12500__;
  assign new_new_n12509__ = ~new_new_n12507__ & ~new_new_n12508__;
  assign new_new_n12510__ = ~new_new_n12495__ & ~new_new_n12509__;
  assign new_new_n12511__ = ~new_new_n12494__ & ~new_new_n12510__;
  assign new_new_n12512__ = ~new_new_n12240__ & new_new_n12511__;
  assign new_new_n12513__ = ~new_new_n12239__ & ~new_new_n12512__;
  assign new_new_n12514__ = ~new_new_n11832__ & ~new_new_n11833__;
  assign new_new_n12515__ = ~new_new_n11837__ & new_new_n12514__;
  assign new_new_n12516__ = new_new_n11837__ & ~new_new_n12514__;
  assign new_new_n12517__ = ~new_new_n12515__ & ~new_new_n12516__;
  assign new_new_n12518__ = ~new_new_n12513__ & ~new_new_n12517__;
  assign new_new_n12519__ = new_new_n12513__ & new_new_n12517__;
  assign new_new_n12520__ = ~new_new_n2313__ & new_new_n10702__;
  assign new_new_n12521__ = new_new_n2420__ & new_new_n10697__;
  assign new_new_n12522__ = new_new_n6751__ & ~new_new_n10697__;
  assign new_new_n12523__ = new_new_n10694__ & ~new_new_n12521__;
  assign new_new_n12524__ = ~new_new_n12522__ & new_new_n12523__;
  assign new_new_n12525__ = ~new_new_n12520__ & ~new_new_n12524__;
  assign new_new_n12526__ = ~new_new_n2572__ & new_new_n10709__;
  assign new_new_n12527__ = pi08 & ~new_new_n12526__;
  assign new_new_n12528__ = ~new_new_n2572__ & new_new_n10712__;
  assign new_new_n12529__ = ~pi08 & ~new_new_n12528__;
  assign new_new_n12530__ = pi05 & ~new_new_n12529__;
  assign new_new_n12531__ = ~new_new_n12527__ & ~new_new_n12530__;
  assign new_new_n12532__ = new_new_n12525__ & ~new_new_n12531__;
  assign new_new_n12533__ = ~pi08 & ~new_new_n12525__;
  assign new_new_n12534__ = ~new_new_n12532__ & ~new_new_n12533__;
  assign new_new_n12535__ = ~new_new_n12519__ & new_new_n12534__;
  assign new_new_n12536__ = ~new_new_n12518__ & ~new_new_n12535__;
  assign new_new_n12537__ = ~new_new_n12206__ & ~new_new_n12536__;
  assign new_new_n12538__ = new_new_n12206__ & new_new_n12536__;
  assign new_new_n12539__ = ~new_new_n2313__ & ~new_new_n11409__;
  assign new_new_n12540__ = ~new_new_n2224__ & new_new_n10698__;
  assign new_new_n12541__ = ~new_new_n2420__ & new_new_n10702__;
  assign new_new_n12542__ = new_new_n6521__ & new_new_n11378__;
  assign new_new_n12543__ = ~new_new_n12539__ & ~new_new_n12540__;
  assign new_new_n12544__ = ~new_new_n12541__ & new_new_n12543__;
  assign new_new_n12545__ = ~new_new_n12542__ & new_new_n12544__;
  assign new_new_n12546__ = ~pi08 & ~new_new_n12545__;
  assign new_new_n12547__ = pi08 & new_new_n12545__;
  assign new_new_n12548__ = ~new_new_n12546__ & ~new_new_n12547__;
  assign new_new_n12549__ = ~new_new_n12538__ & new_new_n12548__;
  assign new_new_n12550__ = ~new_new_n12537__ & ~new_new_n12549__;
  assign new_new_n12551__ = ~new_new_n12202__ & ~new_new_n12550__;
  assign new_new_n12552__ = new_new_n12202__ & new_new_n12550__;
  assign new_new_n12553__ = ~new_new_n2024__ & new_new_n10698__;
  assign new_new_n12554__ = ~new_new_n2224__ & new_new_n10702__;
  assign new_new_n12555__ = ~new_new_n2420__ & ~new_new_n11409__;
  assign new_new_n12556__ = new_new_n7313__ & new_new_n11378__;
  assign new_new_n12557__ = ~new_new_n12553__ & ~new_new_n12554__;
  assign new_new_n12558__ = ~new_new_n12555__ & new_new_n12557__;
  assign new_new_n12559__ = ~new_new_n12556__ & new_new_n12558__;
  assign new_new_n12560__ = pi08 & ~new_new_n12559__;
  assign new_new_n12561__ = ~pi08 & new_new_n12559__;
  assign new_new_n12562__ = ~new_new_n12560__ & ~new_new_n12561__;
  assign new_new_n12563__ = ~new_new_n12552__ & ~new_new_n12562__;
  assign new_new_n12564__ = ~new_new_n12551__ & ~new_new_n12563__;
  assign new_new_n12565__ = new_new_n12187__ & new_new_n12564__;
  assign new_new_n12566__ = ~new_new_n12187__ & ~new_new_n12564__;
  assign new_new_n12567__ = ~new_new_n2224__ & ~new_new_n11409__;
  assign new_new_n12568__ = ~new_new_n2024__ & new_new_n10702__;
  assign new_new_n12569__ = ~new_new_n2130__ & new_new_n10698__;
  assign new_new_n12570__ = ~new_new_n6036__ & new_new_n11378__;
  assign new_new_n12571__ = ~new_new_n12567__ & ~new_new_n12568__;
  assign new_new_n12572__ = ~new_new_n12569__ & new_new_n12571__;
  assign new_new_n12573__ = ~new_new_n12570__ & new_new_n12572__;
  assign new_new_n12574__ = ~pi08 & new_new_n12573__;
  assign new_new_n12575__ = pi08 & ~new_new_n12573__;
  assign new_new_n12576__ = ~new_new_n12574__ & ~new_new_n12575__;
  assign new_new_n12577__ = ~new_new_n12566__ & new_new_n12576__;
  assign new_new_n12578__ = ~new_new_n12565__ & ~new_new_n12577__;
  assign new_new_n12579__ = ~new_new_n12183__ & new_new_n12578__;
  assign new_new_n12580__ = new_new_n12183__ & ~new_new_n12578__;
  assign new_new_n12581__ = ~new_new_n2024__ & ~new_new_n11409__;
  assign new_new_n12582__ = ~new_new_n2130__ & new_new_n10702__;
  assign new_new_n12583__ = ~new_new_n3535__ & new_new_n10698__;
  assign new_new_n12584__ = new_new_n6854__ & new_new_n11378__;
  assign new_new_n12585__ = ~new_new_n12581__ & ~new_new_n12582__;
  assign new_new_n12586__ = ~new_new_n12583__ & new_new_n12585__;
  assign new_new_n12587__ = ~new_new_n12584__ & new_new_n12586__;
  assign new_new_n12588__ = pi08 & ~new_new_n12587__;
  assign new_new_n12589__ = ~pi08 & new_new_n12587__;
  assign new_new_n12590__ = ~new_new_n12588__ & ~new_new_n12589__;
  assign new_new_n12591__ = ~new_new_n12580__ & ~new_new_n12590__;
  assign new_new_n12592__ = ~new_new_n12579__ & ~new_new_n12591__;
  assign new_new_n12593__ = ~new_new_n12179__ & new_new_n12592__;
  assign new_new_n12594__ = new_new_n12179__ & ~new_new_n12592__;
  assign new_new_n12595__ = ~new_new_n1823__ & new_new_n10698__;
  assign new_new_n12596__ = ~new_new_n3535__ & new_new_n10702__;
  assign new_new_n12597__ = ~new_new_n2130__ & ~new_new_n11409__;
  assign new_new_n12598__ = new_new_n7274__ & new_new_n11378__;
  assign new_new_n12599__ = ~new_new_n12595__ & ~new_new_n12596__;
  assign new_new_n12600__ = ~new_new_n12597__ & new_new_n12599__;
  assign new_new_n12601__ = ~new_new_n12598__ & new_new_n12600__;
  assign new_new_n12602__ = pi08 & new_new_n12601__;
  assign new_new_n12603__ = ~pi08 & ~new_new_n12601__;
  assign new_new_n12604__ = ~new_new_n12602__ & ~new_new_n12603__;
  assign new_new_n12605__ = ~new_new_n12594__ & ~new_new_n12604__;
  assign new_new_n12606__ = ~new_new_n12593__ & ~new_new_n12605__;
  assign new_new_n12607__ = ~new_new_n12158__ & new_new_n12606__;
  assign new_new_n12608__ = new_new_n12158__ & ~new_new_n12606__;
  assign new_new_n12609__ = ~new_new_n11160__ & ~new_new_n11908__;
  assign new_new_n12610__ = new_new_n11160__ & new_new_n11908__;
  assign new_new_n12611__ = ~new_new_n12609__ & ~new_new_n12610__;
  assign new_new_n12612__ = new_new_n11162__ & ~new_new_n11586__;
  assign new_new_n12613__ = ~new_new_n11162__ & new_new_n11586__;
  assign new_new_n12614__ = ~new_new_n12612__ & ~new_new_n12613__;
  assign new_new_n12615__ = new_new_n12611__ & new_new_n12614__;
  assign new_new_n12616__ = ~new_new_n12611__ & ~new_new_n12614__;
  assign new_new_n12617__ = ~new_new_n12615__ & ~new_new_n12616__;
  assign new_new_n12618__ = ~new_new_n12608__ & ~new_new_n12617__;
  assign new_new_n12619__ = ~new_new_n12607__ & ~new_new_n12618__;
  assign new_new_n12620__ = new_new_n12140__ & ~new_new_n12619__;
  assign new_new_n12621__ = ~new_new_n12140__ & new_new_n12619__;
  assign new_new_n12622__ = ~new_new_n1823__ & ~new_new_n11409__;
  assign new_new_n12623__ = ~new_new_n1902__ & new_new_n10702__;
  assign new_new_n12624__ = ~new_new_n1660__ & new_new_n10698__;
  assign new_new_n12625__ = ~new_new_n5274__ & new_new_n11378__;
  assign new_new_n12626__ = ~new_new_n12622__ & ~new_new_n12623__;
  assign new_new_n12627__ = ~new_new_n12624__ & new_new_n12626__;
  assign new_new_n12628__ = ~new_new_n12625__ & new_new_n12627__;
  assign new_new_n12629__ = pi08 & ~new_new_n12628__;
  assign new_new_n12630__ = ~pi08 & new_new_n12628__;
  assign new_new_n12631__ = ~new_new_n12629__ & ~new_new_n12630__;
  assign new_new_n12632__ = ~new_new_n12621__ & ~new_new_n12631__;
  assign new_new_n12633__ = ~new_new_n12620__ & ~new_new_n12632__;
  assign new_new_n12634__ = new_new_n12146__ & ~new_new_n12633__;
  assign new_new_n12635__ = ~new_new_n1737__ & new_new_n10698__;
  assign new_new_n12636__ = ~new_new_n1902__ & ~new_new_n11409__;
  assign new_new_n12637__ = ~new_new_n1660__ & new_new_n10702__;
  assign new_new_n12638__ = ~new_new_n12635__ & ~new_new_n12636__;
  assign new_new_n12639__ = ~new_new_n12637__ & new_new_n12638__;
  assign new_new_n12640__ = new_new_n5688__ & new_new_n10694__;
  assign new_new_n12641__ = pi08 & ~new_new_n12640__;
  assign new_new_n12642__ = new_new_n5688__ & new_new_n11498__;
  assign new_new_n12643__ = ~new_new_n12641__ & ~new_new_n12642__;
  assign new_new_n12644__ = new_new_n12639__ & ~new_new_n12643__;
  assign new_new_n12645__ = ~pi08 & ~new_new_n12639__;
  assign new_new_n12646__ = ~new_new_n12644__ & ~new_new_n12645__;
  assign new_new_n12647__ = ~new_new_n12634__ & ~new_new_n12646__;
  assign new_new_n12648__ = new_new_n12126__ & new_new_n12130__;
  assign new_new_n12649__ = ~new_new_n12146__ & new_new_n12633__;
  assign new_new_n12650__ = ~new_new_n12648__ & ~new_new_n12649__;
  assign new_new_n12651__ = ~new_new_n12647__ & new_new_n12650__;
  assign new_new_n12652__ = ~new_new_n12131__ & ~new_new_n12651__;
  assign new_new_n12653__ = ~new_new_n5671__ & new_new_n11378__;
  assign new_new_n12654__ = ~new_new_n1737__ & ~new_new_n11409__;
  assign new_new_n12655__ = ~new_new_n1466__ & new_new_n10702__;
  assign new_new_n12656__ = ~new_new_n12654__ & ~new_new_n12655__;
  assign new_new_n12657__ = ~new_new_n12653__ & new_new_n12656__;
  assign new_new_n12658__ = ~new_new_n1556__ & new_new_n10694__;
  assign new_new_n12659__ = ~pi08 & ~new_new_n12658__;
  assign new_new_n12660__ = ~new_new_n1556__ & new_new_n11498__;
  assign new_new_n12661__ = ~new_new_n12659__ & ~new_new_n12660__;
  assign new_new_n12662__ = new_new_n12657__ & ~new_new_n12661__;
  assign new_new_n12663__ = pi08 & ~new_new_n12657__;
  assign new_new_n12664__ = ~new_new_n12662__ & ~new_new_n12663__;
  assign new_new_n12665__ = ~new_new_n12652__ & ~new_new_n12664__;
  assign new_new_n12666__ = new_new_n12652__ & new_new_n12664__;
  assign new_new_n12667__ = ~new_new_n11954__ & ~new_new_n11955__;
  assign new_new_n12668__ = new_new_n11967__ & ~new_new_n12667__;
  assign new_new_n12669__ = ~new_new_n11967__ & new_new_n12667__;
  assign new_new_n12670__ = ~new_new_n12668__ & ~new_new_n12669__;
  assign new_new_n12671__ = ~new_new_n12666__ & ~new_new_n12670__;
  assign new_new_n12672__ = ~new_new_n12665__ & ~new_new_n12671__;
  assign new_new_n12673__ = ~new_new_n11982__ & ~new_new_n11983__;
  assign new_new_n12674__ = ~new_new_n11987__ & new_new_n12673__;
  assign new_new_n12675__ = new_new_n11987__ & ~new_new_n12673__;
  assign new_new_n12676__ = ~new_new_n12674__ & ~new_new_n12675__;
  assign new_new_n12677__ = new_new_n12672__ & ~new_new_n12676__;
  assign new_new_n12678__ = ~new_new_n12672__ & new_new_n12676__;
  assign new_new_n12679__ = ~new_new_n1466__ & ~new_new_n11409__;
  assign new_new_n12680__ = ~new_new_n1556__ & new_new_n10702__;
  assign new_new_n12681__ = ~new_new_n1325__ & new_new_n10698__;
  assign new_new_n12682__ = new_new_n5048__ & new_new_n11378__;
  assign new_new_n12683__ = ~new_new_n12679__ & ~new_new_n12680__;
  assign new_new_n12684__ = ~new_new_n12681__ & new_new_n12683__;
  assign new_new_n12685__ = ~new_new_n12682__ & new_new_n12684__;
  assign new_new_n12686__ = ~pi08 & ~new_new_n12685__;
  assign new_new_n12687__ = pi08 & new_new_n12685__;
  assign new_new_n12688__ = ~new_new_n12686__ & ~new_new_n12687__;
  assign new_new_n12689__ = ~new_new_n12678__ & ~new_new_n12688__;
  assign new_new_n12690__ = ~new_new_n12677__ & ~new_new_n12689__;
  assign new_new_n12691__ = ~new_new_n12113__ & ~new_new_n12690__;
  assign new_new_n12692__ = ~new_new_n12112__ & ~new_new_n12691__;
  assign new_new_n12693__ = ~new_new_n12010__ & ~new_new_n12011__;
  assign new_new_n12694__ = ~new_new_n12023__ & new_new_n12693__;
  assign new_new_n12695__ = new_new_n12023__ & ~new_new_n12693__;
  assign new_new_n12696__ = ~new_new_n12694__ & ~new_new_n12695__;
  assign new_new_n12697__ = new_new_n12692__ & ~new_new_n12696__;
  assign new_new_n12698__ = ~new_new_n12692__ & new_new_n12696__;
  assign new_new_n12699__ = ~new_new_n1061__ & new_new_n10698__;
  assign new_new_n12700__ = ~new_new_n1325__ & ~new_new_n11409__;
  assign new_new_n12701__ = ~new_new_n3618__ & new_new_n10702__;
  assign new_new_n12702__ = ~new_new_n12699__ & ~new_new_n12700__;
  assign new_new_n12703__ = ~new_new_n12701__ & new_new_n12702__;
  assign new_new_n12704__ = new_new_n4926__ & new_new_n11378__;
  assign new_new_n12705__ = new_new_n12703__ & ~new_new_n12704__;
  assign new_new_n12706__ = pi08 & ~new_new_n12705__;
  assign new_new_n12707__ = ~pi08 & new_new_n12705__;
  assign new_new_n12708__ = ~new_new_n12706__ & ~new_new_n12707__;
  assign new_new_n12709__ = ~new_new_n12698__ & ~new_new_n12708__;
  assign new_new_n12710__ = ~new_new_n12697__ & ~new_new_n12709__;
  assign new_new_n12711__ = ~new_new_n12091__ & new_new_n12710__;
  assign new_new_n12712__ = new_new_n12091__ & ~new_new_n12710__;
  assign new_new_n12713__ = ~new_new_n1207__ & new_new_n10698__;
  assign new_new_n12714__ = ~new_new_n3618__ & ~new_new_n11409__;
  assign new_new_n12715__ = ~new_new_n1061__ & new_new_n10702__;
  assign new_new_n12716__ = ~new_new_n12713__ & ~new_new_n12714__;
  assign new_new_n12717__ = ~new_new_n12715__ & new_new_n12716__;
  assign new_new_n12718__ = ~new_new_n5235__ & new_new_n10694__;
  assign new_new_n12719__ = pi08 & ~new_new_n12718__;
  assign new_new_n12720__ = ~new_new_n5235__ & new_new_n11498__;
  assign new_new_n12721__ = ~new_new_n12719__ & ~new_new_n12720__;
  assign new_new_n12722__ = new_new_n12717__ & ~new_new_n12721__;
  assign new_new_n12723__ = ~pi08 & ~new_new_n12717__;
  assign new_new_n12724__ = ~new_new_n12722__ & ~new_new_n12723__;
  assign new_new_n12725__ = ~new_new_n12712__ & ~new_new_n12724__;
  assign new_new_n12726__ = ~new_new_n12711__ & ~new_new_n12725__;
  assign new_new_n12727__ = ~new_new_n12087__ & new_new_n12726__;
  assign new_new_n12728__ = new_new_n12087__ & ~new_new_n12726__;
  assign new_new_n12729__ = ~new_new_n12727__ & ~new_new_n12728__;
  assign new_new_n12730__ = ~new_new_n1061__ & ~new_new_n11409__;
  assign new_new_n12731__ = ~new_new_n868__ & new_new_n10698__;
  assign new_new_n12732__ = ~new_new_n1207__ & new_new_n10702__;
  assign new_new_n12733__ = ~new_new_n12730__ & ~new_new_n12731__;
  assign new_new_n12734__ = ~new_new_n12732__ & new_new_n12733__;
  assign new_new_n12735__ = ~new_new_n4550__ & new_new_n10694__;
  assign new_new_n12736__ = pi08 & ~new_new_n12735__;
  assign new_new_n12737__ = ~new_new_n4550__ & new_new_n11498__;
  assign new_new_n12738__ = ~new_new_n12736__ & ~new_new_n12737__;
  assign new_new_n12739__ = new_new_n12734__ & ~new_new_n12738__;
  assign new_new_n12740__ = ~pi08 & ~new_new_n12734__;
  assign new_new_n12741__ = ~new_new_n12739__ & ~new_new_n12740__;
  assign new_new_n12742__ = new_new_n12729__ & new_new_n12741__;
  assign new_new_n12743__ = ~new_new_n12727__ & ~new_new_n12742__;
  assign new_new_n12744__ = ~new_new_n12044__ & ~new_new_n12045__;
  assign new_new_n12745__ = ~new_new_n12055__ & new_new_n12744__;
  assign new_new_n12746__ = new_new_n12055__ & ~new_new_n12744__;
  assign new_new_n12747__ = ~new_new_n12745__ & ~new_new_n12746__;
  assign new_new_n12748__ = ~new_new_n12743__ & new_new_n12747__;
  assign new_new_n12749__ = new_new_n12743__ & ~new_new_n12747__;
  assign new_new_n12750__ = ~new_new_n868__ & new_new_n10702__;
  assign new_new_n12751__ = ~new_new_n1207__ & ~new_new_n11409__;
  assign new_new_n12752__ = ~new_new_n4032__ & ~new_new_n10697__;
  assign new_new_n12753__ = new_new_n3720__ & ~new_new_n12752__;
  assign new_new_n12754__ = ~new_new_n3720__ & new_new_n12752__;
  assign new_new_n12755__ = new_new_n10694__ & ~new_new_n12753__;
  assign new_new_n12756__ = ~new_new_n12754__ & new_new_n12755__;
  assign new_new_n12757__ = ~new_new_n12750__ & ~new_new_n12751__;
  assign new_new_n12758__ = ~new_new_n12756__ & new_new_n12757__;
  assign new_new_n12759__ = pi08 & ~new_new_n12758__;
  assign new_new_n12760__ = ~pi08 & new_new_n12758__;
  assign new_new_n12761__ = ~new_new_n12759__ & ~new_new_n12760__;
  assign new_new_n12762__ = ~new_new_n12749__ & ~new_new_n12761__;
  assign new_new_n12763__ = ~new_new_n12748__ & ~new_new_n12762__;
  assign new_new_n12764__ = ~new_new_n12058__ & ~new_new_n12059__;
  assign new_new_n12765__ = new_new_n12069__ & new_new_n12764__;
  assign new_new_n12766__ = ~new_new_n12069__ & ~new_new_n12764__;
  assign new_new_n12767__ = ~new_new_n12765__ & ~new_new_n12766__;
  assign new_new_n12768__ = ~new_new_n12763__ & ~new_new_n12767__;
  assign new_new_n12769__ = new_new_n12763__ & new_new_n12767__;
  assign new_new_n12770__ = ~new_new_n3720__ & new_new_n10702__;
  assign new_new_n12771__ = new_new_n4036__ & ~new_new_n10697__;
  assign new_new_n12772__ = new_new_n910__ & ~new_new_n12771__;
  assign new_new_n12773__ = ~new_new_n910__ & new_new_n12771__;
  assign new_new_n12774__ = new_new_n10694__ & ~new_new_n12772__;
  assign new_new_n12775__ = ~new_new_n12773__ & new_new_n12774__;
  assign new_new_n12776__ = ~new_new_n12770__ & ~new_new_n12775__;
  assign new_new_n12777__ = ~new_new_n868__ & new_new_n10709__;
  assign new_new_n12778__ = pi08 & ~new_new_n12777__;
  assign new_new_n12779__ = ~new_new_n868__ & new_new_n10712__;
  assign new_new_n12780__ = ~pi08 & ~new_new_n12779__;
  assign new_new_n12781__ = pi05 & ~new_new_n12780__;
  assign new_new_n12782__ = ~new_new_n12778__ & ~new_new_n12781__;
  assign new_new_n12783__ = new_new_n12776__ & ~new_new_n12782__;
  assign new_new_n12784__ = ~pi08 & ~new_new_n12776__;
  assign new_new_n12785__ = ~new_new_n12783__ & ~new_new_n12784__;
  assign new_new_n12786__ = ~new_new_n12769__ & new_new_n12785__;
  assign new_new_n12787__ = ~new_new_n12768__ & ~new_new_n12786__;
  assign new_new_n12788__ = ~new_new_n12083__ & ~new_new_n12787__;
  assign new_new_n12789__ = ~new_new_n12082__ & ~new_new_n12788__;
  assign new_new_n12790__ = ~new_new_n12082__ & ~new_new_n12083__;
  assign new_new_n12791__ = new_new_n12787__ & ~new_new_n12790__;
  assign new_new_n12792__ = ~new_new_n12787__ & new_new_n12790__;
  assign new_new_n12793__ = ~new_new_n12791__ & ~new_new_n12792__;
  assign new_new_n12794__ = pi02 & new_new_n3768__;
  assign new_new_n12795__ = ~pi02 & ~new_new_n3768__;
  assign new_new_n12796__ = ~new_new_n12794__ & ~new_new_n12795__;
  assign new_new_n12797__ = pi01 & ~new_new_n12796__;
  assign new_new_n12798__ = ~pi01 & pi02;
  assign new_new_n12799__ = new_new_n583__ & new_new_n12798__;
  assign new_new_n12800__ = ~new_new_n12797__ & ~new_new_n12799__;
  assign new_new_n12801__ = ~pi00 & ~new_new_n12800__;
  assign new_new_n12802__ = pi01 & new_new_n466__;
  assign new_new_n12803__ = ~pi01 & ~new_new_n466__;
  assign new_new_n12804__ = ~new_new_n12802__ & ~new_new_n12803__;
  assign new_new_n12805__ = new_new_n4169__ & new_new_n12804__;
  assign new_new_n12806__ = pi02 & ~new_new_n466__;
  assign new_new_n12807__ = ~pi02 & new_new_n466__;
  assign new_new_n12808__ = ~new_new_n12806__ & ~new_new_n12807__;
  assign new_new_n12809__ = ~new_new_n4169__ & ~new_new_n12808__;
  assign new_new_n12810__ = pi00 & ~new_new_n12805__;
  assign new_new_n12811__ = ~new_new_n12809__ & new_new_n12810__;
  assign new_new_n12812__ = ~new_new_n12801__ & ~new_new_n12811__;
  assign new_new_n12813__ = pi01 & ~new_new_n583__;
  assign new_new_n12814__ = ~pi01 & ~new_new_n691__;
  assign new_new_n12815__ = pi02 & ~new_new_n12814__;
  assign new_new_n12816__ = ~new_new_n12813__ & ~new_new_n12815__;
  assign new_new_n12817__ = pi02 & new_new_n12813__;
  assign new_new_n12818__ = ~pi00 & ~new_new_n12817__;
  assign new_new_n12819__ = ~new_new_n12816__ & new_new_n12818__;
  assign new_new_n12820__ = pi01 & new_new_n3768__;
  assign new_new_n12821__ = ~pi01 & ~new_new_n3768__;
  assign new_new_n12822__ = ~new_new_n12820__ & ~new_new_n12821__;
  assign new_new_n12823__ = new_new_n4141__ & new_new_n12822__;
  assign new_new_n12824__ = ~new_new_n4141__ & new_new_n12796__;
  assign new_new_n12825__ = pi00 & ~new_new_n12823__;
  assign new_new_n12826__ = ~new_new_n12824__ & new_new_n12825__;
  assign new_new_n12827__ = ~new_new_n12819__ & ~new_new_n12826__;
  assign new_new_n12828__ = pi02 & new_new_n11467__;
  assign new_new_n12829__ = ~pi05 & ~new_new_n12828__;
  assign new_new_n12830__ = ~pi02 & new_new_n11466__;
  assign new_new_n12831__ = pi05 & ~new_new_n12830__;
  assign new_new_n12832__ = ~new_new_n12829__ & ~new_new_n12831__;
  assign new_new_n12833__ = ~new_new_n868__ & new_new_n12832__;
  assign new_new_n12834__ = ~new_new_n3720__ & new_new_n11475__;
  assign new_new_n12835__ = ~new_new_n12833__ & ~new_new_n12834__;
  assign new_new_n12836__ = ~new_new_n5129__ & new_new_n11469__;
  assign new_new_n12837__ = pi05 & ~new_new_n12836__;
  assign new_new_n12838__ = ~pi04 & new_new_n910__;
  assign new_new_n12839__ = pi04 & ~new_new_n910__;
  assign new_new_n12840__ = ~new_new_n11482__ & ~new_new_n12838__;
  assign new_new_n12841__ = ~new_new_n12839__ & new_new_n12840__;
  assign new_new_n12842__ = new_new_n4036__ & new_new_n12841__;
  assign new_new_n12843__ = ~new_new_n12837__ & ~new_new_n12842__;
  assign new_new_n12844__ = new_new_n12835__ & ~new_new_n12843__;
  assign new_new_n12845__ = new_new_n5116__ & new_new_n11469__;
  assign new_new_n12846__ = new_new_n12835__ & ~new_new_n12845__;
  assign new_new_n12847__ = ~pi05 & ~new_new_n12846__;
  assign new_new_n12848__ = ~new_new_n12844__ & ~new_new_n12847__;
  assign new_new_n12849__ = ~new_new_n1207__ & new_new_n11471__;
  assign new_new_n12850__ = ~new_new_n11478__ & ~new_new_n11482__;
  assign new_new_n12851__ = ~new_new_n3720__ & new_new_n12850__;
  assign new_new_n12852__ = ~new_new_n868__ & new_new_n11475__;
  assign new_new_n12853__ = ~new_new_n12849__ & ~new_new_n12851__;
  assign new_new_n12854__ = ~new_new_n12852__ & new_new_n12853__;
  assign new_new_n12855__ = pi05 & ~new_new_n12854__;
  assign new_new_n12856__ = ~pi04 & ~new_new_n11482__;
  assign new_new_n12857__ = ~new_new_n5927__ & new_new_n12856__;
  assign new_new_n12858__ = ~new_new_n5927__ & new_new_n11469__;
  assign new_new_n12859__ = ~pi05 & ~new_new_n12858__;
  assign new_new_n12860__ = ~new_new_n12857__ & ~new_new_n12859__;
  assign new_new_n12861__ = new_new_n12854__ & ~new_new_n12860__;
  assign new_new_n12862__ = ~new_new_n12855__ & ~new_new_n12861__;
  assign new_new_n12863__ = ~new_new_n12112__ & ~new_new_n12113__;
  assign new_new_n12864__ = ~new_new_n12690__ & new_new_n12863__;
  assign new_new_n12865__ = new_new_n12690__ & ~new_new_n12863__;
  assign new_new_n12866__ = ~new_new_n12864__ & ~new_new_n12865__;
  assign new_new_n12867__ = ~new_new_n1207__ & new_new_n12850__;
  assign new_new_n12868__ = ~new_new_n3618__ & new_new_n11471__;
  assign new_new_n12869__ = ~new_new_n1061__ & new_new_n11475__;
  assign new_new_n12870__ = ~new_new_n12867__ & ~new_new_n12868__;
  assign new_new_n12871__ = ~new_new_n12869__ & new_new_n12870__;
  assign new_new_n12872__ = ~pi05 & ~new_new_n12871__;
  assign new_new_n12873__ = pi04 & ~new_new_n11482__;
  assign new_new_n12874__ = ~new_new_n5235__ & new_new_n12873__;
  assign new_new_n12875__ = ~new_new_n5235__ & new_new_n11469__;
  assign new_new_n12876__ = pi05 & ~new_new_n12875__;
  assign new_new_n12877__ = ~new_new_n12874__ & ~new_new_n12876__;
  assign new_new_n12878__ = new_new_n12871__ & ~new_new_n12877__;
  assign new_new_n12879__ = ~new_new_n12872__ & ~new_new_n12878__;
  assign new_new_n12880__ = ~new_new_n12665__ & ~new_new_n12666__;
  assign new_new_n12881__ = ~new_new_n12670__ & new_new_n12880__;
  assign new_new_n12882__ = new_new_n12670__ & ~new_new_n12880__;
  assign new_new_n12883__ = ~new_new_n12881__ & ~new_new_n12882__;
  assign new_new_n12884__ = ~new_new_n1325__ & new_new_n11475__;
  assign new_new_n12885__ = new_new_n8344__ & new_new_n11478__;
  assign new_new_n12886__ = ~new_new_n3618__ & ~new_new_n11478__;
  assign new_new_n12887__ = ~new_new_n5981__ & ~new_new_n12886__;
  assign new_new_n12888__ = ~new_new_n12885__ & new_new_n12887__;
  assign new_new_n12889__ = new_new_n11469__ & ~new_new_n12888__;
  assign new_new_n12890__ = ~new_new_n12884__ & ~new_new_n12889__;
  assign new_new_n12891__ = ~pi05 & ~new_new_n12890__;
  assign new_new_n12892__ = ~new_new_n1556__ & new_new_n12828__;
  assign new_new_n12893__ = ~new_new_n1556__ & new_new_n12830__;
  assign new_new_n12894__ = pi05 & ~new_new_n12893__;
  assign new_new_n12895__ = ~new_new_n12892__ & ~new_new_n12894__;
  assign new_new_n12896__ = new_new_n12890__ & ~new_new_n12895__;
  assign new_new_n12897__ = ~new_new_n12891__ & ~new_new_n12896__;
  assign new_new_n12898__ = ~new_new_n12131__ & new_new_n12651__;
  assign new_new_n12899__ = new_new_n12131__ & ~new_new_n12146__;
  assign new_new_n12900__ = ~new_new_n12634__ & ~new_new_n12649__;
  assign new_new_n12901__ = new_new_n12648__ & new_new_n12900__;
  assign new_new_n12902__ = ~new_new_n12899__ & ~new_new_n12901__;
  assign new_new_n12903__ = new_new_n12646__ & ~new_new_n12900__;
  assign new_new_n12904__ = ~new_new_n12646__ & new_new_n12900__;
  assign new_new_n12905__ = ~new_new_n12903__ & ~new_new_n12904__;
  assign new_new_n12906__ = ~new_new_n12902__ & ~new_new_n12905__;
  assign new_new_n12907__ = new_new_n12131__ & ~new_new_n12646__;
  assign new_new_n12908__ = ~new_new_n12146__ & new_new_n12648__;
  assign new_new_n12909__ = ~new_new_n12907__ & ~new_new_n12908__;
  assign new_new_n12910__ = new_new_n12633__ & ~new_new_n12909__;
  assign new_new_n12911__ = ~new_new_n12898__ & ~new_new_n12910__;
  assign new_new_n12912__ = ~new_new_n12906__ & new_new_n12911__;
  assign new_new_n12913__ = new_new_n12897__ & new_new_n12912__;
  assign new_new_n12914__ = ~new_new_n12897__ & ~new_new_n12912__;
  assign new_new_n12915__ = ~new_new_n12620__ & ~new_new_n12621__;
  assign new_new_n12916__ = new_new_n12631__ & new_new_n12915__;
  assign new_new_n12917__ = ~new_new_n12631__ & ~new_new_n12915__;
  assign new_new_n12918__ = ~new_new_n12916__ & ~new_new_n12917__;
  assign new_new_n12919__ = ~new_new_n12607__ & ~new_new_n12608__;
  assign new_new_n12920__ = ~new_new_n11587__ & ~new_new_n11588__;
  assign new_new_n12921__ = new_new_n11908__ & ~new_new_n12920__;
  assign new_new_n12922__ = ~new_new_n11908__ & new_new_n12920__;
  assign new_new_n12923__ = ~new_new_n12921__ & ~new_new_n12922__;
  assign new_new_n12924__ = new_new_n12919__ & new_new_n12923__;
  assign new_new_n12925__ = ~new_new_n12919__ & ~new_new_n12923__;
  assign new_new_n12926__ = ~new_new_n12924__ & ~new_new_n12925__;
  assign new_new_n12927__ = ~new_new_n1660__ & new_new_n11475__;
  assign new_new_n12928__ = ~new_new_n1902__ & new_new_n11471__;
  assign new_new_n12929__ = ~new_new_n1737__ & new_new_n12850__;
  assign new_new_n12930__ = ~new_new_n12927__ & ~new_new_n12928__;
  assign new_new_n12931__ = ~new_new_n12929__ & new_new_n12930__;
  assign new_new_n12932__ = pi05 & ~new_new_n12931__;
  assign new_new_n12933__ = new_new_n5688__ & new_new_n12856__;
  assign new_new_n12934__ = new_new_n5688__ & new_new_n11469__;
  assign new_new_n12935__ = ~pi05 & ~new_new_n12934__;
  assign new_new_n12936__ = ~new_new_n12933__ & ~new_new_n12935__;
  assign new_new_n12937__ = new_new_n12931__ & ~new_new_n12936__;
  assign new_new_n12938__ = ~new_new_n12932__ & ~new_new_n12937__;
  assign new_new_n12939__ = ~new_new_n12579__ & ~new_new_n12580__;
  assign new_new_n12940__ = new_new_n12590__ & new_new_n12939__;
  assign new_new_n12941__ = ~new_new_n12590__ & ~new_new_n12939__;
  assign new_new_n12942__ = ~new_new_n12940__ & ~new_new_n12941__;
  assign new_new_n12943__ = ~new_new_n1823__ & new_new_n11475__;
  assign new_new_n12944__ = new_new_n6487__ & new_new_n11478__;
  assign new_new_n12945__ = new_new_n1902__ & ~new_new_n11478__;
  assign new_new_n12946__ = ~new_new_n11482__ & ~new_new_n12945__;
  assign new_new_n12947__ = ~new_new_n12944__ & new_new_n12946__;
  assign new_new_n12948__ = ~new_new_n12943__ & ~new_new_n12947__;
  assign new_new_n12949__ = ~pi05 & ~new_new_n12948__;
  assign new_new_n12950__ = ~new_new_n3535__ & new_new_n12830__;
  assign new_new_n12951__ = pi05 & ~new_new_n12950__;
  assign new_new_n12952__ = ~new_new_n3535__ & new_new_n12828__;
  assign new_new_n12953__ = ~new_new_n12951__ & ~new_new_n12952__;
  assign new_new_n12954__ = new_new_n12948__ & ~new_new_n12953__;
  assign new_new_n12955__ = ~new_new_n12949__ & ~new_new_n12954__;
  assign new_new_n12956__ = ~new_new_n12551__ & ~new_new_n12552__;
  assign new_new_n12957__ = new_new_n12562__ & ~new_new_n12956__;
  assign new_new_n12958__ = ~new_new_n12562__ & new_new_n12956__;
  assign new_new_n12959__ = ~new_new_n12957__ & ~new_new_n12958__;
  assign new_new_n12960__ = ~new_new_n2130__ & new_new_n12850__;
  assign new_new_n12961__ = ~new_new_n2224__ & new_new_n11471__;
  assign new_new_n12962__ = ~new_new_n2024__ & new_new_n11475__;
  assign new_new_n12963__ = ~new_new_n12960__ & ~new_new_n12961__;
  assign new_new_n12964__ = ~new_new_n12962__ & new_new_n12963__;
  assign new_new_n12965__ = ~pi05 & ~new_new_n12964__;
  assign new_new_n12966__ = ~new_new_n6036__ & new_new_n12873__;
  assign new_new_n12967__ = ~new_new_n6036__ & new_new_n11469__;
  assign new_new_n12968__ = pi05 & ~new_new_n12967__;
  assign new_new_n12969__ = ~new_new_n12966__ & ~new_new_n12968__;
  assign new_new_n12970__ = new_new_n12964__ & ~new_new_n12969__;
  assign new_new_n12971__ = ~new_new_n12965__ & ~new_new_n12970__;
  assign new_new_n12972__ = ~new_new_n12239__ & ~new_new_n12240__;
  assign new_new_n12973__ = new_new_n12511__ & new_new_n12972__;
  assign new_new_n12974__ = ~new_new_n12511__ & ~new_new_n12972__;
  assign new_new_n12975__ = ~new_new_n12973__ & ~new_new_n12974__;
  assign new_new_n12976__ = ~new_new_n2313__ & new_new_n11471__;
  assign new_new_n12977__ = ~new_new_n2420__ & new_new_n11475__;
  assign new_new_n12978__ = new_new_n2224__ & ~new_new_n11478__;
  assign new_new_n12979__ = ~new_new_n6521__ & new_new_n11478__;
  assign new_new_n12980__ = ~new_new_n11482__ & ~new_new_n12978__;
  assign new_new_n12981__ = ~new_new_n12979__ & new_new_n12980__;
  assign new_new_n12982__ = ~new_new_n12976__ & ~new_new_n12977__;
  assign new_new_n12983__ = ~new_new_n12981__ & new_new_n12982__;
  assign new_new_n12984__ = ~pi05 & ~new_new_n12983__;
  assign new_new_n12985__ = pi05 & new_new_n12983__;
  assign new_new_n12986__ = ~new_new_n12984__ & ~new_new_n12985__;
  assign new_new_n12987__ = ~new_new_n2313__ & new_new_n11475__;
  assign new_new_n12988__ = new_new_n6751__ & new_new_n11478__;
  assign new_new_n12989__ = new_new_n2420__ & ~new_new_n11478__;
  assign new_new_n12990__ = ~new_new_n11482__ & ~new_new_n12989__;
  assign new_new_n12991__ = ~new_new_n12988__ & new_new_n12990__;
  assign new_new_n12992__ = ~new_new_n12987__ & ~new_new_n12991__;
  assign new_new_n12993__ = ~pi05 & ~new_new_n12992__;
  assign new_new_n12994__ = ~new_new_n2572__ & new_new_n12830__;
  assign new_new_n12995__ = pi05 & ~new_new_n12994__;
  assign new_new_n12996__ = ~new_new_n2572__ & new_new_n12828__;
  assign new_new_n12997__ = ~new_new_n12995__ & ~new_new_n12996__;
  assign new_new_n12998__ = new_new_n12992__ & ~new_new_n12997__;
  assign new_new_n12999__ = ~new_new_n12993__ & ~new_new_n12998__;
  assign new_new_n13000__ = ~new_new_n2572__ & new_new_n12850__;
  assign new_new_n13001__ = ~new_new_n2636__ & new_new_n11471__;
  assign new_new_n13002__ = ~new_new_n2497__ & new_new_n11475__;
  assign new_new_n13003__ = ~new_new_n13000__ & ~new_new_n13001__;
  assign new_new_n13004__ = ~new_new_n13002__ & new_new_n13003__;
  assign new_new_n13005__ = pi05 & ~new_new_n13004__;
  assign new_new_n13006__ = new_new_n6804__ & new_new_n12856__;
  assign new_new_n13007__ = new_new_n6804__ & new_new_n11469__;
  assign new_new_n13008__ = ~pi05 & ~new_new_n13007__;
  assign new_new_n13009__ = ~new_new_n13006__ & ~new_new_n13008__;
  assign new_new_n13010__ = new_new_n13004__ & ~new_new_n13009__;
  assign new_new_n13011__ = ~new_new_n13005__ & ~new_new_n13010__;
  assign new_new_n13012__ = ~new_new_n2737__ & new_new_n12832__;
  assign new_new_n13013__ = ~new_new_n2636__ & new_new_n11475__;
  assign new_new_n13014__ = ~new_new_n13012__ & ~new_new_n13013__;
  assign new_new_n13015__ = new_new_n7772__ & new_new_n11469__;
  assign new_new_n13016__ = new_new_n13014__ & ~new_new_n13015__;
  assign new_new_n13017__ = pi05 & ~new_new_n13016__;
  assign new_new_n13018__ = ~new_new_n9126__ & new_new_n11469__;
  assign new_new_n13019__ = ~pi05 & ~new_new_n13018__;
  assign new_new_n13020__ = pi04 & new_new_n2497__;
  assign new_new_n13021__ = ~pi04 & ~new_new_n2497__;
  assign new_new_n13022__ = ~new_new_n11482__ & ~new_new_n13020__;
  assign new_new_n13023__ = ~new_new_n13021__ & new_new_n13022__;
  assign new_new_n13024__ = ~new_new_n6797__ & new_new_n13023__;
  assign new_new_n13025__ = ~new_new_n13019__ & ~new_new_n13024__;
  assign new_new_n13026__ = new_new_n13014__ & ~new_new_n13025__;
  assign new_new_n13027__ = ~new_new_n13017__ & ~new_new_n13026__;
  assign new_new_n13028__ = ~new_new_n12368__ & ~new_new_n12369__;
  assign new_new_n13029__ = ~new_new_n12379__ & new_new_n13028__;
  assign new_new_n13030__ = new_new_n12379__ & ~new_new_n13028__;
  assign new_new_n13031__ = ~new_new_n13029__ & ~new_new_n13030__;
  assign new_new_n13032__ = new_new_n13027__ & ~new_new_n13031__;
  assign new_new_n13033__ = ~new_new_n13027__ & new_new_n13031__;
  assign new_new_n13034__ = ~new_new_n2737__ & new_new_n11475__;
  assign new_new_n13035__ = new_new_n7814__ & new_new_n11478__;
  assign new_new_n13036__ = new_new_n2636__ & ~new_new_n11478__;
  assign new_new_n13037__ = ~new_new_n11482__ & ~new_new_n13036__;
  assign new_new_n13038__ = ~new_new_n13035__ & new_new_n13037__;
  assign new_new_n13039__ = ~new_new_n13034__ & ~new_new_n13038__;
  assign new_new_n13040__ = ~new_new_n2886__ & new_new_n11466__;
  assign new_new_n13041__ = pi05 & ~new_new_n13040__;
  assign new_new_n13042__ = ~new_new_n2886__ & new_new_n11467__;
  assign new_new_n13043__ = ~pi05 & ~new_new_n13042__;
  assign new_new_n13044__ = pi02 & ~new_new_n13043__;
  assign new_new_n13045__ = ~new_new_n13041__ & ~new_new_n13044__;
  assign new_new_n13046__ = new_new_n13039__ & ~new_new_n13045__;
  assign new_new_n13047__ = ~pi05 & ~new_new_n13039__;
  assign new_new_n13048__ = ~new_new_n13046__ & ~new_new_n13047__;
  assign new_new_n13049__ = ~new_new_n12338__ & ~new_new_n12339__;
  assign new_new_n13050__ = new_new_n12351__ & ~new_new_n13049__;
  assign new_new_n13051__ = ~new_new_n12351__ & new_new_n13049__;
  assign new_new_n13052__ = ~new_new_n13050__ & ~new_new_n13051__;
  assign new_new_n13053__ = new_new_n12264__ & new_new_n12318__;
  assign new_new_n13054__ = ~new_new_n12319__ & ~new_new_n13053__;
  assign new_new_n13055__ = new_new_n12323__ & ~new_new_n13054__;
  assign new_new_n13056__ = new_new_n12319__ & ~new_new_n12325__;
  assign new_new_n13057__ = new_new_n12328__ & ~new_new_n13056__;
  assign new_new_n13058__ = pi11 & new_new_n12325__;
  assign new_new_n13059__ = new_new_n12318__ & new_new_n13058__;
  assign new_new_n13060__ = ~new_new_n13055__ & ~new_new_n13059__;
  assign new_new_n13061__ = ~new_new_n13057__ & new_new_n13060__;
  assign new_new_n13062__ = ~new_new_n12271__ & ~new_new_n12273__;
  assign new_new_n13063__ = ~new_new_n10694__ & new_new_n13062__;
  assign new_new_n13064__ = pi08 & ~new_new_n13063__;
  assign new_new_n13065__ = ~new_new_n12278__ & new_new_n13064__;
  assign new_new_n13066__ = ~new_new_n12289__ & new_new_n13065__;
  assign new_new_n13067__ = new_new_n12289__ & ~new_new_n13065__;
  assign new_new_n13068__ = ~new_new_n13066__ & ~new_new_n13067__;
  assign new_new_n13069__ = new_new_n11478__ & ~new_new_n11482__;
  assign new_new_n13070__ = ~new_new_n8637__ & new_new_n13069__;
  assign new_new_n13071__ = ~new_new_n3164__ & new_new_n12850__;
  assign new_new_n13072__ = ~new_new_n3055__ & new_new_n11471__;
  assign new_new_n13073__ = ~new_new_n3254__ & new_new_n11475__;
  assign new_new_n13074__ = ~new_new_n13071__ & ~new_new_n13072__;
  assign new_new_n13075__ = ~new_new_n13073__ & new_new_n13074__;
  assign new_new_n13076__ = ~new_new_n13070__ & new_new_n13075__;
  assign new_new_n13077__ = ~new_new_n3055__ & new_new_n11469__;
  assign new_new_n13078__ = new_new_n3356__ & ~new_new_n13077__;
  assign new_new_n13079__ = ~new_new_n11470__ & ~new_new_n13078__;
  assign new_new_n13080__ = pi04 & new_new_n10726__;
  assign new_new_n13081__ = ~pi04 & new_new_n10731__;
  assign new_new_n13082__ = ~new_new_n13080__ & ~new_new_n13081__;
  assign new_new_n13083__ = new_new_n7682__ & new_new_n13069__;
  assign new_new_n13084__ = new_new_n13082__ & ~new_new_n13083__;
  assign new_new_n13085__ = ~new_new_n3055__ & ~new_new_n13084__;
  assign new_new_n13086__ = ~new_new_n3254__ & ~new_new_n11482__;
  assign new_new_n13087__ = ~new_new_n3356__ & new_new_n11471__;
  assign new_new_n13088__ = ~new_new_n13086__ & ~new_new_n13087__;
  assign new_new_n13089__ = ~new_new_n3055__ & new_new_n11478__;
  assign new_new_n13090__ = new_new_n3356__ & new_new_n13089__;
  assign new_new_n13091__ = ~new_new_n13088__ & ~new_new_n13090__;
  assign new_new_n13092__ = ~new_new_n13085__ & ~new_new_n13091__;
  assign new_new_n13093__ = pi05 & ~new_new_n13079__;
  assign new_new_n13094__ = new_new_n13092__ & new_new_n13093__;
  assign new_new_n13095__ = new_new_n13076__ & new_new_n13094__;
  assign new_new_n13096__ = pi06 & ~new_new_n13076__;
  assign new_new_n13097__ = pi05 & new_new_n13076__;
  assign new_new_n13098__ = ~new_new_n13096__ & ~new_new_n13097__;
  assign new_new_n13099__ = ~new_new_n3356__ & ~new_new_n9701__;
  assign new_new_n13100__ = ~new_new_n13098__ & new_new_n13099__;
  assign new_new_n13101__ = ~new_new_n13095__ & ~new_new_n13100__;
  assign new_new_n13102__ = ~new_new_n3055__ & ~new_new_n9697__;
  assign new_new_n13103__ = new_new_n10701__ & ~new_new_n13102__;
  assign new_new_n13104__ = ~new_new_n3356__ & new_new_n13102__;
  assign new_new_n13105__ = ~new_new_n9701__ & ~new_new_n13104__;
  assign new_new_n13106__ = pi07 & ~new_new_n13105__;
  assign new_new_n13107__ = ~new_new_n12278__ & ~new_new_n13103__;
  assign new_new_n13108__ = ~new_new_n13106__ & new_new_n13107__;
  assign new_new_n13109__ = ~new_new_n13101__ & new_new_n13108__;
  assign new_new_n13110__ = new_new_n13101__ & ~new_new_n13108__;
  assign new_new_n13111__ = new_new_n11482__ & new_new_n13082__;
  assign new_new_n13112__ = ~new_new_n3254__ & new_new_n13111__;
  assign new_new_n13113__ = ~new_new_n7570__ & new_new_n11469__;
  assign new_new_n13114__ = ~new_new_n13112__ & ~new_new_n13113__;
  assign new_new_n13115__ = new_new_n11478__ & ~new_new_n13114__;
  assign new_new_n13116__ = ~new_new_n3126__ & new_new_n12850__;
  assign new_new_n13117__ = ~new_new_n3164__ & new_new_n11475__;
  assign new_new_n13118__ = ~new_new_n13116__ & ~new_new_n13117__;
  assign new_new_n13119__ = ~new_new_n13115__ & new_new_n13118__;
  assign new_new_n13120__ = pi05 & ~new_new_n13119__;
  assign new_new_n13121__ = ~pi05 & new_new_n13119__;
  assign new_new_n13122__ = ~new_new_n13120__ & ~new_new_n13121__;
  assign new_new_n13123__ = ~new_new_n13110__ & new_new_n13122__;
  assign new_new_n13124__ = ~new_new_n13109__ & ~new_new_n13123__;
  assign new_new_n13125__ = new_new_n13068__ & ~new_new_n13124__;
  assign new_new_n13126__ = ~new_new_n13068__ & new_new_n13124__;
  assign new_new_n13127__ = ~new_new_n2960__ & new_new_n12850__;
  assign new_new_n13128__ = ~new_new_n3164__ & new_new_n11471__;
  assign new_new_n13129__ = ~new_new_n3126__ & new_new_n11475__;
  assign new_new_n13130__ = ~new_new_n13128__ & ~new_new_n13129__;
  assign new_new_n13131__ = ~new_new_n13127__ & new_new_n13130__;
  assign new_new_n13132__ = pi05 & ~new_new_n13131__;
  assign new_new_n13133__ = ~new_new_n7468__ & new_new_n12856__;
  assign new_new_n13134__ = ~new_new_n7468__ & new_new_n11469__;
  assign new_new_n13135__ = ~pi05 & ~new_new_n13134__;
  assign new_new_n13136__ = ~new_new_n13133__ & ~new_new_n13135__;
  assign new_new_n13137__ = new_new_n13131__ & ~new_new_n13136__;
  assign new_new_n13138__ = ~new_new_n13132__ & ~new_new_n13137__;
  assign new_new_n13139__ = ~new_new_n13126__ & new_new_n13138__;
  assign new_new_n13140__ = ~new_new_n13125__ & ~new_new_n13139__;
  assign new_new_n13141__ = new_new_n7391__ & new_new_n13069__;
  assign new_new_n13142__ = ~new_new_n3126__ & new_new_n11471__;
  assign new_new_n13143__ = ~new_new_n3460__ & new_new_n12850__;
  assign new_new_n13144__ = ~new_new_n2960__ & new_new_n11475__;
  assign new_new_n13145__ = ~new_new_n13142__ & ~new_new_n13143__;
  assign new_new_n13146__ = ~new_new_n13144__ & new_new_n13145__;
  assign new_new_n13147__ = ~new_new_n13141__ & new_new_n13146__;
  assign new_new_n13148__ = ~new_new_n13140__ & ~new_new_n13147__;
  assign new_new_n13149__ = new_new_n13140__ & new_new_n13147__;
  assign new_new_n13150__ = ~new_new_n13148__ & ~new_new_n13149__;
  assign new_new_n13151__ = pi05 & ~new_new_n13150__;
  assign new_new_n13152__ = ~pi05 & new_new_n13150__;
  assign new_new_n13153__ = ~new_new_n13151__ & ~new_new_n13152__;
  assign new_new_n13154__ = ~new_new_n13140__ & new_new_n13153__;
  assign new_new_n13155__ = pi09 & new_new_n12291__;
  assign new_new_n13156__ = pi08 & ~new_new_n12291__;
  assign new_new_n13157__ = new_new_n3356__ & ~new_new_n13156__;
  assign new_new_n13158__ = ~new_new_n13155__ & ~new_new_n13157__;
  assign new_new_n13159__ = new_new_n12298__ & ~new_new_n13158__;
  assign new_new_n13160__ = new_new_n3356__ & ~new_new_n12298__;
  assign new_new_n13161__ = new_new_n13156__ & new_new_n13160__;
  assign new_new_n13162__ = ~pi09 & new_new_n12298__;
  assign new_new_n13163__ = ~new_new_n12300__ & ~new_new_n13162__;
  assign new_new_n13164__ = ~new_new_n3356__ & ~new_new_n12299__;
  assign new_new_n13165__ = ~new_new_n13163__ & new_new_n13164__;
  assign new_new_n13166__ = ~new_new_n13161__ & ~new_new_n13165__;
  assign new_new_n13167__ = ~new_new_n13159__ & new_new_n13166__;
  assign new_new_n13168__ = ~new_new_n13153__ & new_new_n13167__;
  assign new_new_n13169__ = ~new_new_n13154__ & ~new_new_n13168__;
  assign new_new_n13170__ = ~new_new_n12305__ & ~new_new_n12306__;
  assign new_new_n13171__ = ~new_new_n12316__ & new_new_n13170__;
  assign new_new_n13172__ = new_new_n12316__ & ~new_new_n13170__;
  assign new_new_n13173__ = ~new_new_n13171__ & ~new_new_n13172__;
  assign new_new_n13174__ = ~new_new_n13169__ & ~new_new_n13173__;
  assign new_new_n13175__ = new_new_n13169__ & new_new_n13173__;
  assign new_new_n13176__ = ~new_new_n2960__ & new_new_n11471__;
  assign new_new_n13177__ = ~new_new_n2848__ & new_new_n12850__;
  assign new_new_n13178__ = ~new_new_n3460__ & new_new_n11475__;
  assign new_new_n13179__ = ~new_new_n13177__ & ~new_new_n13178__;
  assign new_new_n13180__ = ~new_new_n13176__ & new_new_n13179__;
  assign new_new_n13181__ = pi05 & ~new_new_n13180__;
  assign new_new_n13182__ = ~new_new_n7065__ & new_new_n12856__;
  assign new_new_n13183__ = ~new_new_n7065__ & new_new_n11469__;
  assign new_new_n13184__ = ~pi05 & ~new_new_n13183__;
  assign new_new_n13185__ = ~new_new_n13182__ & ~new_new_n13184__;
  assign new_new_n13186__ = new_new_n13180__ & ~new_new_n13185__;
  assign new_new_n13187__ = ~new_new_n13181__ & ~new_new_n13186__;
  assign new_new_n13188__ = ~new_new_n13175__ & new_new_n13187__;
  assign new_new_n13189__ = ~new_new_n13174__ & ~new_new_n13188__;
  assign new_new_n13190__ = ~new_new_n13061__ & ~new_new_n13189__;
  assign new_new_n13191__ = new_new_n13061__ & new_new_n13189__;
  assign new_new_n13192__ = ~new_new_n3460__ & new_new_n11471__;
  assign new_new_n13193__ = ~new_new_n2848__ & new_new_n11475__;
  assign new_new_n13194__ = new_new_n2886__ & ~new_new_n11478__;
  assign new_new_n13195__ = new_new_n8574__ & new_new_n11478__;
  assign new_new_n13196__ = ~new_new_n11482__ & ~new_new_n13194__;
  assign new_new_n13197__ = ~new_new_n13195__ & new_new_n13196__;
  assign new_new_n13198__ = ~new_new_n13192__ & ~new_new_n13193__;
  assign new_new_n13199__ = ~new_new_n13197__ & new_new_n13198__;
  assign new_new_n13200__ = ~pi05 & ~new_new_n13199__;
  assign new_new_n13201__ = pi05 & new_new_n13199__;
  assign new_new_n13202__ = ~new_new_n13200__ & ~new_new_n13201__;
  assign new_new_n13203__ = ~new_new_n13191__ & ~new_new_n13202__;
  assign new_new_n13204__ = ~new_new_n13190__ & ~new_new_n13203__;
  assign new_new_n13205__ = new_new_n13052__ & ~new_new_n13204__;
  assign new_new_n13206__ = ~new_new_n13052__ & new_new_n13204__;
  assign new_new_n13207__ = ~new_new_n2848__ & new_new_n11471__;
  assign new_new_n13208__ = ~new_new_n2886__ & new_new_n11475__;
  assign new_new_n13209__ = new_new_n7378__ & new_new_n11478__;
  assign new_new_n13210__ = new_new_n2737__ & ~new_new_n11478__;
  assign new_new_n13211__ = ~new_new_n11482__ & ~new_new_n13210__;
  assign new_new_n13212__ = ~new_new_n13209__ & new_new_n13211__;
  assign new_new_n13213__ = ~new_new_n13207__ & ~new_new_n13208__;
  assign new_new_n13214__ = ~new_new_n13212__ & new_new_n13213__;
  assign new_new_n13215__ = ~pi05 & ~new_new_n13214__;
  assign new_new_n13216__ = pi05 & new_new_n13214__;
  assign new_new_n13217__ = ~new_new_n13215__ & ~new_new_n13216__;
  assign new_new_n13218__ = ~new_new_n13206__ & ~new_new_n13217__;
  assign new_new_n13219__ = ~new_new_n13205__ & ~new_new_n13218__;
  assign new_new_n13220__ = new_new_n13048__ & new_new_n13219__;
  assign new_new_n13221__ = ~new_new_n13048__ & ~new_new_n13219__;
  assign new_new_n13222__ = ~new_new_n7065__ & new_new_n10694__;
  assign new_new_n13223__ = pi07 & ~new_new_n12252__;
  assign new_new_n13224__ = ~pi07 & new_new_n12252__;
  assign new_new_n13225__ = ~new_new_n13223__ & ~new_new_n13224__;
  assign new_new_n13226__ = new_new_n13222__ & ~new_new_n13225__;
  assign new_new_n13227__ = pi08 & new_new_n12252__;
  assign new_new_n13228__ = ~pi08 & ~new_new_n12252__;
  assign new_new_n13229__ = ~new_new_n13227__ & ~new_new_n13228__;
  assign new_new_n13230__ = ~new_new_n13222__ & new_new_n13229__;
  assign new_new_n13231__ = ~new_new_n13226__ & ~new_new_n13230__;
  assign new_new_n13232__ = new_new_n12360__ & ~new_new_n13231__;
  assign new_new_n13233__ = ~new_new_n12360__ & ~new_new_n13229__;
  assign new_new_n13234__ = ~new_new_n13232__ & ~new_new_n13233__;
  assign new_new_n13235__ = ~new_new_n12353__ & ~new_new_n13234__;
  assign new_new_n13236__ = new_new_n12353__ & new_new_n13234__;
  assign new_new_n13237__ = ~new_new_n13235__ & ~new_new_n13236__;
  assign new_new_n13238__ = ~new_new_n13221__ & ~new_new_n13237__;
  assign new_new_n13239__ = ~new_new_n13220__ & ~new_new_n13238__;
  assign new_new_n13240__ = ~new_new_n13033__ & new_new_n13239__;
  assign new_new_n13241__ = ~new_new_n13032__ & ~new_new_n13240__;
  assign new_new_n13242__ = new_new_n13011__ & ~new_new_n13241__;
  assign new_new_n13243__ = ~new_new_n13011__ & new_new_n13241__;
  assign new_new_n13244__ = ~new_new_n12394__ & ~new_new_n12405__;
  assign new_new_n13245__ = new_new_n12404__ & ~new_new_n13244__;
  assign new_new_n13246__ = ~new_new_n12404__ & new_new_n13244__;
  assign new_new_n13247__ = ~new_new_n13245__ & ~new_new_n13246__;
  assign new_new_n13248__ = ~new_new_n13243__ & ~new_new_n13247__;
  assign new_new_n13249__ = ~new_new_n13242__ & ~new_new_n13248__;
  assign new_new_n13250__ = ~new_new_n12430__ & ~new_new_n12431__;
  assign new_new_n13251__ = new_new_n12437__ & ~new_new_n13250__;
  assign new_new_n13252__ = ~new_new_n12437__ & new_new_n13250__;
  assign new_new_n13253__ = ~new_new_n13251__ & ~new_new_n13252__;
  assign new_new_n13254__ = ~new_new_n13249__ & new_new_n13253__;
  assign new_new_n13255__ = new_new_n13249__ & ~new_new_n13253__;
  assign new_new_n13256__ = ~new_new_n7236__ & new_new_n13069__;
  assign new_new_n13257__ = ~new_new_n2313__ & new_new_n12850__;
  assign new_new_n13258__ = ~new_new_n2497__ & new_new_n11471__;
  assign new_new_n13259__ = ~new_new_n2572__ & new_new_n11475__;
  assign new_new_n13260__ = ~new_new_n13257__ & ~new_new_n13258__;
  assign new_new_n13261__ = ~new_new_n13259__ & new_new_n13260__;
  assign new_new_n13262__ = ~new_new_n13256__ & new_new_n13261__;
  assign new_new_n13263__ = pi05 & ~new_new_n13262__;
  assign new_new_n13264__ = ~pi05 & new_new_n13262__;
  assign new_new_n13265__ = ~new_new_n13263__ & ~new_new_n13264__;
  assign new_new_n13266__ = ~new_new_n13255__ & new_new_n13265__;
  assign new_new_n13267__ = ~new_new_n13254__ & ~new_new_n13266__;
  assign new_new_n13268__ = ~new_new_n12999__ & ~new_new_n13267__;
  assign new_new_n13269__ = new_new_n12999__ & new_new_n13267__;
  assign new_new_n13270__ = ~new_new_n12469__ & ~new_new_n12470__;
  assign new_new_n13271__ = new_new_n12486__ & ~new_new_n13270__;
  assign new_new_n13272__ = ~new_new_n12486__ & new_new_n13270__;
  assign new_new_n13273__ = ~new_new_n13271__ & ~new_new_n13272__;
  assign new_new_n13274__ = ~new_new_n13269__ & new_new_n13273__;
  assign new_new_n13275__ = ~new_new_n13268__ & ~new_new_n13274__;
  assign new_new_n13276__ = ~new_new_n12986__ & ~new_new_n13275__;
  assign new_new_n13277__ = new_new_n12986__ & new_new_n13275__;
  assign new_new_n13278__ = ~new_new_n12494__ & ~new_new_n12495__;
  assign new_new_n13279__ = new_new_n12509__ & ~new_new_n13278__;
  assign new_new_n13280__ = ~new_new_n12509__ & new_new_n13278__;
  assign new_new_n13281__ = ~new_new_n13279__ & ~new_new_n13280__;
  assign new_new_n13282__ = ~new_new_n13277__ & new_new_n13281__;
  assign new_new_n13283__ = ~new_new_n13276__ & ~new_new_n13282__;
  assign new_new_n13284__ = ~new_new_n12975__ & ~new_new_n13283__;
  assign new_new_n13285__ = new_new_n12975__ & new_new_n13283__;
  assign new_new_n13286__ = ~new_new_n2024__ & new_new_n12850__;
  assign new_new_n13287__ = ~new_new_n2224__ & new_new_n11475__;
  assign new_new_n13288__ = ~new_new_n2420__ & new_new_n11471__;
  assign new_new_n13289__ = new_new_n7313__ & new_new_n13069__;
  assign new_new_n13290__ = ~new_new_n13286__ & ~new_new_n13287__;
  assign new_new_n13291__ = ~new_new_n13288__ & new_new_n13290__;
  assign new_new_n13292__ = ~new_new_n13289__ & new_new_n13291__;
  assign new_new_n13293__ = pi05 & ~new_new_n13292__;
  assign new_new_n13294__ = ~pi05 & new_new_n13292__;
  assign new_new_n13295__ = ~new_new_n13293__ & ~new_new_n13294__;
  assign new_new_n13296__ = ~new_new_n13285__ & new_new_n13295__;
  assign new_new_n13297__ = ~new_new_n13284__ & ~new_new_n13296__;
  assign new_new_n13298__ = ~new_new_n12971__ & ~new_new_n13297__;
  assign new_new_n13299__ = new_new_n12971__ & new_new_n13297__;
  assign new_new_n13300__ = ~new_new_n12518__ & ~new_new_n12519__;
  assign new_new_n13301__ = new_new_n12534__ & new_new_n13300__;
  assign new_new_n13302__ = ~new_new_n12534__ & ~new_new_n13300__;
  assign new_new_n13303__ = ~new_new_n13301__ & ~new_new_n13302__;
  assign new_new_n13304__ = ~new_new_n13299__ & ~new_new_n13303__;
  assign new_new_n13305__ = ~new_new_n13298__ & ~new_new_n13304__;
  assign new_new_n13306__ = pi08 & ~new_new_n12545__;
  assign new_new_n13307__ = ~pi08 & new_new_n12545__;
  assign new_new_n13308__ = ~new_new_n13306__ & ~new_new_n13307__;
  assign new_new_n13309__ = new_new_n12206__ & ~new_new_n12536__;
  assign new_new_n13310__ = ~new_new_n12206__ & new_new_n12536__;
  assign new_new_n13311__ = ~new_new_n13309__ & ~new_new_n13310__;
  assign new_new_n13312__ = new_new_n13308__ & new_new_n13311__;
  assign new_new_n13313__ = ~new_new_n13308__ & ~new_new_n13311__;
  assign new_new_n13314__ = ~new_new_n13312__ & ~new_new_n13313__;
  assign new_new_n13315__ = new_new_n13305__ & new_new_n13314__;
  assign new_new_n13316__ = ~new_new_n13305__ & ~new_new_n13314__;
  assign new_new_n13317__ = ~new_new_n3535__ & new_new_n12850__;
  assign new_new_n13318__ = ~new_new_n2130__ & new_new_n11475__;
  assign new_new_n13319__ = ~new_new_n2024__ & new_new_n11471__;
  assign new_new_n13320__ = new_new_n6854__ & new_new_n13069__;
  assign new_new_n13321__ = ~new_new_n13317__ & ~new_new_n13318__;
  assign new_new_n13322__ = ~new_new_n13319__ & new_new_n13321__;
  assign new_new_n13323__ = ~new_new_n13320__ & new_new_n13322__;
  assign new_new_n13324__ = pi05 & ~new_new_n13323__;
  assign new_new_n13325__ = ~pi05 & new_new_n13323__;
  assign new_new_n13326__ = ~new_new_n13324__ & ~new_new_n13325__;
  assign new_new_n13327__ = ~new_new_n13316__ & ~new_new_n13326__;
  assign new_new_n13328__ = ~new_new_n13315__ & ~new_new_n13327__;
  assign new_new_n13329__ = new_new_n12959__ & ~new_new_n13328__;
  assign new_new_n13330__ = ~new_new_n12959__ & new_new_n13328__;
  assign new_new_n13331__ = ~new_new_n2130__ & new_new_n12832__;
  assign new_new_n13332__ = ~new_new_n3535__ & new_new_n11475__;
  assign new_new_n13333__ = ~new_new_n13331__ & ~new_new_n13332__;
  assign new_new_n13334__ = new_new_n6553__ & new_new_n11469__;
  assign new_new_n13335__ = new_new_n13333__ & ~new_new_n13334__;
  assign new_new_n13336__ = pi05 & ~new_new_n13335__;
  assign new_new_n13337__ = ~new_new_n5520__ & new_new_n11469__;
  assign new_new_n13338__ = ~pi05 & ~new_new_n13337__;
  assign new_new_n13339__ = pi04 & new_new_n1823__;
  assign new_new_n13340__ = ~pi04 & ~new_new_n1823__;
  assign new_new_n13341__ = ~new_new_n11482__ & ~new_new_n13339__;
  assign new_new_n13342__ = ~new_new_n13340__ & new_new_n13341__;
  assign new_new_n13343__ = new_new_n5501__ & new_new_n13342__;
  assign new_new_n13344__ = ~new_new_n13338__ & ~new_new_n13343__;
  assign new_new_n13345__ = new_new_n13333__ & ~new_new_n13344__;
  assign new_new_n13346__ = ~new_new_n13336__ & ~new_new_n13345__;
  assign new_new_n13347__ = ~new_new_n13330__ & ~new_new_n13346__;
  assign new_new_n13348__ = ~new_new_n13329__ & ~new_new_n13347__;
  assign new_new_n13349__ = ~new_new_n12955__ & new_new_n13348__;
  assign new_new_n13350__ = new_new_n12955__ & ~new_new_n13348__;
  assign new_new_n13351__ = ~new_new_n12565__ & ~new_new_n12566__;
  assign new_new_n13352__ = new_new_n12576__ & ~new_new_n13351__;
  assign new_new_n13353__ = ~new_new_n12576__ & new_new_n13351__;
  assign new_new_n13354__ = ~new_new_n13352__ & ~new_new_n13353__;
  assign new_new_n13355__ = ~new_new_n13350__ & ~new_new_n13354__;
  assign new_new_n13356__ = ~new_new_n13349__ & ~new_new_n13355__;
  assign new_new_n13357__ = new_new_n12942__ & ~new_new_n13356__;
  assign new_new_n13358__ = ~new_new_n12942__ & new_new_n13356__;
  assign new_new_n13359__ = ~new_new_n1660__ & new_new_n12850__;
  assign new_new_n13360__ = ~new_new_n1823__ & new_new_n13111__;
  assign new_new_n13361__ = ~new_new_n5274__ & new_new_n11469__;
  assign new_new_n13362__ = ~new_new_n13360__ & ~new_new_n13361__;
  assign new_new_n13363__ = new_new_n11478__ & ~new_new_n13362__;
  assign new_new_n13364__ = ~new_new_n1902__ & new_new_n11475__;
  assign new_new_n13365__ = ~new_new_n13359__ & ~new_new_n13364__;
  assign new_new_n13366__ = ~new_new_n13363__ & new_new_n13365__;
  assign new_new_n13367__ = ~pi05 & ~new_new_n13366__;
  assign new_new_n13368__ = pi05 & new_new_n13366__;
  assign new_new_n13369__ = ~new_new_n13367__ & ~new_new_n13368__;
  assign new_new_n13370__ = ~new_new_n13358__ & ~new_new_n13369__;
  assign new_new_n13371__ = ~new_new_n13357__ & ~new_new_n13370__;
  assign new_new_n13372__ = ~new_new_n12938__ & new_new_n13371__;
  assign new_new_n13373__ = new_new_n12938__ & ~new_new_n13371__;
  assign new_new_n13374__ = ~new_new_n12179__ & ~new_new_n12604__;
  assign new_new_n13375__ = new_new_n12179__ & new_new_n12604__;
  assign new_new_n13376__ = ~new_new_n13374__ & ~new_new_n13375__;
  assign new_new_n13377__ = new_new_n12592__ & new_new_n13376__;
  assign new_new_n13378__ = ~new_new_n12592__ & ~new_new_n13376__;
  assign new_new_n13379__ = ~new_new_n13377__ & ~new_new_n13378__;
  assign new_new_n13380__ = ~new_new_n13373__ & ~new_new_n13379__;
  assign new_new_n13381__ = ~new_new_n13372__ & ~new_new_n13380__;
  assign new_new_n13382__ = ~new_new_n12926__ & new_new_n13381__;
  assign new_new_n13383__ = new_new_n12926__ & ~new_new_n13381__;
  assign new_new_n13384__ = ~new_new_n1466__ & new_new_n12850__;
  assign new_new_n13385__ = ~new_new_n1737__ & new_new_n11475__;
  assign new_new_n13386__ = ~new_new_n1660__ & new_new_n11471__;
  assign new_new_n13387__ = ~new_new_n6410__ & new_new_n13069__;
  assign new_new_n13388__ = ~new_new_n13384__ & ~new_new_n13385__;
  assign new_new_n13389__ = ~new_new_n13386__ & new_new_n13388__;
  assign new_new_n13390__ = ~new_new_n13387__ & new_new_n13389__;
  assign new_new_n13391__ = ~pi05 & ~new_new_n13390__;
  assign new_new_n13392__ = pi05 & new_new_n13390__;
  assign new_new_n13393__ = ~new_new_n13391__ & ~new_new_n13392__;
  assign new_new_n13394__ = ~new_new_n13383__ & ~new_new_n13393__;
  assign new_new_n13395__ = ~new_new_n13382__ & ~new_new_n13394__;
  assign new_new_n13396__ = ~new_new_n12918__ & new_new_n13395__;
  assign new_new_n13397__ = new_new_n12918__ & ~new_new_n13395__;
  assign new_new_n13398__ = ~new_new_n1737__ & new_new_n13111__;
  assign new_new_n13399__ = ~new_new_n5671__ & new_new_n11469__;
  assign new_new_n13400__ = ~new_new_n13398__ & ~new_new_n13399__;
  assign new_new_n13401__ = new_new_n11478__ & ~new_new_n13400__;
  assign new_new_n13402__ = ~new_new_n1466__ & new_new_n11475__;
  assign new_new_n13403__ = ~new_new_n13401__ & ~new_new_n13402__;
  assign new_new_n13404__ = ~pi05 & ~new_new_n13403__;
  assign new_new_n13405__ = ~new_new_n1556__ & new_new_n12856__;
  assign new_new_n13406__ = ~new_new_n1556__ & new_new_n11469__;
  assign new_new_n13407__ = pi05 & ~new_new_n13406__;
  assign new_new_n13408__ = ~new_new_n13405__ & ~new_new_n13407__;
  assign new_new_n13409__ = new_new_n13403__ & ~new_new_n13408__;
  assign new_new_n13410__ = ~new_new_n13404__ & ~new_new_n13409__;
  assign new_new_n13411__ = ~new_new_n13397__ & new_new_n13410__;
  assign new_new_n13412__ = ~new_new_n13396__ & ~new_new_n13411__;
  assign new_new_n13413__ = new_new_n12905__ & new_new_n13412__;
  assign new_new_n13414__ = ~new_new_n12905__ & ~new_new_n13412__;
  assign new_new_n13415__ = ~new_new_n1466__ & new_new_n11471__;
  assign new_new_n13416__ = ~new_new_n1325__ & new_new_n12850__;
  assign new_new_n13417__ = ~new_new_n1556__ & new_new_n11475__;
  assign new_new_n13418__ = ~new_new_n13415__ & ~new_new_n13416__;
  assign new_new_n13419__ = ~new_new_n13417__ & new_new_n13418__;
  assign new_new_n13420__ = pi05 & ~new_new_n13419__;
  assign new_new_n13421__ = new_new_n5048__ & new_new_n12856__;
  assign new_new_n13422__ = new_new_n5048__ & new_new_n11469__;
  assign new_new_n13423__ = ~pi05 & ~new_new_n13422__;
  assign new_new_n13424__ = ~new_new_n13421__ & ~new_new_n13423__;
  assign new_new_n13425__ = new_new_n13419__ & ~new_new_n13424__;
  assign new_new_n13426__ = ~new_new_n13420__ & ~new_new_n13425__;
  assign new_new_n13427__ = ~new_new_n13414__ & new_new_n13426__;
  assign new_new_n13428__ = ~new_new_n12914__ & ~new_new_n13413__;
  assign new_new_n13429__ = ~new_new_n13427__ & new_new_n13428__;
  assign new_new_n13430__ = ~new_new_n12913__ & ~new_new_n13429__;
  assign new_new_n13431__ = ~new_new_n12883__ & new_new_n13430__;
  assign new_new_n13432__ = new_new_n12883__ & ~new_new_n13430__;
  assign new_new_n13433__ = ~new_new_n1061__ & new_new_n12850__;
  assign new_new_n13434__ = ~new_new_n3618__ & new_new_n11475__;
  assign new_new_n13435__ = ~new_new_n1325__ & new_new_n11471__;
  assign new_new_n13436__ = new_new_n4926__ & new_new_n13069__;
  assign new_new_n13437__ = ~new_new_n13433__ & ~new_new_n13434__;
  assign new_new_n13438__ = ~new_new_n13435__ & new_new_n13437__;
  assign new_new_n13439__ = ~new_new_n13436__ & new_new_n13438__;
  assign new_new_n13440__ = pi05 & ~new_new_n13439__;
  assign new_new_n13441__ = ~pi05 & new_new_n13439__;
  assign new_new_n13442__ = ~new_new_n13440__ & ~new_new_n13441__;
  assign new_new_n13443__ = ~new_new_n13432__ & new_new_n13442__;
  assign new_new_n13444__ = ~new_new_n13431__ & ~new_new_n13443__;
  assign new_new_n13445__ = ~new_new_n12879__ & ~new_new_n13444__;
  assign new_new_n13446__ = new_new_n12879__ & new_new_n13444__;
  assign new_new_n13447__ = ~new_new_n12677__ & ~new_new_n12678__;
  assign new_new_n13448__ = new_new_n12688__ & new_new_n13447__;
  assign new_new_n13449__ = ~new_new_n12688__ & ~new_new_n13447__;
  assign new_new_n13450__ = ~new_new_n13448__ & ~new_new_n13449__;
  assign new_new_n13451__ = ~new_new_n13446__ & ~new_new_n13450__;
  assign new_new_n13452__ = ~new_new_n13445__ & ~new_new_n13451__;
  assign new_new_n13453__ = new_new_n12866__ & ~new_new_n13452__;
  assign new_new_n13454__ = ~new_new_n12866__ & new_new_n13452__;
  assign new_new_n13455__ = ~new_new_n868__ & new_new_n12850__;
  assign new_new_n13456__ = ~new_new_n1061__ & new_new_n11471__;
  assign new_new_n13457__ = ~new_new_n1207__ & new_new_n11475__;
  assign new_new_n13458__ = ~new_new_n13455__ & ~new_new_n13456__;
  assign new_new_n13459__ = ~new_new_n13457__ & new_new_n13458__;
  assign new_new_n13460__ = ~pi05 & ~new_new_n13459__;
  assign new_new_n13461__ = ~new_new_n4550__ & new_new_n12873__;
  assign new_new_n13462__ = ~new_new_n4550__ & new_new_n11469__;
  assign new_new_n13463__ = pi05 & ~new_new_n13462__;
  assign new_new_n13464__ = ~new_new_n13461__ & ~new_new_n13463__;
  assign new_new_n13465__ = new_new_n13459__ & ~new_new_n13464__;
  assign new_new_n13466__ = ~new_new_n13460__ & ~new_new_n13465__;
  assign new_new_n13467__ = ~new_new_n13454__ & ~new_new_n13466__;
  assign new_new_n13468__ = ~new_new_n13453__ & ~new_new_n13467__;
  assign new_new_n13469__ = new_new_n12862__ & ~new_new_n13468__;
  assign new_new_n13470__ = ~new_new_n12862__ & new_new_n13468__;
  assign new_new_n13471__ = new_new_n4926__ & new_new_n10694__;
  assign new_new_n13472__ = pi08 & new_new_n12696__;
  assign new_new_n13473__ = ~pi08 & ~new_new_n12696__;
  assign new_new_n13474__ = ~new_new_n13472__ & ~new_new_n13473__;
  assign new_new_n13475__ = ~new_new_n13471__ & ~new_new_n13474__;
  assign new_new_n13476__ = pi07 & new_new_n12696__;
  assign new_new_n13477__ = ~pi07 & ~new_new_n12696__;
  assign new_new_n13478__ = ~new_new_n13476__ & ~new_new_n13477__;
  assign new_new_n13479__ = new_new_n13471__ & ~new_new_n13478__;
  assign new_new_n13480__ = ~new_new_n13475__ & ~new_new_n13479__;
  assign new_new_n13481__ = new_new_n12703__ & ~new_new_n13480__;
  assign new_new_n13482__ = ~new_new_n12703__ & new_new_n13474__;
  assign new_new_n13483__ = ~new_new_n13481__ & ~new_new_n13482__;
  assign new_new_n13484__ = ~new_new_n12692__ & new_new_n13483__;
  assign new_new_n13485__ = new_new_n12692__ & ~new_new_n13483__;
  assign new_new_n13486__ = ~new_new_n13484__ & ~new_new_n13485__;
  assign new_new_n13487__ = ~new_new_n13470__ & new_new_n13486__;
  assign new_new_n13488__ = ~new_new_n13469__ & ~new_new_n13487__;
  assign new_new_n13489__ = new_new_n12848__ & new_new_n13488__;
  assign new_new_n13490__ = ~new_new_n12848__ & ~new_new_n13488__;
  assign new_new_n13491__ = ~new_new_n13489__ & ~new_new_n13490__;
  assign new_new_n13492__ = ~new_new_n12711__ & ~new_new_n12712__;
  assign new_new_n13493__ = ~new_new_n12724__ & new_new_n13492__;
  assign new_new_n13494__ = new_new_n12724__ & ~new_new_n13492__;
  assign new_new_n13495__ = ~new_new_n13493__ & ~new_new_n13494__;
  assign new_new_n13496__ = new_new_n13491__ & ~new_new_n13495__;
  assign new_new_n13497__ = ~new_new_n13491__ & new_new_n13495__;
  assign new_new_n13498__ = ~new_new_n13496__ & ~new_new_n13497__;
  assign new_new_n13499__ = new_new_n12827__ & new_new_n13498__;
  assign new_new_n13500__ = ~new_new_n12827__ & ~new_new_n13498__;
  assign new_new_n13501__ = pi02 & ~new_new_n4039__;
  assign new_new_n13502__ = pi01 & new_new_n4039__;
  assign new_new_n13503__ = ~new_new_n13501__ & ~new_new_n13502__;
  assign new_new_n13504__ = new_new_n691__ & ~new_new_n13503__;
  assign new_new_n13505__ = ~new_new_n691__ & new_new_n13503__;
  assign new_new_n13506__ = pi00 & ~new_new_n13504__;
  assign new_new_n13507__ = ~new_new_n13505__ & new_new_n13506__;
  assign new_new_n13508__ = pi01 & ~pi02;
  assign new_new_n13509__ = ~new_new_n910__ & new_new_n13508__;
  assign new_new_n13510__ = ~pi01 & ~new_new_n3720__;
  assign new_new_n13511__ = pi01 & ~new_new_n910__;
  assign new_new_n13512__ = pi02 & ~new_new_n13510__;
  assign new_new_n13513__ = ~new_new_n13511__ & new_new_n13512__;
  assign new_new_n13514__ = ~pi00 & ~new_new_n13509__;
  assign new_new_n13515__ = ~new_new_n13513__ & new_new_n13514__;
  assign new_new_n13516__ = ~new_new_n13507__ & ~new_new_n13515__;
  assign new_new_n13517__ = ~new_new_n3720__ & new_new_n13508__;
  assign new_new_n13518__ = pi01 & ~new_new_n3720__;
  assign new_new_n13519__ = ~pi01 & ~new_new_n868__;
  assign new_new_n13520__ = pi02 & ~new_new_n13518__;
  assign new_new_n13521__ = ~new_new_n13519__ & new_new_n13520__;
  assign new_new_n13522__ = ~pi00 & ~new_new_n13517__;
  assign new_new_n13523__ = ~new_new_n13521__ & new_new_n13522__;
  assign new_new_n13524__ = pi02 & ~new_new_n4036__;
  assign new_new_n13525__ = pi01 & new_new_n4036__;
  assign new_new_n13526__ = ~new_new_n13524__ & ~new_new_n13525__;
  assign new_new_n13527__ = new_new_n910__ & ~new_new_n13526__;
  assign new_new_n13528__ = ~new_new_n910__ & new_new_n13526__;
  assign new_new_n13529__ = pi00 & ~new_new_n13527__;
  assign new_new_n13530__ = ~new_new_n13528__ & new_new_n13529__;
  assign new_new_n13531__ = ~new_new_n13523__ & ~new_new_n13530__;
  assign new_new_n13532__ = ~new_new_n13445__ & ~new_new_n13446__;
  assign new_new_n13533__ = ~new_new_n13450__ & new_new_n13532__;
  assign new_new_n13534__ = new_new_n13450__ & ~new_new_n13532__;
  assign new_new_n13535__ = ~new_new_n13533__ & ~new_new_n13534__;
  assign new_new_n13536__ = ~new_new_n13531__ & ~new_new_n13535__;
  assign new_new_n13537__ = new_new_n13531__ & new_new_n13535__;
  assign new_new_n13538__ = ~pi02 & ~new_new_n868__;
  assign new_new_n13539__ = pi01 & new_new_n868__;
  assign new_new_n13540__ = ~new_new_n13538__ & ~new_new_n13539__;
  assign new_new_n13541__ = ~new_new_n4550__ & ~new_new_n13540__;
  assign new_new_n13542__ = pi02 & new_new_n868__;
  assign new_new_n13543__ = ~new_new_n13519__ & ~new_new_n13542__;
  assign new_new_n13544__ = new_new_n4550__ & ~new_new_n13543__;
  assign new_new_n13545__ = pi00 & ~new_new_n13541__;
  assign new_new_n13546__ = ~new_new_n13544__ & new_new_n13545__;
  assign new_new_n13547__ = ~new_new_n1207__ & new_new_n13508__;
  assign new_new_n13548__ = ~pi01 & ~new_new_n1061__;
  assign new_new_n13549__ = pi01 & ~new_new_n1207__;
  assign new_new_n13550__ = pi02 & ~new_new_n13548__;
  assign new_new_n13551__ = ~new_new_n13549__ & new_new_n13550__;
  assign new_new_n13552__ = ~pi00 & ~new_new_n13547__;
  assign new_new_n13553__ = ~new_new_n13551__ & new_new_n13552__;
  assign new_new_n13554__ = ~new_new_n13546__ & ~new_new_n13553__;
  assign new_new_n13555__ = ~new_new_n1061__ & new_new_n13508__;
  assign new_new_n13556__ = pi01 & new_new_n1061__;
  assign new_new_n13557__ = ~pi01 & new_new_n3618__;
  assign new_new_n13558__ = ~new_new_n13556__ & ~new_new_n13557__;
  assign new_new_n13559__ = pi02 & ~new_new_n13558__;
  assign new_new_n13560__ = ~pi00 & ~new_new_n13555__;
  assign new_new_n13561__ = ~new_new_n13559__ & new_new_n13560__;
  assign new_new_n13562__ = ~pi01 & new_new_n1207__;
  assign new_new_n13563__ = pi02 & ~new_new_n1207__;
  assign new_new_n13564__ = ~new_new_n13562__ & ~new_new_n13563__;
  assign new_new_n13565__ = ~new_new_n5235__ & new_new_n13564__;
  assign new_new_n13566__ = ~pi02 & new_new_n1207__;
  assign new_new_n13567__ = ~new_new_n13549__ & ~new_new_n13566__;
  assign new_new_n13568__ = new_new_n5235__ & new_new_n13567__;
  assign new_new_n13569__ = pi00 & ~new_new_n13565__;
  assign new_new_n13570__ = ~new_new_n13568__ & new_new_n13569__;
  assign new_new_n13571__ = ~new_new_n13561__ & ~new_new_n13570__;
  assign new_new_n13572__ = ~new_new_n3618__ & new_new_n13508__;
  assign new_new_n13573__ = pi01 & new_new_n3618__;
  assign new_new_n13574__ = ~pi01 & new_new_n1325__;
  assign new_new_n13575__ = ~new_new_n13573__ & ~new_new_n13574__;
  assign new_new_n13576__ = pi02 & ~new_new_n13575__;
  assign new_new_n13577__ = ~new_new_n13572__ & ~new_new_n13576__;
  assign new_new_n13578__ = ~pi00 & ~new_new_n13577__;
  assign new_new_n13579__ = ~new_new_n3553__ & ~new_new_n3618__;
  assign new_new_n13580__ = ~new_new_n5982__ & ~new_new_n13579__;
  assign new_new_n13581__ = ~new_new_n13548__ & ~new_new_n13556__;
  assign new_new_n13582__ = new_new_n13580__ & new_new_n13581__;
  assign new_new_n13583__ = ~pi02 & ~new_new_n1061__;
  assign new_new_n13584__ = pi02 & new_new_n1061__;
  assign new_new_n13585__ = ~new_new_n13583__ & ~new_new_n13584__;
  assign new_new_n13586__ = ~new_new_n13580__ & new_new_n13585__;
  assign new_new_n13587__ = pi00 & ~new_new_n13582__;
  assign new_new_n13588__ = ~new_new_n13586__ & new_new_n13587__;
  assign new_new_n13589__ = ~new_new_n13578__ & ~new_new_n13588__;
  assign new_new_n13590__ = pi02 & ~new_new_n4921__;
  assign new_new_n13591__ = pi01 & new_new_n4921__;
  assign new_new_n13592__ = ~new_new_n13590__ & ~new_new_n13591__;
  assign new_new_n13593__ = ~new_new_n3618__ & new_new_n13592__;
  assign new_new_n13594__ = new_new_n3618__ & ~new_new_n13592__;
  assign new_new_n13595__ = pi00 & ~new_new_n13593__;
  assign new_new_n13596__ = ~new_new_n13594__ & new_new_n13595__;
  assign new_new_n13597__ = ~new_new_n1325__ & new_new_n13508__;
  assign new_new_n13598__ = ~pi01 & ~new_new_n1556__;
  assign new_new_n13599__ = pi01 & ~new_new_n1325__;
  assign new_new_n13600__ = pi02 & ~new_new_n13598__;
  assign new_new_n13601__ = ~new_new_n13599__ & new_new_n13600__;
  assign new_new_n13602__ = ~pi00 & ~new_new_n13597__;
  assign new_new_n13603__ = ~new_new_n13601__ & new_new_n13602__;
  assign new_new_n13604__ = ~new_new_n13596__ & ~new_new_n13603__;
  assign new_new_n13605__ = ~new_new_n13382__ & ~new_new_n13383__;
  assign new_new_n13606__ = new_new_n13393__ & new_new_n13605__;
  assign new_new_n13607__ = ~new_new_n13393__ & ~new_new_n13605__;
  assign new_new_n13608__ = ~new_new_n13606__ & ~new_new_n13607__;
  assign new_new_n13609__ = new_new_n13604__ & ~new_new_n13608__;
  assign new_new_n13610__ = ~new_new_n13604__ & new_new_n13608__;
  assign new_new_n13611__ = ~new_new_n1556__ & new_new_n13508__;
  assign new_new_n13612__ = ~pi01 & new_new_n1466__;
  assign new_new_n13613__ = pi01 & new_new_n1556__;
  assign new_new_n13614__ = ~new_new_n13612__ & ~new_new_n13613__;
  assign new_new_n13615__ = pi02 & ~new_new_n13614__;
  assign new_new_n13616__ = ~pi00 & ~new_new_n13611__;
  assign new_new_n13617__ = ~new_new_n13615__ & new_new_n13616__;
  assign new_new_n13618__ = ~pi02 & new_new_n1325__;
  assign new_new_n13619__ = ~new_new_n13599__ & ~new_new_n13618__;
  assign new_new_n13620__ = ~new_new_n5048__ & new_new_n13619__;
  assign new_new_n13621__ = pi02 & ~new_new_n1325__;
  assign new_new_n13622__ = ~new_new_n13574__ & ~new_new_n13621__;
  assign new_new_n13623__ = new_new_n5048__ & new_new_n13622__;
  assign new_new_n13624__ = pi00 & ~new_new_n13620__;
  assign new_new_n13625__ = ~new_new_n13623__ & new_new_n13624__;
  assign new_new_n13626__ = ~new_new_n13372__ & ~new_new_n13373__;
  assign new_new_n13627__ = ~new_new_n12592__ & new_new_n13376__;
  assign new_new_n13628__ = new_new_n12592__ & ~new_new_n13376__;
  assign new_new_n13629__ = ~new_new_n13627__ & ~new_new_n13628__;
  assign new_new_n13630__ = new_new_n13626__ & new_new_n13629__;
  assign new_new_n13631__ = ~new_new_n13626__ & ~new_new_n13629__;
  assign new_new_n13632__ = ~new_new_n13630__ & ~new_new_n13631__;
  assign new_new_n13633__ = ~pi02 & new_new_n5671__;
  assign new_new_n13634__ = pi02 & ~new_new_n1556__;
  assign new_new_n13635__ = pi01 & ~new_new_n13634__;
  assign new_new_n13636__ = ~new_new_n13633__ & new_new_n13635__;
  assign new_new_n13637__ = ~pi02 & new_new_n1556__;
  assign new_new_n13638__ = pi02 & ~new_new_n5671__;
  assign new_new_n13639__ = ~pi01 & ~new_new_n13637__;
  assign new_new_n13640__ = ~new_new_n13638__ & new_new_n13639__;
  assign new_new_n13641__ = ~new_new_n13636__ & ~new_new_n13640__;
  assign new_new_n13642__ = pi00 & ~new_new_n13641__;
  assign new_new_n13643__ = pi02 & new_new_n1737__;
  assign new_new_n13644__ = ~pi01 & ~new_new_n13643__;
  assign new_new_n13645__ = pi02 & ~new_new_n1466__;
  assign new_new_n13646__ = ~pi02 & new_new_n1466__;
  assign new_new_n13647__ = ~new_new_n13645__ & ~new_new_n13646__;
  assign new_new_n13648__ = pi01 & ~new_new_n13647__;
  assign new_new_n13649__ = ~pi00 & ~new_new_n13644__;
  assign new_new_n13650__ = ~new_new_n13648__ & new_new_n13649__;
  assign new_new_n13651__ = ~new_new_n13642__ & ~new_new_n13650__;
  assign new_new_n13652__ = ~new_new_n13357__ & ~new_new_n13358__;
  assign new_new_n13653__ = ~new_new_n13369__ & new_new_n13652__;
  assign new_new_n13654__ = new_new_n13369__ & ~new_new_n13652__;
  assign new_new_n13655__ = ~new_new_n13653__ & ~new_new_n13654__;
  assign new_new_n13656__ = new_new_n13651__ & ~new_new_n13655__;
  assign new_new_n13657__ = ~new_new_n13651__ & new_new_n13655__;
  assign new_new_n13658__ = new_new_n12187__ & ~new_new_n12564__;
  assign new_new_n13659__ = ~new_new_n12187__ & new_new_n12564__;
  assign new_new_n13660__ = ~new_new_n13658__ & ~new_new_n13659__;
  assign new_new_n13661__ = new_new_n13348__ & new_new_n13660__;
  assign new_new_n13662__ = ~new_new_n13348__ & ~new_new_n13660__;
  assign new_new_n13663__ = ~new_new_n13661__ & ~new_new_n13662__;
  assign new_new_n13664__ = new_new_n12576__ & ~new_new_n13663__;
  assign new_new_n13665__ = ~new_new_n12576__ & new_new_n13663__;
  assign new_new_n13666__ = ~new_new_n13664__ & ~new_new_n13665__;
  assign new_new_n13667__ = new_new_n12955__ & new_new_n13666__;
  assign new_new_n13668__ = ~new_new_n12955__ & ~new_new_n13666__;
  assign new_new_n13669__ = pi01 & new_new_n1737__;
  assign new_new_n13670__ = ~pi01 & new_new_n1660__;
  assign new_new_n13671__ = ~new_new_n13669__ & ~new_new_n13670__;
  assign new_new_n13672__ = pi02 & ~new_new_n13671__;
  assign new_new_n13673__ = ~new_new_n1737__ & new_new_n13508__;
  assign new_new_n13674__ = ~new_new_n13672__ & ~new_new_n13673__;
  assign new_new_n13675__ = ~pi00 & ~new_new_n13674__;
  assign new_new_n13676__ = pi01 & ~new_new_n1466__;
  assign new_new_n13677__ = ~new_new_n13612__ & ~new_new_n13676__;
  assign new_new_n13678__ = new_new_n5664__ & ~new_new_n13677__;
  assign new_new_n13679__ = ~new_new_n5664__ & ~new_new_n13647__;
  assign new_new_n13680__ = pi00 & ~new_new_n13678__;
  assign new_new_n13681__ = ~new_new_n13679__ & new_new_n13680__;
  assign new_new_n13682__ = ~new_new_n13675__ & ~new_new_n13681__;
  assign new_new_n13683__ = ~pi01 & ~new_new_n1737__;
  assign new_new_n13684__ = ~new_new_n13643__ & ~new_new_n13683__;
  assign new_new_n13685__ = ~new_new_n5688__ & ~new_new_n13684__;
  assign new_new_n13686__ = ~pi02 & ~new_new_n1737__;
  assign new_new_n13687__ = ~new_new_n13669__ & ~new_new_n13686__;
  assign new_new_n13688__ = new_new_n5688__ & ~new_new_n13687__;
  assign new_new_n13689__ = pi00 & ~new_new_n13685__;
  assign new_new_n13690__ = ~new_new_n13688__ & new_new_n13689__;
  assign new_new_n13691__ = ~new_new_n1660__ & new_new_n13508__;
  assign new_new_n13692__ = ~pi01 & ~new_new_n1902__;
  assign new_new_n13693__ = pi01 & ~new_new_n1660__;
  assign new_new_n13694__ = pi02 & ~new_new_n13692__;
  assign new_new_n13695__ = ~new_new_n13693__ & new_new_n13694__;
  assign new_new_n13696__ = ~pi00 & ~new_new_n13691__;
  assign new_new_n13697__ = ~new_new_n13695__ & new_new_n13696__;
  assign new_new_n13698__ = ~new_new_n13690__ & ~new_new_n13697__;
  assign new_new_n13699__ = ~pi01 & ~new_new_n5274__;
  assign new_new_n13700__ = ~pi02 & new_new_n5274__;
  assign new_new_n13701__ = new_new_n1660__ & ~new_new_n13699__;
  assign new_new_n13702__ = ~new_new_n13700__ & new_new_n13701__;
  assign new_new_n13703__ = pi01 & new_new_n5274__;
  assign new_new_n13704__ = pi02 & ~new_new_n5274__;
  assign new_new_n13705__ = ~new_new_n1660__ & ~new_new_n13703__;
  assign new_new_n13706__ = ~new_new_n13704__ & new_new_n13705__;
  assign new_new_n13707__ = ~new_new_n13702__ & ~new_new_n13706__;
  assign new_new_n13708__ = pi00 & ~new_new_n13707__;
  assign new_new_n13709__ = pi02 & new_new_n1823__;
  assign new_new_n13710__ = ~pi01 & ~new_new_n13709__;
  assign new_new_n13711__ = pi02 & ~new_new_n1902__;
  assign new_new_n13712__ = ~pi02 & new_new_n1902__;
  assign new_new_n13713__ = ~new_new_n13711__ & ~new_new_n13712__;
  assign new_new_n13714__ = pi01 & ~new_new_n13713__;
  assign new_new_n13715__ = ~pi00 & ~new_new_n13710__;
  assign new_new_n13716__ = ~new_new_n13714__ & new_new_n13715__;
  assign new_new_n13717__ = ~new_new_n13708__ & ~new_new_n13716__;
  assign new_new_n13718__ = ~new_new_n13315__ & ~new_new_n13316__;
  assign new_new_n13719__ = new_new_n13326__ & ~new_new_n13718__;
  assign new_new_n13720__ = ~new_new_n13326__ & new_new_n13718__;
  assign new_new_n13721__ = ~new_new_n13719__ & ~new_new_n13720__;
  assign new_new_n13722__ = new_new_n13717__ & new_new_n13721__;
  assign new_new_n13723__ = ~new_new_n13717__ & ~new_new_n13721__;
  assign new_new_n13724__ = ~new_new_n6484__ & ~new_new_n13713__;
  assign new_new_n13725__ = pi01 & new_new_n1902__;
  assign new_new_n13726__ = ~new_new_n13692__ & ~new_new_n13725__;
  assign new_new_n13727__ = new_new_n6484__ & new_new_n13726__;
  assign new_new_n13728__ = pi00 & ~new_new_n13724__;
  assign new_new_n13729__ = ~new_new_n13727__ & new_new_n13728__;
  assign new_new_n13730__ = pi01 & ~new_new_n1823__;
  assign new_new_n13731__ = pi02 & new_new_n13730__;
  assign new_new_n13732__ = ~pi01 & ~new_new_n3535__;
  assign new_new_n13733__ = pi02 & ~new_new_n13732__;
  assign new_new_n13734__ = ~new_new_n13730__ & ~new_new_n13733__;
  assign new_new_n13735__ = ~pi00 & ~new_new_n13731__;
  assign new_new_n13736__ = ~new_new_n13734__ & new_new_n13735__;
  assign new_new_n13737__ = ~new_new_n13298__ & ~new_new_n13299__;
  assign new_new_n13738__ = ~new_new_n13303__ & new_new_n13737__;
  assign new_new_n13739__ = new_new_n13303__ & ~new_new_n13737__;
  assign new_new_n13740__ = ~new_new_n13738__ & ~new_new_n13739__;
  assign new_new_n13741__ = pi02 & ~new_new_n5501__;
  assign new_new_n13742__ = pi01 & new_new_n5501__;
  assign new_new_n13743__ = ~new_new_n13741__ & ~new_new_n13742__;
  assign new_new_n13744__ = ~new_new_n1823__ & new_new_n13743__;
  assign new_new_n13745__ = new_new_n1823__ & ~new_new_n13743__;
  assign new_new_n13746__ = pi00 & ~new_new_n13744__;
  assign new_new_n13747__ = ~new_new_n13745__ & new_new_n13746__;
  assign new_new_n13748__ = ~new_new_n3535__ & new_new_n13508__;
  assign new_new_n13749__ = pi01 & ~new_new_n3535__;
  assign new_new_n13750__ = ~pi01 & ~new_new_n2130__;
  assign new_new_n13751__ = pi02 & ~new_new_n13749__;
  assign new_new_n13752__ = ~new_new_n13750__ & new_new_n13751__;
  assign new_new_n13753__ = ~pi00 & ~new_new_n13748__;
  assign new_new_n13754__ = ~new_new_n13752__ & new_new_n13753__;
  assign new_new_n13755__ = ~new_new_n13747__ & ~new_new_n13754__;
  assign new_new_n13756__ = ~new_new_n13284__ & ~new_new_n13285__;
  assign new_new_n13757__ = ~new_new_n13295__ & new_new_n13756__;
  assign new_new_n13758__ = new_new_n13295__ & ~new_new_n13756__;
  assign new_new_n13759__ = ~new_new_n13757__ & ~new_new_n13758__;
  assign new_new_n13760__ = ~new_new_n13755__ & new_new_n13759__;
  assign new_new_n13761__ = new_new_n13755__ & ~new_new_n13759__;
  assign new_new_n13762__ = new_new_n12488__ & ~new_new_n12983__;
  assign new_new_n13763__ = ~new_new_n12488__ & new_new_n12983__;
  assign new_new_n13764__ = ~new_new_n13762__ & ~new_new_n13763__;
  assign new_new_n13765__ = pi05 & ~new_new_n12493__;
  assign new_new_n13766__ = ~pi05 & new_new_n12493__;
  assign new_new_n13767__ = ~new_new_n13765__ & ~new_new_n13766__;
  assign new_new_n13768__ = new_new_n12509__ & new_new_n13767__;
  assign new_new_n13769__ = ~new_new_n12509__ & ~new_new_n13767__;
  assign new_new_n13770__ = ~new_new_n13768__ & ~new_new_n13769__;
  assign new_new_n13771__ = new_new_n13275__ & ~new_new_n13770__;
  assign new_new_n13772__ = ~new_new_n13275__ & new_new_n13770__;
  assign new_new_n13773__ = ~new_new_n13771__ & ~new_new_n13772__;
  assign new_new_n13774__ = new_new_n13764__ & new_new_n13773__;
  assign new_new_n13775__ = ~new_new_n13764__ & ~new_new_n13773__;
  assign new_new_n13776__ = pi01 & new_new_n2130__;
  assign new_new_n13777__ = ~pi01 & new_new_n2024__;
  assign new_new_n13778__ = ~new_new_n13776__ & ~new_new_n13777__;
  assign new_new_n13779__ = pi02 & ~new_new_n13778__;
  assign new_new_n13780__ = ~new_new_n2130__ & new_new_n13508__;
  assign new_new_n13781__ = ~new_new_n13779__ & ~new_new_n13780__;
  assign new_new_n13782__ = ~pi00 & ~new_new_n13781__;
  assign new_new_n13783__ = pi02 & ~new_new_n5500__;
  assign new_new_n13784__ = pi01 & new_new_n6852__;
  assign new_new_n13785__ = ~new_new_n13783__ & ~new_new_n13784__;
  assign new_new_n13786__ = ~new_new_n3535__ & ~new_new_n13785__;
  assign new_new_n13787__ = ~new_new_n5498__ & ~new_new_n5501__;
  assign new_new_n13788__ = pi01 & new_new_n13787__;
  assign new_new_n13789__ = pi02 & ~new_new_n13787__;
  assign new_new_n13790__ = new_new_n3535__ & ~new_new_n13788__;
  assign new_new_n13791__ = ~new_new_n13789__ & new_new_n13790__;
  assign new_new_n13792__ = pi00 & ~new_new_n13786__;
  assign new_new_n13793__ = ~new_new_n13791__ & new_new_n13792__;
  assign new_new_n13794__ = ~new_new_n13782__ & ~new_new_n13793__;
  assign new_new_n13795__ = ~pi02 & ~new_new_n2130__;
  assign new_new_n13796__ = ~new_new_n13776__ & ~new_new_n13795__;
  assign new_new_n13797__ = ~new_new_n6036__ & ~new_new_n13796__;
  assign new_new_n13798__ = pi02 & new_new_n2130__;
  assign new_new_n13799__ = ~new_new_n13750__ & ~new_new_n13798__;
  assign new_new_n13800__ = new_new_n6036__ & ~new_new_n13799__;
  assign new_new_n13801__ = pi00 & ~new_new_n13797__;
  assign new_new_n13802__ = ~new_new_n13800__ & new_new_n13801__;
  assign new_new_n13803__ = ~new_new_n2024__ & new_new_n13508__;
  assign new_new_n13804__ = ~pi01 & ~new_new_n2224__;
  assign new_new_n13805__ = pi01 & ~new_new_n2024__;
  assign new_new_n13806__ = pi02 & ~new_new_n13804__;
  assign new_new_n13807__ = ~new_new_n13805__ & new_new_n13806__;
  assign new_new_n13808__ = ~pi00 & ~new_new_n13803__;
  assign new_new_n13809__ = ~new_new_n13807__ & new_new_n13808__;
  assign new_new_n13810__ = ~new_new_n13802__ & ~new_new_n13809__;
  assign new_new_n13811__ = ~new_new_n13268__ & ~new_new_n13269__;
  assign new_new_n13812__ = new_new_n13273__ & new_new_n13811__;
  assign new_new_n13813__ = ~new_new_n13273__ & ~new_new_n13811__;
  assign new_new_n13814__ = ~new_new_n13812__ & ~new_new_n13813__;
  assign new_new_n13815__ = ~new_new_n13810__ & ~new_new_n13814__;
  assign new_new_n13816__ = new_new_n13810__ & new_new_n13814__;
  assign new_new_n13817__ = ~new_new_n2420__ & new_new_n13508__;
  assign new_new_n13818__ = pi01 & new_new_n2420__;
  assign new_new_n13819__ = ~pi01 & new_new_n2313__;
  assign new_new_n13820__ = ~new_new_n13818__ & ~new_new_n13819__;
  assign new_new_n13821__ = pi02 & ~new_new_n13820__;
  assign new_new_n13822__ = ~new_new_n13817__ & ~new_new_n13821__;
  assign new_new_n13823__ = ~pi00 & ~new_new_n13822__;
  assign new_new_n13824__ = ~pi02 & ~new_new_n2224__;
  assign new_new_n13825__ = ~new_new_n3476__ & ~new_new_n6512__;
  assign new_new_n13826__ = pi02 & new_new_n2224__;
  assign new_new_n13827__ = ~new_new_n13824__ & ~new_new_n13826__;
  assign new_new_n13828__ = ~new_new_n13825__ & new_new_n13827__;
  assign new_new_n13829__ = pi01 & new_new_n2224__;
  assign new_new_n13830__ = ~new_new_n13804__ & ~new_new_n13829__;
  assign new_new_n13831__ = new_new_n13825__ & new_new_n13830__;
  assign new_new_n13832__ = pi00 & ~new_new_n13828__;
  assign new_new_n13833__ = ~new_new_n13831__ & new_new_n13832__;
  assign new_new_n13834__ = ~new_new_n13823__ & ~new_new_n13833__;
  assign new_new_n13835__ = ~new_new_n13242__ & ~new_new_n13243__;
  assign new_new_n13836__ = ~new_new_n13247__ & new_new_n13835__;
  assign new_new_n13837__ = new_new_n13247__ & ~new_new_n13835__;
  assign new_new_n13838__ = ~new_new_n13836__ & ~new_new_n13837__;
  assign new_new_n13839__ = ~new_new_n13834__ & new_new_n13838__;
  assign new_new_n13840__ = new_new_n13834__ & ~new_new_n13838__;
  assign new_new_n13841__ = ~new_new_n13032__ & ~new_new_n13033__;
  assign new_new_n13842__ = new_new_n13239__ & new_new_n13841__;
  assign new_new_n13843__ = ~new_new_n13239__ & ~new_new_n13841__;
  assign new_new_n13844__ = ~new_new_n2313__ & new_new_n13508__;
  assign new_new_n13845__ = ~pi01 & ~new_new_n2572__;
  assign new_new_n13846__ = pi01 & ~new_new_n2313__;
  assign new_new_n13847__ = pi02 & ~new_new_n13845__;
  assign new_new_n13848__ = ~new_new_n13846__ & new_new_n13847__;
  assign new_new_n13849__ = ~pi00 & ~new_new_n13844__;
  assign new_new_n13850__ = ~new_new_n13848__ & new_new_n13849__;
  assign new_new_n13851__ = pi02 & ~new_new_n6748__;
  assign new_new_n13852__ = pi01 & new_new_n6748__;
  assign new_new_n13853__ = ~new_new_n13851__ & ~new_new_n13852__;
  assign new_new_n13854__ = new_new_n2420__ & ~new_new_n13853__;
  assign new_new_n13855__ = ~new_new_n2420__ & new_new_n13853__;
  assign new_new_n13856__ = pi00 & ~new_new_n13854__;
  assign new_new_n13857__ = ~new_new_n13855__ & new_new_n13856__;
  assign new_new_n13858__ = ~new_new_n13850__ & ~new_new_n13857__;
  assign new_new_n13859__ = ~new_new_n2572__ & new_new_n13508__;
  assign new_new_n13860__ = ~pi01 & new_new_n2497__;
  assign new_new_n13861__ = pi01 & new_new_n2572__;
  assign new_new_n13862__ = ~new_new_n13860__ & ~new_new_n13861__;
  assign new_new_n13863__ = pi02 & ~new_new_n13862__;
  assign new_new_n13864__ = ~pi00 & ~new_new_n13859__;
  assign new_new_n13865__ = ~new_new_n13863__ & new_new_n13864__;
  assign new_new_n13866__ = pi02 & ~new_new_n2313__;
  assign new_new_n13867__ = ~new_new_n13819__ & ~new_new_n13866__;
  assign new_new_n13868__ = ~new_new_n7236__ & new_new_n13867__;
  assign new_new_n13869__ = ~pi02 & new_new_n2313__;
  assign new_new_n13870__ = ~new_new_n13846__ & ~new_new_n13869__;
  assign new_new_n13871__ = new_new_n7236__ & new_new_n13870__;
  assign new_new_n13872__ = pi00 & ~new_new_n13868__;
  assign new_new_n13873__ = ~new_new_n13871__ & new_new_n13872__;
  assign new_new_n13874__ = ~new_new_n13865__ & ~new_new_n13873__;
  assign new_new_n13875__ = pi01 & ~new_new_n2497__;
  assign new_new_n13876__ = ~new_new_n2636__ & new_new_n12798__;
  assign new_new_n13877__ = ~new_new_n13875__ & ~new_new_n13876__;
  assign new_new_n13878__ = ~pi00 & ~new_new_n13877__;
  assign new_new_n13879__ = pi00 & new_new_n10874__;
  assign new_new_n13880__ = ~new_new_n13878__ & ~new_new_n13879__;
  assign new_new_n13881__ = ~pi02 & ~new_new_n13880__;
  assign new_new_n13882__ = pi00 & ~new_new_n6802__;
  assign new_new_n13883__ = pi02 & ~new_new_n13878__;
  assign new_new_n13884__ = ~new_new_n13882__ & new_new_n13883__;
  assign new_new_n13885__ = ~new_new_n13845__ & ~new_new_n13861__;
  assign new_new_n13886__ = pi00 & ~new_new_n13885__;
  assign new_new_n13887__ = new_new_n6801__ & new_new_n13886__;
  assign new_new_n13888__ = ~new_new_n13884__ & ~new_new_n13887__;
  assign new_new_n13889__ = ~new_new_n13881__ & new_new_n13888__;
  assign new_new_n13890__ = ~new_new_n13205__ & ~new_new_n13206__;
  assign new_new_n13891__ = ~new_new_n13217__ & new_new_n13890__;
  assign new_new_n13892__ = new_new_n13217__ & ~new_new_n13890__;
  assign new_new_n13893__ = ~new_new_n13891__ & ~new_new_n13892__;
  assign new_new_n13894__ = new_new_n13889__ & ~new_new_n13893__;
  assign new_new_n13895__ = ~new_new_n13889__ & new_new_n13893__;
  assign new_new_n13896__ = pi00 & new_new_n9126__;
  assign new_new_n13897__ = pi01 & ~new_new_n2636__;
  assign new_new_n13898__ = ~new_new_n2737__ & new_new_n12798__;
  assign new_new_n13899__ = ~pi00 & ~new_new_n13897__;
  assign new_new_n13900__ = ~new_new_n13898__ & new_new_n13899__;
  assign new_new_n13901__ = ~new_new_n13896__ & ~new_new_n13900__;
  assign new_new_n13902__ = ~pi02 & ~new_new_n13901__;
  assign new_new_n13903__ = pi00 & ~new_new_n7772__;
  assign new_new_n13904__ = pi02 & ~new_new_n13900__;
  assign new_new_n13905__ = ~new_new_n13903__ & new_new_n13904__;
  assign new_new_n13906__ = ~new_new_n13860__ & ~new_new_n13875__;
  assign new_new_n13907__ = pi00 & ~new_new_n13906__;
  assign new_new_n13908__ = ~new_new_n6797__ & new_new_n13907__;
  assign new_new_n13909__ = ~new_new_n13905__ & ~new_new_n13908__;
  assign new_new_n13910__ = ~new_new_n13902__ & new_new_n13909__;
  assign new_new_n13911__ = ~new_new_n13190__ & ~new_new_n13191__;
  assign new_new_n13912__ = ~new_new_n13202__ & new_new_n13911__;
  assign new_new_n13913__ = new_new_n13202__ & ~new_new_n13911__;
  assign new_new_n13914__ = ~new_new_n13912__ & ~new_new_n13913__;
  assign new_new_n13915__ = ~new_new_n13910__ & ~new_new_n13914__;
  assign new_new_n13916__ = new_new_n13910__ & new_new_n13914__;
  assign new_new_n13917__ = pi01 & new_new_n2737__;
  assign new_new_n13918__ = ~pi01 & new_new_n2886__;
  assign new_new_n13919__ = ~new_new_n13917__ & ~new_new_n13918__;
  assign new_new_n13920__ = pi02 & ~new_new_n13919__;
  assign new_new_n13921__ = ~pi02 & ~new_new_n2737__;
  assign new_new_n13922__ = pi01 & new_new_n13921__;
  assign new_new_n13923__ = ~new_new_n13920__ & ~new_new_n13922__;
  assign new_new_n13924__ = ~pi00 & ~new_new_n13923__;
  assign new_new_n13925__ = ~pi01 & new_new_n2636__;
  assign new_new_n13926__ = ~new_new_n13897__ & ~new_new_n13925__;
  assign new_new_n13927__ = new_new_n7811__ & ~new_new_n13926__;
  assign new_new_n13928__ = ~pi02 & ~new_new_n2636__;
  assign new_new_n13929__ = pi02 & new_new_n2636__;
  assign new_new_n13930__ = ~new_new_n13928__ & ~new_new_n13929__;
  assign new_new_n13931__ = ~new_new_n7811__ & new_new_n13930__;
  assign new_new_n13932__ = pi00 & ~new_new_n13927__;
  assign new_new_n13933__ = ~new_new_n13931__ & new_new_n13932__;
  assign new_new_n13934__ = ~new_new_n13924__ & ~new_new_n13933__;
  assign new_new_n13935__ = ~new_new_n13917__ & ~new_new_n13921__;
  assign new_new_n13936__ = ~new_new_n7378__ & ~new_new_n13935__;
  assign new_new_n13937__ = ~pi02 & new_new_n2737__;
  assign new_new_n13938__ = pi01 & ~new_new_n2737__;
  assign new_new_n13939__ = ~new_new_n13937__ & ~new_new_n13938__;
  assign new_new_n13940__ = new_new_n7378__ & new_new_n13939__;
  assign new_new_n13941__ = pi00 & ~new_new_n13936__;
  assign new_new_n13942__ = ~new_new_n13940__ & new_new_n13941__;
  assign new_new_n13943__ = ~new_new_n2886__ & new_new_n13508__;
  assign new_new_n13944__ = pi01 & ~new_new_n2886__;
  assign new_new_n13945__ = ~pi01 & ~new_new_n2848__;
  assign new_new_n13946__ = pi02 & ~new_new_n13944__;
  assign new_new_n13947__ = ~new_new_n13945__ & new_new_n13946__;
  assign new_new_n13948__ = ~pi00 & ~new_new_n13943__;
  assign new_new_n13949__ = ~new_new_n13947__ & new_new_n13948__;
  assign new_new_n13950__ = ~new_new_n13942__ & ~new_new_n13949__;
  assign new_new_n13951__ = ~pi02 & ~new_new_n2848__;
  assign new_new_n13952__ = pi01 & new_new_n13951__;
  assign new_new_n13953__ = ~pi01 & ~new_new_n3460__;
  assign new_new_n13954__ = pi01 & ~new_new_n2848__;
  assign new_new_n13955__ = pi02 & ~new_new_n13953__;
  assign new_new_n13956__ = ~new_new_n13954__ & new_new_n13955__;
  assign new_new_n13957__ = ~pi00 & ~new_new_n13952__;
  assign new_new_n13958__ = ~new_new_n13956__ & new_new_n13957__;
  assign new_new_n13959__ = pi02 & ~new_new_n2886__;
  assign new_new_n13960__ = ~new_new_n13918__ & ~new_new_n13959__;
  assign new_new_n13961__ = ~new_new_n8574__ & new_new_n13960__;
  assign new_new_n13962__ = ~pi02 & new_new_n2886__;
  assign new_new_n13963__ = ~new_new_n13944__ & ~new_new_n13962__;
  assign new_new_n13964__ = new_new_n8574__ & new_new_n13963__;
  assign new_new_n13965__ = pi00 & ~new_new_n13961__;
  assign new_new_n13966__ = ~new_new_n13964__ & new_new_n13965__;
  assign new_new_n13967__ = ~new_new_n13958__ & ~new_new_n13966__;
  assign new_new_n13968__ = new_new_n2960__ & ~new_new_n7055__;
  assign new_new_n13969__ = pi02 & new_new_n2848__;
  assign new_new_n13970__ = ~new_new_n2960__ & ~new_new_n13969__;
  assign new_new_n13971__ = ~new_new_n13968__ & ~new_new_n13970__;
  assign new_new_n13972__ = new_new_n3361__ & new_new_n13971__;
  assign new_new_n13973__ = new_new_n2960__ & new_new_n3460__;
  assign new_new_n13974__ = ~new_new_n3460__ & ~new_new_n13969__;
  assign new_new_n13975__ = ~new_new_n7711__ & ~new_new_n13973__;
  assign new_new_n13976__ = ~new_new_n13974__ & new_new_n13975__;
  assign new_new_n13977__ = ~new_new_n3361__ & new_new_n13976__;
  assign new_new_n13978__ = ~new_new_n13951__ & ~new_new_n13972__;
  assign new_new_n13979__ = ~new_new_n13977__ & new_new_n13978__;
  assign new_new_n13980__ = pi00 & ~new_new_n13979__;
  assign new_new_n13981__ = pi00 & ~new_new_n7711__;
  assign new_new_n13982__ = pi02 & new_new_n2960__;
  assign new_new_n13983__ = ~new_new_n13981__ & new_new_n13982__;
  assign new_new_n13984__ = ~new_new_n13980__ & ~new_new_n13983__;
  assign new_new_n13985__ = ~pi01 & ~new_new_n13984__;
  assign new_new_n13986__ = ~pi00 & pi02;
  assign new_new_n13987__ = new_new_n3460__ & new_new_n13986__;
  assign new_new_n13988__ = ~new_new_n2848__ & ~new_new_n2960__;
  assign new_new_n13989__ = pi00 & ~new_new_n13988__;
  assign new_new_n13990__ = ~pi02 & ~new_new_n3460__;
  assign new_new_n13991__ = ~new_new_n13989__ & new_new_n13990__;
  assign new_new_n13992__ = pi02 & ~new_new_n3361__;
  assign new_new_n13993__ = new_new_n2960__ & ~new_new_n7711__;
  assign new_new_n13994__ = ~new_new_n13992__ & new_new_n13993__;
  assign new_new_n13995__ = new_new_n7058__ & new_new_n13994__;
  assign new_new_n13996__ = new_new_n3361__ & new_new_n13951__;
  assign new_new_n13997__ = ~new_new_n8567__ & ~new_new_n13996__;
  assign new_new_n13998__ = new_new_n3460__ & ~new_new_n13997__;
  assign new_new_n13999__ = ~new_new_n13969__ & ~new_new_n13995__;
  assign new_new_n14000__ = ~new_new_n13998__ & new_new_n13999__;
  assign new_new_n14001__ = pi00 & ~new_new_n14000__;
  assign new_new_n14002__ = ~new_new_n13987__ & ~new_new_n13991__;
  assign new_new_n14003__ = ~new_new_n14001__ & new_new_n14002__;
  assign new_new_n14004__ = pi01 & ~new_new_n14003__;
  assign new_new_n14005__ = ~new_new_n13985__ & ~new_new_n14004__;
  assign new_new_n14006__ = ~new_new_n13109__ & ~new_new_n13110__;
  assign new_new_n14007__ = new_new_n13122__ & new_new_n14006__;
  assign new_new_n14008__ = ~new_new_n13122__ & ~new_new_n14006__;
  assign new_new_n14009__ = ~new_new_n14007__ & ~new_new_n14008__;
  assign new_new_n14010__ = new_new_n14005__ & ~new_new_n14009__;
  assign new_new_n14011__ = ~new_new_n14005__ & new_new_n14009__;
  assign new_new_n14012__ = pi00 & new_new_n13953__;
  assign new_new_n14013__ = ~pi00 & ~new_new_n2960__;
  assign new_new_n14014__ = ~new_new_n2960__ & ~new_new_n3460__;
  assign new_new_n14015__ = pi00 & new_new_n2960__;
  assign new_new_n14016__ = new_new_n3460__ & new_new_n14015__;
  assign new_new_n14017__ = ~new_new_n14014__ & ~new_new_n14016__;
  assign new_new_n14018__ = ~new_new_n3361__ & ~new_new_n14017__;
  assign new_new_n14019__ = ~new_new_n14013__ & ~new_new_n14018__;
  assign new_new_n14020__ = pi01 & ~new_new_n14019__;
  assign new_new_n14021__ = pi01 & new_new_n3460__;
  assign new_new_n14022__ = ~new_new_n14015__ & ~new_new_n14021__;
  assign new_new_n14023__ = ~new_new_n13973__ & ~new_new_n14022__;
  assign new_new_n14024__ = new_new_n3361__ & new_new_n14023__;
  assign new_new_n14025__ = ~new_new_n14012__ & ~new_new_n14024__;
  assign new_new_n14026__ = ~new_new_n14020__ & new_new_n14025__;
  assign new_new_n14027__ = ~pi02 & ~new_new_n14026__;
  assign new_new_n14028__ = pi01 & new_new_n2960__;
  assign new_new_n14029__ = ~new_new_n13973__ & ~new_new_n14014__;
  assign new_new_n14030__ = ~new_new_n14028__ & new_new_n14029__;
  assign new_new_n14031__ = ~new_new_n3361__ & new_new_n14030__;
  assign new_new_n14032__ = ~new_new_n14021__ & ~new_new_n14031__;
  assign new_new_n14033__ = pi00 & ~new_new_n14032__;
  assign new_new_n14034__ = ~pi01 & new_new_n14014__;
  assign new_new_n14035__ = ~new_new_n14016__ & ~new_new_n14034__;
  assign new_new_n14036__ = new_new_n3361__ & ~new_new_n14035__;
  assign new_new_n14037__ = ~pi01 & new_new_n3126__;
  assign new_new_n14038__ = ~new_new_n14028__ & ~new_new_n14037__;
  assign new_new_n14039__ = ~pi00 & ~new_new_n14038__;
  assign new_new_n14040__ = ~new_new_n14036__ & ~new_new_n14039__;
  assign new_new_n14041__ = ~new_new_n14033__ & new_new_n14040__;
  assign new_new_n14042__ = pi02 & ~new_new_n14041__;
  assign new_new_n14043__ = ~new_new_n14027__ & ~new_new_n14042__;
  assign new_new_n14044__ = ~pi01 & new_new_n3164__;
  assign new_new_n14045__ = pi01 & new_new_n3126__;
  assign new_new_n14046__ = ~new_new_n14044__ & ~new_new_n14045__;
  assign new_new_n14047__ = pi02 & ~new_new_n14046__;
  assign new_new_n14048__ = ~new_new_n3126__ & new_new_n13508__;
  assign new_new_n14049__ = ~new_new_n14047__ & ~new_new_n14048__;
  assign new_new_n14050__ = ~pi00 & ~new_new_n14049__;
  assign new_new_n14051__ = ~pi01 & ~new_new_n7468__;
  assign new_new_n14052__ = ~pi02 & new_new_n7468__;
  assign new_new_n14053__ = new_new_n2960__ & ~new_new_n14051__;
  assign new_new_n14054__ = ~new_new_n14052__ & new_new_n14053__;
  assign new_new_n14055__ = pi01 & new_new_n7468__;
  assign new_new_n14056__ = pi02 & ~new_new_n7468__;
  assign new_new_n14057__ = ~new_new_n2960__ & ~new_new_n14055__;
  assign new_new_n14058__ = ~new_new_n14056__ & new_new_n14057__;
  assign new_new_n14059__ = ~new_new_n14054__ & ~new_new_n14058__;
  assign new_new_n14060__ = pi00 & ~new_new_n14059__;
  assign new_new_n14061__ = ~new_new_n14050__ & ~new_new_n14060__;
  assign new_new_n14062__ = pi01 & ~new_new_n3164__;
  assign new_new_n14063__ = ~pi01 & ~new_new_n3254__;
  assign new_new_n14064__ = pi02 & ~new_new_n14062__;
  assign new_new_n14065__ = ~new_new_n14063__ & new_new_n14064__;
  assign new_new_n14066__ = ~new_new_n3164__ & new_new_n13508__;
  assign new_new_n14067__ = ~new_new_n14065__ & ~new_new_n14066__;
  assign new_new_n14068__ = ~pi00 & ~new_new_n14067__;
  assign new_new_n14069__ = ~pi01 & ~new_new_n7570__;
  assign new_new_n14070__ = ~pi02 & new_new_n7570__;
  assign new_new_n14071__ = new_new_n3126__ & ~new_new_n14069__;
  assign new_new_n14072__ = ~new_new_n14070__ & new_new_n14071__;
  assign new_new_n14073__ = pi01 & new_new_n7570__;
  assign new_new_n14074__ = pi02 & ~new_new_n7570__;
  assign new_new_n14075__ = ~new_new_n3126__ & ~new_new_n14073__;
  assign new_new_n14076__ = ~new_new_n14074__ & new_new_n14075__;
  assign new_new_n14077__ = ~new_new_n14072__ & ~new_new_n14076__;
  assign new_new_n14078__ = pi00 & ~new_new_n14077__;
  assign new_new_n14079__ = ~new_new_n14068__ & ~new_new_n14078__;
  assign new_new_n14080__ = pi00 & ~new_new_n7682__;
  assign new_new_n14081__ = pi01 & ~new_new_n3254__;
  assign new_new_n14082__ = pi03 & ~new_new_n3356__;
  assign new_new_n14083__ = pi02 & new_new_n3055__;
  assign new_new_n14084__ = ~new_new_n14081__ & new_new_n14083__;
  assign new_new_n14085__ = ~new_new_n14082__ & new_new_n14084__;
  assign new_new_n14086__ = ~new_new_n14080__ & new_new_n14085__;
  assign new_new_n14087__ = ~new_new_n14079__ & new_new_n14086__;
  assign new_new_n14088__ = pi00 & new_new_n11469__;
  assign new_new_n14089__ = ~new_new_n3254__ & ~new_new_n11480__;
  assign new_new_n14090__ = new_new_n3254__ & ~new_new_n11481__;
  assign new_new_n14091__ = pi01 & ~new_new_n14089__;
  assign new_new_n14092__ = ~new_new_n14090__ & new_new_n14091__;
  assign new_new_n14093__ = ~new_new_n14088__ & ~new_new_n14092__;
  assign new_new_n14094__ = ~new_new_n3055__ & ~new_new_n10726__;
  assign new_new_n14095__ = new_new_n11473__ & ~new_new_n14094__;
  assign new_new_n14096__ = ~new_new_n3356__ & new_new_n14094__;
  assign new_new_n14097__ = ~new_new_n10731__ & ~new_new_n14096__;
  assign new_new_n14098__ = pi04 & ~new_new_n14097__;
  assign new_new_n14099__ = ~new_new_n13078__ & ~new_new_n14095__;
  assign new_new_n14100__ = ~new_new_n14098__ & new_new_n14099__;
  assign new_new_n14101__ = new_new_n14079__ & ~new_new_n14100__;
  assign new_new_n14102__ = ~new_new_n3356__ & ~new_new_n14093__;
  assign new_new_n14103__ = ~new_new_n14101__ & new_new_n14102__;
  assign new_new_n14104__ = ~new_new_n14087__ & ~new_new_n14103__;
  assign new_new_n14105__ = pi02 & ~new_new_n3164__;
  assign new_new_n14106__ = ~new_new_n14044__ & ~new_new_n14105__;
  assign new_new_n14107__ = ~new_new_n8637__ & new_new_n14106__;
  assign new_new_n14108__ = ~pi02 & new_new_n3164__;
  assign new_new_n14109__ = ~new_new_n14062__ & ~new_new_n14108__;
  assign new_new_n14110__ = new_new_n8637__ & new_new_n14109__;
  assign new_new_n14111__ = pi00 & ~new_new_n14107__;
  assign new_new_n14112__ = ~new_new_n14110__ & new_new_n14111__;
  assign new_new_n14113__ = ~new_new_n14104__ & ~new_new_n14112__;
  assign new_new_n14114__ = new_new_n14079__ & ~new_new_n14086__;
  assign new_new_n14115__ = new_new_n14100__ & ~new_new_n14114__;
  assign new_new_n14116__ = ~new_new_n14113__ & ~new_new_n14115__;
  assign new_new_n14117__ = pi05 & ~new_new_n11470__;
  assign new_new_n14118__ = ~new_new_n13078__ & new_new_n14117__;
  assign new_new_n14119__ = ~new_new_n13092__ & ~new_new_n14118__;
  assign new_new_n14120__ = ~new_new_n9017__ & new_new_n14117__;
  assign new_new_n14121__ = new_new_n13092__ & new_new_n14120__;
  assign new_new_n14122__ = ~new_new_n14119__ & ~new_new_n14121__;
  assign new_new_n14123__ = new_new_n14116__ & new_new_n14122__;
  assign new_new_n14124__ = ~new_new_n14061__ & ~new_new_n14123__;
  assign new_new_n14125__ = ~new_new_n14116__ & ~new_new_n14122__;
  assign new_new_n14126__ = ~new_new_n14124__ & ~new_new_n14125__;
  assign new_new_n14127__ = new_new_n14043__ & new_new_n14126__;
  assign new_new_n14128__ = ~new_new_n14043__ & ~new_new_n14126__;
  assign new_new_n14129__ = pi06 & new_new_n13094__;
  assign new_new_n14130__ = pi05 & ~new_new_n13094__;
  assign new_new_n14131__ = new_new_n3356__ & ~new_new_n14130__;
  assign new_new_n14132__ = ~new_new_n14129__ & ~new_new_n14131__;
  assign new_new_n14133__ = new_new_n13076__ & ~new_new_n14132__;
  assign new_new_n14134__ = new_new_n3356__ & ~new_new_n13076__;
  assign new_new_n14135__ = new_new_n14130__ & new_new_n14134__;
  assign new_new_n14136__ = ~pi06 & new_new_n13076__;
  assign new_new_n14137__ = ~new_new_n13096__ & ~new_new_n14136__;
  assign new_new_n14138__ = ~new_new_n3356__ & ~new_new_n13095__;
  assign new_new_n14139__ = ~new_new_n14137__ & new_new_n14138__;
  assign new_new_n14140__ = ~new_new_n14135__ & ~new_new_n14139__;
  assign new_new_n14141__ = ~new_new_n14133__ & new_new_n14140__;
  assign new_new_n14142__ = ~new_new_n14128__ & ~new_new_n14141__;
  assign new_new_n14143__ = ~new_new_n14127__ & ~new_new_n14142__;
  assign new_new_n14144__ = ~new_new_n14011__ & ~new_new_n14143__;
  assign new_new_n14145__ = ~new_new_n14010__ & ~new_new_n14144__;
  assign new_new_n14146__ = new_new_n13967__ & new_new_n14145__;
  assign new_new_n14147__ = ~new_new_n13967__ & ~new_new_n14145__;
  assign new_new_n14148__ = ~new_new_n13125__ & ~new_new_n13126__;
  assign new_new_n14149__ = new_new_n13138__ & ~new_new_n14148__;
  assign new_new_n14150__ = ~new_new_n13138__ & new_new_n14148__;
  assign new_new_n14151__ = ~new_new_n14149__ & ~new_new_n14150__;
  assign new_new_n14152__ = ~new_new_n14147__ & ~new_new_n14151__;
  assign new_new_n14153__ = ~new_new_n14146__ & ~new_new_n14152__;
  assign new_new_n14154__ = new_new_n13950__ & ~new_new_n14153__;
  assign new_new_n14155__ = ~new_new_n13950__ & new_new_n14153__;
  assign new_new_n14156__ = new_new_n13153__ & ~new_new_n13167__;
  assign new_new_n14157__ = ~new_new_n13168__ & ~new_new_n14156__;
  assign new_new_n14158__ = ~new_new_n14155__ & new_new_n14157__;
  assign new_new_n14159__ = ~new_new_n14154__ & ~new_new_n14158__;
  assign new_new_n14160__ = new_new_n13934__ & new_new_n14159__;
  assign new_new_n14161__ = ~new_new_n13934__ & ~new_new_n14159__;
  assign new_new_n14162__ = ~new_new_n13174__ & ~new_new_n13175__;
  assign new_new_n14163__ = new_new_n13187__ & ~new_new_n14162__;
  assign new_new_n14164__ = ~new_new_n13187__ & new_new_n14162__;
  assign new_new_n14165__ = ~new_new_n14163__ & ~new_new_n14164__;
  assign new_new_n14166__ = ~new_new_n14161__ & new_new_n14165__;
  assign new_new_n14167__ = ~new_new_n14160__ & ~new_new_n14166__;
  assign new_new_n14168__ = ~new_new_n13916__ & ~new_new_n14167__;
  assign new_new_n14169__ = ~new_new_n13915__ & ~new_new_n14168__;
  assign new_new_n14170__ = ~new_new_n13895__ & ~new_new_n14169__;
  assign new_new_n14171__ = ~new_new_n13894__ & ~new_new_n14170__;
  assign new_new_n14172__ = ~new_new_n13874__ & ~new_new_n14171__;
  assign new_new_n14173__ = new_new_n13874__ & new_new_n14171__;
  assign new_new_n14174__ = ~new_new_n13048__ & new_new_n13234__;
  assign new_new_n14175__ = new_new_n13048__ & ~new_new_n13234__;
  assign new_new_n14176__ = ~new_new_n14174__ & ~new_new_n14175__;
  assign new_new_n14177__ = new_new_n13219__ & ~new_new_n14176__;
  assign new_new_n14178__ = ~new_new_n13219__ & new_new_n14176__;
  assign new_new_n14179__ = ~new_new_n14177__ & ~new_new_n14178__;
  assign new_new_n14180__ = new_new_n12353__ & new_new_n14179__;
  assign new_new_n14181__ = ~new_new_n12353__ & ~new_new_n14179__;
  assign new_new_n14182__ = ~new_new_n14180__ & ~new_new_n14181__;
  assign new_new_n14183__ = ~new_new_n14173__ & ~new_new_n14182__;
  assign new_new_n14184__ = ~new_new_n14172__ & ~new_new_n14183__;
  assign new_new_n14185__ = ~new_new_n13858__ & ~new_new_n14184__;
  assign new_new_n14186__ = ~new_new_n13842__ & ~new_new_n13843__;
  assign new_new_n14187__ = ~new_new_n14185__ & new_new_n14186__;
  assign new_new_n14188__ = new_new_n13858__ & new_new_n14184__;
  assign new_new_n14189__ = ~new_new_n14187__ & ~new_new_n14188__;
  assign new_new_n14190__ = ~new_new_n13840__ & ~new_new_n14189__;
  assign new_new_n14191__ = ~new_new_n2224__ & new_new_n13508__;
  assign new_new_n14192__ = ~pi01 & new_new_n2420__;
  assign new_new_n14193__ = ~new_new_n13829__ & ~new_new_n14192__;
  assign new_new_n14194__ = pi02 & ~new_new_n14193__;
  assign new_new_n14195__ = ~pi00 & ~new_new_n14191__;
  assign new_new_n14196__ = ~new_new_n14194__ & new_new_n14195__;
  assign new_new_n14197__ = ~pi02 & new_new_n2024__;
  assign new_new_n14198__ = ~new_new_n13805__ & ~new_new_n14197__;
  assign new_new_n14199__ = ~new_new_n7313__ & new_new_n14198__;
  assign new_new_n14200__ = pi02 & ~new_new_n2024__;
  assign new_new_n14201__ = ~new_new_n13777__ & ~new_new_n14200__;
  assign new_new_n14202__ = new_new_n7313__ & new_new_n14201__;
  assign new_new_n14203__ = pi00 & ~new_new_n14199__;
  assign new_new_n14204__ = ~new_new_n14202__ & new_new_n14203__;
  assign new_new_n14205__ = ~new_new_n14196__ & ~new_new_n14204__;
  assign new_new_n14206__ = ~new_new_n13254__ & ~new_new_n13255__;
  assign new_new_n14207__ = ~new_new_n13265__ & ~new_new_n14206__;
  assign new_new_n14208__ = new_new_n13265__ & new_new_n14206__;
  assign new_new_n14209__ = ~new_new_n14207__ & ~new_new_n14208__;
  assign new_new_n14210__ = new_new_n14205__ & new_new_n14209__;
  assign new_new_n14211__ = ~new_new_n13839__ & ~new_new_n14190__;
  assign new_new_n14212__ = ~new_new_n14210__ & new_new_n14211__;
  assign new_new_n14213__ = ~new_new_n14205__ & ~new_new_n14209__;
  assign new_new_n14214__ = ~new_new_n14212__ & ~new_new_n14213__;
  assign new_new_n14215__ = ~new_new_n13816__ & ~new_new_n14214__;
  assign new_new_n14216__ = ~new_new_n13815__ & ~new_new_n14215__;
  assign new_new_n14217__ = ~new_new_n13794__ & new_new_n14216__;
  assign new_new_n14218__ = ~new_new_n13774__ & ~new_new_n13775__;
  assign new_new_n14219__ = ~new_new_n14217__ & new_new_n14218__;
  assign new_new_n14220__ = new_new_n13794__ & ~new_new_n14216__;
  assign new_new_n14221__ = ~new_new_n14219__ & ~new_new_n14220__;
  assign new_new_n14222__ = ~new_new_n13761__ & ~new_new_n14221__;
  assign new_new_n14223__ = ~new_new_n13760__ & ~new_new_n14222__;
  assign new_new_n14224__ = new_new_n13740__ & new_new_n14223__;
  assign new_new_n14225__ = ~new_new_n13729__ & ~new_new_n13736__;
  assign new_new_n14226__ = ~new_new_n14224__ & new_new_n14225__;
  assign new_new_n14227__ = ~new_new_n13740__ & ~new_new_n14223__;
  assign new_new_n14228__ = ~new_new_n14226__ & ~new_new_n14227__;
  assign new_new_n14229__ = ~new_new_n13723__ & ~new_new_n14228__;
  assign new_new_n14230__ = ~new_new_n13722__ & ~new_new_n14229__;
  assign new_new_n14231__ = new_new_n13698__ & new_new_n14230__;
  assign new_new_n14232__ = ~new_new_n13698__ & ~new_new_n14230__;
  assign new_new_n14233__ = ~new_new_n13329__ & ~new_new_n13330__;
  assign new_new_n14234__ = new_new_n13346__ & ~new_new_n14233__;
  assign new_new_n14235__ = ~new_new_n13346__ & new_new_n14233__;
  assign new_new_n14236__ = ~new_new_n14234__ & ~new_new_n14235__;
  assign new_new_n14237__ = ~new_new_n14232__ & ~new_new_n14236__;
  assign new_new_n14238__ = ~new_new_n14231__ & ~new_new_n14237__;
  assign new_new_n14239__ = ~new_new_n13682__ & ~new_new_n14238__;
  assign new_new_n14240__ = ~new_new_n13667__ & ~new_new_n13668__;
  assign new_new_n14241__ = ~new_new_n14239__ & new_new_n14240__;
  assign new_new_n14242__ = new_new_n13682__ & new_new_n14238__;
  assign new_new_n14243__ = ~new_new_n14241__ & ~new_new_n14242__;
  assign new_new_n14244__ = ~new_new_n13657__ & ~new_new_n14243__;
  assign new_new_n14245__ = ~new_new_n13656__ & ~new_new_n14244__;
  assign new_new_n14246__ = new_new_n13632__ & ~new_new_n14245__;
  assign new_new_n14247__ = ~new_new_n13617__ & ~new_new_n13625__;
  assign new_new_n14248__ = ~new_new_n14246__ & new_new_n14247__;
  assign new_new_n14249__ = ~new_new_n13632__ & new_new_n14245__;
  assign new_new_n14250__ = ~new_new_n14248__ & ~new_new_n14249__;
  assign new_new_n14251__ = ~new_new_n13610__ & ~new_new_n14250__;
  assign new_new_n14252__ = ~new_new_n13609__ & ~new_new_n14251__;
  assign new_new_n14253__ = new_new_n13589__ & new_new_n14252__;
  assign new_new_n14254__ = ~new_new_n13589__ & ~new_new_n14252__;
  assign new_new_n14255__ = ~new_new_n13396__ & ~new_new_n13397__;
  assign new_new_n14256__ = new_new_n13410__ & ~new_new_n14255__;
  assign new_new_n14257__ = ~new_new_n13410__ & new_new_n14255__;
  assign new_new_n14258__ = ~new_new_n14256__ & ~new_new_n14257__;
  assign new_new_n14259__ = ~new_new_n14254__ & ~new_new_n14258__;
  assign new_new_n14260__ = ~new_new_n14253__ & ~new_new_n14259__;
  assign new_new_n14261__ = ~new_new_n13571__ & ~new_new_n14260__;
  assign new_new_n14262__ = new_new_n13554__ & ~new_new_n14261__;
  assign new_new_n14263__ = ~new_new_n13413__ & new_new_n13427__;
  assign new_new_n14264__ = ~new_new_n14262__ & ~new_new_n14263__;
  assign new_new_n14265__ = new_new_n13571__ & new_new_n14260__;
  assign new_new_n14266__ = ~new_new_n13413__ & ~new_new_n13414__;
  assign new_new_n14267__ = ~new_new_n13426__ & ~new_new_n14266__;
  assign new_new_n14268__ = new_new_n13554__ & ~new_new_n14267__;
  assign new_new_n14269__ = ~new_new_n14265__ & ~new_new_n14268__;
  assign new_new_n14270__ = ~new_new_n14264__ & ~new_new_n14269__;
  assign new_new_n14271__ = ~new_new_n12913__ & ~new_new_n12914__;
  assign new_new_n14272__ = ~new_new_n13413__ & new_new_n14271__;
  assign new_new_n14273__ = new_new_n13413__ & ~new_new_n14271__;
  assign new_new_n14274__ = ~new_new_n14272__ & ~new_new_n14273__;
  assign new_new_n14275__ = ~new_new_n14270__ & new_new_n14274__;
  assign new_new_n14276__ = ~new_new_n14261__ & ~new_new_n14267__;
  assign new_new_n14277__ = ~new_new_n13554__ & ~new_new_n14265__;
  assign new_new_n14278__ = ~new_new_n14276__ & new_new_n14277__;
  assign new_new_n14279__ = new_new_n13554__ & new_new_n14265__;
  assign new_new_n14280__ = new_new_n14263__ & new_new_n14271__;
  assign new_new_n14281__ = ~new_new_n14279__ & new_new_n14280__;
  assign new_new_n14282__ = ~new_new_n14278__ & ~new_new_n14281__;
  assign new_new_n14283__ = ~new_new_n14275__ & new_new_n14282__;
  assign new_new_n14284__ = ~new_new_n13431__ & ~new_new_n13432__;
  assign new_new_n14285__ = new_new_n13442__ & new_new_n14284__;
  assign new_new_n14286__ = ~new_new_n13442__ & ~new_new_n14284__;
  assign new_new_n14287__ = ~new_new_n14285__ & ~new_new_n14286__;
  assign new_new_n14288__ = ~new_new_n14283__ & ~new_new_n14287__;
  assign new_new_n14289__ = new_new_n14283__ & new_new_n14287__;
  assign new_new_n14290__ = ~pi02 & new_new_n4032__;
  assign new_new_n14291__ = ~pi01 & ~new_new_n4032__;
  assign new_new_n14292__ = ~new_new_n14290__ & ~new_new_n14291__;
  assign new_new_n14293__ = ~new_new_n3720__ & ~new_new_n14292__;
  assign new_new_n14294__ = new_new_n3720__ & new_new_n14292__;
  assign new_new_n14295__ = pi00 & ~new_new_n14293__;
  assign new_new_n14296__ = ~new_new_n14294__ & new_new_n14295__;
  assign new_new_n14297__ = ~new_new_n13539__ & ~new_new_n13562__;
  assign new_new_n14298__ = pi02 & ~new_new_n14297__;
  assign new_new_n14299__ = ~new_new_n868__ & new_new_n13508__;
  assign new_new_n14300__ = ~pi00 & ~new_new_n14299__;
  assign new_new_n14301__ = ~new_new_n14298__ & new_new_n14300__;
  assign new_new_n14302__ = ~new_new_n14296__ & ~new_new_n14301__;
  assign new_new_n14303__ = ~new_new_n14289__ & ~new_new_n14302__;
  assign new_new_n14304__ = ~new_new_n14288__ & ~new_new_n14303__;
  assign new_new_n14305__ = ~new_new_n13537__ & ~new_new_n14304__;
  assign new_new_n14306__ = ~new_new_n13536__ & ~new_new_n14305__;
  assign new_new_n14307__ = ~new_new_n13516__ & ~new_new_n14306__;
  assign new_new_n14308__ = new_new_n13516__ & new_new_n14306__;
  assign new_new_n14309__ = ~new_new_n13453__ & ~new_new_n13454__;
  assign new_new_n14310__ = ~new_new_n13466__ & new_new_n14309__;
  assign new_new_n14311__ = new_new_n13466__ & ~new_new_n14309__;
  assign new_new_n14312__ = ~new_new_n14310__ & ~new_new_n14311__;
  assign new_new_n14313__ = ~new_new_n14308__ & ~new_new_n14312__;
  assign new_new_n14314__ = ~new_new_n14307__ & ~new_new_n14313__;
  assign new_new_n14315__ = ~new_new_n13469__ & ~new_new_n13470__;
  assign new_new_n14316__ = new_new_n13486__ & new_new_n14315__;
  assign new_new_n14317__ = ~new_new_n13486__ & ~new_new_n14315__;
  assign new_new_n14318__ = ~new_new_n14316__ & ~new_new_n14317__;
  assign new_new_n14319__ = ~new_new_n14314__ & ~new_new_n14318__;
  assign new_new_n14320__ = new_new_n14314__ & new_new_n14318__;
  assign new_new_n14321__ = ~pi02 & ~new_new_n3742__;
  assign new_new_n14322__ = ~pi01 & new_new_n3742__;
  assign new_new_n14323__ = new_new_n583__ & ~new_new_n14321__;
  assign new_new_n14324__ = ~new_new_n14322__ & new_new_n14323__;
  assign new_new_n14325__ = pi02 & new_new_n3742__;
  assign new_new_n14326__ = pi01 & ~new_new_n3742__;
  assign new_new_n14327__ = ~new_new_n583__ & ~new_new_n14325__;
  assign new_new_n14328__ = ~new_new_n14326__ & new_new_n14327__;
  assign new_new_n14329__ = ~new_new_n14324__ & ~new_new_n14328__;
  assign new_new_n14330__ = pi00 & ~new_new_n14329__;
  assign new_new_n14331__ = pi01 & ~new_new_n691__;
  assign new_new_n14332__ = ~pi01 & ~new_new_n910__;
  assign new_new_n14333__ = pi02 & ~new_new_n14332__;
  assign new_new_n14334__ = ~new_new_n14331__ & ~new_new_n14333__;
  assign new_new_n14335__ = pi02 & new_new_n14331__;
  assign new_new_n14336__ = ~pi00 & ~new_new_n14335__;
  assign new_new_n14337__ = ~new_new_n14334__ & new_new_n14336__;
  assign new_new_n14338__ = ~new_new_n14330__ & ~new_new_n14337__;
  assign new_new_n14339__ = ~new_new_n14320__ & new_new_n14338__;
  assign new_new_n14340__ = ~new_new_n14319__ & ~new_new_n14339__;
  assign new_new_n14341__ = ~new_new_n13500__ & ~new_new_n14340__;
  assign new_new_n14342__ = ~new_new_n13499__ & ~new_new_n14341__;
  assign new_new_n14343__ = ~new_new_n12812__ & new_new_n14342__;
  assign new_new_n14344__ = new_new_n12812__ & ~new_new_n14342__;
  assign new_new_n14345__ = ~new_new_n13489__ & new_new_n13495__;
  assign new_new_n14346__ = ~new_new_n13490__ & ~new_new_n14345__;
  assign new_new_n14347__ = ~new_new_n3720__ & new_new_n11471__;
  assign new_new_n14348__ = ~new_new_n691__ & new_new_n12850__;
  assign new_new_n14349__ = ~new_new_n910__ & new_new_n11475__;
  assign new_new_n14350__ = ~new_new_n14347__ & ~new_new_n14348__;
  assign new_new_n14351__ = ~new_new_n14349__ & new_new_n14350__;
  assign new_new_n14352__ = pi05 & ~new_new_n14351__;
  assign new_new_n14353__ = new_new_n4042__ & new_new_n12856__;
  assign new_new_n14354__ = new_new_n4042__ & new_new_n11469__;
  assign new_new_n14355__ = ~pi05 & ~new_new_n14354__;
  assign new_new_n14356__ = ~new_new_n14353__ & ~new_new_n14355__;
  assign new_new_n14357__ = new_new_n14351__ & ~new_new_n14356__;
  assign new_new_n14358__ = ~new_new_n14352__ & ~new_new_n14357__;
  assign new_new_n14359__ = new_new_n12729__ & ~new_new_n14358__;
  assign new_new_n14360__ = ~new_new_n12729__ & new_new_n14358__;
  assign new_new_n14361__ = ~new_new_n14359__ & ~new_new_n14360__;
  assign new_new_n14362__ = new_new_n12741__ & new_new_n14361__;
  assign new_new_n14363__ = ~new_new_n12741__ & ~new_new_n14361__;
  assign new_new_n14364__ = ~new_new_n14362__ & ~new_new_n14363__;
  assign new_new_n14365__ = ~new_new_n14346__ & new_new_n14364__;
  assign new_new_n14366__ = new_new_n14346__ & ~new_new_n14364__;
  assign new_new_n14367__ = ~new_new_n14365__ & ~new_new_n14366__;
  assign new_new_n14368__ = ~new_new_n14344__ & new_new_n14367__;
  assign new_new_n14369__ = ~new_new_n14343__ & ~new_new_n14368__;
  assign new_new_n14370__ = ~new_new_n12729__ & ~new_new_n12741__;
  assign new_new_n14371__ = ~new_new_n12742__ & ~new_new_n14370__;
  assign new_new_n14372__ = new_new_n14346__ & new_new_n14371__;
  assign new_new_n14373__ = new_new_n14358__ & ~new_new_n14372__;
  assign new_new_n14374__ = ~new_new_n14346__ & ~new_new_n14371__;
  assign new_new_n14375__ = ~new_new_n14373__ & ~new_new_n14374__;
  assign new_new_n14376__ = new_new_n14369__ & new_new_n14375__;
  assign new_new_n14377__ = ~new_new_n12748__ & ~new_new_n12749__;
  assign new_new_n14378__ = ~new_new_n12761__ & new_new_n14377__;
  assign new_new_n14379__ = new_new_n12761__ & ~new_new_n14377__;
  assign new_new_n14380__ = ~new_new_n14378__ & ~new_new_n14379__;
  assign new_new_n14381__ = pi01 & ~new_new_n466__;
  assign new_new_n14382__ = ~pi00 & ~pi02;
  assign new_new_n14383__ = new_new_n14381__ & new_new_n14382__;
  assign new_new_n14384__ = ~new_new_n3744__ & ~new_new_n4168__;
  assign new_new_n14385__ = new_new_n3768__ & ~new_new_n14381__;
  assign new_new_n14386__ = ~new_new_n12795__ & ~new_new_n14385__;
  assign new_new_n14387__ = ~new_new_n14384__ & ~new_new_n14386__;
  assign new_new_n14388__ = ~new_new_n3768__ & new_new_n12802__;
  assign new_new_n14389__ = ~new_new_n12806__ & ~new_new_n14388__;
  assign new_new_n14390__ = new_new_n14384__ & new_new_n14389__;
  assign new_new_n14391__ = pi00 & ~new_new_n14387__;
  assign new_new_n14392__ = ~new_new_n14390__ & new_new_n14391__;
  assign new_new_n14393__ = ~pi00 & ~pi01;
  assign new_new_n14394__ = ~new_new_n466__ & ~new_new_n14393__;
  assign new_new_n14395__ = pi02 & ~new_new_n12821__;
  assign new_new_n14396__ = ~new_new_n14394__ & new_new_n14395__;
  assign new_new_n14397__ = ~new_new_n14383__ & ~new_new_n14396__;
  assign new_new_n14398__ = ~new_new_n14392__ & new_new_n14397__;
  assign new_new_n14399__ = ~new_new_n14380__ & ~new_new_n14398__;
  assign new_new_n14400__ = new_new_n14380__ & new_new_n14398__;
  assign new_new_n14401__ = ~new_new_n910__ & new_new_n13111__;
  assign new_new_n14402__ = new_new_n3742__ & new_new_n11469__;
  assign new_new_n14403__ = ~new_new_n14401__ & ~new_new_n14402__;
  assign new_new_n14404__ = new_new_n11478__ & ~new_new_n14403__;
  assign new_new_n14405__ = ~new_new_n691__ & new_new_n11475__;
  assign new_new_n14406__ = ~new_new_n14404__ & ~new_new_n14405__;
  assign new_new_n14407__ = ~pi05 & ~new_new_n14406__;
  assign new_new_n14408__ = ~new_new_n583__ & new_new_n12856__;
  assign new_new_n14409__ = ~new_new_n583__ & new_new_n11469__;
  assign new_new_n14410__ = pi05 & ~new_new_n14409__;
  assign new_new_n14411__ = ~new_new_n14408__ & ~new_new_n14410__;
  assign new_new_n14412__ = new_new_n14406__ & ~new_new_n14411__;
  assign new_new_n14413__ = ~new_new_n14407__ & ~new_new_n14412__;
  assign new_new_n14414__ = ~new_new_n14400__ & ~new_new_n14413__;
  assign new_new_n14415__ = ~new_new_n14399__ & ~new_new_n14414__;
  assign new_new_n14416__ = ~new_new_n14376__ & ~new_new_n14415__;
  assign new_new_n14417__ = ~new_new_n12768__ & ~new_new_n12769__;
  assign new_new_n14418__ = ~new_new_n12785__ & new_new_n14417__;
  assign new_new_n14419__ = new_new_n12785__ & ~new_new_n14417__;
  assign new_new_n14420__ = ~new_new_n14418__ & ~new_new_n14419__;
  assign new_new_n14421__ = ~new_new_n691__ & new_new_n11471__;
  assign new_new_n14422__ = ~new_new_n583__ & new_new_n11475__;
  assign new_new_n14423__ = ~new_new_n3768__ & new_new_n12850__;
  assign new_new_n14424__ = ~new_new_n4144__ & new_new_n13069__;
  assign new_new_n14425__ = ~new_new_n14422__ & ~new_new_n14423__;
  assign new_new_n14426__ = ~new_new_n14424__ & new_new_n14425__;
  assign new_new_n14427__ = ~new_new_n14421__ & new_new_n14426__;
  assign new_new_n14428__ = ~pi05 & ~new_new_n14427__;
  assign new_new_n14429__ = new_new_n691__ & ~new_new_n12850__;
  assign new_new_n14430__ = new_new_n11471__ & ~new_new_n14429__;
  assign new_new_n14431__ = pi05 & ~new_new_n14430__;
  assign new_new_n14432__ = new_new_n14426__ & new_new_n14431__;
  assign new_new_n14433__ = ~new_new_n14428__ & ~new_new_n14432__;
  assign new_new_n14434__ = ~new_new_n14420__ & new_new_n14433__;
  assign new_new_n14435__ = new_new_n14420__ & ~new_new_n14433__;
  assign new_new_n14436__ = ~new_new_n14434__ & ~new_new_n14435__;
  assign new_new_n14437__ = pi00 & new_new_n3768__;
  assign new_new_n14438__ = ~new_new_n14384__ & new_new_n14437__;
  assign new_new_n14439__ = new_new_n12803__ & ~new_new_n14438__;
  assign new_new_n14440__ = pi02 & ~new_new_n14439__;
  assign new_new_n14441__ = pi00 & pi01;
  assign new_new_n14442__ = new_new_n6950__ & new_new_n14441__;
  assign new_new_n14443__ = ~new_new_n14440__ & ~new_new_n14442__;
  assign new_new_n14444__ = ~new_new_n14436__ & new_new_n14443__;
  assign new_new_n14445__ = new_new_n14436__ & ~new_new_n14443__;
  assign new_new_n14446__ = ~new_new_n14444__ & ~new_new_n14445__;
  assign new_new_n14447__ = ~new_new_n14416__ & ~new_new_n14446__;
  assign new_new_n14448__ = ~new_new_n14369__ & ~new_new_n14375__;
  assign new_new_n14449__ = new_new_n14400__ & new_new_n14413__;
  assign new_new_n14450__ = new_new_n14399__ & ~new_new_n14413__;
  assign new_new_n14451__ = ~new_new_n14446__ & ~new_new_n14450__;
  assign new_new_n14452__ = ~new_new_n14449__ & ~new_new_n14451__;
  assign new_new_n14453__ = ~new_new_n14448__ & ~new_new_n14452__;
  assign new_new_n14454__ = new_new_n14376__ & new_new_n14415__;
  assign new_new_n14455__ = ~new_new_n14453__ & ~new_new_n14454__;
  assign new_new_n14456__ = ~new_new_n14447__ & new_new_n14455__;
  assign new_new_n14457__ = new_new_n12793__ & ~new_new_n14456__;
  assign new_new_n14458__ = ~new_new_n12793__ & new_new_n14456__;
  assign new_new_n14459__ = ~new_new_n14434__ & ~new_new_n14443__;
  assign new_new_n14460__ = ~new_new_n14435__ & ~new_new_n14459__;
  assign new_new_n14461__ = ~new_new_n14458__ & new_new_n14460__;
  assign new_new_n14462__ = ~new_new_n14457__ & ~new_new_n14461__;
  assign new_new_n14463__ = ~new_new_n12789__ & ~new_new_n14462__;
  assign new_new_n14464__ = ~new_new_n12073__ & ~new_new_n12078__;
  assign new_new_n14465__ = ~new_new_n12072__ & ~new_new_n14464__;
  assign new_new_n14466__ = new_new_n10690__ & ~new_new_n11393__;
  assign new_new_n14467__ = ~new_new_n10690__ & new_new_n11393__;
  assign new_new_n14468__ = ~new_new_n14466__ & ~new_new_n14467__;
  assign new_new_n14469__ = ~new_new_n11391__ & ~new_new_n11392__;
  assign new_new_n14470__ = new_new_n14468__ & ~new_new_n14469__;
  assign new_new_n14471__ = ~new_new_n14468__ & new_new_n14469__;
  assign new_new_n14472__ = ~new_new_n14470__ & ~new_new_n14471__;
  assign new_new_n14473__ = ~new_new_n14465__ & new_new_n14472__;
  assign new_new_n14474__ = new_new_n14465__ & ~new_new_n14472__;
  assign new_new_n14475__ = new_new_n466__ & ~new_new_n11482__;
  assign new_new_n14476__ = new_new_n14384__ & new_new_n14475__;
  assign new_new_n14477__ = ~new_new_n13111__ & ~new_new_n14476__;
  assign new_new_n14478__ = ~new_new_n3768__ & ~new_new_n14477__;
  assign new_new_n14479__ = ~new_new_n466__ & ~new_new_n11482__;
  assign new_new_n14480__ = new_new_n4168__ & new_new_n14479__;
  assign new_new_n14481__ = ~new_new_n14478__ & ~new_new_n14480__;
  assign new_new_n14482__ = new_new_n11478__ & ~new_new_n14481__;
  assign new_new_n14483__ = ~new_new_n466__ & new_new_n11475__;
  assign new_new_n14484__ = ~new_new_n14482__ & ~new_new_n14483__;
  assign new_new_n14485__ = ~pi05 & new_new_n14484__;
  assign new_new_n14486__ = pi05 & ~new_new_n14484__;
  assign new_new_n14487__ = ~new_new_n14485__ & ~new_new_n14486__;
  assign new_new_n14488__ = ~new_new_n14474__ & new_new_n14487__;
  assign new_new_n14489__ = ~new_new_n14473__ & ~new_new_n14488__;
  assign new_new_n14490__ = ~new_new_n14463__ & ~new_new_n14489__;
  assign new_new_n14491__ = ~new_new_n11399__ & ~new_new_n11402__;
  assign new_new_n14492__ = new_new_n11401__ & ~new_new_n14491__;
  assign new_new_n14493__ = ~new_new_n11401__ & new_new_n14491__;
  assign new_new_n14494__ = ~new_new_n14492__ & ~new_new_n14493__;
  assign new_new_n14495__ = ~new_new_n14490__ & new_new_n14494__;
  assign new_new_n14496__ = new_new_n14473__ & new_new_n14487__;
  assign new_new_n14497__ = new_new_n12789__ & new_new_n14462__;
  assign new_new_n14498__ = new_new_n14474__ & ~new_new_n14487__;
  assign new_new_n14499__ = ~new_new_n14494__ & ~new_new_n14498__;
  assign new_new_n14500__ = ~new_new_n14496__ & ~new_new_n14499__;
  assign new_new_n14501__ = ~new_new_n14497__ & new_new_n14500__;
  assign new_new_n14502__ = new_new_n14463__ & new_new_n14489__;
  assign new_new_n14503__ = ~new_new_n14501__ & ~new_new_n14502__;
  assign new_new_n14504__ = ~new_new_n14495__ & new_new_n14503__;
  assign new_new_n14505__ = ~new_new_n11423__ & ~new_new_n11424__;
  assign new_new_n14506__ = new_new_n11436__ & ~new_new_n14505__;
  assign new_new_n14507__ = ~new_new_n11436__ & new_new_n14505__;
  assign new_new_n14508__ = ~new_new_n14506__ & ~new_new_n14507__;
  assign new_new_n14509__ = ~new_new_n14504__ & ~new_new_n14508__;
  assign new_new_n14510__ = new_new_n11448__ & ~new_new_n14509__;
  assign new_new_n14511__ = new_new_n11465__ & ~new_new_n14510__;
  assign new_new_n14512__ = new_new_n14504__ & new_new_n14508__;
  assign new_new_n14513__ = ~new_new_n11448__ & ~new_new_n14512__;
  assign new_new_n14514__ = ~new_new_n11450__ & ~new_new_n14513__;
  assign new_new_n14515__ = ~new_new_n14511__ & new_new_n14514__;
  assign new_new_n14516__ = ~new_new_n11405__ & ~new_new_n11448__;
  assign new_new_n14517__ = ~new_new_n11465__ & ~new_new_n14509__;
  assign new_new_n14518__ = ~new_new_n14512__ & ~new_new_n14517__;
  assign new_new_n14519__ = ~new_new_n14516__ & ~new_new_n14518__;
  assign new_new_n14520__ = ~new_new_n11449__ & ~new_new_n14515__;
  assign new_new_n14521__ = ~new_new_n14519__ & new_new_n14520__;
  assign new_new_n14522__ = new_new_n11416__ & ~new_new_n11444__;
  assign new_new_n14523__ = ~new_new_n11443__ & ~new_new_n14522__;
  assign new_new_n14524__ = ~new_new_n14521__ & ~new_new_n14523__;
  assign new_new_n14525__ = new_new_n14521__ & new_new_n14523__;
  assign new_new_n14526__ = ~new_new_n9693__ & ~new_new_n9707__;
  assign new_new_n14527__ = ~new_new_n9706__ & new_new_n14526__;
  assign new_new_n14528__ = new_new_n9706__ & ~new_new_n14526__;
  assign new_new_n14529__ = ~new_new_n14527__ & ~new_new_n14528__;
  assign new_new_n14530__ = ~new_new_n14525__ & ~new_new_n14529__;
  assign new_new_n14531__ = ~new_new_n14524__ & ~new_new_n14530__;
  assign new_new_n14532__ = ~new_new_n9709__ & new_new_n14531__;
  assign new_new_n14533__ = ~new_new_n9685__ & new_new_n9689__;
  assign new_new_n14534__ = ~new_new_n9686__ & ~new_new_n14533__;
  assign new_new_n14535__ = ~new_new_n8507__ & ~new_new_n8508__;
  assign new_new_n14536__ = new_new_n8836__ & ~new_new_n14535__;
  assign new_new_n14537__ = ~new_new_n8836__ & new_new_n14535__;
  assign new_new_n14538__ = ~new_new_n14536__ & ~new_new_n14537__;
  assign new_new_n14539__ = new_new_n14534__ & new_new_n14538__;
  assign new_new_n14540__ = ~new_new_n14534__ & ~new_new_n14538__;
  assign new_new_n14541__ = new_new_n4172__ & new_new_n8470__;
  assign new_new_n14542__ = ~new_new_n3768__ & new_new_n8474__;
  assign new_new_n14543__ = ~new_new_n583__ & ~new_new_n8479__;
  assign new_new_n14544__ = ~new_new_n14542__ & ~new_new_n14543__;
  assign new_new_n14545__ = ~new_new_n14541__ & new_new_n14544__;
  assign new_new_n14546__ = ~new_new_n466__ & new_new_n8469__;
  assign new_new_n14547__ = pi11 & ~new_new_n14546__;
  assign new_new_n14548__ = ~new_new_n466__ & new_new_n11368__;
  assign new_new_n14549__ = ~new_new_n14547__ & ~new_new_n14548__;
  assign new_new_n14550__ = new_new_n14545__ & ~new_new_n14549__;
  assign new_new_n14551__ = ~pi11 & ~new_new_n14545__;
  assign new_new_n14552__ = ~new_new_n14550__ & ~new_new_n14551__;
  assign new_new_n14553__ = ~new_new_n14540__ & ~new_new_n14552__;
  assign new_new_n14554__ = ~new_new_n14539__ & ~new_new_n14553__;
  assign new_new_n14555__ = ~new_new_n14532__ & ~new_new_n14554__;
  assign new_new_n14556__ = ~new_new_n8839__ & ~new_new_n8840__;
  assign new_new_n14557__ = ~new_new_n8848__ & new_new_n14556__;
  assign new_new_n14558__ = new_new_n8848__ & ~new_new_n14556__;
  assign new_new_n14559__ = ~new_new_n14557__ & ~new_new_n14558__;
  assign new_new_n14560__ = ~new_new_n14555__ & new_new_n14559__;
  assign new_new_n14561__ = new_new_n9709__ & ~new_new_n14531__;
  assign new_new_n14562__ = new_new_n14540__ & new_new_n14552__;
  assign new_new_n14563__ = new_new_n14539__ & ~new_new_n14552__;
  assign new_new_n14564__ = new_new_n14559__ & ~new_new_n14563__;
  assign new_new_n14565__ = ~new_new_n14562__ & ~new_new_n14564__;
  assign new_new_n14566__ = ~new_new_n14561__ & ~new_new_n14565__;
  assign new_new_n14567__ = new_new_n14532__ & new_new_n14554__;
  assign new_new_n14568__ = ~new_new_n14566__ & ~new_new_n14567__;
  assign new_new_n14569__ = ~new_new_n14560__ & new_new_n14568__;
  assign new_new_n14570__ = ~new_new_n8850__ & new_new_n14569__;
  assign new_new_n14571__ = new_new_n8850__ & ~new_new_n14569__;
  assign new_new_n14572__ = ~new_new_n8298__ & ~new_new_n8312__;
  assign new_new_n14573__ = new_new_n8311__ & new_new_n14572__;
  assign new_new_n14574__ = ~new_new_n8311__ & ~new_new_n14572__;
  assign new_new_n14575__ = ~new_new_n14573__ & ~new_new_n14574__;
  assign new_new_n14576__ = ~new_new_n14571__ & new_new_n14575__;
  assign new_new_n14577__ = ~new_new_n14570__ & ~new_new_n14576__;
  assign new_new_n14578__ = ~new_new_n8465__ & new_new_n14577__;
  assign new_new_n14579__ = ~new_new_n8461__ & ~new_new_n14578__;
  assign new_new_n14580__ = new_new_n8317__ & new_new_n14579__;
  assign new_new_n14581__ = new_new_n8465__ & ~new_new_n14577__;
  assign new_new_n14582__ = ~new_new_n14579__ & ~new_new_n14581__;
  assign new_new_n14583__ = new_new_n8444__ & ~new_new_n14582__;
  assign new_new_n14584__ = ~new_new_n8317__ & ~new_new_n8460__;
  assign new_new_n14585__ = ~new_new_n8444__ & ~new_new_n14581__;
  assign new_new_n14586__ = ~new_new_n8318__ & ~new_new_n14584__;
  assign new_new_n14587__ = ~new_new_n14585__ & new_new_n14586__;
  assign new_new_n14588__ = ~new_new_n14580__ & ~new_new_n14587__;
  assign new_new_n14589__ = ~new_new_n14583__ & new_new_n14588__;
  assign new_new_n14590__ = pi14 & ~new_new_n8456__;
  assign new_new_n14591__ = ~new_new_n6981__ & ~new_new_n10770__;
  assign new_new_n14592__ = ~new_new_n466__ & new_new_n14591__;
  assign new_new_n14593__ = ~new_new_n14590__ & ~new_new_n14592__;
  assign new_new_n14594__ = ~new_new_n4168__ & ~new_new_n8456__;
  assign new_new_n14595__ = pi14 & new_new_n4168__;
  assign new_new_n14596__ = ~new_new_n6983__ & ~new_new_n14594__;
  assign new_new_n14597__ = ~new_new_n14595__ & new_new_n14596__;
  assign new_new_n14598__ = ~new_new_n14593__ & ~new_new_n14597__;
  assign new_new_n14599__ = ~new_new_n3768__ & new_new_n7935__;
  assign new_new_n14600__ = ~new_new_n691__ & new_new_n6964__;
  assign new_new_n14601__ = ~new_new_n583__ & new_new_n6968__;
  assign new_new_n14602__ = ~new_new_n14599__ & ~new_new_n14600__;
  assign new_new_n14603__ = ~new_new_n14601__ & new_new_n14602__;
  assign new_new_n14604__ = ~new_new_n4144__ & new_new_n6958__;
  assign new_new_n14605__ = pi17 & ~new_new_n14604__;
  assign new_new_n14606__ = ~new_new_n4144__ & new_new_n7942__;
  assign new_new_n14607__ = ~new_new_n14605__ & ~new_new_n14606__;
  assign new_new_n14608__ = new_new_n14603__ & ~new_new_n14607__;
  assign new_new_n14609__ = ~pi17 & ~new_new_n14603__;
  assign new_new_n14610__ = ~new_new_n14608__ & ~new_new_n14609__;
  assign new_new_n14611__ = ~new_new_n6921__ & ~new_new_n6922__;
  assign new_new_n14612__ = new_new_n6928__ & new_new_n14611__;
  assign new_new_n14613__ = ~new_new_n6928__ & ~new_new_n14611__;
  assign new_new_n14614__ = ~new_new_n14612__ & ~new_new_n14613__;
  assign new_new_n14615__ = ~new_new_n14610__ & ~new_new_n14614__;
  assign new_new_n14616__ = new_new_n14610__ & new_new_n14614__;
  assign new_new_n14617__ = ~new_new_n14615__ & ~new_new_n14616__;
  assign new_new_n14618__ = ~new_new_n8432__ & ~new_new_n8435__;
  assign new_new_n14619__ = ~new_new_n8431__ & ~new_new_n14618__;
  assign new_new_n14620__ = new_new_n14617__ & ~new_new_n14619__;
  assign new_new_n14621__ = ~new_new_n14617__ & new_new_n14619__;
  assign new_new_n14622__ = ~new_new_n14620__ & ~new_new_n14621__;
  assign new_new_n14623__ = new_new_n14598__ & ~new_new_n14622__;
  assign new_new_n14624__ = ~new_new_n14598__ & new_new_n14622__;
  assign new_new_n14625__ = ~new_new_n14623__ & ~new_new_n14624__;
  assign new_new_n14626__ = ~new_new_n8413__ & new_new_n8438__;
  assign new_new_n14627__ = ~new_new_n8412__ & ~new_new_n14626__;
  assign new_new_n14628__ = new_new_n14625__ & ~new_new_n14627__;
  assign new_new_n14629__ = ~new_new_n14625__ & new_new_n14627__;
  assign new_new_n14630__ = ~new_new_n14628__ & ~new_new_n14629__;
  assign new_new_n14631__ = ~new_new_n14589__ & ~new_new_n14630__;
  assign new_new_n14632__ = new_new_n14589__ & new_new_n14630__;
  assign new_new_n14633__ = ~new_new_n8395__ & ~new_new_n8441__;
  assign new_new_n14634__ = ~new_new_n8396__ & ~new_new_n14633__;
  assign new_new_n14635__ = ~new_new_n14632__ & ~new_new_n14634__;
  assign new_new_n14636__ = ~new_new_n14631__ & ~new_new_n14635__;
  assign new_new_n14637__ = ~new_new_n6947__ & new_new_n14636__;
  assign new_new_n14638__ = ~new_new_n6699__ & new_new_n6977__;
  assign new_new_n14639__ = ~new_new_n6978__ & ~new_new_n14638__;
  assign new_new_n14640__ = new_new_n14637__ & ~new_new_n14639__;
  assign new_new_n14641__ = ~new_new_n14624__ & new_new_n14627__;
  assign new_new_n14642__ = ~new_new_n14623__ & ~new_new_n14641__;
  assign new_new_n14643__ = ~new_new_n14616__ & new_new_n14619__;
  assign new_new_n14644__ = ~new_new_n14615__ & ~new_new_n14643__;
  assign new_new_n14645__ = new_new_n14642__ & new_new_n14644__;
  assign new_new_n14646__ = ~new_new_n3768__ & new_new_n6968__;
  assign new_new_n14647__ = ~new_new_n583__ & new_new_n6964__;
  assign new_new_n14648__ = ~new_new_n466__ & new_new_n7935__;
  assign new_new_n14649__ = ~new_new_n14646__ & ~new_new_n14647__;
  assign new_new_n14650__ = ~new_new_n14648__ & new_new_n14649__;
  assign new_new_n14651__ = new_new_n4172__ & new_new_n6958__;
  assign new_new_n14652__ = ~pi17 & ~new_new_n14651__;
  assign new_new_n14653__ = new_new_n4172__ & new_new_n8160__;
  assign new_new_n14654__ = ~new_new_n14652__ & ~new_new_n14653__;
  assign new_new_n14655__ = new_new_n14650__ & ~new_new_n14654__;
  assign new_new_n14656__ = pi17 & ~new_new_n14650__;
  assign new_new_n14657__ = ~new_new_n14655__ & ~new_new_n14656__;
  assign new_new_n14658__ = ~new_new_n14645__ & new_new_n14657__;
  assign new_new_n14659__ = ~new_new_n14637__ & new_new_n14639__;
  assign new_new_n14660__ = ~new_new_n14642__ & ~new_new_n14644__;
  assign new_new_n14661__ = ~new_new_n14658__ & ~new_new_n14660__;
  assign new_new_n14662__ = ~new_new_n14659__ & new_new_n14661__;
  assign new_new_n14663__ = new_new_n14657__ & new_new_n14660__;
  assign new_new_n14664__ = new_new_n14645__ & ~new_new_n14657__;
  assign new_new_n14665__ = new_new_n14639__ & ~new_new_n14664__;
  assign new_new_n14666__ = new_new_n6947__ & ~new_new_n14636__;
  assign new_new_n14667__ = ~new_new_n14663__ & ~new_new_n14665__;
  assign new_new_n14668__ = ~new_new_n14666__ & new_new_n14667__;
  assign new_new_n14669__ = ~new_new_n14640__ & ~new_new_n14668__;
  assign new_new_n14670__ = ~new_new_n14662__ & new_new_n14669__;
  assign new_new_n14671__ = new_new_n6980__ & ~new_new_n14670__;
  assign new_new_n14672__ = ~new_new_n6647__ & ~new_new_n6696__;
  assign new_new_n14673__ = ~new_new_n6646__ & ~new_new_n14672__;
  assign new_new_n14674__ = ~new_new_n3720__ & new_new_n5183__;
  assign new_new_n14675__ = ~new_new_n868__ & new_new_n5191__;
  assign new_new_n14676__ = ~new_new_n14674__ & ~new_new_n14675__;
  assign new_new_n14677__ = new_new_n5116__ & new_new_n5195__;
  assign new_new_n14678__ = new_new_n14676__ & ~new_new_n14677__;
  assign new_new_n14679__ = pi23 & ~new_new_n14678__;
  assign new_new_n14680__ = ~new_new_n5129__ & new_new_n5195__;
  assign new_new_n14681__ = ~pi23 & ~new_new_n14680__;
  assign new_new_n14682__ = pi22 & new_new_n910__;
  assign new_new_n14683__ = ~pi22 & ~new_new_n910__;
  assign new_new_n14684__ = new_new_n5195__ & ~new_new_n14682__;
  assign new_new_n14685__ = ~new_new_n14683__ & new_new_n14684__;
  assign new_new_n14686__ = new_new_n4036__ & new_new_n14685__;
  assign new_new_n14687__ = ~new_new_n14681__ & ~new_new_n14686__;
  assign new_new_n14688__ = new_new_n14676__ & ~new_new_n14687__;
  assign new_new_n14689__ = ~new_new_n14679__ & ~new_new_n14688__;
  assign new_new_n14690__ = ~new_new_n5681__ & ~new_new_n5682__;
  assign new_new_n14691__ = new_new_n5740__ & new_new_n14690__;
  assign new_new_n14692__ = ~new_new_n5740__ & ~new_new_n14690__;
  assign new_new_n14693__ = ~new_new_n14691__ & ~new_new_n14692__;
  assign new_new_n14694__ = ~new_new_n14689__ & new_new_n14693__;
  assign new_new_n14695__ = new_new_n14689__ & ~new_new_n14693__;
  assign new_new_n14696__ = ~new_new_n14694__ & ~new_new_n14695__;
  assign new_new_n14697__ = ~new_new_n6660__ & ~new_new_n6668__;
  assign new_new_n14698__ = ~new_new_n6667__ & ~new_new_n14697__;
  assign new_new_n14699__ = new_new_n14696__ & ~new_new_n14698__;
  assign new_new_n14700__ = ~new_new_n14696__ & new_new_n14698__;
  assign new_new_n14701__ = ~new_new_n14699__ & ~new_new_n14700__;
  assign new_new_n14702__ = ~new_new_n3768__ & new_new_n6634__;
  assign new_new_n14703__ = ~new_new_n691__ & ~new_new_n6625__;
  assign new_new_n14704__ = ~new_new_n583__ & new_new_n6629__;
  assign new_new_n14705__ = ~new_new_n14702__ & ~new_new_n14703__;
  assign new_new_n14706__ = ~new_new_n14704__ & new_new_n14705__;
  assign new_new_n14707__ = ~new_new_n4144__ & new_new_n6631__;
  assign new_new_n14708__ = pi20 & ~new_new_n14707__;
  assign new_new_n14709__ = ~new_new_n4144__ & new_new_n6640__;
  assign new_new_n14710__ = ~new_new_n14708__ & ~new_new_n14709__;
  assign new_new_n14711__ = new_new_n14706__ & ~new_new_n14710__;
  assign new_new_n14712__ = ~pi20 & ~new_new_n14706__;
  assign new_new_n14713__ = ~new_new_n14711__ & ~new_new_n14712__;
  assign new_new_n14714__ = new_new_n14701__ & new_new_n14713__;
  assign new_new_n14715__ = ~new_new_n14701__ & ~new_new_n14713__;
  assign new_new_n14716__ = ~new_new_n14714__ & ~new_new_n14715__;
  assign new_new_n14717__ = ~new_new_n6660__ & ~new_new_n6669__;
  assign new_new_n14718__ = new_new_n6660__ & new_new_n6669__;
  assign new_new_n14719__ = ~new_new_n14717__ & ~new_new_n14718__;
  assign new_new_n14720__ = ~new_new_n6691__ & ~new_new_n14719__;
  assign new_new_n14721__ = ~new_new_n6692__ & ~new_new_n14720__;
  assign new_new_n14722__ = new_new_n14716__ & new_new_n14721__;
  assign new_new_n14723__ = ~new_new_n14716__ & ~new_new_n14721__;
  assign new_new_n14724__ = ~new_new_n14722__ & ~new_new_n14723__;
  assign new_new_n14725__ = new_new_n14673__ & ~new_new_n14724__;
  assign new_new_n14726__ = ~new_new_n14673__ & new_new_n14724__;
  assign new_new_n14727__ = ~pi16 & ~new_new_n466__;
  assign new_new_n14728__ = pi17 & ~new_new_n14727__;
  assign new_new_n14729__ = ~new_new_n6953__ & ~new_new_n6956__;
  assign new_new_n14730__ = ~new_new_n466__ & new_new_n14729__;
  assign new_new_n14731__ = ~new_new_n14728__ & ~new_new_n14730__;
  assign new_new_n14732__ = ~new_new_n4168__ & ~new_new_n14727__;
  assign new_new_n14733__ = pi17 & new_new_n4168__;
  assign new_new_n14734__ = ~new_new_n6957__ & ~new_new_n14732__;
  assign new_new_n14735__ = ~new_new_n14733__ & new_new_n14734__;
  assign new_new_n14736__ = ~new_new_n14731__ & ~new_new_n14735__;
  assign new_new_n14737__ = ~new_new_n14726__ & ~new_new_n14736__;
  assign new_new_n14738__ = ~new_new_n14725__ & ~new_new_n14737__;
  assign new_new_n14739__ = ~new_new_n14671__ & new_new_n14738__;
  assign new_new_n14740__ = ~new_new_n3768__ & new_new_n6629__;
  assign new_new_n14741__ = ~new_new_n466__ & new_new_n6634__;
  assign new_new_n14742__ = ~new_new_n583__ & ~new_new_n6625__;
  assign new_new_n14743__ = new_new_n4172__ & new_new_n6936__;
  assign new_new_n14744__ = ~new_new_n14740__ & ~new_new_n14741__;
  assign new_new_n14745__ = ~new_new_n14742__ & new_new_n14744__;
  assign new_new_n14746__ = ~new_new_n14743__ & new_new_n14745__;
  assign new_new_n14747__ = pi20 & ~new_new_n14746__;
  assign new_new_n14748__ = ~pi20 & new_new_n14746__;
  assign new_new_n14749__ = ~new_new_n14747__ & ~new_new_n14748__;
  assign new_new_n14750__ = ~new_new_n14694__ & ~new_new_n14699__;
  assign new_new_n14751__ = new_new_n4042__ & new_new_n5215__;
  assign new_new_n14752__ = ~new_new_n691__ & new_new_n5213__;
  assign new_new_n14753__ = ~new_new_n3720__ & new_new_n5191__;
  assign new_new_n14754__ = ~new_new_n910__ & new_new_n5183__;
  assign new_new_n14755__ = ~new_new_n14752__ & ~new_new_n14753__;
  assign new_new_n14756__ = ~new_new_n14754__ & new_new_n14755__;
  assign new_new_n14757__ = ~new_new_n14751__ & new_new_n14756__;
  assign new_new_n14758__ = ~pi23 & ~new_new_n14757__;
  assign new_new_n14759__ = pi23 & new_new_n14757__;
  assign new_new_n14760__ = ~new_new_n14758__ & ~new_new_n14759__;
  assign new_new_n14761__ = new_new_n14750__ & ~new_new_n14760__;
  assign new_new_n14762__ = ~new_new_n14750__ & new_new_n14760__;
  assign new_new_n14763__ = ~new_new_n14761__ & ~new_new_n14762__;
  assign new_new_n14764__ = ~new_new_n5860__ & ~new_new_n5871__;
  assign new_new_n14765__ = new_new_n5870__ & new_new_n14764__;
  assign new_new_n14766__ = ~new_new_n5870__ & ~new_new_n14764__;
  assign new_new_n14767__ = ~new_new_n14765__ & ~new_new_n14766__;
  assign new_new_n14768__ = ~new_new_n14763__ & new_new_n14767__;
  assign new_new_n14769__ = new_new_n14763__ & ~new_new_n14767__;
  assign new_new_n14770__ = ~new_new_n14768__ & ~new_new_n14769__;
  assign new_new_n14771__ = ~new_new_n14714__ & new_new_n14721__;
  assign new_new_n14772__ = ~new_new_n14715__ & ~new_new_n14771__;
  assign new_new_n14773__ = ~new_new_n14770__ & ~new_new_n14772__;
  assign new_new_n14774__ = new_new_n14770__ & new_new_n14772__;
  assign new_new_n14775__ = ~new_new_n14773__ & ~new_new_n14774__;
  assign new_new_n14776__ = new_new_n14749__ & ~new_new_n14775__;
  assign new_new_n14777__ = ~new_new_n14749__ & new_new_n14775__;
  assign new_new_n14778__ = ~new_new_n14776__ & ~new_new_n14777__;
  assign new_new_n14779__ = ~new_new_n14739__ & new_new_n14778__;
  assign new_new_n14780__ = new_new_n14726__ & new_new_n14736__;
  assign new_new_n14781__ = ~new_new_n6980__ & new_new_n14670__;
  assign new_new_n14782__ = new_new_n14725__ & ~new_new_n14736__;
  assign new_new_n14783__ = ~new_new_n14778__ & ~new_new_n14782__;
  assign new_new_n14784__ = ~new_new_n14780__ & ~new_new_n14783__;
  assign new_new_n14785__ = ~new_new_n14781__ & new_new_n14784__;
  assign new_new_n14786__ = new_new_n14671__ & ~new_new_n14738__;
  assign new_new_n14787__ = ~new_new_n14785__ & ~new_new_n14786__;
  assign new_new_n14788__ = ~new_new_n14779__ & new_new_n14787__;
  assign new_new_n14789__ = new_new_n5966__ & new_new_n14788__;
  assign new_new_n14790__ = ~new_new_n583__ & new_new_n5183__;
  assign new_new_n14791__ = new_new_n3768__ & ~new_new_n5212__;
  assign new_new_n14792__ = new_new_n4144__ & new_new_n5212__;
  assign new_new_n14793__ = new_new_n5195__ & ~new_new_n14791__;
  assign new_new_n14794__ = ~new_new_n14792__ & new_new_n14793__;
  assign new_new_n14795__ = ~new_new_n14790__ & ~new_new_n14794__;
  assign new_new_n14796__ = ~new_new_n691__ & new_new_n5185__;
  assign new_new_n14797__ = pi23 & ~new_new_n14796__;
  assign new_new_n14798__ = ~new_new_n691__ & new_new_n5188__;
  assign new_new_n14799__ = ~pi23 & ~new_new_n14798__;
  assign new_new_n14800__ = pi20 & ~new_new_n14799__;
  assign new_new_n14801__ = ~new_new_n14797__ & ~new_new_n14800__;
  assign new_new_n14802__ = new_new_n14795__ & ~new_new_n14801__;
  assign new_new_n14803__ = ~pi23 & ~new_new_n14795__;
  assign new_new_n14804__ = ~new_new_n14802__ & ~new_new_n14803__;
  assign new_new_n14805__ = ~new_new_n5913__ & new_new_n5931__;
  assign new_new_n14806__ = new_new_n5913__ & ~new_new_n5931__;
  assign new_new_n14807__ = ~new_new_n5911__ & ~new_new_n5941__;
  assign new_new_n14808__ = new_new_n5911__ & new_new_n5941__;
  assign new_new_n14809__ = ~new_new_n14807__ & ~new_new_n14808__;
  assign new_new_n14810__ = ~new_new_n5945__ & ~new_new_n14809__;
  assign new_new_n14811__ = new_new_n5945__ & new_new_n14809__;
  assign new_new_n14812__ = ~new_new_n14806__ & ~new_new_n14810__;
  assign new_new_n14813__ = ~new_new_n14811__ & new_new_n14812__;
  assign new_new_n14814__ = ~new_new_n14805__ & ~new_new_n14813__;
  assign new_new_n14815__ = new_new_n5896__ & new_new_n5941__;
  assign new_new_n14816__ = ~new_new_n5908__ & ~new_new_n5942__;
  assign new_new_n14817__ = new_new_n5908__ & new_new_n5942__;
  assign new_new_n14818__ = ~new_new_n4452__ & ~new_new_n14817__;
  assign new_new_n14819__ = ~new_new_n14816__ & ~new_new_n14818__;
  assign new_new_n14820__ = new_new_n14815__ & new_new_n14819__;
  assign new_new_n14821__ = new_new_n4452__ & ~new_new_n5056__;
  assign new_new_n14822__ = ~new_new_n4452__ & new_new_n5056__;
  assign new_new_n14823__ = ~new_new_n14821__ & ~new_new_n14822__;
  assign new_new_n14824__ = new_new_n5020__ & new_new_n14823__;
  assign new_new_n14825__ = ~new_new_n5020__ & ~new_new_n14823__;
  assign new_new_n14826__ = ~new_new_n14824__ & ~new_new_n14825__;
  assign new_new_n14827__ = ~new_new_n5896__ & ~new_new_n5941__;
  assign new_new_n14828__ = ~new_new_n14816__ & ~new_new_n14817__;
  assign new_new_n14829__ = new_new_n5945__ & ~new_new_n14828__;
  assign new_new_n14830__ = ~new_new_n14815__ & ~new_new_n14827__;
  assign new_new_n14831__ = ~new_new_n14829__ & new_new_n14830__;
  assign new_new_n14832__ = ~new_new_n14819__ & new_new_n14827__;
  assign new_new_n14833__ = ~new_new_n14820__ & new_new_n14826__;
  assign new_new_n14834__ = ~new_new_n14831__ & ~new_new_n14832__;
  assign new_new_n14835__ = new_new_n14833__ & new_new_n14834__;
  assign new_new_n14836__ = ~new_new_n5908__ & new_new_n5941__;
  assign new_new_n14837__ = new_new_n5896__ & new_new_n14836__;
  assign new_new_n14838__ = ~new_new_n5942__ & new_new_n14837__;
  assign new_new_n14839__ = new_new_n14817__ & new_new_n14827__;
  assign new_new_n14840__ = new_new_n5908__ & new_new_n14827__;
  assign new_new_n14841__ = ~new_new_n5908__ & ~new_new_n14827__;
  assign new_new_n14842__ = ~new_new_n14815__ & ~new_new_n14841__;
  assign new_new_n14843__ = new_new_n5942__ & new_new_n14842__;
  assign new_new_n14844__ = new_new_n4452__ & ~new_new_n14840__;
  assign new_new_n14845__ = ~new_new_n14843__ & new_new_n14844__;
  assign new_new_n14846__ = ~new_new_n5942__ & ~new_new_n14842__;
  assign new_new_n14847__ = ~new_new_n4452__ & ~new_new_n14837__;
  assign new_new_n14848__ = ~new_new_n14846__ & new_new_n14847__;
  assign new_new_n14849__ = ~new_new_n14845__ & ~new_new_n14848__;
  assign new_new_n14850__ = ~new_new_n14826__ & ~new_new_n14839__;
  assign new_new_n14851__ = ~new_new_n14838__ & new_new_n14850__;
  assign new_new_n14852__ = ~new_new_n14849__ & new_new_n14851__;
  assign new_new_n14853__ = ~new_new_n14835__ & ~new_new_n14852__;
  assign new_new_n14854__ = ~new_new_n333__ & ~new_new_n868__;
  assign new_new_n14855__ = new_new_n873__ & ~new_new_n3720__;
  assign new_new_n14856__ = ~new_new_n14854__ & ~new_new_n14855__;
  assign new_new_n14857__ = pi25 & new_new_n4036__;
  assign new_new_n14858__ = ~new_new_n110__ & ~new_new_n5127__;
  assign new_new_n14859__ = ~new_new_n5129__ & ~new_new_n14857__;
  assign new_new_n14860__ = new_new_n14858__ & new_new_n14859__;
  assign new_new_n14861__ = new_new_n14856__ & ~new_new_n14860__;
  assign new_new_n14862__ = pi26 & ~new_new_n14861__;
  assign new_new_n14863__ = new_new_n910__ & ~new_new_n14857__;
  assign new_new_n14864__ = pi25 & new_new_n5127__;
  assign new_new_n14865__ = ~new_new_n110__ & ~new_new_n14863__;
  assign new_new_n14866__ = ~new_new_n14864__ & new_new_n14865__;
  assign new_new_n14867__ = ~pi26 & new_new_n14856__;
  assign new_new_n14868__ = ~new_new_n14866__ & new_new_n14867__;
  assign new_new_n14869__ = ~new_new_n14862__ & ~new_new_n14868__;
  assign new_new_n14870__ = ~new_new_n14853__ & ~new_new_n14869__;
  assign new_new_n14871__ = new_new_n14853__ & new_new_n14869__;
  assign new_new_n14872__ = ~new_new_n14870__ & ~new_new_n14871__;
  assign new_new_n14873__ = ~new_new_n1061__ & new_new_n4212__;
  assign new_new_n14874__ = ~new_new_n3618__ & ~new_new_n4818__;
  assign new_new_n14875__ = ~new_new_n1207__ & new_new_n4815__;
  assign new_new_n14876__ = ~new_new_n14873__ & ~new_new_n14874__;
  assign new_new_n14877__ = ~new_new_n14875__ & new_new_n14876__;
  assign new_new_n14878__ = new_new_n4214__ & ~new_new_n5235__;
  assign new_new_n14879__ = ~pi29 & ~new_new_n14878__;
  assign new_new_n14880__ = ~new_new_n5235__ & new_new_n5732__;
  assign new_new_n14881__ = ~new_new_n14879__ & ~new_new_n14880__;
  assign new_new_n14882__ = new_new_n14877__ & ~new_new_n14881__;
  assign new_new_n14883__ = pi29 & ~new_new_n14877__;
  assign new_new_n14884__ = ~new_new_n14882__ & ~new_new_n14883__;
  assign new_new_n14885__ = new_new_n14872__ & ~new_new_n14884__;
  assign new_new_n14886__ = ~new_new_n14872__ & new_new_n14884__;
  assign new_new_n14887__ = ~new_new_n14885__ & ~new_new_n14886__;
  assign new_new_n14888__ = new_new_n14814__ & new_new_n14887__;
  assign new_new_n14889__ = ~new_new_n14814__ & ~new_new_n14887__;
  assign new_new_n14890__ = ~new_new_n14888__ & ~new_new_n14889__;
  assign new_new_n14891__ = ~new_new_n14804__ & ~new_new_n14890__;
  assign new_new_n14892__ = new_new_n14804__ & new_new_n14890__;
  assign new_new_n14893__ = ~new_new_n14891__ & ~new_new_n14892__;
  assign new_new_n14894__ = pi19 & ~new_new_n466__;
  assign new_new_n14895__ = ~pi20 & ~new_new_n14894__;
  assign new_new_n14896__ = pi19 & pi20;
  assign new_new_n14897__ = ~new_new_n6619__ & ~new_new_n14896__;
  assign new_new_n14898__ = ~new_new_n466__ & new_new_n14897__;
  assign new_new_n14899__ = ~new_new_n14895__ & ~new_new_n14898__;
  assign new_new_n14900__ = ~new_new_n4168__ & ~new_new_n14894__;
  assign new_new_n14901__ = ~pi20 & new_new_n4168__;
  assign new_new_n14902__ = ~new_new_n6622__ & ~new_new_n14900__;
  assign new_new_n14903__ = ~new_new_n14901__ & new_new_n14902__;
  assign new_new_n14904__ = ~new_new_n14899__ & ~new_new_n14903__;
  assign new_new_n14905__ = ~new_new_n5958__ & ~new_new_n5966__;
  assign new_new_n14906__ = ~new_new_n5959__ & ~new_new_n14905__;
  assign new_new_n14907__ = ~new_new_n14904__ & ~new_new_n14906__;
  assign new_new_n14908__ = new_new_n14904__ & new_new_n14906__;
  assign new_new_n14909__ = ~new_new_n14907__ & ~new_new_n14908__;
  assign new_new_n14910__ = new_new_n14893__ & ~new_new_n14909__;
  assign new_new_n14911__ = ~new_new_n14893__ & new_new_n14909__;
  assign new_new_n14912__ = ~new_new_n14910__ & ~new_new_n14911__;
  assign new_new_n14913__ = new_new_n14789__ & new_new_n14912__;
  assign new_new_n14914__ = ~new_new_n14789__ & ~new_new_n14912__;
  assign new_new_n14915__ = new_new_n14749__ & ~new_new_n14774__;
  assign new_new_n14916__ = ~new_new_n14773__ & ~new_new_n14915__;
  assign new_new_n14917__ = ~new_new_n14761__ & ~new_new_n14767__;
  assign new_new_n14918__ = ~new_new_n14762__ & ~new_new_n14917__;
  assign new_new_n14919__ = new_new_n14916__ & ~new_new_n14918__;
  assign new_new_n14920__ = new_new_n6936__ & new_new_n6952__;
  assign new_new_n14921__ = ~new_new_n3768__ & ~new_new_n6625__;
  assign new_new_n14922__ = ~new_new_n466__ & new_new_n6629__;
  assign new_new_n14923__ = ~new_new_n14921__ & ~new_new_n14922__;
  assign new_new_n14924__ = ~new_new_n14920__ & new_new_n14923__;
  assign new_new_n14925__ = ~pi20 & new_new_n14924__;
  assign new_new_n14926__ = pi20 & ~new_new_n14924__;
  assign new_new_n14927__ = ~new_new_n14925__ & ~new_new_n14926__;
  assign new_new_n14928__ = ~new_new_n14916__ & new_new_n14918__;
  assign new_new_n14929__ = ~new_new_n5966__ & ~new_new_n14788__;
  assign new_new_n14930__ = new_new_n14912__ & ~new_new_n14929__;
  assign new_new_n14931__ = ~new_new_n14927__ & ~new_new_n14928__;
  assign new_new_n14932__ = ~new_new_n14930__ & new_new_n14931__;
  assign new_new_n14933__ = ~new_new_n14914__ & ~new_new_n14919__;
  assign new_new_n14934__ = ~new_new_n14932__ & new_new_n14933__;
  assign new_new_n14935__ = ~new_new_n14912__ & ~new_new_n14928__;
  assign new_new_n14936__ = new_new_n14927__ & ~new_new_n14935__;
  assign new_new_n14937__ = ~new_new_n14929__ & new_new_n14936__;
  assign new_new_n14938__ = ~new_new_n14913__ & ~new_new_n14937__;
  assign new_new_n14939__ = ~new_new_n14934__ & new_new_n14938__;
  assign new_new_n14940__ = ~new_new_n5207__ & new_new_n14939__;
  assign new_new_n14941__ = new_new_n5215__ & new_new_n6952__;
  assign new_new_n14942__ = ~new_new_n3768__ & new_new_n5191__;
  assign new_new_n14943__ = ~new_new_n466__ & new_new_n5183__;
  assign new_new_n14944__ = ~new_new_n14942__ & ~new_new_n14943__;
  assign new_new_n14945__ = ~new_new_n14941__ & new_new_n14944__;
  assign new_new_n14946__ = pi23 & ~new_new_n14945__;
  assign new_new_n14947__ = ~pi23 & new_new_n14945__;
  assign new_new_n14948__ = ~new_new_n14946__ & ~new_new_n14947__;
  assign new_new_n14949__ = ~new_new_n333__ & ~new_new_n910__;
  assign new_new_n14950__ = ~new_new_n691__ & new_new_n873__;
  assign new_new_n14951__ = ~new_new_n583__ & new_new_n3311__;
  assign new_new_n14952__ = ~new_new_n14950__ & ~new_new_n14951__;
  assign new_new_n14953__ = ~new_new_n14949__ & new_new_n14952__;
  assign new_new_n14954__ = ~pi26 & ~new_new_n14953__;
  assign new_new_n14955__ = new_new_n512__ & new_new_n3742__;
  assign new_new_n14956__ = new_new_n801__ & new_new_n3742__;
  assign new_new_n14957__ = pi26 & ~new_new_n14956__;
  assign new_new_n14958__ = ~new_new_n14955__ & ~new_new_n14957__;
  assign new_new_n14959__ = new_new_n14953__ & ~new_new_n14958__;
  assign new_new_n14960__ = ~new_new_n14954__ & ~new_new_n14959__;
  assign new_new_n14961__ = ~new_new_n4385__ & ~new_new_n5068__;
  assign new_new_n14962__ = new_new_n4385__ & new_new_n5068__;
  assign new_new_n14963__ = ~new_new_n14961__ & ~new_new_n14962__;
  assign new_new_n14964__ = ~new_new_n5020__ & ~new_new_n14821__;
  assign new_new_n14965__ = ~new_new_n14822__ & ~new_new_n14964__;
  assign new_new_n14966__ = pi20 & ~new_new_n5056__;
  assign new_new_n14967__ = ~pi20 & new_new_n5056__;
  assign new_new_n14968__ = ~new_new_n14966__ & ~new_new_n14967__;
  assign new_new_n14969__ = new_new_n14965__ & new_new_n14968__;
  assign new_new_n14970__ = ~new_new_n14965__ & ~new_new_n14968__;
  assign new_new_n14971__ = ~new_new_n14969__ & ~new_new_n14970__;
  assign new_new_n14972__ = new_new_n14963__ & new_new_n14971__;
  assign new_new_n14973__ = ~new_new_n4353__ & new_new_n4385__;
  assign new_new_n14974__ = ~new_new_n14963__ & ~new_new_n14973__;
  assign new_new_n14975__ = ~new_new_n14971__ & new_new_n14974__;
  assign new_new_n14976__ = ~new_new_n14972__ & ~new_new_n14975__;
  assign new_new_n14977__ = new_new_n5908__ & ~new_new_n5941__;
  assign new_new_n14978__ = ~new_new_n14826__ & new_new_n14977__;
  assign new_new_n14979__ = new_new_n14826__ & ~new_new_n14977__;
  assign new_new_n14980__ = new_new_n5896__ & ~new_new_n5942__;
  assign new_new_n14981__ = ~new_new_n5896__ & new_new_n5942__;
  assign new_new_n14982__ = ~new_new_n14826__ & ~new_new_n14836__;
  assign new_new_n14983__ = ~new_new_n4452__ & ~new_new_n14981__;
  assign new_new_n14984__ = ~new_new_n14982__ & new_new_n14983__;
  assign new_new_n14985__ = ~new_new_n14979__ & ~new_new_n14980__;
  assign new_new_n14986__ = ~new_new_n14984__ & new_new_n14985__;
  assign new_new_n14987__ = new_new_n14826__ & ~new_new_n14981__;
  assign new_new_n14988__ = new_new_n4452__ & ~new_new_n14987__;
  assign new_new_n14989__ = ~new_new_n14836__ & new_new_n14988__;
  assign new_new_n14990__ = ~new_new_n14978__ & ~new_new_n14989__;
  assign new_new_n14991__ = ~new_new_n14986__ & new_new_n14990__;
  assign new_new_n14992__ = new_new_n14976__ & ~new_new_n14991__;
  assign new_new_n14993__ = ~new_new_n14976__ & new_new_n14991__;
  assign new_new_n14994__ = ~new_new_n4550__ & new_new_n4813__;
  assign new_new_n14995__ = ~new_new_n868__ & new_new_n4815__;
  assign new_new_n14996__ = ~new_new_n1061__ & ~new_new_n4818__;
  assign new_new_n14997__ = ~new_new_n1207__ & new_new_n4212__;
  assign new_new_n14998__ = ~new_new_n14995__ & ~new_new_n14996__;
  assign new_new_n14999__ = ~new_new_n14997__ & new_new_n14998__;
  assign new_new_n15000__ = ~new_new_n14994__ & new_new_n14999__;
  assign new_new_n15001__ = ~new_new_n14992__ & ~new_new_n14993__;
  assign new_new_n15002__ = pi29 & ~new_new_n15001__;
  assign new_new_n15003__ = ~pi29 & new_new_n15001__;
  assign new_new_n15004__ = ~new_new_n15002__ & ~new_new_n15003__;
  assign new_new_n15005__ = new_new_n15000__ & new_new_n15004__;
  assign new_new_n15006__ = ~new_new_n15000__ & ~new_new_n15004__;
  assign new_new_n15007__ = ~new_new_n15005__ & ~new_new_n15006__;
  assign new_new_n15008__ = ~new_new_n14993__ & ~new_new_n15007__;
  assign new_new_n15009__ = ~new_new_n14992__ & ~new_new_n15008__;
  assign new_new_n15010__ = new_new_n14960__ & new_new_n15009__;
  assign new_new_n15011__ = ~new_new_n14960__ & ~new_new_n15009__;
  assign new_new_n15012__ = ~new_new_n15010__ & ~new_new_n15011__;
  assign new_new_n15013__ = ~new_new_n5086__ & ~new_new_n5087__;
  assign new_new_n15014__ = new_new_n5103__ & new_new_n15013__;
  assign new_new_n15015__ = ~new_new_n5103__ & ~new_new_n15013__;
  assign new_new_n15016__ = ~new_new_n15014__ & ~new_new_n15015__;
  assign new_new_n15017__ = new_new_n15012__ & ~new_new_n15016__;
  assign new_new_n15018__ = ~new_new_n15012__ & new_new_n15016__;
  assign new_new_n15019__ = ~new_new_n15017__ & ~new_new_n15018__;
  assign new_new_n15020__ = ~new_new_n333__ & ~new_new_n3720__;
  assign new_new_n15021__ = ~new_new_n691__ & new_new_n3311__;
  assign new_new_n15022__ = new_new_n873__ & ~new_new_n910__;
  assign new_new_n15023__ = ~new_new_n15020__ & ~new_new_n15021__;
  assign new_new_n15024__ = ~new_new_n15022__ & new_new_n15023__;
  assign new_new_n15025__ = ~pi26 & ~new_new_n15024__;
  assign new_new_n15026__ = new_new_n512__ & new_new_n4042__;
  assign new_new_n15027__ = new_new_n801__ & new_new_n4042__;
  assign new_new_n15028__ = pi26 & ~new_new_n15027__;
  assign new_new_n15029__ = ~new_new_n15026__ & ~new_new_n15028__;
  assign new_new_n15030__ = new_new_n15024__ & ~new_new_n15029__;
  assign new_new_n15031__ = ~new_new_n15025__ & ~new_new_n15030__;
  assign new_new_n15032__ = ~new_new_n15007__ & new_new_n15031__;
  assign new_new_n15033__ = new_new_n15007__ & ~new_new_n15031__;
  assign new_new_n15034__ = ~new_new_n14871__ & ~new_new_n14884__;
  assign new_new_n15035__ = ~new_new_n14870__ & ~new_new_n15034__;
  assign new_new_n15036__ = ~new_new_n15033__ & ~new_new_n15035__;
  assign new_new_n15037__ = ~new_new_n15032__ & ~new_new_n15036__;
  assign new_new_n15038__ = new_new_n15019__ & new_new_n15037__;
  assign new_new_n15039__ = ~new_new_n15019__ & ~new_new_n15037__;
  assign new_new_n15040__ = ~new_new_n15038__ & ~new_new_n15039__;
  assign new_new_n15041__ = new_new_n14948__ & ~new_new_n15040__;
  assign new_new_n15042__ = ~new_new_n14948__ & new_new_n15040__;
  assign new_new_n15043__ = ~new_new_n15041__ & ~new_new_n15042__;
  assign new_new_n15044__ = new_new_n14940__ & new_new_n15043__;
  assign new_new_n15045__ = ~new_new_n14888__ & ~new_new_n14892__;
  assign new_new_n15046__ = ~new_new_n14893__ & ~new_new_n14908__;
  assign new_new_n15047__ = ~new_new_n14907__ & ~new_new_n15046__;
  assign new_new_n15048__ = ~new_new_n15045__ & new_new_n15047__;
  assign new_new_n15049__ = ~new_new_n15043__ & ~new_new_n15048__;
  assign new_new_n15050__ = new_new_n15045__ & ~new_new_n15047__;
  assign new_new_n15051__ = new_new_n15043__ & ~new_new_n15050__;
  assign new_new_n15052__ = ~new_new_n15032__ & ~new_new_n15033__;
  assign new_new_n15053__ = new_new_n15035__ & new_new_n15052__;
  assign new_new_n15054__ = ~new_new_n15035__ & ~new_new_n15052__;
  assign new_new_n15055__ = ~new_new_n15053__ & ~new_new_n15054__;
  assign new_new_n15056__ = ~new_new_n15051__ & new_new_n15055__;
  assign new_new_n15057__ = new_new_n5207__ & ~new_new_n14939__;
  assign new_new_n15058__ = ~new_new_n15049__ & ~new_new_n15056__;
  assign new_new_n15059__ = ~new_new_n15057__ & new_new_n15058__;
  assign new_new_n15060__ = ~new_new_n15048__ & new_new_n15055__;
  assign new_new_n15061__ = ~new_new_n14940__ & ~new_new_n15043__;
  assign new_new_n15062__ = ~new_new_n15050__ & ~new_new_n15060__;
  assign new_new_n15063__ = ~new_new_n15061__ & new_new_n15062__;
  assign new_new_n15064__ = ~new_new_n15044__ & ~new_new_n15059__;
  assign new_new_n15065__ = ~new_new_n15063__ & new_new_n15064__;
  assign new_new_n15066__ = ~new_new_n14948__ & ~new_new_n15038__;
  assign new_new_n15067__ = ~new_new_n15039__ & ~new_new_n15066__;
  assign new_new_n15068__ = ~new_new_n15065__ & ~new_new_n15067__;
  assign new_new_n15069__ = ~new_new_n15011__ & new_new_n15016__;
  assign new_new_n15070__ = ~new_new_n15010__ & ~new_new_n15069__;
  assign new_new_n15071__ = ~new_new_n5137__ & ~new_new_n5138__;
  assign new_new_n15072__ = new_new_n5148__ & new_new_n15071__;
  assign new_new_n15073__ = ~new_new_n5148__ & ~new_new_n15071__;
  assign new_new_n15074__ = ~new_new_n15072__ & ~new_new_n15073__;
  assign new_new_n15075__ = ~new_new_n15070__ & ~new_new_n15074__;
  assign new_new_n15076__ = new_new_n15070__ & new_new_n15074__;
  assign new_new_n15077__ = pi23 & ~new_new_n5201__;
  assign new_new_n15078__ = ~new_new_n5179__ & ~new_new_n5210__;
  assign new_new_n15079__ = ~new_new_n466__ & new_new_n15078__;
  assign new_new_n15080__ = ~new_new_n15077__ & ~new_new_n15079__;
  assign new_new_n15081__ = ~new_new_n4168__ & ~new_new_n5201__;
  assign new_new_n15082__ = pi23 & new_new_n4168__;
  assign new_new_n15083__ = ~new_new_n5181__ & ~new_new_n15081__;
  assign new_new_n15084__ = ~new_new_n15082__ & new_new_n15083__;
  assign new_new_n15085__ = ~new_new_n15080__ & ~new_new_n15084__;
  assign new_new_n15086__ = ~new_new_n15076__ & ~new_new_n15085__;
  assign new_new_n15087__ = ~new_new_n15075__ & ~new_new_n15086__;
  assign new_new_n15088__ = ~new_new_n15068__ & new_new_n15087__;
  assign new_new_n15089__ = ~new_new_n5151__ & ~new_new_n5152__;
  assign new_new_n15090__ = new_new_n5176__ & ~new_new_n15089__;
  assign new_new_n15091__ = ~new_new_n5176__ & new_new_n15089__;
  assign new_new_n15092__ = ~new_new_n15090__ & ~new_new_n15091__;
  assign new_new_n15093__ = ~new_new_n15088__ & new_new_n15092__;
  assign new_new_n15094__ = new_new_n15065__ & new_new_n15067__;
  assign new_new_n15095__ = new_new_n15076__ & new_new_n15085__;
  assign new_new_n15096__ = new_new_n15075__ & ~new_new_n15085__;
  assign new_new_n15097__ = ~new_new_n15092__ & ~new_new_n15096__;
  assign new_new_n15098__ = ~new_new_n15095__ & ~new_new_n15097__;
  assign new_new_n15099__ = ~new_new_n15094__ & new_new_n15098__;
  assign new_new_n15100__ = new_new_n15068__ & ~new_new_n15087__;
  assign new_new_n15101__ = ~new_new_n15099__ & ~new_new_n15100__;
  assign new_new_n15102__ = ~new_new_n15093__ & new_new_n15101__;
  assign new_new_n15103__ = new_new_n5178__ & new_new_n15102__;
  assign new_new_n15104__ = ~new_new_n4900__ & new_new_n6952__;
  assign new_new_n15105__ = ~new_new_n333__ & ~new_new_n3768__;
  assign new_new_n15106__ = ~new_new_n466__ & new_new_n873__;
  assign new_new_n15107__ = ~new_new_n15105__ & ~new_new_n15106__;
  assign new_new_n15108__ = ~new_new_n15104__ & new_new_n15107__;
  assign new_new_n15109__ = ~pi26 & new_new_n15108__;
  assign new_new_n15110__ = pi26 & ~new_new_n15108__;
  assign new_new_n15111__ = ~new_new_n15109__ & ~new_new_n15110__;
  assign new_new_n15112__ = new_new_n5166__ & new_new_n5170__;
  assign new_new_n15113__ = ~new_new_n5154__ & ~new_new_n15112__;
  assign new_new_n15114__ = ~new_new_n5166__ & ~new_new_n5170__;
  assign new_new_n15115__ = ~new_new_n15113__ & ~new_new_n15114__;
  assign new_new_n15116__ = ~new_new_n15111__ & new_new_n15115__;
  assign new_new_n15117__ = new_new_n15111__ & ~new_new_n15115__;
  assign new_new_n15118__ = ~new_new_n4673__ & ~new_new_n4677__;
  assign new_new_n15119__ = new_new_n4648__ & new_new_n4790__;
  assign new_new_n15120__ = ~new_new_n4648__ & ~new_new_n4790__;
  assign new_new_n15121__ = ~new_new_n15119__ & ~new_new_n15120__;
  assign new_new_n15122__ = ~new_new_n15118__ & new_new_n15121__;
  assign new_new_n15123__ = ~new_new_n1959__ & new_new_n4672__;
  assign new_new_n15124__ = new_new_n15118__ & ~new_new_n15123__;
  assign new_new_n15125__ = ~new_new_n15121__ & new_new_n15124__;
  assign new_new_n15126__ = ~new_new_n15122__ & ~new_new_n15125__;
  assign new_new_n15127__ = ~new_new_n15117__ & ~new_new_n15126__;
  assign new_new_n15128__ = ~new_new_n15116__ & ~new_new_n15127__;
  assign new_new_n15129__ = ~new_new_n15103__ & ~new_new_n15128__;
  assign new_new_n15130__ = pi29 & new_new_n4811__;
  assign new_new_n15131__ = new_new_n4144__ & new_new_n15130__;
  assign new_new_n15132__ = pi29 & new_new_n5732__;
  assign new_new_n15133__ = ~pi29 & ~new_new_n4811__;
  assign new_new_n15134__ = ~new_new_n15130__ & ~new_new_n15133__;
  assign new_new_n15135__ = new_new_n4822__ & ~new_new_n15132__;
  assign new_new_n15136__ = ~new_new_n15134__ & new_new_n15135__;
  assign new_new_n15137__ = ~new_new_n4811__ & ~new_new_n4822__;
  assign new_new_n15138__ = new_new_n4814__ & ~new_new_n15130__;
  assign new_new_n15139__ = ~new_new_n15137__ & new_new_n15138__;
  assign new_new_n15140__ = ~new_new_n15131__ & ~new_new_n15136__;
  assign new_new_n15141__ = ~new_new_n15139__ & new_new_n15140__;
  assign new_new_n15142__ = new_new_n4787__ & ~new_new_n15141__;
  assign new_new_n15143__ = ~new_new_n4787__ & ~new_new_n4823__;
  assign new_new_n15144__ = ~new_new_n15134__ & new_new_n15143__;
  assign new_new_n15145__ = new_new_n4787__ & new_new_n4822__;
  assign new_new_n15146__ = ~new_new_n15143__ & ~new_new_n15145__;
  assign new_new_n15147__ = new_new_n15134__ & new_new_n15146__;
  assign new_new_n15148__ = ~new_new_n15144__ & ~new_new_n15147__;
  assign new_new_n15149__ = ~new_new_n15142__ & new_new_n15148__;
  assign new_new_n15150__ = ~new_new_n15129__ & new_new_n15149__;
  assign new_new_n15151__ = ~new_new_n5178__ & ~new_new_n15102__;
  assign new_new_n15152__ = new_new_n15117__ & new_new_n15126__;
  assign new_new_n15153__ = new_new_n15116__ & ~new_new_n15126__;
  assign new_new_n15154__ = new_new_n15149__ & ~new_new_n15153__;
  assign new_new_n15155__ = ~new_new_n15152__ & ~new_new_n15154__;
  assign new_new_n15156__ = ~new_new_n15151__ & ~new_new_n15155__;
  assign new_new_n15157__ = new_new_n15103__ & new_new_n15128__;
  assign new_new_n15158__ = ~new_new_n15156__ & ~new_new_n15157__;
  assign new_new_n15159__ = ~new_new_n15150__ & new_new_n15158__;
  assign new_new_n15160__ = ~new_new_n4897__ & ~new_new_n15159__;
  assign new_new_n15161__ = ~new_new_n4126__ & ~new_new_n4181__;
  assign new_new_n15162__ = new_new_n4059__ & ~new_new_n15161__;
  assign new_new_n15163__ = ~new_new_n4059__ & new_new_n15161__;
  assign new_new_n15164__ = ~new_new_n15162__ & ~new_new_n15163__;
  assign new_new_n15165__ = ~new_new_n4210__ & ~new_new_n4221__;
  assign new_new_n15166__ = new_new_n5126__ & new_new_n15165__;
  assign new_new_n15167__ = ~new_new_n5126__ & ~new_new_n15165__;
  assign new_new_n15168__ = ~new_new_n15166__ & ~new_new_n15167__;
  assign new_new_n15169__ = ~new_new_n466__ & new_new_n15168__;
  assign new_new_n15170__ = ~new_new_n4212__ & ~new_new_n4215__;
  assign new_new_n15171__ = ~new_new_n3768__ & new_new_n15170__;
  assign new_new_n15172__ = ~new_new_n15169__ & ~new_new_n15171__;
  assign new_new_n15173__ = ~pi29 & new_new_n15172__;
  assign new_new_n15174__ = pi29 & ~new_new_n15172__;
  assign new_new_n15175__ = ~new_new_n15173__ & ~new_new_n15174__;
  assign new_new_n15176__ = new_new_n4889__ & ~new_new_n15175__;
  assign new_new_n15177__ = ~new_new_n4889__ & new_new_n15175__;
  assign new_new_n15178__ = ~new_new_n15176__ & ~new_new_n15177__;
  assign new_new_n15179__ = new_new_n15164__ & new_new_n15178__;
  assign new_new_n15180__ = ~new_new_n15164__ & ~new_new_n15178__;
  assign new_new_n15181__ = ~new_new_n15179__ & ~new_new_n15180__;
  assign new_new_n15182__ = ~new_new_n15160__ & ~new_new_n15181__;
  assign new_new_n15183__ = ~new_new_n4845__ & ~new_new_n15182__;
  assign new_new_n15184__ = ~new_new_n4777__ & new_new_n15183__;
  assign new_new_n15185__ = new_new_n4897__ & new_new_n15159__;
  assign new_new_n15186__ = ~new_new_n4845__ & new_new_n15181__;
  assign new_new_n15187__ = new_new_n4777__ & ~new_new_n15186__;
  assign new_new_n15188__ = ~new_new_n15185__ & ~new_new_n15187__;
  assign new_new_n15189__ = ~new_new_n15160__ & ~new_new_n15188__;
  assign new_new_n15190__ = new_new_n15181__ & ~new_new_n15189__;
  assign new_new_n15191__ = ~new_new_n15183__ & ~new_new_n15188__;
  assign new_new_n15192__ = ~new_new_n4833__ & new_new_n4844__;
  assign new_new_n15193__ = ~new_new_n15191__ & new_new_n15192__;
  assign new_new_n15194__ = ~new_new_n15184__ & ~new_new_n15190__;
  assign new_new_n15195__ = ~new_new_n15193__ & new_new_n15194__;
  assign new_new_n15196__ = new_new_n4208__ & new_new_n15195__;
  assign new_new_n15197__ = ~new_new_n4208__ & ~new_new_n15195__;
  assign new_new_n15198__ = ~new_new_n15164__ & ~new_new_n15177__;
  assign new_new_n15199__ = ~new_new_n15176__ & ~new_new_n15198__;
  assign new_new_n15200__ = ~new_new_n15197__ & ~new_new_n15199__;
  assign new_new_n15201__ = ~new_new_n15196__ & ~new_new_n15200__;
  assign new_new_n15202__ = ~new_new_n3824__ & ~new_new_n4193__;
  assign new_new_n15203__ = ~new_new_n4195__ & ~new_new_n15202__;
  assign new_new_n15204__ = new_new_n15201__ & new_new_n15203__;
  assign new_new_n15205__ = ~new_new_n15201__ & ~new_new_n15203__;
  assign new_new_n15206__ = ~new_new_n15204__ & ~new_new_n15205__;
  assign new_new_n15207__ = new_new_n4167__ & new_new_n4177__;
  assign new_new_n15208__ = ~new_new_n3888__ & new_new_n15207__;
  assign new_new_n15209__ = ~new_new_n4179__ & ~new_new_n15208__;
  assign new_new_n15210__ = new_new_n15206__ & new_new_n15209__;
  assign new_new_n15211__ = new_new_n3888__ & ~new_new_n15207__;
  assign new_new_n15212__ = ~new_new_n4178__ & ~new_new_n15211__;
  assign new_new_n15213__ = new_new_n15204__ & ~new_new_n15212__;
  assign new_new_n15214__ = new_new_n15205__ & new_new_n15212__;
  assign new_new_n15215__ = ~new_new_n15213__ & ~new_new_n15214__;
  assign new_new_n15216__ = ~new_new_n15210__ & new_new_n15215__;
  assign new_new_n15217__ = ~new_new_n3884__ & ~new_new_n15216__;
  assign new_new_n15218__ = new_new_n4167__ & new_new_n15203__;
  assign new_new_n15219__ = new_new_n15201__ & new_new_n15218__;
  assign new_new_n15220__ = new_new_n4177__ & new_new_n15219__;
  assign new_new_n15221__ = ~new_new_n4167__ & ~new_new_n15203__;
  assign new_new_n15222__ = ~new_new_n15201__ & new_new_n15221__;
  assign new_new_n15223__ = new_new_n4177__ & ~new_new_n15222__;
  assign new_new_n15224__ = ~new_new_n15201__ & ~new_new_n15218__;
  assign new_new_n15225__ = ~new_new_n15221__ & ~new_new_n15224__;
  assign new_new_n15226__ = new_new_n3888__ & ~new_new_n15223__;
  assign new_new_n15227__ = ~new_new_n15225__ & new_new_n15226__;
  assign new_new_n15228__ = new_new_n4177__ & new_new_n15225__;
  assign new_new_n15229__ = ~new_new_n15219__ & ~new_new_n15228__;
  assign new_new_n15230__ = ~new_new_n3888__ & ~new_new_n15229__;
  assign new_new_n15231__ = ~new_new_n4177__ & ~new_new_n15201__;
  assign new_new_n15232__ = new_new_n15221__ & new_new_n15231__;
  assign new_new_n15233__ = ~new_new_n15220__ & ~new_new_n15232__;
  assign new_new_n15234__ = ~new_new_n15227__ & new_new_n15233__;
  assign new_new_n15235__ = ~new_new_n15230__ & new_new_n15234__;
  assign new_new_n15236__ = new_new_n3884__ & ~new_new_n15235__;
  assign new_new_n15237__ = ~new_new_n15217__ & ~new_new_n15236__;
  assign new_new_n15238__ = ~new_new_n4178__ & ~new_new_n15207__;
  assign new_new_n15239__ = new_new_n3888__ & ~new_new_n15238__;
  assign new_new_n15240__ = ~new_new_n3888__ & new_new_n15238__;
  assign new_new_n15241__ = ~new_new_n15239__ & ~new_new_n15240__;
  assign new_new_n15242__ = new_new_n15206__ & new_new_n15241__;
  assign new_new_n15243__ = ~new_new_n15206__ & ~new_new_n15241__;
  assign new_new_n15244__ = ~new_new_n15242__ & ~new_new_n15243__;
  assign new_new_n15245__ = ~new_new_n15196__ & ~new_new_n15197__;
  assign new_new_n15246__ = new_new_n15199__ & ~new_new_n15245__;
  assign new_new_n15247__ = ~new_new_n15199__ & new_new_n15245__;
  assign new_new_n15248__ = ~new_new_n15246__ & ~new_new_n15247__;
  assign new_new_n15249__ = ~new_new_n15244__ & new_new_n15248__;
  assign new_new_n15250__ = new_new_n15128__ & ~new_new_n15151__;
  assign new_new_n15251__ = ~new_new_n15129__ & ~new_new_n15250__;
  assign new_new_n15252__ = ~new_new_n15103__ & ~new_new_n15151__;
  assign new_new_n15253__ = ~new_new_n15152__ & ~new_new_n15153__;
  assign new_new_n15254__ = new_new_n15252__ & new_new_n15253__;
  assign new_new_n15255__ = ~new_new_n15251__ & ~new_new_n15254__;
  assign new_new_n15256__ = ~new_new_n15149__ & ~new_new_n15255__;
  assign new_new_n15257__ = new_new_n15103__ & ~new_new_n15115__;
  assign new_new_n15258__ = new_new_n15111__ & new_new_n15257__;
  assign new_new_n15259__ = ~new_new_n15103__ & new_new_n15115__;
  assign new_new_n15260__ = new_new_n15111__ & ~new_new_n15151__;
  assign new_new_n15261__ = ~new_new_n15259__ & new_new_n15260__;
  assign new_new_n15262__ = ~new_new_n15257__ & ~new_new_n15261__;
  assign new_new_n15263__ = new_new_n15126__ & ~new_new_n15262__;
  assign new_new_n15264__ = ~new_new_n15117__ & new_new_n15151__;
  assign new_new_n15265__ = ~new_new_n15111__ & new_new_n15259__;
  assign new_new_n15266__ = ~new_new_n15264__ & ~new_new_n15265__;
  assign new_new_n15267__ = ~new_new_n15126__ & ~new_new_n15266__;
  assign new_new_n15268__ = new_new_n15116__ & new_new_n15151__;
  assign new_new_n15269__ = ~new_new_n15258__ & ~new_new_n15268__;
  assign new_new_n15270__ = ~new_new_n15263__ & new_new_n15269__;
  assign new_new_n15271__ = ~new_new_n15267__ & new_new_n15270__;
  assign new_new_n15272__ = new_new_n15149__ & ~new_new_n15271__;
  assign new_new_n15273__ = ~new_new_n15256__ & ~new_new_n15272__;
  assign new_new_n15274__ = new_new_n4844__ & ~new_new_n4897__;
  assign new_new_n15275__ = ~new_new_n4844__ & new_new_n4897__;
  assign new_new_n15276__ = ~new_new_n15274__ & ~new_new_n15275__;
  assign new_new_n15277__ = new_new_n4833__ & new_new_n15159__;
  assign new_new_n15278__ = ~new_new_n4833__ & ~new_new_n15159__;
  assign new_new_n15279__ = ~new_new_n15277__ & ~new_new_n15278__;
  assign new_new_n15280__ = ~new_new_n4777__ & new_new_n15279__;
  assign new_new_n15281__ = new_new_n4777__ & ~new_new_n15279__;
  assign new_new_n15282__ = ~new_new_n15280__ & ~new_new_n15281__;
  assign new_new_n15283__ = new_new_n15276__ & new_new_n15282__;
  assign new_new_n15284__ = ~new_new_n15276__ & ~new_new_n15282__;
  assign new_new_n15285__ = ~new_new_n15283__ & ~new_new_n15284__;
  assign new_new_n15286__ = ~new_new_n15248__ & new_new_n15285__;
  assign new_new_n15287__ = new_new_n4777__ & new_new_n15275__;
  assign new_new_n15288__ = ~new_new_n4777__ & new_new_n15274__;
  assign new_new_n15289__ = ~new_new_n15287__ & ~new_new_n15288__;
  assign new_new_n15290__ = new_new_n15279__ & new_new_n15289__;
  assign new_new_n15291__ = new_new_n4777__ & ~new_new_n15274__;
  assign new_new_n15292__ = ~new_new_n15275__ & ~new_new_n15291__;
  assign new_new_n15293__ = new_new_n15278__ & ~new_new_n15292__;
  assign new_new_n15294__ = new_new_n15277__ & new_new_n15292__;
  assign new_new_n15295__ = ~new_new_n15293__ & ~new_new_n15294__;
  assign new_new_n15296__ = ~new_new_n15290__ & new_new_n15295__;
  assign new_new_n15297__ = ~new_new_n15181__ & ~new_new_n15296__;
  assign new_new_n15298__ = ~new_new_n4833__ & new_new_n15160__;
  assign new_new_n15299__ = new_new_n4844__ & new_new_n15298__;
  assign new_new_n15300__ = ~new_new_n4833__ & ~new_new_n15185__;
  assign new_new_n15301__ = ~new_new_n15160__ & ~new_new_n15300__;
  assign new_new_n15302__ = ~new_new_n4844__ & new_new_n15301__;
  assign new_new_n15303__ = new_new_n4833__ & new_new_n15185__;
  assign new_new_n15304__ = ~new_new_n15302__ & ~new_new_n15303__;
  assign new_new_n15305__ = new_new_n4777__ & ~new_new_n15304__;
  assign new_new_n15306__ = ~new_new_n4844__ & ~new_new_n15298__;
  assign new_new_n15307__ = ~new_new_n4777__ & ~new_new_n15301__;
  assign new_new_n15308__ = ~new_new_n15306__ & new_new_n15307__;
  assign new_new_n15309__ = new_new_n4845__ & new_new_n15185__;
  assign new_new_n15310__ = ~new_new_n15299__ & ~new_new_n15309__;
  assign new_new_n15311__ = ~new_new_n15308__ & new_new_n15310__;
  assign new_new_n15312__ = ~new_new_n15305__ & new_new_n15311__;
  assign new_new_n15313__ = new_new_n15181__ & ~new_new_n15312__;
  assign new_new_n15314__ = ~new_new_n15297__ & ~new_new_n15313__;
  assign new_new_n15315__ = ~new_new_n15116__ & ~new_new_n15117__;
  assign new_new_n15316__ = ~new_new_n15252__ & new_new_n15315__;
  assign new_new_n15317__ = new_new_n15252__ & ~new_new_n15315__;
  assign new_new_n15318__ = ~new_new_n15316__ & ~new_new_n15317__;
  assign new_new_n15319__ = new_new_n15126__ & new_new_n15318__;
  assign new_new_n15320__ = ~new_new_n15126__ & ~new_new_n15318__;
  assign new_new_n15321__ = ~new_new_n15319__ & ~new_new_n15320__;
  assign new_new_n15322__ = ~new_new_n15314__ & ~new_new_n15321__;
  assign new_new_n15323__ = ~new_new_n15286__ & ~new_new_n15322__;
  assign new_new_n15324__ = ~new_new_n15273__ & ~new_new_n15323__;
  assign new_new_n15325__ = ~new_new_n15248__ & ~new_new_n15314__;
  assign new_new_n15326__ = new_new_n15070__ & new_new_n15094__;
  assign new_new_n15327__ = ~new_new_n15070__ & ~new_new_n15094__;
  assign new_new_n15328__ = ~new_new_n15068__ & new_new_n15074__;
  assign new_new_n15329__ = ~new_new_n15327__ & new_new_n15328__;
  assign new_new_n15330__ = ~new_new_n15326__ & ~new_new_n15329__;
  assign new_new_n15331__ = new_new_n15085__ & ~new_new_n15330__;
  assign new_new_n15332__ = new_new_n15076__ & new_new_n15094__;
  assign new_new_n15333__ = new_new_n15068__ & new_new_n15075__;
  assign new_new_n15334__ = new_new_n15068__ & ~new_new_n15076__;
  assign new_new_n15335__ = new_new_n15075__ & ~new_new_n15094__;
  assign new_new_n15336__ = ~new_new_n15334__ & ~new_new_n15335__;
  assign new_new_n15337__ = ~new_new_n15085__ & ~new_new_n15336__;
  assign new_new_n15338__ = new_new_n15092__ & ~new_new_n15332__;
  assign new_new_n15339__ = ~new_new_n15333__ & new_new_n15338__;
  assign new_new_n15340__ = ~new_new_n15337__ & new_new_n15339__;
  assign new_new_n15341__ = ~new_new_n15331__ & new_new_n15340__;
  assign new_new_n15342__ = ~new_new_n15087__ & ~new_new_n15094__;
  assign new_new_n15343__ = ~new_new_n15088__ & ~new_new_n15342__;
  assign new_new_n15344__ = ~new_new_n15068__ & ~new_new_n15094__;
  assign new_new_n15345__ = ~new_new_n15095__ & ~new_new_n15096__;
  assign new_new_n15346__ = new_new_n15344__ & new_new_n15345__;
  assign new_new_n15347__ = ~new_new_n15092__ & ~new_new_n15343__;
  assign new_new_n15348__ = ~new_new_n15346__ & new_new_n15347__;
  assign new_new_n15349__ = ~new_new_n15341__ & ~new_new_n15348__;
  assign new_new_n15350__ = new_new_n15321__ & new_new_n15349__;
  assign new_new_n15351__ = ~new_new_n14939__ & ~new_new_n15047__;
  assign new_new_n15352__ = new_new_n14939__ & new_new_n15047__;
  assign new_new_n15353__ = ~new_new_n15351__ & ~new_new_n15352__;
  assign new_new_n15354__ = new_new_n5207__ & new_new_n15045__;
  assign new_new_n15355__ = ~new_new_n5207__ & ~new_new_n15045__;
  assign new_new_n15356__ = ~new_new_n15354__ & ~new_new_n15355__;
  assign new_new_n15357__ = new_new_n15353__ & ~new_new_n15356__;
  assign new_new_n15358__ = ~new_new_n15353__ & new_new_n15356__;
  assign new_new_n15359__ = ~new_new_n15357__ & ~new_new_n15358__;
  assign new_new_n15360__ = new_new_n15055__ & new_new_n15359__;
  assign new_new_n15361__ = ~new_new_n15055__ & ~new_new_n15359__;
  assign new_new_n15362__ = ~new_new_n15360__ & ~new_new_n15361__;
  assign new_new_n15363__ = new_new_n15055__ & new_new_n15354__;
  assign new_new_n15364__ = ~new_new_n15055__ & new_new_n15355__;
  assign new_new_n15365__ = ~new_new_n15363__ & ~new_new_n15364__;
  assign new_new_n15366__ = new_new_n15353__ & new_new_n15365__;
  assign new_new_n15367__ = new_new_n15055__ & ~new_new_n15355__;
  assign new_new_n15368__ = ~new_new_n15354__ & ~new_new_n15367__;
  assign new_new_n15369__ = new_new_n15352__ & ~new_new_n15368__;
  assign new_new_n15370__ = new_new_n15351__ & new_new_n15368__;
  assign new_new_n15371__ = ~new_new_n15369__ & ~new_new_n15370__;
  assign new_new_n15372__ = ~new_new_n15366__ & new_new_n15371__;
  assign new_new_n15373__ = ~new_new_n15043__ & ~new_new_n15372__;
  assign new_new_n15374__ = ~new_new_n14939__ & new_new_n15050__;
  assign new_new_n15375__ = new_new_n5207__ & new_new_n15374__;
  assign new_new_n15376__ = new_new_n14939__ & ~new_new_n15050__;
  assign new_new_n15377__ = ~new_new_n15048__ & ~new_new_n15376__;
  assign new_new_n15378__ = new_new_n5207__ & new_new_n15377__;
  assign new_new_n15379__ = ~new_new_n15374__ & ~new_new_n15378__;
  assign new_new_n15380__ = new_new_n15055__ & ~new_new_n15379__;
  assign new_new_n15381__ = new_new_n14939__ & new_new_n15048__;
  assign new_new_n15382__ = new_new_n5207__ & ~new_new_n15381__;
  assign new_new_n15383__ = ~new_new_n15055__ & ~new_new_n15377__;
  assign new_new_n15384__ = ~new_new_n15382__ & new_new_n15383__;
  assign new_new_n15385__ = new_new_n14940__ & new_new_n15048__;
  assign new_new_n15386__ = ~new_new_n15375__ & ~new_new_n15385__;
  assign new_new_n15387__ = ~new_new_n15384__ & new_new_n15386__;
  assign new_new_n15388__ = ~new_new_n15380__ & new_new_n15387__;
  assign new_new_n15389__ = new_new_n15043__ & ~new_new_n15388__;
  assign new_new_n15390__ = ~new_new_n15373__ & ~new_new_n15389__;
  assign new_new_n15391__ = new_new_n15349__ & ~new_new_n15390__;
  assign new_new_n15392__ = ~new_new_n15075__ & ~new_new_n15076__;
  assign new_new_n15393__ = new_new_n15085__ & ~new_new_n15392__;
  assign new_new_n15394__ = ~new_new_n15085__ & new_new_n15392__;
  assign new_new_n15395__ = ~new_new_n15393__ & ~new_new_n15394__;
  assign new_new_n15396__ = new_new_n15344__ & new_new_n15395__;
  assign new_new_n15397__ = ~new_new_n15344__ & ~new_new_n15395__;
  assign new_new_n15398__ = ~new_new_n15396__ & ~new_new_n15397__;
  assign new_new_n15399__ = new_new_n15321__ & new_new_n15398__;
  assign new_new_n15400__ = new_new_n14788__ & ~new_new_n14916__;
  assign new_new_n15401__ = new_new_n14918__ & new_new_n15400__;
  assign new_new_n15402__ = new_new_n5966__ & new_new_n15401__;
  assign new_new_n15403__ = ~new_new_n14788__ & new_new_n14916__;
  assign new_new_n15404__ = ~new_new_n14918__ & new_new_n15403__;
  assign new_new_n15405__ = ~new_new_n14788__ & ~new_new_n14928__;
  assign new_new_n15406__ = ~new_new_n14919__ & ~new_new_n15405__;
  assign new_new_n15407__ = ~new_new_n5966__ & ~new_new_n15406__;
  assign new_new_n15408__ = ~new_new_n14927__ & ~new_new_n15404__;
  assign new_new_n15409__ = ~new_new_n15407__ & new_new_n15408__;
  assign new_new_n15410__ = new_new_n5966__ & new_new_n15406__;
  assign new_new_n15411__ = new_new_n14927__ & ~new_new_n15401__;
  assign new_new_n15412__ = ~new_new_n15410__ & new_new_n15411__;
  assign new_new_n15413__ = ~new_new_n15409__ & ~new_new_n15412__;
  assign new_new_n15414__ = ~new_new_n5966__ & ~new_new_n14918__;
  assign new_new_n15415__ = new_new_n15403__ & new_new_n15414__;
  assign new_new_n15416__ = ~new_new_n14912__ & ~new_new_n15415__;
  assign new_new_n15417__ = ~new_new_n15402__ & new_new_n15416__;
  assign new_new_n15418__ = ~new_new_n15413__ & new_new_n15417__;
  assign new_new_n15419__ = new_new_n5966__ & new_new_n14918__;
  assign new_new_n15420__ = ~new_new_n14927__ & ~new_new_n15419__;
  assign new_new_n15421__ = ~new_new_n15414__ & ~new_new_n15420__;
  assign new_new_n15422__ = new_new_n15403__ & new_new_n15421__;
  assign new_new_n15423__ = ~new_new_n14927__ & new_new_n15414__;
  assign new_new_n15424__ = ~new_new_n15400__ & ~new_new_n15403__;
  assign new_new_n15425__ = new_new_n14927__ & new_new_n15419__;
  assign new_new_n15426__ = ~new_new_n15423__ & ~new_new_n15425__;
  assign new_new_n15427__ = new_new_n15424__ & new_new_n15426__;
  assign new_new_n15428__ = new_new_n15400__ & ~new_new_n15421__;
  assign new_new_n15429__ = new_new_n14912__ & ~new_new_n15422__;
  assign new_new_n15430__ = ~new_new_n15428__ & new_new_n15429__;
  assign new_new_n15431__ = ~new_new_n15427__ & new_new_n15430__;
  assign new_new_n15432__ = ~new_new_n15418__ & ~new_new_n15431__;
  assign new_new_n15433__ = ~new_new_n15414__ & ~new_new_n15419__;
  assign new_new_n15434__ = new_new_n14927__ & ~new_new_n15433__;
  assign new_new_n15435__ = ~new_new_n14927__ & new_new_n15433__;
  assign new_new_n15436__ = ~new_new_n15434__ & ~new_new_n15435__;
  assign new_new_n15437__ = new_new_n15424__ & new_new_n15436__;
  assign new_new_n15438__ = ~new_new_n15424__ & ~new_new_n15436__;
  assign new_new_n15439__ = ~new_new_n15437__ & ~new_new_n15438__;
  assign new_new_n15440__ = ~new_new_n15432__ & ~new_new_n15439__;
  assign new_new_n15441__ = ~new_new_n14738__ & ~new_new_n14781__;
  assign new_new_n15442__ = ~new_new_n14739__ & ~new_new_n15441__;
  assign new_new_n15443__ = ~new_new_n14671__ & ~new_new_n14781__;
  assign new_new_n15444__ = ~new_new_n14780__ & ~new_new_n14782__;
  assign new_new_n15445__ = new_new_n15443__ & new_new_n15444__;
  assign new_new_n15446__ = ~new_new_n15442__ & ~new_new_n15445__;
  assign new_new_n15447__ = ~new_new_n14778__ & ~new_new_n15446__;
  assign new_new_n15448__ = new_new_n14726__ & new_new_n14781__;
  assign new_new_n15449__ = new_new_n14724__ & new_new_n14781__;
  assign new_new_n15450__ = ~new_new_n14724__ & ~new_new_n14781__;
  assign new_new_n15451__ = ~new_new_n14671__ & ~new_new_n14673__;
  assign new_new_n15452__ = ~new_new_n15450__ & new_new_n15451__;
  assign new_new_n15453__ = ~new_new_n15449__ & ~new_new_n15452__;
  assign new_new_n15454__ = new_new_n14736__ & ~new_new_n15453__;
  assign new_new_n15455__ = new_new_n14671__ & new_new_n14725__;
  assign new_new_n15456__ = new_new_n14671__ & ~new_new_n14726__;
  assign new_new_n15457__ = new_new_n14725__ & ~new_new_n14781__;
  assign new_new_n15458__ = ~new_new_n15456__ & ~new_new_n15457__;
  assign new_new_n15459__ = ~new_new_n14736__ & ~new_new_n15458__;
  assign new_new_n15460__ = ~new_new_n15448__ & ~new_new_n15455__;
  assign new_new_n15461__ = ~new_new_n15459__ & new_new_n15460__;
  assign new_new_n15462__ = ~new_new_n15454__ & new_new_n15461__;
  assign new_new_n15463__ = new_new_n14778__ & ~new_new_n15462__;
  assign new_new_n15464__ = ~new_new_n15447__ & ~new_new_n15463__;
  assign new_new_n15465__ = ~new_new_n14725__ & ~new_new_n14726__;
  assign new_new_n15466__ = new_new_n14736__ & ~new_new_n15465__;
  assign new_new_n15467__ = ~new_new_n14736__ & new_new_n15465__;
  assign new_new_n15468__ = ~new_new_n15466__ & ~new_new_n15467__;
  assign new_new_n15469__ = new_new_n15443__ & new_new_n15468__;
  assign new_new_n15470__ = ~new_new_n15443__ & ~new_new_n15468__;
  assign new_new_n15471__ = ~new_new_n15469__ & ~new_new_n15470__;
  assign new_new_n15472__ = ~new_new_n15439__ & ~new_new_n15471__;
  assign new_new_n15473__ = ~new_new_n15464__ & ~new_new_n15472__;
  assign new_new_n15474__ = ~new_new_n15440__ & new_new_n15473__;
  assign new_new_n15475__ = new_new_n15432__ & new_new_n15439__;
  assign new_new_n15476__ = ~new_new_n6947__ & new_new_n14644__;
  assign new_new_n15477__ = new_new_n6947__ & ~new_new_n14644__;
  assign new_new_n15478__ = ~new_new_n15476__ & ~new_new_n15477__;
  assign new_new_n15479__ = ~new_new_n14636__ & ~new_new_n14642__;
  assign new_new_n15480__ = new_new_n14636__ & new_new_n14642__;
  assign new_new_n15481__ = ~new_new_n15479__ & ~new_new_n15480__;
  assign new_new_n15482__ = new_new_n15478__ & ~new_new_n15481__;
  assign new_new_n15483__ = ~new_new_n15478__ & new_new_n15481__;
  assign new_new_n15484__ = ~new_new_n15482__ & ~new_new_n15483__;
  assign new_new_n15485__ = new_new_n14657__ & new_new_n15484__;
  assign new_new_n15486__ = ~new_new_n14657__ & ~new_new_n15484__;
  assign new_new_n15487__ = ~new_new_n15485__ & ~new_new_n15486__;
  assign new_new_n15488__ = new_new_n8316__ & new_new_n8465__;
  assign new_new_n15489__ = new_new_n8460__ & new_new_n15488__;
  assign new_new_n15490__ = new_new_n8314__ & ~new_new_n14577__;
  assign new_new_n15491__ = ~new_new_n8314__ & new_new_n14577__;
  assign new_new_n15492__ = ~new_new_n15490__ & ~new_new_n15491__;
  assign new_new_n15493__ = ~new_new_n8316__ & ~new_new_n8465__;
  assign new_new_n15494__ = ~new_new_n8460__ & new_new_n15493__;
  assign new_new_n15495__ = ~new_new_n15489__ & ~new_new_n15494__;
  assign new_new_n15496__ = new_new_n15492__ & new_new_n15495__;
  assign new_new_n15497__ = ~new_new_n8460__ & ~new_new_n15488__;
  assign new_new_n15498__ = ~new_new_n15493__ & ~new_new_n15497__;
  assign new_new_n15499__ = new_new_n15490__ & ~new_new_n15498__;
  assign new_new_n15500__ = new_new_n15491__ & new_new_n15498__;
  assign new_new_n15501__ = ~new_new_n15499__ & ~new_new_n15500__;
  assign new_new_n15502__ = ~new_new_n15496__ & new_new_n15501__;
  assign new_new_n15503__ = new_new_n8444__ & ~new_new_n15502__;
  assign new_new_n15504__ = ~new_new_n8314__ & new_new_n14578__;
  assign new_new_n15505__ = ~new_new_n8316__ & new_new_n15504__;
  assign new_new_n15506__ = ~new_new_n8465__ & ~new_new_n15490__;
  assign new_new_n15507__ = ~new_new_n15491__ & ~new_new_n15506__;
  assign new_new_n15508__ = ~new_new_n8316__ & ~new_new_n15507__;
  assign new_new_n15509__ = ~new_new_n15504__ & ~new_new_n15508__;
  assign new_new_n15510__ = ~new_new_n8460__ & ~new_new_n15509__;
  assign new_new_n15511__ = new_new_n8316__ & new_new_n15507__;
  assign new_new_n15512__ = new_new_n8314__ & new_new_n14581__;
  assign new_new_n15513__ = ~new_new_n15511__ & ~new_new_n15512__;
  assign new_new_n15514__ = new_new_n8460__ & ~new_new_n15513__;
  assign new_new_n15515__ = new_new_n15488__ & new_new_n15490__;
  assign new_new_n15516__ = ~new_new_n15505__ & ~new_new_n15515__;
  assign new_new_n15517__ = ~new_new_n15510__ & new_new_n15516__;
  assign new_new_n15518__ = ~new_new_n15514__ & new_new_n15517__;
  assign new_new_n15519__ = ~new_new_n8444__ & ~new_new_n15518__;
  assign new_new_n15520__ = ~new_new_n15503__ & ~new_new_n15519__;
  assign new_new_n15521__ = ~new_new_n14631__ & ~new_new_n14632__;
  assign new_new_n15522__ = new_new_n14634__ & ~new_new_n15521__;
  assign new_new_n15523__ = ~new_new_n14634__ & new_new_n15521__;
  assign new_new_n15524__ = ~new_new_n15522__ & ~new_new_n15523__;
  assign new_new_n15525__ = new_new_n15520__ & new_new_n15524__;
  assign new_new_n15526__ = new_new_n15487__ & ~new_new_n15525__;
  assign new_new_n15527__ = ~new_new_n15488__ & ~new_new_n15493__;
  assign new_new_n15528__ = ~new_new_n8460__ & new_new_n15492__;
  assign new_new_n15529__ = new_new_n8460__ & ~new_new_n15492__;
  assign new_new_n15530__ = ~new_new_n15528__ & ~new_new_n15529__;
  assign new_new_n15531__ = new_new_n15527__ & new_new_n15530__;
  assign new_new_n15532__ = ~new_new_n15527__ & ~new_new_n15530__;
  assign new_new_n15533__ = ~new_new_n15531__ & ~new_new_n15532__;
  assign new_new_n15534__ = new_new_n15520__ & ~new_new_n15533__;
  assign new_new_n15535__ = ~new_new_n15524__ & ~new_new_n15534__;
  assign new_new_n15536__ = ~new_new_n15526__ & ~new_new_n15535__;
  assign new_new_n15537__ = new_new_n14554__ & ~new_new_n14561__;
  assign new_new_n15538__ = ~new_new_n14555__ & ~new_new_n15537__;
  assign new_new_n15539__ = ~new_new_n14532__ & ~new_new_n14561__;
  assign new_new_n15540__ = ~new_new_n14562__ & ~new_new_n14563__;
  assign new_new_n15541__ = new_new_n15539__ & new_new_n15540__;
  assign new_new_n15542__ = ~new_new_n15538__ & ~new_new_n15541__;
  assign new_new_n15543__ = ~new_new_n14559__ & ~new_new_n15542__;
  assign new_new_n15544__ = new_new_n14534__ & new_new_n14561__;
  assign new_new_n15545__ = new_new_n14538__ & new_new_n15544__;
  assign new_new_n15546__ = ~new_new_n14534__ & ~new_new_n14561__;
  assign new_new_n15547__ = ~new_new_n14532__ & new_new_n14538__;
  assign new_new_n15548__ = ~new_new_n15546__ & new_new_n15547__;
  assign new_new_n15549__ = ~new_new_n15544__ & ~new_new_n15548__;
  assign new_new_n15550__ = ~new_new_n14552__ & ~new_new_n15549__;
  assign new_new_n15551__ = new_new_n14532__ & new_new_n14540__;
  assign new_new_n15552__ = new_new_n14532__ & ~new_new_n14539__;
  assign new_new_n15553__ = ~new_new_n14538__ & new_new_n15546__;
  assign new_new_n15554__ = ~new_new_n15552__ & ~new_new_n15553__;
  assign new_new_n15555__ = new_new_n14552__ & ~new_new_n15554__;
  assign new_new_n15556__ = ~new_new_n15545__ & ~new_new_n15551__;
  assign new_new_n15557__ = ~new_new_n15550__ & new_new_n15556__;
  assign new_new_n15558__ = ~new_new_n15555__ & new_new_n15557__;
  assign new_new_n15559__ = new_new_n14559__ & ~new_new_n15558__;
  assign new_new_n15560__ = ~new_new_n15543__ & ~new_new_n15559__;
  assign new_new_n15561__ = ~new_new_n14524__ & ~new_new_n14525__;
  assign new_new_n15562__ = new_new_n14529__ & ~new_new_n15561__;
  assign new_new_n15563__ = ~new_new_n14529__ & new_new_n15561__;
  assign new_new_n15564__ = ~new_new_n15562__ & ~new_new_n15563__;
  assign new_new_n15565__ = ~new_new_n15560__ & ~new_new_n15564__;
  assign new_new_n15566__ = ~new_new_n14539__ & ~new_new_n14540__;
  assign new_new_n15567__ = new_new_n15539__ & ~new_new_n15566__;
  assign new_new_n15568__ = ~new_new_n15539__ & new_new_n15566__;
  assign new_new_n15569__ = ~new_new_n15567__ & ~new_new_n15568__;
  assign new_new_n15570__ = new_new_n14552__ & new_new_n15569__;
  assign new_new_n15571__ = ~new_new_n14552__ & ~new_new_n15569__;
  assign new_new_n15572__ = ~new_new_n15570__ & ~new_new_n15571__;
  assign new_new_n15573__ = ~new_new_n15565__ & new_new_n15572__;
  assign new_new_n15574__ = new_new_n15560__ & new_new_n15564__;
  assign new_new_n15575__ = ~new_new_n14463__ & ~new_new_n14497__;
  assign new_new_n15576__ = ~new_new_n14473__ & ~new_new_n14474__;
  assign new_new_n15577__ = new_new_n14487__ & ~new_new_n15576__;
  assign new_new_n15578__ = ~new_new_n14487__ & new_new_n15576__;
  assign new_new_n15579__ = ~new_new_n15577__ & ~new_new_n15578__;
  assign new_new_n15580__ = new_new_n15575__ & new_new_n15579__;
  assign new_new_n15581__ = ~new_new_n15575__ & ~new_new_n15579__;
  assign new_new_n15582__ = ~new_new_n15580__ & ~new_new_n15581__;
  assign new_new_n15583__ = ~new_new_n11404__ & ~new_new_n14504__;
  assign new_new_n15584__ = ~new_new_n11405__ & ~new_new_n15583__;
  assign new_new_n15585__ = new_new_n10723__ & ~new_new_n14508__;
  assign new_new_n15586__ = ~new_new_n14512__ & ~new_new_n15585__;
  assign new_new_n15587__ = ~new_new_n15584__ & ~new_new_n15586__;
  assign new_new_n15588__ = new_new_n10723__ & new_new_n15583__;
  assign new_new_n15589__ = new_new_n11404__ & new_new_n14504__;
  assign new_new_n15590__ = new_new_n10723__ & ~new_new_n15589__;
  assign new_new_n15591__ = ~new_new_n15583__ & ~new_new_n15590__;
  assign new_new_n15592__ = ~new_new_n14508__ & ~new_new_n15591__;
  assign new_new_n15593__ = new_new_n11465__ & ~new_new_n15588__;
  assign new_new_n15594__ = ~new_new_n15592__ & new_new_n15593__;
  assign new_new_n15595__ = ~new_new_n10723__ & new_new_n15589__;
  assign new_new_n15596__ = new_new_n14508__ & new_new_n15591__;
  assign new_new_n15597__ = ~new_new_n11465__ & ~new_new_n15595__;
  assign new_new_n15598__ = ~new_new_n15596__ & new_new_n15597__;
  assign new_new_n15599__ = ~new_new_n15594__ & ~new_new_n15598__;
  assign new_new_n15600__ = ~new_new_n11448__ & ~new_new_n15587__;
  assign new_new_n15601__ = ~new_new_n15599__ & new_new_n15600__;
  assign new_new_n15602__ = ~new_new_n10723__ & new_new_n14508__;
  assign new_new_n15603__ = ~new_new_n11465__ & ~new_new_n15585__;
  assign new_new_n15604__ = ~new_new_n15602__ & ~new_new_n15603__;
  assign new_new_n15605__ = new_new_n15589__ & new_new_n15604__;
  assign new_new_n15606__ = ~new_new_n15583__ & ~new_new_n15589__;
  assign new_new_n15607__ = ~new_new_n11465__ & new_new_n15602__;
  assign new_new_n15608__ = new_new_n11465__ & new_new_n15585__;
  assign new_new_n15609__ = ~new_new_n15607__ & ~new_new_n15608__;
  assign new_new_n15610__ = new_new_n15606__ & new_new_n15609__;
  assign new_new_n15611__ = new_new_n15583__ & ~new_new_n15604__;
  assign new_new_n15612__ = new_new_n11448__ & ~new_new_n15605__;
  assign new_new_n15613__ = ~new_new_n15611__ & new_new_n15612__;
  assign new_new_n15614__ = ~new_new_n15610__ & new_new_n15613__;
  assign new_new_n15615__ = ~new_new_n15601__ & ~new_new_n15614__;
  assign new_new_n15616__ = ~new_new_n14465__ & new_new_n14497__;
  assign new_new_n15617__ = new_new_n14465__ & ~new_new_n14497__;
  assign new_new_n15618__ = ~new_new_n14463__ & new_new_n14472__;
  assign new_new_n15619__ = ~new_new_n15617__ & new_new_n15618__;
  assign new_new_n15620__ = ~new_new_n15616__ & ~new_new_n15619__;
  assign new_new_n15621__ = new_new_n14487__ & ~new_new_n15620__;
  assign new_new_n15622__ = new_new_n14473__ & new_new_n14497__;
  assign new_new_n15623__ = new_new_n14463__ & new_new_n14474__;
  assign new_new_n15624__ = new_new_n14463__ & ~new_new_n14473__;
  assign new_new_n15625__ = new_new_n14474__ & ~new_new_n14497__;
  assign new_new_n15626__ = ~new_new_n15624__ & ~new_new_n15625__;
  assign new_new_n15627__ = ~new_new_n14487__ & ~new_new_n15626__;
  assign new_new_n15628__ = new_new_n14494__ & ~new_new_n15622__;
  assign new_new_n15629__ = ~new_new_n15623__ & new_new_n15628__;
  assign new_new_n15630__ = ~new_new_n15627__ & new_new_n15629__;
  assign new_new_n15631__ = ~new_new_n15621__ & new_new_n15630__;
  assign new_new_n15632__ = new_new_n14489__ & ~new_new_n14497__;
  assign new_new_n15633__ = ~new_new_n14490__ & ~new_new_n15632__;
  assign new_new_n15634__ = ~new_new_n14496__ & ~new_new_n14498__;
  assign new_new_n15635__ = new_new_n15575__ & new_new_n15634__;
  assign new_new_n15636__ = ~new_new_n14494__ & ~new_new_n15633__;
  assign new_new_n15637__ = ~new_new_n15635__ & new_new_n15636__;
  assign new_new_n15638__ = ~new_new_n15631__ & ~new_new_n15637__;
  assign new_new_n15639__ = ~new_new_n15615__ & ~new_new_n15638__;
  assign new_new_n15640__ = ~new_new_n14343__ & ~new_new_n14344__;
  assign new_new_n15641__ = new_new_n14367__ & new_new_n15640__;
  assign new_new_n15642__ = ~new_new_n14367__ & ~new_new_n15640__;
  assign new_new_n15643__ = ~new_new_n15641__ & ~new_new_n15642__;
  assign new_new_n15644__ = ~new_new_n14457__ & ~new_new_n14458__;
  assign new_new_n15645__ = ~new_new_n14460__ & ~new_new_n15644__;
  assign new_new_n15646__ = new_new_n14460__ & new_new_n15644__;
  assign new_new_n15647__ = ~new_new_n15645__ & ~new_new_n15646__;
  assign new_new_n15648__ = ~new_new_n15582__ & ~new_new_n15647__;
  assign new_new_n15649__ = ~new_new_n14376__ & ~new_new_n14448__;
  assign new_new_n15650__ = ~new_new_n14399__ & ~new_new_n14400__;
  assign new_new_n15651__ = new_new_n14413__ & ~new_new_n15650__;
  assign new_new_n15652__ = ~new_new_n14413__ & new_new_n15650__;
  assign new_new_n15653__ = ~new_new_n15651__ & ~new_new_n15652__;
  assign new_new_n15654__ = new_new_n15649__ & new_new_n15653__;
  assign new_new_n15655__ = ~new_new_n15649__ & ~new_new_n15653__;
  assign new_new_n15656__ = ~new_new_n15654__ & ~new_new_n15655__;
  assign new_new_n15657__ = new_new_n15648__ & new_new_n15656__;
  assign new_new_n15658__ = ~new_new_n13499__ & ~new_new_n13500__;
  assign new_new_n15659__ = new_new_n14340__ & ~new_new_n15658__;
  assign new_new_n15660__ = ~new_new_n14340__ & new_new_n15658__;
  assign new_new_n15661__ = ~new_new_n15659__ & ~new_new_n15660__;
  assign new_new_n15662__ = new_new_n15643__ & new_new_n15661__;
  assign new_new_n15663__ = ~new_new_n15643__ & ~new_new_n15661__;
  assign new_new_n15664__ = ~new_new_n15662__ & ~new_new_n15663__;
  assign new_new_n15665__ = ~new_new_n14319__ & ~new_new_n14320__;
  assign new_new_n15666__ = ~new_new_n14338__ & new_new_n15665__;
  assign new_new_n15667__ = new_new_n14338__ & ~new_new_n15665__;
  assign new_new_n15668__ = ~new_new_n15666__ & ~new_new_n15667__;
  assign new_new_n15669__ = ~new_new_n15661__ & ~new_new_n15668__;
  assign new_new_n15670__ = ~new_new_n14307__ & ~new_new_n14308__;
  assign new_new_n15671__ = ~new_new_n14312__ & new_new_n15670__;
  assign new_new_n15672__ = new_new_n14312__ & ~new_new_n15670__;
  assign new_new_n15673__ = ~new_new_n15671__ & ~new_new_n15672__;
  assign new_new_n15674__ = new_new_n15668__ & ~new_new_n15673__;
  assign new_new_n15675__ = new_new_n15643__ & new_new_n15674__;
  assign new_new_n15676__ = ~new_new_n15669__ & ~new_new_n15675__;
  assign new_new_n15677__ = ~new_new_n15664__ & new_new_n15676__;
  assign new_new_n15678__ = ~new_new_n15656__ & ~new_new_n15677__;
  assign new_new_n15679__ = new_new_n15661__ & new_new_n15673__;
  assign new_new_n15680__ = new_new_n15668__ & ~new_new_n15679__;
  assign new_new_n15681__ = new_new_n15643__ & ~new_new_n15680__;
  assign new_new_n15682__ = new_new_n15661__ & ~new_new_n15673__;
  assign new_new_n15683__ = new_new_n15668__ & ~new_new_n15682__;
  assign new_new_n15684__ = ~new_new_n15681__ & ~new_new_n15683__;
  assign new_new_n15685__ = ~new_new_n15664__ & ~new_new_n15684__;
  assign new_new_n15686__ = new_new_n15656__ & new_new_n15685__;
  assign new_new_n15687__ = ~new_new_n15678__ & ~new_new_n15686__;
  assign new_new_n15688__ = new_new_n14415__ & ~new_new_n14448__;
  assign new_new_n15689__ = ~new_new_n14416__ & ~new_new_n15688__;
  assign new_new_n15690__ = ~new_new_n14449__ & ~new_new_n14450__;
  assign new_new_n15691__ = new_new_n15649__ & new_new_n15690__;
  assign new_new_n15692__ = new_new_n14446__ & ~new_new_n15689__;
  assign new_new_n15693__ = ~new_new_n15691__ & new_new_n15692__;
  assign new_new_n15694__ = new_new_n14376__ & new_new_n14400__;
  assign new_new_n15695__ = new_new_n14376__ & new_new_n14380__;
  assign new_new_n15696__ = ~new_new_n14376__ & ~new_new_n14380__;
  assign new_new_n15697__ = new_new_n14398__ & ~new_new_n14448__;
  assign new_new_n15698__ = ~new_new_n15696__ & new_new_n15697__;
  assign new_new_n15699__ = ~new_new_n15695__ & ~new_new_n15698__;
  assign new_new_n15700__ = new_new_n14413__ & ~new_new_n15699__;
  assign new_new_n15701__ = ~new_new_n14400__ & new_new_n14448__;
  assign new_new_n15702__ = ~new_new_n14398__ & new_new_n15696__;
  assign new_new_n15703__ = ~new_new_n15701__ & ~new_new_n15702__;
  assign new_new_n15704__ = ~new_new_n14413__ & ~new_new_n15703__;
  assign new_new_n15705__ = new_new_n14399__ & new_new_n14448__;
  assign new_new_n15706__ = ~new_new_n14446__ & ~new_new_n15694__;
  assign new_new_n15707__ = ~new_new_n15705__ & new_new_n15706__;
  assign new_new_n15708__ = ~new_new_n15700__ & new_new_n15707__;
  assign new_new_n15709__ = ~new_new_n15704__ & new_new_n15708__;
  assign new_new_n15710__ = ~new_new_n15693__ & ~new_new_n15709__;
  assign new_new_n15711__ = new_new_n15582__ & new_new_n15647__;
  assign new_new_n15712__ = ~new_new_n15710__ & new_new_n15711__;
  assign new_new_n15713__ = ~new_new_n15687__ & new_new_n15712__;
  assign new_new_n15714__ = ~new_new_n15657__ & ~new_new_n15713__;
  assign new_new_n15715__ = new_new_n15643__ & ~new_new_n15714__;
  assign new_new_n15716__ = ~new_new_n15582__ & new_new_n15647__;
  assign new_new_n15717__ = new_new_n15687__ & new_new_n15716__;
  assign new_new_n15718__ = new_new_n15582__ & ~new_new_n15647__;
  assign new_new_n15719__ = new_new_n15710__ & new_new_n15718__;
  assign new_new_n15720__ = ~new_new_n15717__ & ~new_new_n15719__;
  assign new_new_n15721__ = ~new_new_n15656__ & ~new_new_n15720__;
  assign new_new_n15722__ = ~new_new_n15647__ & ~new_new_n15710__;
  assign new_new_n15723__ = new_new_n15647__ & new_new_n15710__;
  assign new_new_n15724__ = ~new_new_n15722__ & ~new_new_n15723__;
  assign new_new_n15725__ = ~new_new_n15582__ & ~new_new_n15724__;
  assign new_new_n15726__ = new_new_n15648__ & ~new_new_n15687__;
  assign new_new_n15727__ = ~new_new_n15712__ & ~new_new_n15726__;
  assign new_new_n15728__ = new_new_n15656__ & ~new_new_n15727__;
  assign new_new_n15729__ = ~new_new_n15656__ & new_new_n15716__;
  assign new_new_n15730__ = new_new_n15687__ & new_new_n15719__;
  assign new_new_n15731__ = ~new_new_n15729__ & ~new_new_n15730__;
  assign new_new_n15732__ = ~new_new_n15643__ & ~new_new_n15731__;
  assign new_new_n15733__ = ~new_new_n15721__ & ~new_new_n15725__;
  assign new_new_n15734__ = ~new_new_n15728__ & new_new_n15733__;
  assign new_new_n15735__ = ~new_new_n15715__ & ~new_new_n15732__;
  assign new_new_n15736__ = new_new_n15734__ & new_new_n15735__;
  assign new_new_n15737__ = ~new_new_n15585__ & ~new_new_n15602__;
  assign new_new_n15738__ = new_new_n11465__ & ~new_new_n15606__;
  assign new_new_n15739__ = ~new_new_n11465__ & new_new_n15606__;
  assign new_new_n15740__ = ~new_new_n15738__ & ~new_new_n15739__;
  assign new_new_n15741__ = new_new_n15737__ & new_new_n15740__;
  assign new_new_n15742__ = ~new_new_n15737__ & ~new_new_n15740__;
  assign new_new_n15743__ = ~new_new_n15741__ & ~new_new_n15742__;
  assign new_new_n15744__ = new_new_n15736__ & new_new_n15743__;
  assign new_new_n15745__ = ~new_new_n15639__ & ~new_new_n15744__;
  assign new_new_n15746__ = ~new_new_n15582__ & ~new_new_n15745__;
  assign new_new_n15747__ = ~new_new_n15582__ & new_new_n15743__;
  assign new_new_n15748__ = ~new_new_n15638__ & new_new_n15736__;
  assign new_new_n15749__ = ~new_new_n15615__ & new_new_n15748__;
  assign new_new_n15750__ = ~new_new_n15747__ & ~new_new_n15749__;
  assign new_new_n15751__ = ~new_new_n15647__ & ~new_new_n15750__;
  assign new_new_n15752__ = new_new_n15615__ & new_new_n15638__;
  assign new_new_n15753__ = new_new_n15743__ & ~new_new_n15752__;
  assign new_new_n15754__ = ~new_new_n15746__ & ~new_new_n15753__;
  assign new_new_n15755__ = ~new_new_n15751__ & new_new_n15754__;
  assign new_new_n15756__ = new_new_n15574__ & ~new_new_n15755__;
  assign new_new_n15757__ = new_new_n15572__ & ~new_new_n15755__;
  assign new_new_n15758__ = ~new_new_n15574__ & ~new_new_n15757__;
  assign new_new_n15759__ = ~new_new_n15615__ & ~new_new_n15758__;
  assign new_new_n15760__ = ~new_new_n15573__ & ~new_new_n15756__;
  assign new_new_n15761__ = ~new_new_n15759__ & new_new_n15760__;
  assign new_new_n15762__ = ~new_new_n15533__ & new_new_n15560__;
  assign new_new_n15763__ = ~new_new_n15761__ & new_new_n15762__;
  assign new_new_n15764__ = ~new_new_n14570__ & ~new_new_n14571__;
  assign new_new_n15765__ = new_new_n14575__ & new_new_n15764__;
  assign new_new_n15766__ = ~new_new_n14575__ & ~new_new_n15764__;
  assign new_new_n15767__ = ~new_new_n15765__ & ~new_new_n15766__;
  assign new_new_n15768__ = new_new_n15533__ & ~new_new_n15560__;
  assign new_new_n15769__ = new_new_n15761__ & new_new_n15768__;
  assign new_new_n15770__ = new_new_n15767__ & ~new_new_n15769__;
  assign new_new_n15771__ = ~new_new_n15763__ & ~new_new_n15770__;
  assign new_new_n15772__ = new_new_n15524__ & ~new_new_n15533__;
  assign new_new_n15773__ = ~new_new_n15771__ & new_new_n15772__;
  assign new_new_n15774__ = ~new_new_n15536__ & ~new_new_n15773__;
  assign new_new_n15775__ = new_new_n15487__ & new_new_n15774__;
  assign new_new_n15776__ = new_new_n15471__ & new_new_n15775__;
  assign new_new_n15777__ = new_new_n15520__ & ~new_new_n15771__;
  assign new_new_n15778__ = ~new_new_n15487__ & new_new_n15777__;
  assign new_new_n15779__ = new_new_n15774__ & ~new_new_n15778__;
  assign new_new_n15780__ = ~new_new_n15487__ & ~new_new_n15779__;
  assign new_new_n15781__ = ~new_new_n15471__ & new_new_n15780__;
  assign new_new_n15782__ = new_new_n14657__ & new_new_n15477__;
  assign new_new_n15783__ = ~new_new_n14657__ & new_new_n15476__;
  assign new_new_n15784__ = ~new_new_n15782__ & ~new_new_n15783__;
  assign new_new_n15785__ = new_new_n15481__ & new_new_n15784__;
  assign new_new_n15786__ = ~new_new_n14657__ & ~new_new_n15477__;
  assign new_new_n15787__ = ~new_new_n15476__ & ~new_new_n15786__;
  assign new_new_n15788__ = new_new_n15479__ & ~new_new_n15787__;
  assign new_new_n15789__ = new_new_n15480__ & new_new_n15787__;
  assign new_new_n15790__ = new_new_n14639__ & ~new_new_n15788__;
  assign new_new_n15791__ = ~new_new_n15789__ & new_new_n15790__;
  assign new_new_n15792__ = ~new_new_n15785__ & new_new_n15791__;
  assign new_new_n15793__ = new_new_n14636__ & new_new_n14645__;
  assign new_new_n15794__ = ~new_new_n6947__ & new_new_n15793__;
  assign new_new_n15795__ = ~new_new_n14636__ & ~new_new_n14645__;
  assign new_new_n15796__ = ~new_new_n14660__ & ~new_new_n15795__;
  assign new_new_n15797__ = ~new_new_n6947__ & new_new_n15796__;
  assign new_new_n15798__ = ~new_new_n15793__ & ~new_new_n15797__;
  assign new_new_n15799__ = ~new_new_n14657__ & ~new_new_n15798__;
  assign new_new_n15800__ = ~new_new_n14636__ & new_new_n14660__;
  assign new_new_n15801__ = ~new_new_n6947__ & ~new_new_n15800__;
  assign new_new_n15802__ = new_new_n14657__ & ~new_new_n15796__;
  assign new_new_n15803__ = ~new_new_n15801__ & new_new_n15802__;
  assign new_new_n15804__ = new_new_n15477__ & new_new_n15479__;
  assign new_new_n15805__ = ~new_new_n14639__ & ~new_new_n15794__;
  assign new_new_n15806__ = ~new_new_n15804__ & new_new_n15805__;
  assign new_new_n15807__ = ~new_new_n15803__ & new_new_n15806__;
  assign new_new_n15808__ = ~new_new_n15799__ & new_new_n15807__;
  assign new_new_n15809__ = ~new_new_n15792__ & ~new_new_n15808__;
  assign new_new_n15810__ = ~new_new_n15781__ & new_new_n15809__;
  assign new_new_n15811__ = ~new_new_n15776__ & ~new_new_n15810__;
  assign new_new_n15812__ = new_new_n15439__ & ~new_new_n15811__;
  assign new_new_n15813__ = ~new_new_n15432__ & ~new_new_n15812__;
  assign new_new_n15814__ = new_new_n15464__ & new_new_n15471__;
  assign new_new_n15815__ = ~new_new_n15464__ & ~new_new_n15471__;
  assign new_new_n15816__ = ~new_new_n15814__ & ~new_new_n15815__;
  assign new_new_n15817__ = new_new_n15811__ & ~new_new_n15816__;
  assign new_new_n15818__ = ~new_new_n15811__ & new_new_n15816__;
  assign new_new_n15819__ = ~new_new_n15817__ & ~new_new_n15818__;
  assign new_new_n15820__ = new_new_n15464__ & ~new_new_n15812__;
  assign new_new_n15821__ = ~new_new_n15813__ & new_new_n15819__;
  assign new_new_n15822__ = ~new_new_n15820__ & new_new_n15821__;
  assign new_new_n15823__ = ~new_new_n15474__ & ~new_new_n15475__;
  assign new_new_n15824__ = ~new_new_n15822__ & new_new_n15823__;
  assign new_new_n15825__ = ~new_new_n15432__ & new_new_n15824__;
  assign new_new_n15826__ = new_new_n15362__ & ~new_new_n15825__;
  assign new_new_n15827__ = new_new_n15432__ & ~new_new_n15824__;
  assign new_new_n15828__ = ~new_new_n15362__ & ~new_new_n15827__;
  assign new_new_n15829__ = ~new_new_n15826__ & ~new_new_n15828__;
  assign new_new_n15830__ = new_new_n15399__ & ~new_new_n15829__;
  assign new_new_n15831__ = ~new_new_n15391__ & ~new_new_n15830__;
  assign new_new_n15832__ = new_new_n15362__ & ~new_new_n15831__;
  assign new_new_n15833__ = new_new_n15349__ & new_new_n15829__;
  assign new_new_n15834__ = ~new_new_n15399__ & ~new_new_n15833__;
  assign new_new_n15835__ = ~new_new_n15390__ & ~new_new_n15834__;
  assign new_new_n15836__ = new_new_n15349__ & new_new_n15398__;
  assign new_new_n15837__ = ~new_new_n15835__ & ~new_new_n15836__;
  assign new_new_n15838__ = ~new_new_n15832__ & new_new_n15837__;
  assign new_new_n15839__ = ~new_new_n15350__ & new_new_n15838__;
  assign new_new_n15840__ = ~new_new_n15273__ & ~new_new_n15314__;
  assign new_new_n15841__ = new_new_n15286__ & ~new_new_n15321__;
  assign new_new_n15842__ = ~new_new_n15840__ & ~new_new_n15841__;
  assign new_new_n15843__ = new_new_n15839__ & ~new_new_n15842__;
  assign new_new_n15844__ = new_new_n15285__ & ~new_new_n15314__;
  assign new_new_n15845__ = ~new_new_n15325__ & ~new_new_n15844__;
  assign new_new_n15846__ = ~new_new_n15324__ & new_new_n15845__;
  assign new_new_n15847__ = ~new_new_n15843__ & new_new_n15846__;
  assign new_new_n15848__ = new_new_n15248__ & new_new_n15847__;
  assign new_new_n15849__ = ~new_new_n15244__ & ~new_new_n15847__;
  assign new_new_n15850__ = ~new_new_n15848__ & ~new_new_n15849__;
  assign new_new_n15851__ = ~new_new_n15249__ & ~new_new_n15850__;
  assign new_new_n15852__ = ~new_new_n15237__ & ~new_new_n15851__;
  assign new_new_n15853__ = ~new_new_n94__ & ~new_new_n125__;
  assign new_new_n15854__ = ~new_new_n15249__ & new_new_n15853__;
  assign new_new_n15855__ = new_new_n15852__ & ~new_new_n15854__;
  assign new_new_n15856__ = new_new_n15244__ & new_new_n15847__;
  assign new_new_n15857__ = new_new_n15237__ & new_new_n15856__;
  assign new_new_n15858__ = ~new_new_n161__ & ~new_new_n15857__;
  assign new_new_n15859__ = ~new_new_n71__ & new_new_n15248__;
  assign new_new_n15860__ = ~new_new_n15858__ & new_new_n15859__;
  assign new_new_n15861__ = new_new_n15237__ & ~new_new_n15847__;
  assign new_new_n15862__ = ~new_new_n15248__ & new_new_n15861__;
  assign new_new_n15863__ = ~new_new_n71__ & ~new_new_n15862__;
  assign new_new_n15864__ = ~new_new_n161__ & ~new_new_n15244__;
  assign new_new_n15865__ = ~new_new_n15863__ & new_new_n15864__;
  assign new_new_n15866__ = ~new_new_n15855__ & ~new_new_n15860__;
  assign new_new_n15867__ = ~new_new_n15865__ & new_new_n15866__;
  assign new_new_n15868__ = pi31 & ~new_new_n15867__;
  assign new_new_n15869__ = new_new_n161__ & new_new_n15244__;
  assign new_new_n15870__ = new_new_n765__ & new_new_n15237__;
  assign new_new_n15871__ = ~pi31 & ~new_new_n15869__;
  assign new_new_n15872__ = ~new_new_n15870__ & new_new_n15871__;
  assign new_new_n15873__ = ~new_new_n15868__ & ~new_new_n15872__;
  assign new_new_n15874__ = new_new_n418__ & ~new_new_n15873__;
  assign new_new_n15875__ = ~new_new_n3853__ & new_new_n3881__;
  assign new_new_n15876__ = ~new_new_n3854__ & ~new_new_n15875__;
  assign new_new_n15877__ = ~new_new_n76__ & ~new_new_n168__;
  assign new_new_n15878__ = ~new_new_n320__ & ~new_new_n438__;
  assign new_new_n15879__ = new_new_n15877__ & new_new_n15878__;
  assign new_new_n15880__ = ~new_new_n655__ & new_new_n15879__;
  assign new_new_n15881__ = ~new_new_n437__ & new_new_n15880__;
  assign new_new_n15882__ = new_new_n3831__ & new_new_n15881__;
  assign new_new_n15883__ = new_new_n3764__ & new_new_n15882__;
  assign new_new_n15884__ = new_new_n3881__ & new_new_n15883__;
  assign new_new_n15885__ = ~new_new_n3881__ & ~new_new_n15883__;
  assign new_new_n15886__ = ~new_new_n15884__ & ~new_new_n15885__;
  assign new_new_n15887__ = ~new_new_n3884__ & new_new_n15218__;
  assign new_new_n15888__ = ~new_new_n3884__ & ~new_new_n15231__;
  assign new_new_n15889__ = new_new_n3888__ & ~new_new_n15888__;
  assign new_new_n15890__ = new_new_n4177__ & new_new_n15201__;
  assign new_new_n15891__ = new_new_n3884__ & ~new_new_n15890__;
  assign new_new_n15892__ = ~new_new_n15221__ & ~new_new_n15891__;
  assign new_new_n15893__ = ~new_new_n15889__ & new_new_n15892__;
  assign new_new_n15894__ = new_new_n3884__ & ~new_new_n15218__;
  assign new_new_n15895__ = ~new_new_n3888__ & ~new_new_n15231__;
  assign new_new_n15896__ = ~new_new_n15890__ & ~new_new_n15895__;
  assign new_new_n15897__ = ~new_new_n15894__ & ~new_new_n15896__;
  assign new_new_n15898__ = ~new_new_n15887__ & ~new_new_n15893__;
  assign new_new_n15899__ = ~new_new_n15897__ & new_new_n15898__;
  assign new_new_n15900__ = new_new_n15886__ & ~new_new_n15899__;
  assign new_new_n15901__ = ~new_new_n15886__ & new_new_n15899__;
  assign new_new_n15902__ = ~new_new_n15900__ & ~new_new_n15901__;
  assign new_new_n15903__ = new_new_n15876__ & new_new_n15902__;
  assign new_new_n15904__ = ~new_new_n15876__ & ~new_new_n15902__;
  assign new_new_n15905__ = ~new_new_n15903__ & ~new_new_n15904__;
  assign new_new_n15906__ = ~pi31 & ~new_new_n15905__;
  assign new_new_n15907__ = ~new_new_n15237__ & new_new_n15905__;
  assign new_new_n15908__ = new_new_n15237__ & ~new_new_n15905__;
  assign new_new_n15909__ = ~new_new_n15907__ & ~new_new_n15908__;
  assign new_new_n15910__ = new_new_n15244__ & ~new_new_n15848__;
  assign new_new_n15911__ = ~new_new_n15244__ & new_new_n15847__;
  assign new_new_n15912__ = new_new_n15237__ & ~new_new_n15249__;
  assign new_new_n15913__ = ~new_new_n15911__ & new_new_n15912__;
  assign new_new_n15914__ = ~new_new_n15910__ & ~new_new_n15913__;
  assign new_new_n15915__ = new_new_n15909__ & ~new_new_n15914__;
  assign new_new_n15916__ = ~new_new_n15909__ & new_new_n15914__;
  assign new_new_n15917__ = ~new_new_n15915__ & ~new_new_n15916__;
  assign new_new_n15918__ = pi31 & new_new_n15917__;
  assign new_new_n15919__ = new_new_n765__ & ~new_new_n15906__;
  assign new_new_n15920__ = ~new_new_n15918__ & new_new_n15919__;
  assign new_new_n15921__ = ~new_new_n4148__ & new_new_n15853__;
  assign new_new_n15922__ = new_new_n15237__ & new_new_n15921__;
  assign new_new_n15923__ = ~new_new_n15920__ & ~new_new_n15922__;
  assign new_new_n15924__ = new_new_n15874__ & new_new_n15923__;
  assign new_new_n15925__ = ~new_new_n418__ & new_new_n15873__;
  assign new_new_n15926__ = ~new_new_n15923__ & new_new_n15925__;
  assign new_new_n15927__ = new_new_n15923__ & ~new_new_n15925__;
  assign new_new_n15928__ = ~pi26 & ~new_new_n303__;
  assign new_new_n15929__ = ~new_new_n2759__ & ~new_new_n15928__;
  assign new_new_n15930__ = ~new_new_n91__ & new_new_n165__;
  assign new_new_n15931__ = ~new_new_n88__ & ~new_new_n718__;
  assign new_new_n15932__ = ~new_new_n15930__ & new_new_n15931__;
  assign new_new_n15933__ = ~new_new_n424__ & new_new_n15932__;
  assign new_new_n15934__ = ~new_new_n1372__ & new_new_n15933__;
  assign new_new_n15935__ = ~new_new_n76__ & new_new_n674__;
  assign new_new_n15936__ = new_new_n15934__ & new_new_n15935__;
  assign new_new_n15937__ = new_new_n503__ & new_new_n15936__;
  assign new_new_n15938__ = new_new_n575__ & new_new_n15937__;
  assign new_new_n15939__ = ~new_new_n15929__ & new_new_n15938__;
  assign new_new_n15940__ = new_new_n15929__ & ~new_new_n15938__;
  assign new_new_n15941__ = ~new_new_n15939__ & ~new_new_n15940__;
  assign new_new_n15942__ = ~new_new_n15927__ & ~new_new_n15941__;
  assign new_new_n15943__ = ~new_new_n200__ & ~new_new_n482__;
  assign new_new_n15944__ = ~new_new_n816__ & new_new_n15943__;
  assign new_new_n15945__ = new_new_n1368__ & new_new_n15944__;
  assign new_new_n15946__ = new_new_n589__ & new_new_n592__;
  assign new_new_n15947__ = ~new_new_n676__ & new_new_n15946__;
  assign new_new_n15948__ = new_new_n7607__ & new_new_n15945__;
  assign new_new_n15949__ = new_new_n15947__ & new_new_n15948__;
  assign new_new_n15950__ = ~new_new_n88__ & ~new_new_n441__;
  assign new_new_n15951__ = ~new_new_n692__ & new_new_n15950__;
  assign new_new_n15952__ = ~new_new_n198__ & new_new_n3258__;
  assign new_new_n15953__ = new_new_n5699__ & new_new_n15952__;
  assign new_new_n15954__ = new_new_n354__ & new_new_n15951__;
  assign new_new_n15955__ = ~new_new_n837__ & new_new_n15954__;
  assign new_new_n15956__ = new_new_n15953__ & new_new_n15955__;
  assign new_new_n15957__ = new_new_n187__ & new_new_n15956__;
  assign new_new_n15958__ = new_new_n889__ & new_new_n15949__;
  assign new_new_n15959__ = new_new_n15957__ & new_new_n15958__;
  assign new_new_n15960__ = new_new_n3685__ & new_new_n15959__;
  assign new_new_n15961__ = ~new_new_n15926__ & ~new_new_n15960__;
  assign new_new_n15962__ = ~new_new_n15942__ & new_new_n15961__;
  assign new_new_n15963__ = ~new_new_n15874__ & ~new_new_n15923__;
  assign new_new_n15964__ = ~new_new_n15941__ & new_new_n15960__;
  assign new_new_n15965__ = ~new_new_n15963__ & new_new_n15964__;
  assign new_new_n15966__ = ~new_new_n15924__ & ~new_new_n15965__;
  assign new_new_n15967__ = ~new_new_n15962__ & new_new_n15966__;
  assign new_new_n15968__ = new_new_n70__ & ~new_new_n15967__;
  assign new_new_n15969__ = ~new_new_n70__ & new_new_n15967__;
  assign new_new_n15970__ = ~new_new_n15968__ & ~new_new_n15969__;
  assign new_new_n15971__ = pi30 & new_new_n15905__;
  assign new_new_n15972__ = ~new_new_n15883__ & ~new_new_n15899__;
  assign new_new_n15973__ = ~new_new_n3852__ & ~new_new_n15972__;
  assign new_new_n15974__ = new_new_n15883__ & new_new_n15899__;
  assign new_new_n15975__ = new_new_n3852__ & ~new_new_n15974__;
  assign new_new_n15976__ = new_new_n3881__ & ~new_new_n15973__;
  assign new_new_n15977__ = ~new_new_n15975__ & new_new_n15976__;
  assign new_new_n15978__ = new_new_n165__ & new_new_n9357__;
  assign new_new_n15979__ = ~new_new_n718__ & ~new_new_n1372__;
  assign new_new_n15980__ = ~new_new_n192__ & new_new_n15979__;
  assign new_new_n15981__ = new_new_n210__ & ~new_new_n321__;
  assign new_new_n15982__ = ~new_new_n15978__ & new_new_n15981__;
  assign new_new_n15983__ = new_new_n628__ & new_new_n15980__;
  assign new_new_n15984__ = new_new_n15982__ & new_new_n15983__;
  assign new_new_n15985__ = new_new_n806__ & new_new_n15984__;
  assign new_new_n15986__ = new_new_n578__ & new_new_n15985__;
  assign new_new_n15987__ = new_new_n3881__ & ~new_new_n15883__;
  assign new_new_n15988__ = ~new_new_n15986__ & ~new_new_n15987__;
  assign new_new_n15989__ = ~new_new_n15972__ & new_new_n15988__;
  assign new_new_n15990__ = ~new_new_n15977__ & ~new_new_n15989__;
  assign new_new_n15991__ = ~new_new_n3772__ & ~new_new_n15990__;
  assign new_new_n15992__ = new_new_n3772__ & new_new_n15972__;
  assign new_new_n15993__ = ~new_new_n3854__ & ~new_new_n15972__;
  assign new_new_n15994__ = ~new_new_n3881__ & ~new_new_n15974__;
  assign new_new_n15995__ = ~new_new_n15993__ & new_new_n15994__;
  assign new_new_n15996__ = ~new_new_n15992__ & ~new_new_n15995__;
  assign new_new_n15997__ = new_new_n15986__ & ~new_new_n15996__;
  assign new_new_n15998__ = ~new_new_n15991__ & ~new_new_n15997__;
  assign new_new_n15999__ = new_new_n765__ & ~new_new_n15998__;
  assign new_new_n16000__ = ~new_new_n15971__ & ~new_new_n15999__;
  assign new_new_n16001__ = ~pi31 & ~new_new_n16000__;
  assign new_new_n16002__ = new_new_n15909__ & new_new_n15998__;
  assign new_new_n16003__ = ~new_new_n15905__ & new_new_n15998__;
  assign new_new_n16004__ = ~new_new_n15244__ & new_new_n16003__;
  assign new_new_n16005__ = new_new_n15907__ & ~new_new_n15998__;
  assign new_new_n16006__ = new_new_n15847__ & new_new_n16005__;
  assign new_new_n16007__ = ~new_new_n16004__ & ~new_new_n16006__;
  assign new_new_n16008__ = new_new_n15248__ & ~new_new_n16007__;
  assign new_new_n16009__ = new_new_n15847__ & new_new_n16003__;
  assign new_new_n16010__ = ~new_new_n16005__ & ~new_new_n16009__;
  assign new_new_n16011__ = ~new_new_n15244__ & ~new_new_n16010__;
  assign new_new_n16012__ = new_new_n15905__ & new_new_n15998__;
  assign new_new_n16013__ = ~new_new_n15847__ & new_new_n16012__;
  assign new_new_n16014__ = ~new_new_n15905__ & ~new_new_n15998__;
  assign new_new_n16015__ = new_new_n15237__ & new_new_n16014__;
  assign new_new_n16016__ = ~new_new_n16013__ & ~new_new_n16015__;
  assign new_new_n16017__ = new_new_n15244__ & ~new_new_n16016__;
  assign new_new_n16018__ = new_new_n15244__ & new_new_n16012__;
  assign new_new_n16019__ = new_new_n15861__ & new_new_n16014__;
  assign new_new_n16020__ = ~new_new_n16018__ & ~new_new_n16019__;
  assign new_new_n16021__ = ~new_new_n15248__ & ~new_new_n16020__;
  assign new_new_n16022__ = ~new_new_n16008__ & ~new_new_n16011__;
  assign new_new_n16023__ = ~new_new_n16017__ & ~new_new_n16021__;
  assign new_new_n16024__ = new_new_n16022__ & new_new_n16023__;
  assign new_new_n16025__ = ~new_new_n16002__ & new_new_n16024__;
  assign new_new_n16026__ = new_new_n765__ & new_new_n16025__;
  assign new_new_n16027__ = new_new_n71__ & new_new_n15905__;
  assign new_new_n16028__ = ~new_new_n15869__ & ~new_new_n16027__;
  assign new_new_n16029__ = ~new_new_n16026__ & new_new_n16028__;
  assign new_new_n16030__ = pi31 & ~new_new_n16029__;
  assign new_new_n16031__ = ~new_new_n16001__ & ~new_new_n16030__;
  assign new_new_n16032__ = ~new_new_n15939__ & ~new_new_n15960__;
  assign new_new_n16033__ = ~new_new_n15940__ & ~new_new_n16032__;
  assign new_new_n16034__ = ~new_new_n16031__ & ~new_new_n16033__;
  assign new_new_n16035__ = new_new_n16031__ & new_new_n16033__;
  assign new_new_n16036__ = ~new_new_n16034__ & ~new_new_n16035__;
  assign new_new_n16037__ = new_new_n537__ & new_new_n15934__;
  assign new_new_n16038__ = new_new_n462__ & new_new_n16037__;
  assign new_new_n16039__ = ~new_new_n16036__ & new_new_n16038__;
  assign new_new_n16040__ = new_new_n16036__ & ~new_new_n16038__;
  assign new_new_n16041__ = ~new_new_n16039__ & ~new_new_n16040__;
  assign new_new_n16042__ = new_new_n15970__ & ~new_new_n16041__;
  assign new_new_n16043__ = ~new_new_n15970__ & new_new_n16041__;
  assign new_new_n16044__ = ~new_new_n16042__ & ~new_new_n16043__;
  assign new_new_n16045__ = new_new_n4212__ & ~new_new_n15998__;
  assign new_new_n16046__ = ~new_new_n15237__ & ~new_new_n15910__;
  assign new_new_n16047__ = new_new_n15905__ & ~new_new_n16046__;
  assign new_new_n16048__ = new_new_n15998__ & ~new_new_n16047__;
  assign new_new_n16049__ = ~new_new_n15905__ & ~new_new_n15913__;
  assign new_new_n16050__ = ~new_new_n15998__ & ~new_new_n16049__;
  assign new_new_n16051__ = ~new_new_n16048__ & ~new_new_n16050__;
  assign new_new_n16052__ = ~new_new_n4215__ & new_new_n16051__;
  assign new_new_n16053__ = new_new_n15884__ & new_new_n15986__;
  assign new_new_n16054__ = ~new_new_n97__ & ~new_new_n16053__;
  assign new_new_n16055__ = new_new_n15876__ & ~new_new_n16054__;
  assign new_new_n16056__ = new_new_n15899__ & new_new_n16055__;
  assign new_new_n16057__ = new_new_n4214__ & ~new_new_n16056__;
  assign new_new_n16058__ = ~new_new_n16052__ & new_new_n16057__;
  assign new_new_n16059__ = ~new_new_n16045__ & ~new_new_n16058__;
  assign new_new_n16060__ = ~pi29 & new_new_n16059__;
  assign new_new_n16061__ = ~new_new_n15905__ & new_new_n16060__;
  assign new_new_n16062__ = new_new_n161__ & ~new_new_n15314__;
  assign new_new_n16063__ = new_new_n765__ & ~new_new_n15248__;
  assign new_new_n16064__ = ~new_new_n16062__ & ~new_new_n16063__;
  assign new_new_n16065__ = ~pi31 & ~new_new_n16064__;
  assign new_new_n16066__ = new_new_n71__ & new_new_n15314__;
  assign new_new_n16067__ = new_new_n15248__ & new_new_n15314__;
  assign new_new_n16068__ = ~new_new_n15273__ & new_new_n15285__;
  assign new_new_n16069__ = new_new_n15285__ & ~new_new_n15839__;
  assign new_new_n16070__ = ~new_new_n15285__ & new_new_n15839__;
  assign new_new_n16071__ = ~new_new_n16069__ & ~new_new_n16070__;
  assign new_new_n16072__ = ~new_new_n15273__ & new_new_n15839__;
  assign new_new_n16073__ = new_new_n15273__ & ~new_new_n15839__;
  assign new_new_n16074__ = new_new_n15321__ & ~new_new_n16073__;
  assign new_new_n16075__ = ~new_new_n16072__ & ~new_new_n16074__;
  assign new_new_n16076__ = new_new_n16071__ & new_new_n16075__;
  assign new_new_n16077__ = ~new_new_n16071__ & ~new_new_n16075__;
  assign new_new_n16078__ = ~new_new_n16076__ & ~new_new_n16077__;
  assign new_new_n16079__ = new_new_n15285__ & new_new_n16078__;
  assign new_new_n16080__ = ~new_new_n15273__ & ~new_new_n16078__;
  assign new_new_n16081__ = ~new_new_n16079__ & ~new_new_n16080__;
  assign new_new_n16082__ = ~new_new_n16068__ & ~new_new_n16081__;
  assign new_new_n16083__ = new_new_n15325__ & ~new_new_n16082__;
  assign new_new_n16084__ = ~new_new_n161__ & ~new_new_n16067__;
  assign new_new_n16085__ = ~new_new_n16083__ & new_new_n16084__;
  assign new_new_n16086__ = ~new_new_n15285__ & ~new_new_n16085__;
  assign new_new_n16087__ = ~new_new_n161__ & new_new_n15285__;
  assign new_new_n16088__ = ~new_new_n15285__ & ~new_new_n16078__;
  assign new_new_n16089__ = new_new_n15840__ & new_new_n16088__;
  assign new_new_n16090__ = ~new_new_n16087__ & ~new_new_n16089__;
  assign new_new_n16091__ = new_new_n15314__ & ~new_new_n16082__;
  assign new_new_n16092__ = ~new_new_n15248__ & ~new_new_n16091__;
  assign new_new_n16093__ = new_new_n15248__ & new_new_n16091__;
  assign new_new_n16094__ = ~new_new_n16090__ & ~new_new_n16092__;
  assign new_new_n16095__ = ~new_new_n16093__ & new_new_n16094__;
  assign new_new_n16096__ = ~new_new_n16086__ & ~new_new_n16095__;
  assign new_new_n16097__ = ~new_new_n71__ & ~new_new_n16096__;
  assign new_new_n16098__ = pi31 & ~new_new_n16066__;
  assign new_new_n16099__ = ~new_new_n16097__ & new_new_n16098__;
  assign new_new_n16100__ = ~new_new_n16065__ & ~new_new_n16099__;
  assign new_new_n16101__ = new_new_n15273__ & new_new_n15321__;
  assign new_new_n16102__ = ~new_new_n15321__ & ~new_new_n15838__;
  assign new_new_n16103__ = ~new_new_n16072__ & ~new_new_n16102__;
  assign new_new_n16104__ = new_new_n765__ & ~new_new_n16103__;
  assign new_new_n16105__ = ~new_new_n16101__ & ~new_new_n16104__;
  assign new_new_n16106__ = ~new_new_n15285__ & ~new_new_n16105__;
  assign new_new_n16107__ = new_new_n15285__ & ~new_new_n15321__;
  assign new_new_n16108__ = new_new_n15839__ & new_new_n16107__;
  assign new_new_n16109__ = ~new_new_n71__ & ~new_new_n16108__;
  assign new_new_n16110__ = ~new_new_n161__ & new_new_n15273__;
  assign new_new_n16111__ = ~new_new_n16109__ & new_new_n16110__;
  assign new_new_n16112__ = ~new_new_n15273__ & new_new_n16069__;
  assign new_new_n16113__ = ~new_new_n161__ & ~new_new_n16112__;
  assign new_new_n16114__ = ~new_new_n71__ & new_new_n15321__;
  assign new_new_n16115__ = ~new_new_n16113__ & new_new_n16114__;
  assign new_new_n16116__ = pi31 & ~new_new_n16111__;
  assign new_new_n16117__ = ~new_new_n16115__ & new_new_n16116__;
  assign new_new_n16118__ = ~new_new_n16106__ & new_new_n16117__;
  assign new_new_n16119__ = new_new_n161__ & ~new_new_n15273__;
  assign new_new_n16120__ = new_new_n765__ & new_new_n15285__;
  assign new_new_n16121__ = ~new_new_n16119__ & ~new_new_n16120__;
  assign new_new_n16122__ = ~pi31 & ~new_new_n16121__;
  assign new_new_n16123__ = ~new_new_n16118__ & ~new_new_n16122__;
  assign new_new_n16124__ = ~new_new_n673__ & ~new_new_n846__;
  assign new_new_n16125__ = ~new_new_n921__ & new_new_n16124__;
  assign new_new_n16126__ = new_new_n4565__ & new_new_n16125__;
  assign new_new_n16127__ = new_new_n2029__ & new_new_n16126__;
  assign new_new_n16128__ = ~new_new_n483__ & ~new_new_n1176__;
  assign new_new_n16129__ = ~new_new_n212__ & ~new_new_n385__;
  assign new_new_n16130__ = ~new_new_n624__ & ~new_new_n693__;
  assign new_new_n16131__ = ~new_new_n875__ & ~new_new_n1007__;
  assign new_new_n16132__ = new_new_n16130__ & new_new_n16131__;
  assign new_new_n16133__ = ~new_new_n155__ & new_new_n16129__;
  assign new_new_n16134__ = ~new_new_n477__ & new_new_n16133__;
  assign new_new_n16135__ = new_new_n3369__ & new_new_n16132__;
  assign new_new_n16136__ = new_new_n5431__ & new_new_n16128__;
  assign new_new_n16137__ = new_new_n16135__ & new_new_n16136__;
  assign new_new_n16138__ = ~new_new_n1539__ & new_new_n16134__;
  assign new_new_n16139__ = new_new_n16137__ & new_new_n16138__;
  assign new_new_n16140__ = ~new_new_n959__ & ~new_new_n1031__;
  assign new_new_n16141__ = ~new_new_n1151__ & new_new_n16140__;
  assign new_new_n16142__ = ~new_new_n479__ & new_new_n1157__;
  assign new_new_n16143__ = new_new_n2064__ & new_new_n16142__;
  assign new_new_n16144__ = new_new_n4091__ & new_new_n16141__;
  assign new_new_n16145__ = new_new_n7746__ & new_new_n16144__;
  assign new_new_n16146__ = new_new_n16143__ & new_new_n16145__;
  assign new_new_n16147__ = ~new_new_n277__ & ~new_new_n1009__;
  assign new_new_n16148__ = ~new_new_n300__ & ~new_new_n896__;
  assign new_new_n16149__ = ~new_new_n76__ & ~new_new_n164__;
  assign new_new_n16150__ = ~new_new_n321__ & new_new_n16149__;
  assign new_new_n16151__ = new_new_n2712__ & new_new_n16150__;
  assign new_new_n16152__ = new_new_n16148__ & new_new_n16151__;
  assign new_new_n16153__ = ~new_new_n266__ & ~new_new_n939__;
  assign new_new_n16154__ = ~new_new_n1568__ & new_new_n16153__;
  assign new_new_n16155__ = new_new_n1945__ & new_new_n16147__;
  assign new_new_n16156__ = new_new_n16154__ & new_new_n16155__;
  assign new_new_n16157__ = new_new_n2912__ & new_new_n16156__;
  assign new_new_n16158__ = new_new_n16152__ & new_new_n16157__;
  assign new_new_n16159__ = new_new_n16146__ & new_new_n16158__;
  assign new_new_n16160__ = ~new_new_n837__ & new_new_n5412__;
  assign new_new_n16161__ = ~new_new_n213__ & ~new_new_n250__;
  assign new_new_n16162__ = ~new_new_n597__ & ~new_new_n845__;
  assign new_new_n16163__ = new_new_n16161__ & new_new_n16162__;
  assign new_new_n16164__ = ~new_new_n329__ & ~new_new_n566__;
  assign new_new_n16165__ = new_new_n2233__ & new_new_n16164__;
  assign new_new_n16166__ = new_new_n16163__ & new_new_n16165__;
  assign new_new_n16167__ = ~new_new_n130__ & ~new_new_n238__;
  assign new_new_n16168__ = ~new_new_n375__ & ~new_new_n950__;
  assign new_new_n16169__ = ~new_new_n1109__ & new_new_n16168__;
  assign new_new_n16170__ = ~new_new_n255__ & new_new_n16167__;
  assign new_new_n16171__ = ~new_new_n842__ & new_new_n1741__;
  assign new_new_n16172__ = new_new_n4342__ & new_new_n16171__;
  assign new_new_n16173__ = new_new_n16169__ & new_new_n16170__;
  assign new_new_n16174__ = new_new_n4949__ & new_new_n16173__;
  assign new_new_n16175__ = new_new_n16172__ & new_new_n16174__;
  assign new_new_n16176__ = new_new_n16160__ & new_new_n16166__;
  assign new_new_n16177__ = new_new_n16175__ & new_new_n16176__;
  assign new_new_n16178__ = new_new_n16127__ & new_new_n16139__;
  assign new_new_n16179__ = new_new_n16177__ & new_new_n16178__;
  assign new_new_n16180__ = new_new_n3237__ & new_new_n16179__;
  assign new_new_n16181__ = new_new_n16159__ & new_new_n16180__;
  assign new_new_n16182__ = pi17 & new_new_n9800__;
  assign new_new_n16183__ = ~pi17 & new_new_n9797__;
  assign new_new_n16184__ = ~pi20 & ~new_new_n16183__;
  assign new_new_n16185__ = ~new_new_n16182__ & ~new_new_n16184__;
  assign new_new_n16186__ = ~new_new_n16181__ & new_new_n16185__;
  assign new_new_n16187__ = new_new_n16181__ & ~new_new_n16185__;
  assign new_new_n16188__ = ~new_new_n238__ & ~new_new_n783__;
  assign new_new_n16189__ = ~new_new_n838__ & new_new_n16188__;
  assign new_new_n16190__ = ~new_new_n274__ & ~new_new_n631__;
  assign new_new_n16191__ = new_new_n1095__ & new_new_n3010__;
  assign new_new_n16192__ = new_new_n7155__ & new_new_n16191__;
  assign new_new_n16193__ = new_new_n16189__ & new_new_n16190__;
  assign new_new_n16194__ = new_new_n2175__ & new_new_n2548__;
  assign new_new_n16195__ = new_new_n3260__ & new_new_n6066__;
  assign new_new_n16196__ = new_new_n16194__ & new_new_n16195__;
  assign new_new_n16197__ = new_new_n16192__ & new_new_n16193__;
  assign new_new_n16198__ = ~new_new_n1539__ & new_new_n3208__;
  assign new_new_n16199__ = new_new_n4478__ & new_new_n16198__;
  assign new_new_n16200__ = new_new_n16196__ & new_new_n16197__;
  assign new_new_n16201__ = new_new_n3521__ & new_new_n16200__;
  assign new_new_n16202__ = new_new_n16199__ & new_new_n16201__;
  assign new_new_n16203__ = ~new_new_n91__ & ~new_new_n129__;
  assign new_new_n16204__ = new_new_n165__ & ~new_new_n16203__;
  assign new_new_n16205__ = ~new_new_n207__ & ~new_new_n624__;
  assign new_new_n16206__ = ~new_new_n715__ & new_new_n16205__;
  assign new_new_n16207__ = ~new_new_n1008__ & new_new_n1263__;
  assign new_new_n16208__ = ~new_new_n3566__ & ~new_new_n16204__;
  assign new_new_n16209__ = new_new_n16207__ & new_new_n16208__;
  assign new_new_n16210__ = ~new_new_n809__ & new_new_n16206__;
  assign new_new_n16211__ = new_new_n1216__ & new_new_n1331__;
  assign new_new_n16212__ = ~new_new_n1486__ & new_new_n16211__;
  assign new_new_n16213__ = new_new_n16209__ & new_new_n16210__;
  assign new_new_n16214__ = new_new_n7657__ & new_new_n16213__;
  assign new_new_n16215__ = new_new_n1579__ & new_new_n16212__;
  assign new_new_n16216__ = new_new_n16214__ & new_new_n16215__;
  assign new_new_n16217__ = new_new_n3273__ & new_new_n16216__;
  assign new_new_n16218__ = new_new_n2366__ & new_new_n16217__;
  assign new_new_n16219__ = new_new_n16202__ & new_new_n16218__;
  assign new_new_n16220__ = ~new_new_n16187__ & ~new_new_n16219__;
  assign new_new_n16221__ = ~new_new_n16186__ & ~new_new_n16220__;
  assign new_new_n16222__ = ~new_new_n16123__ & ~new_new_n16221__;
  assign new_new_n16223__ = ~new_new_n160__ & ~new_new_n207__;
  assign new_new_n16224__ = ~new_new_n247__ & ~new_new_n374__;
  assign new_new_n16225__ = ~new_new_n675__ & new_new_n16224__;
  assign new_new_n16226__ = ~new_new_n894__ & new_new_n1678__;
  assign new_new_n16227__ = new_new_n1903__ & new_new_n4720__;
  assign new_new_n16228__ = new_new_n4728__ & new_new_n16223__;
  assign new_new_n16229__ = new_new_n16227__ & new_new_n16228__;
  assign new_new_n16230__ = new_new_n16225__ & new_new_n16226__;
  assign new_new_n16231__ = new_new_n2324__ & new_new_n3294__;
  assign new_new_n16232__ = new_new_n4716__ & new_new_n16231__;
  assign new_new_n16233__ = new_new_n16229__ & new_new_n16230__;
  assign new_new_n16234__ = new_new_n16232__ & new_new_n16233__;
  assign new_new_n16235__ = ~new_new_n439__ & new_new_n3398__;
  assign new_new_n16236__ = ~new_new_n828__ & ~new_new_n871__;
  assign new_new_n16237__ = ~new_new_n508__ & ~new_new_n778__;
  assign new_new_n16238__ = ~new_new_n198__ & ~new_new_n884__;
  assign new_new_n16239__ = ~new_new_n82__ & ~new_new_n229__;
  assign new_new_n16240__ = ~new_new_n88__ & ~new_new_n874__;
  assign new_new_n16241__ = new_new_n3195__ & new_new_n16239__;
  assign new_new_n16242__ = new_new_n16240__ & new_new_n16241__;
  assign new_new_n16243__ = new_new_n589__ & new_new_n944__;
  assign new_new_n16244__ = new_new_n984__ & new_new_n1142__;
  assign new_new_n16245__ = new_new_n1680__ & new_new_n3637__;
  assign new_new_n16246__ = new_new_n16236__ & new_new_n16238__;
  assign new_new_n16247__ = new_new_n16245__ & new_new_n16246__;
  assign new_new_n16248__ = new_new_n16243__ & new_new_n16244__;
  assign new_new_n16249__ = new_new_n16235__ & new_new_n16242__;
  assign new_new_n16250__ = new_new_n16237__ & new_new_n16249__;
  assign new_new_n16251__ = new_new_n16247__ & new_new_n16248__;
  assign new_new_n16252__ = new_new_n16250__ & new_new_n16251__;
  assign new_new_n16253__ = new_new_n16234__ & new_new_n16252__;
  assign new_new_n16254__ = new_new_n5410__ & new_new_n16253__;
  assign new_new_n16255__ = new_new_n16159__ & new_new_n16254__;
  assign new_new_n16256__ = new_new_n16222__ & ~new_new_n16255__;
  assign new_new_n16257__ = new_new_n16100__ & ~new_new_n16256__;
  assign new_new_n16258__ = new_new_n16123__ & new_new_n16221__;
  assign new_new_n16259__ = new_new_n16255__ & new_new_n16258__;
  assign new_new_n16260__ = ~new_new_n16100__ & ~new_new_n16259__;
  assign new_new_n16261__ = ~new_new_n816__ & ~new_new_n853__;
  assign new_new_n16262__ = ~new_new_n316__ & new_new_n16261__;
  assign new_new_n16263__ = new_new_n1774__ & new_new_n16262__;
  assign new_new_n16264__ = new_new_n163__ & ~new_new_n1880__;
  assign new_new_n16265__ = ~new_new_n283__ & ~new_new_n508__;
  assign new_new_n16266__ = ~new_new_n16264__ & new_new_n16265__;
  assign new_new_n16267__ = ~new_new_n226__ & ~new_new_n698__;
  assign new_new_n16268__ = ~new_new_n276__ & ~new_new_n595__;
  assign new_new_n16269__ = ~new_new_n894__ & new_new_n16239__;
  assign new_new_n16270__ = new_new_n16268__ & new_new_n16269__;
  assign new_new_n16271__ = new_new_n4322__ & new_new_n16267__;
  assign new_new_n16272__ = new_new_n5457__ & new_new_n6143__;
  assign new_new_n16273__ = new_new_n16271__ & new_new_n16272__;
  assign new_new_n16274__ = new_new_n2092__ & new_new_n16270__;
  assign new_new_n16275__ = new_new_n16273__ & new_new_n16274__;
  assign new_new_n16276__ = new_new_n16263__ & new_new_n16266__;
  assign new_new_n16277__ = new_new_n16275__ & new_new_n16276__;
  assign new_new_n16278__ = new_new_n3325__ & new_new_n16277__;
  assign new_new_n16279__ = new_new_n1941__ & new_new_n16278__;
  assign new_new_n16280__ = new_new_n4715__ & new_new_n16279__;
  assign new_new_n16281__ = ~new_new_n16260__ & new_new_n16280__;
  assign new_new_n16282__ = ~new_new_n209__ & ~new_new_n495__;
  assign new_new_n16283__ = ~new_new_n298__ & ~new_new_n385__;
  assign new_new_n16284__ = ~new_new_n445__ & ~new_new_n632__;
  assign new_new_n16285__ = new_new_n16283__ & new_new_n16284__;
  assign new_new_n16286__ = ~new_new_n263__ & ~new_new_n959__;
  assign new_new_n16287__ = new_new_n1858__ & new_new_n16286__;
  assign new_new_n16288__ = ~new_new_n344__ & new_new_n16285__;
  assign new_new_n16289__ = new_new_n542__ & new_new_n2850__;
  assign new_new_n16290__ = new_new_n3059__ & new_new_n5303__;
  assign new_new_n16291__ = new_new_n16289__ & new_new_n16290__;
  assign new_new_n16292__ = new_new_n16287__ & new_new_n16288__;
  assign new_new_n16293__ = ~new_new_n668__ & new_new_n16292__;
  assign new_new_n16294__ = new_new_n16291__ & new_new_n16293__;
  assign new_new_n16295__ = new_new_n636__ & new_new_n1929__;
  assign new_new_n16296__ = new_new_n16236__ & new_new_n16295__;
  assign new_new_n16297__ = ~new_new_n235__ & ~new_new_n838__;
  assign new_new_n16298__ = ~new_new_n963__ & new_new_n16297__;
  assign new_new_n16299__ = ~new_new_n198__ & ~new_new_n277__;
  assign new_new_n16300__ = ~new_new_n329__ & ~new_new_n747__;
  assign new_new_n16301__ = new_new_n16299__ & new_new_n16300__;
  assign new_new_n16302__ = new_new_n3912__ & new_new_n16298__;
  assign new_new_n16303__ = new_new_n6070__ & new_new_n6211__;
  assign new_new_n16304__ = new_new_n16302__ & new_new_n16303__;
  assign new_new_n16305__ = new_new_n16301__ & new_new_n16304__;
  assign new_new_n16306__ = new_new_n7158__ & new_new_n16296__;
  assign new_new_n16307__ = new_new_n16305__ & new_new_n16306__;
  assign new_new_n16308__ = new_new_n5377__ & new_new_n16307__;
  assign new_new_n16309__ = ~new_new_n260__ & ~new_new_n693__;
  assign new_new_n16310__ = ~new_new_n785__ & new_new_n16309__;
  assign new_new_n16311__ = new_new_n1711__ & new_new_n2342__;
  assign new_new_n16312__ = new_new_n3794__ & new_new_n16311__;
  assign new_new_n16313__ = new_new_n1329__ & new_new_n16310__;
  assign new_new_n16314__ = new_new_n2142__ & new_new_n3419__;
  assign new_new_n16315__ = new_new_n6183__ & new_new_n16314__;
  assign new_new_n16316__ = new_new_n16312__ & new_new_n16313__;
  assign new_new_n16317__ = new_new_n1826__ & new_new_n16316__;
  assign new_new_n16318__ = new_new_n16315__ & new_new_n16317__;
  assign new_new_n16319__ = ~new_new_n346__ & ~new_new_n1515__;
  assign new_new_n16320__ = ~new_new_n721__ & ~new_new_n884__;
  assign new_new_n16321__ = new_new_n1368__ & ~new_new_n4316__;
  assign new_new_n16322__ = new_new_n6149__ & new_new_n16282__;
  assign new_new_n16323__ = new_new_n16321__ & new_new_n16322__;
  assign new_new_n16324__ = new_new_n16319__ & new_new_n16320__;
  assign new_new_n16325__ = new_new_n1114__ & new_new_n4963__;
  assign new_new_n16326__ = new_new_n16324__ & new_new_n16325__;
  assign new_new_n16327__ = new_new_n16237__ & new_new_n16323__;
  assign new_new_n16328__ = new_new_n16326__ & new_new_n16327__;
  assign new_new_n16329__ = new_new_n326__ & new_new_n16328__;
  assign new_new_n16330__ = new_new_n5622__ & new_new_n16329__;
  assign new_new_n16331__ = new_new_n16294__ & new_new_n16318__;
  assign new_new_n16332__ = new_new_n16330__ & new_new_n16331__;
  assign new_new_n16333__ = new_new_n16308__ & new_new_n16332__;
  assign new_new_n16334__ = ~new_new_n5188__ & ~new_new_n16333__;
  assign new_new_n16335__ = ~new_new_n5185__ & new_new_n16333__;
  assign new_new_n16336__ = ~new_new_n5195__ & ~new_new_n16334__;
  assign new_new_n16337__ = ~new_new_n16335__ & new_new_n16336__;
  assign new_new_n16338__ = ~new_new_n5185__ & ~new_new_n16333__;
  assign new_new_n16339__ = ~new_new_n5188__ & new_new_n16333__;
  assign new_new_n16340__ = ~new_new_n5195__ & ~new_new_n16338__;
  assign new_new_n16341__ = ~new_new_n16339__ & new_new_n16340__;
  assign new_new_n16342__ = pi23 & ~new_new_n16333__;
  assign new_new_n16343__ = ~pi23 & new_new_n16333__;
  assign new_new_n16344__ = ~new_new_n16342__ & ~new_new_n16343__;
  assign new_new_n16345__ = ~new_new_n16341__ & new_new_n16344__;
  assign new_new_n16346__ = ~new_new_n16337__ & ~new_new_n16345__;
  assign new_new_n16347__ = ~new_new_n16257__ & new_new_n16346__;
  assign new_new_n16348__ = ~new_new_n16281__ & new_new_n16347__;
  assign new_new_n16349__ = new_new_n16255__ & ~new_new_n16346__;
  assign new_new_n16350__ = ~new_new_n16100__ & new_new_n16222__;
  assign new_new_n16351__ = ~new_new_n16349__ & ~new_new_n16350__;
  assign new_new_n16352__ = new_new_n16100__ & new_new_n16258__;
  assign new_new_n16353__ = new_new_n16349__ & ~new_new_n16352__;
  assign new_new_n16354__ = new_new_n16280__ & ~new_new_n16353__;
  assign new_new_n16355__ = ~new_new_n16351__ & ~new_new_n16354__;
  assign new_new_n16356__ = ~new_new_n16348__ & ~new_new_n16355__;
  assign new_new_n16357__ = new_new_n4815__ & ~new_new_n15998__;
  assign new_new_n16358__ = new_new_n4212__ & new_new_n15905__;
  assign new_new_n16359__ = ~new_new_n4818__ & new_new_n15237__;
  assign new_new_n16360__ = new_new_n4813__ & new_new_n16025__;
  assign new_new_n16361__ = ~new_new_n16358__ & ~new_new_n16359__;
  assign new_new_n16362__ = ~new_new_n16357__ & new_new_n16361__;
  assign new_new_n16363__ = ~new_new_n16360__ & new_new_n16362__;
  assign new_new_n16364__ = pi29 & ~new_new_n16363__;
  assign new_new_n16365__ = ~pi29 & new_new_n16363__;
  assign new_new_n16366__ = ~new_new_n16364__ & ~new_new_n16365__;
  assign new_new_n16367__ = new_new_n16356__ & new_new_n16366__;
  assign new_new_n16368__ = new_new_n16333__ & new_new_n16346__;
  assign new_new_n16369__ = ~new_new_n16349__ & ~new_new_n16368__;
  assign new_new_n16370__ = new_new_n161__ & ~new_new_n15248__;
  assign new_new_n16371__ = new_new_n765__ & new_new_n15244__;
  assign new_new_n16372__ = ~new_new_n16370__ & ~new_new_n16371__;
  assign new_new_n16373__ = ~pi31 & ~new_new_n16372__;
  assign new_new_n16374__ = new_new_n71__ & ~new_new_n15248__;
  assign new_new_n16375__ = ~new_new_n15849__ & ~new_new_n15856__;
  assign new_new_n16376__ = new_new_n15248__ & new_new_n16375__;
  assign new_new_n16377__ = ~new_new_n15248__ & ~new_new_n16375__;
  assign new_new_n16378__ = ~new_new_n16376__ & ~new_new_n16377__;
  assign new_new_n16379__ = new_new_n765__ & new_new_n16378__;
  assign new_new_n16380__ = ~new_new_n16062__ & ~new_new_n16374__;
  assign new_new_n16381__ = ~new_new_n16379__ & new_new_n16380__;
  assign new_new_n16382__ = pi31 & ~new_new_n16381__;
  assign new_new_n16383__ = ~new_new_n16373__ & ~new_new_n16382__;
  assign new_new_n16384__ = new_new_n16369__ & ~new_new_n16383__;
  assign new_new_n16385__ = ~new_new_n15960__ & new_new_n16384__;
  assign new_new_n16386__ = ~new_new_n16367__ & new_new_n16385__;
  assign new_new_n16387__ = ~new_new_n16356__ & ~new_new_n16366__;
  assign new_new_n16388__ = ~new_new_n16369__ & new_new_n16383__;
  assign new_new_n16389__ = new_new_n15960__ & new_new_n16388__;
  assign new_new_n16390__ = ~new_new_n16387__ & new_new_n16389__;
  assign new_new_n16391__ = ~new_new_n16386__ & ~new_new_n16390__;
  assign new_new_n16392__ = ~new_new_n15874__ & ~new_new_n15925__;
  assign new_new_n16393__ = ~new_new_n16366__ & new_new_n16392__;
  assign new_new_n16394__ = new_new_n16366__ & ~new_new_n16392__;
  assign new_new_n16395__ = ~new_new_n16393__ & ~new_new_n16394__;
  assign new_new_n16396__ = ~new_new_n16391__ & new_new_n16395__;
  assign new_new_n16397__ = ~new_new_n16367__ & ~new_new_n16387__;
  assign new_new_n16398__ = ~new_new_n15960__ & ~new_new_n16388__;
  assign new_new_n16399__ = ~new_new_n16384__ & ~new_new_n16398__;
  assign new_new_n16400__ = new_new_n16392__ & ~new_new_n16399__;
  assign new_new_n16401__ = ~new_new_n16392__ & new_new_n16399__;
  assign new_new_n16402__ = ~new_new_n16400__ & ~new_new_n16401__;
  assign new_new_n16403__ = ~new_new_n16397__ & new_new_n16402__;
  assign new_new_n16404__ = ~new_new_n16385__ & ~new_new_n16389__;
  assign new_new_n16405__ = ~new_new_n16395__ & new_new_n16404__;
  assign new_new_n16406__ = new_new_n16397__ & new_new_n16405__;
  assign new_new_n16407__ = ~new_new_n16396__ & ~new_new_n16403__;
  assign new_new_n16408__ = ~new_new_n16406__ & new_new_n16407__;
  assign new_new_n16409__ = ~new_new_n16061__ & ~new_new_n16408__;
  assign new_new_n16410__ = new_new_n15929__ & ~new_new_n16409__;
  assign new_new_n16411__ = ~new_new_n15929__ & ~new_new_n16408__;
  assign new_new_n16412__ = pi29 & ~new_new_n16059__;
  assign new_new_n16413__ = ~new_new_n16060__ & ~new_new_n16412__;
  assign new_new_n16414__ = ~new_new_n3890__ & ~new_new_n16413__;
  assign new_new_n16415__ = ~new_new_n16411__ & new_new_n16414__;
  assign new_new_n16416__ = new_new_n4817__ & new_new_n15905__;
  assign new_new_n16417__ = new_new_n16408__ & new_new_n16416__;
  assign new_new_n16418__ = ~new_new_n16410__ & ~new_new_n16417__;
  assign new_new_n16419__ = ~new_new_n16415__ & new_new_n16418__;
  assign new_new_n16420__ = new_new_n873__ & ~new_new_n15998__;
  assign new_new_n16421__ = new_new_n550__ & new_new_n16051__;
  assign new_new_n16422__ = ~new_new_n110__ & ~new_new_n16056__;
  assign new_new_n16423__ = ~new_new_n16421__ & new_new_n16422__;
  assign new_new_n16424__ = ~new_new_n16420__ & ~new_new_n16423__;
  assign new_new_n16425__ = new_new_n303__ & new_new_n15905__;
  assign new_new_n16426__ = pi26 & ~new_new_n16425__;
  assign new_new_n16427__ = new_new_n145__ & new_new_n15905__;
  assign new_new_n16428__ = ~pi26 & ~new_new_n16427__;
  assign new_new_n16429__ = pi23 & ~new_new_n16428__;
  assign new_new_n16430__ = ~new_new_n16426__ & ~new_new_n16429__;
  assign new_new_n16431__ = new_new_n16424__ & ~new_new_n16430__;
  assign new_new_n16432__ = ~pi26 & ~new_new_n16424__;
  assign new_new_n16433__ = ~new_new_n16431__ & ~new_new_n16432__;
  assign new_new_n16434__ = new_new_n161__ & new_new_n15398__;
  assign new_new_n16435__ = ~new_new_n15321__ & ~new_new_n15829__;
  assign new_new_n16436__ = new_new_n15349__ & ~new_new_n15398__;
  assign new_new_n16437__ = new_new_n16435__ & new_new_n16436__;
  assign new_new_n16438__ = new_new_n15390__ & new_new_n15399__;
  assign new_new_n16439__ = ~new_new_n16437__ & ~new_new_n16438__;
  assign new_new_n16440__ = ~new_new_n15362__ & ~new_new_n16439__;
  assign new_new_n16441__ = ~new_new_n15390__ & ~new_new_n15398__;
  assign new_new_n16442__ = new_new_n15321__ & new_new_n16441__;
  assign new_new_n16443__ = ~new_new_n15349__ & new_new_n15398__;
  assign new_new_n16444__ = new_new_n16435__ & new_new_n16443__;
  assign new_new_n16445__ = ~new_new_n16442__ & ~new_new_n16444__;
  assign new_new_n16446__ = new_new_n15362__ & ~new_new_n16445__;
  assign new_new_n16447__ = new_new_n15390__ & new_new_n15398__;
  assign new_new_n16448__ = ~new_new_n16441__ & ~new_new_n16447__;
  assign new_new_n16449__ = new_new_n15829__ & ~new_new_n16448__;
  assign new_new_n16450__ = ~new_new_n15349__ & ~new_new_n15398__;
  assign new_new_n16451__ = ~new_new_n15836__ & ~new_new_n16450__;
  assign new_new_n16452__ = ~new_new_n16449__ & new_new_n16451__;
  assign new_new_n16453__ = new_new_n15321__ & ~new_new_n16452__;
  assign new_new_n16454__ = new_new_n16448__ & new_new_n16451__;
  assign new_new_n16455__ = ~new_new_n15321__ & new_new_n16454__;
  assign new_new_n16456__ = ~new_new_n16453__ & ~new_new_n16455__;
  assign new_new_n16457__ = ~new_new_n16440__ & new_new_n16456__;
  assign new_new_n16458__ = ~new_new_n16446__ & new_new_n16457__;
  assign new_new_n16459__ = new_new_n765__ & ~new_new_n16458__;
  assign new_new_n16460__ = ~new_new_n16434__ & ~new_new_n16459__;
  assign new_new_n16461__ = pi31 & ~new_new_n16460__;
  assign new_new_n16462__ = pi31 & ~new_new_n15349__;
  assign new_new_n16463__ = new_new_n71__ & ~new_new_n16462__;
  assign new_new_n16464__ = ~new_new_n161__ & ~new_new_n15321__;
  assign new_new_n16465__ = new_new_n161__ & ~new_new_n15349__;
  assign new_new_n16466__ = ~pi31 & ~new_new_n16465__;
  assign new_new_n16467__ = ~new_new_n16464__ & new_new_n16466__;
  assign new_new_n16468__ = ~new_new_n16463__ & ~new_new_n16467__;
  assign new_new_n16469__ = ~new_new_n16461__ & new_new_n16468__;
  assign new_new_n16470__ = ~new_new_n108__ & ~new_new_n585__;
  assign new_new_n16471__ = ~new_new_n940__ & ~new_new_n1073__;
  assign new_new_n16472__ = ~new_new_n127__ & ~new_new_n200__;
  assign new_new_n16473__ = ~new_new_n252__ & ~new_new_n723__;
  assign new_new_n16474__ = new_new_n16472__ & new_new_n16473__;
  assign new_new_n16475__ = ~new_new_n280__ & ~new_new_n317__;
  assign new_new_n16476__ = ~new_new_n329__ & ~new_new_n372__;
  assign new_new_n16477__ = new_new_n3209__ & new_new_n16470__;
  assign new_new_n16478__ = new_new_n16476__ & new_new_n16477__;
  assign new_new_n16479__ = new_new_n16474__ & new_new_n16475__;
  assign new_new_n16480__ = ~new_new_n508__ & new_new_n16471__;
  assign new_new_n16481__ = new_new_n16479__ & new_new_n16480__;
  assign new_new_n16482__ = new_new_n1079__ & new_new_n16478__;
  assign new_new_n16483__ = new_new_n2764__ & new_new_n6090__;
  assign new_new_n16484__ = new_new_n16482__ & new_new_n16483__;
  assign new_new_n16485__ = new_new_n2475__ & new_new_n16481__;
  assign new_new_n16486__ = new_new_n16484__ & new_new_n16485__;
  assign new_new_n16487__ = ~new_new_n247__ & ~new_new_n694__;
  assign new_new_n16488__ = ~new_new_n942__ & new_new_n1285__;
  assign new_new_n16489__ = new_new_n2428__ & new_new_n16488__;
  assign new_new_n16490__ = ~new_new_n388__ & ~new_new_n715__;
  assign new_new_n16491__ = ~new_new_n1031__ & new_new_n16490__;
  assign new_new_n16492__ = ~new_new_n602__ & ~new_new_n816__;
  assign new_new_n16493__ = new_new_n16487__ & new_new_n16492__;
  assign new_new_n16494__ = ~new_new_n254__ & new_new_n16491__;
  assign new_new_n16495__ = new_new_n1096__ & new_new_n1961__;
  assign new_new_n16496__ = new_new_n2377__ & new_new_n2653__;
  assign new_new_n16497__ = new_new_n3911__ & new_new_n16496__;
  assign new_new_n16498__ = new_new_n16494__ & new_new_n16495__;
  assign new_new_n16499__ = new_new_n1771__ & new_new_n16493__;
  assign new_new_n16500__ = new_new_n16498__ & new_new_n16499__;
  assign new_new_n16501__ = new_new_n609__ & new_new_n16497__;
  assign new_new_n16502__ = new_new_n16489__ & new_new_n16501__;
  assign new_new_n16503__ = new_new_n2464__ & new_new_n16500__;
  assign new_new_n16504__ = new_new_n16502__ & new_new_n16503__;
  assign new_new_n16505__ = new_new_n16486__ & new_new_n16504__;
  assign new_new_n16506__ = new_new_n6271__ & new_new_n16505__;
  assign new_new_n16507__ = ~new_new_n16469__ & new_new_n16506__;
  assign new_new_n16508__ = new_new_n16469__ & ~new_new_n16506__;
  assign new_new_n16509__ = ~new_new_n16507__ & ~new_new_n16508__;
  assign new_new_n16510__ = ~new_new_n16181__ & new_new_n16469__;
  assign new_new_n16511__ = new_new_n16181__ & ~new_new_n16469__;
  assign new_new_n16512__ = ~new_new_n16510__ & ~new_new_n16511__;
  assign new_new_n16513__ = ~new_new_n3221__ & new_new_n16469__;
  assign new_new_n16514__ = new_new_n16512__ & ~new_new_n16513__;
  assign new_new_n16515__ = new_new_n161__ & new_new_n16462__;
  assign new_new_n16516__ = ~new_new_n16072__ & ~new_new_n16073__;
  assign new_new_n16517__ = new_new_n15321__ & new_new_n16516__;
  assign new_new_n16518__ = pi31 & ~new_new_n16517__;
  assign new_new_n16519__ = ~pi31 & new_new_n15273__;
  assign new_new_n16520__ = ~new_new_n15853__ & ~new_new_n16519__;
  assign new_new_n16521__ = ~new_new_n16518__ & new_new_n16520__;
  assign new_new_n16522__ = ~new_new_n15853__ & new_new_n16516__;
  assign new_new_n16523__ = new_new_n8646__ & ~new_new_n15321__;
  assign new_new_n16524__ = ~new_new_n16522__ & new_new_n16523__;
  assign new_new_n16525__ = ~new_new_n16515__ & ~new_new_n16524__;
  assign new_new_n16526__ = ~new_new_n16521__ & new_new_n16525__;
  assign new_new_n16527__ = new_new_n16219__ & ~new_new_n16526__;
  assign new_new_n16528__ = ~new_new_n16219__ & new_new_n16526__;
  assign new_new_n16529__ = ~new_new_n16527__ & ~new_new_n16528__;
  assign new_new_n16530__ = ~new_new_n16185__ & new_new_n16529__;
  assign new_new_n16531__ = new_new_n16185__ & ~new_new_n16529__;
  assign new_new_n16532__ = ~new_new_n16530__ & ~new_new_n16531__;
  assign new_new_n16533__ = ~new_new_n16509__ & ~new_new_n16514__;
  assign new_new_n16534__ = new_new_n16532__ & new_new_n16533__;
  assign new_new_n16535__ = ~new_new_n16509__ & ~new_new_n16512__;
  assign new_new_n16536__ = ~new_new_n16532__ & ~new_new_n16535__;
  assign new_new_n16537__ = ~new_new_n16534__ & ~new_new_n16536__;
  assign new_new_n16538__ = new_new_n16507__ & ~new_new_n16537__;
  assign new_new_n16539__ = ~new_new_n16221__ & new_new_n16508__;
  assign new_new_n16540__ = new_new_n16526__ & new_new_n16539__;
  assign new_new_n16541__ = ~new_new_n16538__ & ~new_new_n16540__;
  assign new_new_n16542__ = new_new_n16181__ & ~new_new_n16541__;
  assign new_new_n16543__ = new_new_n16506__ & new_new_n16510__;
  assign new_new_n16544__ = ~new_new_n16221__ & ~new_new_n16469__;
  assign new_new_n16545__ = ~new_new_n16526__ & ~new_new_n16544__;
  assign new_new_n16546__ = ~new_new_n16543__ & new_new_n16545__;
  assign new_new_n16547__ = ~new_new_n16181__ & ~new_new_n16221__;
  assign new_new_n16548__ = ~new_new_n16508__ & new_new_n16547__;
  assign new_new_n16549__ = ~new_new_n16507__ & ~new_new_n16548__;
  assign new_new_n16550__ = new_new_n16526__ & ~new_new_n16549__;
  assign new_new_n16551__ = new_new_n16537__ & ~new_new_n16550__;
  assign new_new_n16552__ = ~new_new_n16546__ & ~new_new_n16551__;
  assign new_new_n16553__ = ~new_new_n16542__ & ~new_new_n16552__;
  assign new_new_n16554__ = ~new_new_n4818__ & ~new_new_n15314__;
  assign new_new_n16555__ = new_new_n4212__ & ~new_new_n15248__;
  assign new_new_n16556__ = new_new_n4815__ & new_new_n15244__;
  assign new_new_n16557__ = ~new_new_n16554__ & ~new_new_n16555__;
  assign new_new_n16558__ = ~new_new_n16556__ & new_new_n16557__;
  assign new_new_n16559__ = new_new_n4214__ & new_new_n16378__;
  assign new_new_n16560__ = ~pi29 & ~new_new_n16559__;
  assign new_new_n16561__ = new_new_n5732__ & new_new_n16378__;
  assign new_new_n16562__ = ~new_new_n16560__ & ~new_new_n16561__;
  assign new_new_n16563__ = new_new_n16558__ & ~new_new_n16562__;
  assign new_new_n16564__ = pi29 & ~new_new_n16558__;
  assign new_new_n16565__ = ~new_new_n16563__ & ~new_new_n16564__;
  assign new_new_n16566__ = ~new_new_n16553__ & ~new_new_n16565__;
  assign new_new_n16567__ = new_new_n16553__ & new_new_n16565__;
  assign new_new_n16568__ = ~new_new_n16222__ & ~new_new_n16258__;
  assign new_new_n16569__ = new_new_n16280__ & ~new_new_n16568__;
  assign new_new_n16570__ = ~new_new_n16280__ & new_new_n16568__;
  assign new_new_n16571__ = ~new_new_n16569__ & ~new_new_n16570__;
  assign new_new_n16572__ = ~new_new_n16567__ & new_new_n16571__;
  assign new_new_n16573__ = ~new_new_n16566__ & ~new_new_n16572__;
  assign new_new_n16574__ = ~new_new_n16433__ & new_new_n16573__;
  assign new_new_n16575__ = new_new_n16433__ & ~new_new_n16573__;
  assign new_new_n16576__ = new_new_n15273__ & new_new_n15314__;
  assign new_new_n16577__ = new_new_n16078__ & new_new_n16576__;
  assign new_new_n16578__ = ~new_new_n71__ & ~new_new_n16577__;
  assign new_new_n16579__ = new_new_n16087__ & ~new_new_n16578__;
  assign new_new_n16580__ = ~new_new_n15285__ & new_new_n15314__;
  assign new_new_n16581__ = ~new_new_n16078__ & new_new_n16580__;
  assign new_new_n16582__ = ~new_new_n161__ & ~new_new_n16581__;
  assign new_new_n16583__ = ~new_new_n71__ & ~new_new_n15273__;
  assign new_new_n16584__ = ~new_new_n16582__ & new_new_n16583__;
  assign new_new_n16585__ = new_new_n15853__ & ~new_new_n16068__;
  assign new_new_n16586__ = ~new_new_n15314__ & ~new_new_n16585__;
  assign new_new_n16587__ = ~new_new_n16082__ & new_new_n16586__;
  assign new_new_n16588__ = ~new_new_n16579__ & ~new_new_n16584__;
  assign new_new_n16589__ = ~new_new_n16587__ & new_new_n16588__;
  assign new_new_n16590__ = pi31 & ~new_new_n16589__;
  assign new_new_n16591__ = new_new_n161__ & new_new_n15285__;
  assign new_new_n16592__ = new_new_n765__ & ~new_new_n15314__;
  assign new_new_n16593__ = ~new_new_n16591__ & ~new_new_n16592__;
  assign new_new_n16594__ = ~pi31 & ~new_new_n16593__;
  assign new_new_n16595__ = ~new_new_n16590__ & ~new_new_n16594__;
  assign new_new_n16596__ = new_new_n4815__ & new_new_n15237__;
  assign new_new_n16597__ = ~new_new_n4818__ & ~new_new_n15248__;
  assign new_new_n16598__ = new_new_n4212__ & new_new_n15244__;
  assign new_new_n16599__ = ~new_new_n16597__ & ~new_new_n16598__;
  assign new_new_n16600__ = ~new_new_n16596__ & new_new_n16599__;
  assign new_new_n16601__ = new_new_n15237__ & ~new_new_n15851__;
  assign new_new_n16602__ = ~new_new_n15237__ & new_new_n15851__;
  assign new_new_n16603__ = ~new_new_n16601__ & ~new_new_n16602__;
  assign new_new_n16604__ = new_new_n4214__ & ~new_new_n16603__;
  assign new_new_n16605__ = pi29 & ~new_new_n16604__;
  assign new_new_n16606__ = new_new_n4825__ & ~new_new_n16603__;
  assign new_new_n16607__ = ~new_new_n16605__ & ~new_new_n16606__;
  assign new_new_n16608__ = new_new_n16600__ & ~new_new_n16607__;
  assign new_new_n16609__ = ~pi29 & ~new_new_n16600__;
  assign new_new_n16610__ = ~new_new_n16608__ & ~new_new_n16609__;
  assign new_new_n16611__ = ~new_new_n16258__ & new_new_n16280__;
  assign new_new_n16612__ = ~new_new_n16222__ & ~new_new_n16280__;
  assign new_new_n16613__ = ~new_new_n16611__ & ~new_new_n16612__;
  assign new_new_n16614__ = new_new_n16255__ & ~new_new_n16613__;
  assign new_new_n16615__ = ~new_new_n16255__ & new_new_n16613__;
  assign new_new_n16616__ = ~new_new_n16614__ & ~new_new_n16615__;
  assign new_new_n16617__ = ~new_new_n16610__ & new_new_n16616__;
  assign new_new_n16618__ = new_new_n16610__ & ~new_new_n16616__;
  assign new_new_n16619__ = ~new_new_n16617__ & ~new_new_n16618__;
  assign new_new_n16620__ = new_new_n16595__ & new_new_n16619__;
  assign new_new_n16621__ = ~new_new_n16595__ & ~new_new_n16619__;
  assign new_new_n16622__ = ~new_new_n16620__ & ~new_new_n16621__;
  assign new_new_n16623__ = ~new_new_n16575__ & ~new_new_n16622__;
  assign new_new_n16624__ = ~new_new_n16574__ & ~new_new_n16623__;
  assign new_new_n16625__ = pi26 & ~new_new_n16624__;
  assign new_new_n16626__ = ~pi26 & new_new_n16624__;
  assign new_new_n16627__ = ~new_new_n16625__ & ~new_new_n16626__;
  assign new_new_n16628__ = new_new_n873__ & ~new_new_n16056__;
  assign new_new_n16629__ = ~new_new_n333__ & ~new_new_n15998__;
  assign new_new_n16630__ = ~new_new_n16048__ & ~new_new_n16056__;
  assign new_new_n16631__ = new_new_n550__ & ~new_new_n16630__;
  assign new_new_n16632__ = new_new_n801__ & ~new_new_n16631__;
  assign new_new_n16633__ = ~new_new_n16628__ & ~new_new_n16629__;
  assign new_new_n16634__ = ~new_new_n16632__ & new_new_n16633__;
  assign new_new_n16635__ = new_new_n4815__ & new_new_n15905__;
  assign new_new_n16636__ = ~new_new_n4818__ & new_new_n15244__;
  assign new_new_n16637__ = new_new_n4212__ & new_new_n15237__;
  assign new_new_n16638__ = new_new_n4813__ & ~new_new_n15917__;
  assign new_new_n16639__ = ~new_new_n16636__ & ~new_new_n16637__;
  assign new_new_n16640__ = ~new_new_n16635__ & new_new_n16639__;
  assign new_new_n16641__ = ~new_new_n16638__ & new_new_n16640__;
  assign new_new_n16642__ = ~pi29 & new_new_n16641__;
  assign new_new_n16643__ = pi29 & ~new_new_n16641__;
  assign new_new_n16644__ = ~new_new_n16642__ & ~new_new_n16643__;
  assign new_new_n16645__ = ~new_new_n16255__ & ~new_new_n16280__;
  assign new_new_n16646__ = ~new_new_n16259__ & ~new_new_n16645__;
  assign new_new_n16647__ = ~new_new_n16612__ & ~new_new_n16646__;
  assign new_new_n16648__ = new_new_n16100__ & ~new_new_n16346__;
  assign new_new_n16649__ = ~new_new_n16100__ & new_new_n16346__;
  assign new_new_n16650__ = ~new_new_n16648__ & ~new_new_n16649__;
  assign new_new_n16651__ = new_new_n16647__ & new_new_n16650__;
  assign new_new_n16652__ = ~new_new_n16647__ & ~new_new_n16650__;
  assign new_new_n16653__ = ~new_new_n16651__ & ~new_new_n16652__;
  assign new_new_n16654__ = ~new_new_n16644__ & ~new_new_n16653__;
  assign new_new_n16655__ = new_new_n16644__ & new_new_n16653__;
  assign new_new_n16656__ = ~new_new_n16654__ & ~new_new_n16655__;
  assign new_new_n16657__ = ~new_new_n16595__ & ~new_new_n16618__;
  assign new_new_n16658__ = ~new_new_n16617__ & ~new_new_n16657__;
  assign new_new_n16659__ = new_new_n16656__ & new_new_n16658__;
  assign new_new_n16660__ = ~new_new_n16656__ & ~new_new_n16658__;
  assign new_new_n16661__ = ~new_new_n16659__ & ~new_new_n16660__;
  assign new_new_n16662__ = new_new_n16634__ & ~new_new_n16661__;
  assign new_new_n16663__ = ~new_new_n16634__ & new_new_n16661__;
  assign new_new_n16664__ = ~new_new_n16662__ & ~new_new_n16663__;
  assign new_new_n16665__ = new_new_n16627__ & new_new_n16664__;
  assign new_new_n16666__ = ~new_new_n16627__ & ~new_new_n16664__;
  assign new_new_n16667__ = ~new_new_n16665__ & ~new_new_n16666__;
  assign new_new_n16668__ = ~new_new_n16574__ & ~new_new_n16575__;
  assign new_new_n16669__ = ~new_new_n16622__ & new_new_n16668__;
  assign new_new_n16670__ = new_new_n16622__ & ~new_new_n16668__;
  assign new_new_n16671__ = ~new_new_n16669__ & ~new_new_n16670__;
  assign new_new_n16672__ = ~new_new_n333__ & new_new_n15237__;
  assign new_new_n16673__ = new_new_n873__ & new_new_n15905__;
  assign new_new_n16674__ = ~new_new_n16672__ & ~new_new_n16673__;
  assign new_new_n16675__ = ~new_new_n110__ & ~new_new_n15998__;
  assign new_new_n16676__ = new_new_n16025__ & new_new_n16675__;
  assign new_new_n16677__ = new_new_n16674__ & ~new_new_n16676__;
  assign new_new_n16678__ = pi26 & ~new_new_n16677__;
  assign new_new_n16679__ = new_new_n15998__ & ~new_new_n16025__;
  assign new_new_n16680__ = new_new_n801__ & ~new_new_n16679__;
  assign new_new_n16681__ = ~pi26 & ~new_new_n16680__;
  assign new_new_n16682__ = new_new_n15998__ & new_new_n16025__;
  assign new_new_n16683__ = ~pi25 & ~new_new_n16682__;
  assign new_new_n16684__ = ~new_new_n15998__ & ~new_new_n16024__;
  assign new_new_n16685__ = pi25 & ~new_new_n16684__;
  assign new_new_n16686__ = ~new_new_n110__ & ~new_new_n16685__;
  assign new_new_n16687__ = ~new_new_n16683__ & new_new_n16686__;
  assign new_new_n16688__ = ~new_new_n16681__ & ~new_new_n16687__;
  assign new_new_n16689__ = new_new_n16674__ & ~new_new_n16688__;
  assign new_new_n16690__ = ~new_new_n16678__ & ~new_new_n16689__;
  assign new_new_n16691__ = ~new_new_n16566__ & ~new_new_n16567__;
  assign new_new_n16692__ = ~new_new_n16571__ & new_new_n16691__;
  assign new_new_n16693__ = new_new_n16571__ & ~new_new_n16691__;
  assign new_new_n16694__ = ~new_new_n16692__ & ~new_new_n16693__;
  assign new_new_n16695__ = new_new_n16690__ & new_new_n16694__;
  assign new_new_n16696__ = ~new_new_n16690__ & ~new_new_n16694__;
  assign new_new_n16697__ = new_new_n4212__ & ~new_new_n15314__;
  assign new_new_n16698__ = ~new_new_n4818__ & new_new_n15285__;
  assign new_new_n16699__ = new_new_n4815__ & ~new_new_n15248__;
  assign new_new_n16700__ = ~new_new_n16697__ & ~new_new_n16698__;
  assign new_new_n16701__ = ~new_new_n16699__ & new_new_n16700__;
  assign new_new_n16702__ = new_new_n15248__ & new_new_n15285__;
  assign new_new_n16703__ = new_new_n15273__ & new_new_n16702__;
  assign new_new_n16704__ = ~new_new_n15285__ & new_new_n15325__;
  assign new_new_n16705__ = ~new_new_n15839__ & new_new_n16704__;
  assign new_new_n16706__ = ~new_new_n16703__ & ~new_new_n16705__;
  assign new_new_n16707__ = new_new_n15321__ & ~new_new_n16706__;
  assign new_new_n16708__ = new_new_n15248__ & ~new_new_n15285__;
  assign new_new_n16709__ = ~new_new_n15273__ & new_new_n16708__;
  assign new_new_n16710__ = new_new_n15286__ & new_new_n15314__;
  assign new_new_n16711__ = new_new_n15839__ & new_new_n16710__;
  assign new_new_n16712__ = ~new_new_n16709__ & ~new_new_n16711__;
  assign new_new_n16713__ = ~new_new_n15321__ & ~new_new_n16712__;
  assign new_new_n16714__ = ~new_new_n15839__ & new_new_n16702__;
  assign new_new_n16715__ = ~new_new_n16704__ & ~new_new_n16714__;
  assign new_new_n16716__ = new_new_n15273__ & ~new_new_n16715__;
  assign new_new_n16717__ = new_new_n15839__ & new_new_n16708__;
  assign new_new_n16718__ = ~new_new_n16710__ & ~new_new_n16717__;
  assign new_new_n16719__ = ~new_new_n15273__ & ~new_new_n16718__;
  assign new_new_n16720__ = ~new_new_n15844__ & ~new_new_n16580__;
  assign new_new_n16721__ = new_new_n15248__ & ~new_new_n16720__;
  assign new_new_n16722__ = ~new_new_n16716__ & ~new_new_n16721__;
  assign new_new_n16723__ = ~new_new_n16719__ & new_new_n16722__;
  assign new_new_n16724__ = ~new_new_n16707__ & ~new_new_n16713__;
  assign new_new_n16725__ = new_new_n16723__ & new_new_n16724__;
  assign new_new_n16726__ = new_new_n4214__ & new_new_n16725__;
  assign new_new_n16727__ = pi29 & ~new_new_n16726__;
  assign new_new_n16728__ = new_new_n4825__ & new_new_n16725__;
  assign new_new_n16729__ = ~new_new_n16727__ & ~new_new_n16728__;
  assign new_new_n16730__ = new_new_n16701__ & ~new_new_n16729__;
  assign new_new_n16731__ = ~pi29 & ~new_new_n16701__;
  assign new_new_n16732__ = ~new_new_n16730__ & ~new_new_n16731__;
  assign new_new_n16733__ = new_new_n161__ & new_new_n15390__;
  assign new_new_n16734__ = new_new_n765__ & ~new_new_n15398__;
  assign new_new_n16735__ = ~new_new_n16733__ & ~new_new_n16734__;
  assign new_new_n16736__ = ~pi31 & ~new_new_n16735__;
  assign new_new_n16737__ = ~pi29 & new_new_n15362__;
  assign new_new_n16738__ = new_new_n16441__ & new_new_n16737__;
  assign new_new_n16739__ = ~new_new_n15398__ & new_new_n15829__;
  assign new_new_n16740__ = new_new_n15398__ & ~new_new_n15829__;
  assign new_new_n16741__ = ~new_new_n16739__ & ~new_new_n16740__;
  assign new_new_n16742__ = ~new_new_n15362__ & ~new_new_n16447__;
  assign new_new_n16743__ = ~new_new_n16741__ & new_new_n16742__;
  assign new_new_n16744__ = ~new_new_n16738__ & ~new_new_n16743__;
  assign new_new_n16745__ = pi30 & ~new_new_n16744__;
  assign new_new_n16746__ = ~pi30 & new_new_n15362__;
  assign new_new_n16747__ = ~new_new_n16740__ & ~new_new_n16746__;
  assign new_new_n16748__ = ~new_new_n15362__ & ~new_new_n15390__;
  assign new_new_n16749__ = ~new_new_n16441__ & ~new_new_n16748__;
  assign new_new_n16750__ = ~new_new_n16747__ & ~new_new_n16749__;
  assign new_new_n16751__ = ~pi30 & ~new_new_n16739__;
  assign new_new_n16752__ = ~new_new_n15362__ & ~new_new_n16751__;
  assign new_new_n16753__ = ~new_new_n16750__ & ~new_new_n16752__;
  assign new_new_n16754__ = pi29 & ~new_new_n16753__;
  assign new_new_n16755__ = new_new_n15398__ & new_new_n15826__;
  assign new_new_n16756__ = ~new_new_n16739__ & ~new_new_n16755__;
  assign new_new_n16757__ = ~new_new_n161__ & ~new_new_n16756__;
  assign new_new_n16758__ = ~new_new_n15362__ & ~new_new_n15398__;
  assign new_new_n16759__ = ~new_new_n71__ & ~new_new_n16758__;
  assign new_new_n16760__ = ~new_new_n16757__ & new_new_n16759__;
  assign new_new_n16761__ = new_new_n15390__ & ~new_new_n16760__;
  assign new_new_n16762__ = ~new_new_n16745__ & ~new_new_n16754__;
  assign new_new_n16763__ = ~new_new_n16761__ & new_new_n16762__;
  assign new_new_n16764__ = pi31 & ~new_new_n16763__;
  assign new_new_n16765__ = ~new_new_n16736__ & ~new_new_n16764__;
  assign new_new_n16766__ = new_new_n71__ & new_new_n15432__;
  assign new_new_n16767__ = new_new_n161__ & new_new_n15439__;
  assign new_new_n16768__ = ~new_new_n15825__ & ~new_new_n15827__;
  assign new_new_n16769__ = new_new_n15362__ & ~new_new_n16768__;
  assign new_new_n16770__ = ~new_new_n15362__ & new_new_n16768__;
  assign new_new_n16771__ = ~new_new_n16769__ & ~new_new_n16770__;
  assign new_new_n16772__ = new_new_n765__ & ~new_new_n16771__;
  assign new_new_n16773__ = ~new_new_n16767__ & ~new_new_n16772__;
  assign new_new_n16774__ = pi31 & ~new_new_n16773__;
  assign new_new_n16775__ = pi29 & ~new_new_n15432__;
  assign new_new_n16776__ = new_new_n15853__ & ~new_new_n16775__;
  assign new_new_n16777__ = ~new_new_n16737__ & ~new_new_n16776__;
  assign new_new_n16778__ = ~new_new_n16746__ & new_new_n16777__;
  assign new_new_n16779__ = ~pi31 & ~new_new_n16778__;
  assign new_new_n16780__ = ~new_new_n16766__ & ~new_new_n16779__;
  assign new_new_n16781__ = ~new_new_n16774__ & new_new_n16780__;
  assign new_new_n16782__ = ~new_new_n783__ & ~new_new_n1515__;
  assign new_new_n16783__ = ~new_new_n300__ & new_new_n16782__;
  assign new_new_n16784__ = new_new_n3193__ & new_new_n3638__;
  assign new_new_n16785__ = new_new_n16783__ & new_new_n16784__;
  assign new_new_n16786__ = new_new_n997__ & new_new_n3280__;
  assign new_new_n16787__ = new_new_n16785__ & new_new_n16786__;
  assign new_new_n16788__ = new_new_n850__ & new_new_n1566__;
  assign new_new_n16789__ = new_new_n16787__ & new_new_n16788__;
  assign new_new_n16790__ = ~new_new_n263__ & ~new_new_n842__;
  assign new_new_n16791__ = ~new_new_n383__ & new_new_n16471__;
  assign new_new_n16792__ = new_new_n16308__ & new_new_n16791__;
  assign new_new_n16793__ = ~new_new_n723__ & ~new_new_n1151__;
  assign new_new_n16794__ = ~new_new_n103__ & ~new_new_n374__;
  assign new_new_n16795__ = ~new_new_n1070__ & new_new_n16794__;
  assign new_new_n16796__ = ~new_new_n321__ & ~new_new_n566__;
  assign new_new_n16797__ = ~new_new_n1064__ & new_new_n1214__;
  assign new_new_n16798__ = ~new_new_n1506__ & new_new_n2158__;
  assign new_new_n16799__ = new_new_n16797__ & new_new_n16798__;
  assign new_new_n16800__ = new_new_n16795__ & new_new_n16796__;
  assign new_new_n16801__ = new_new_n2439__ & new_new_n2992__;
  assign new_new_n16802__ = new_new_n16790__ & new_new_n16793__;
  assign new_new_n16803__ = new_new_n16801__ & new_new_n16802__;
  assign new_new_n16804__ = new_new_n16799__ & new_new_n16800__;
  assign new_new_n16805__ = ~new_new_n1539__ & new_new_n16804__;
  assign new_new_n16806__ = new_new_n3955__ & new_new_n16803__;
  assign new_new_n16807__ = new_new_n16805__ & new_new_n16806__;
  assign new_new_n16808__ = new_new_n16789__ & new_new_n16807__;
  assign new_new_n16809__ = new_new_n3338__ & new_new_n16808__;
  assign new_new_n16810__ = new_new_n16792__ & new_new_n16809__;
  assign new_new_n16811__ = new_new_n16781__ & ~new_new_n16810__;
  assign new_new_n16812__ = ~new_new_n232__ & ~new_new_n826__;
  assign new_new_n16813__ = ~new_new_n896__ & ~new_new_n921__;
  assign new_new_n16814__ = ~new_new_n1008__ & ~new_new_n1009__;
  assign new_new_n16815__ = new_new_n16813__ & new_new_n16814__;
  assign new_new_n16816__ = new_new_n2032__ & new_new_n16815__;
  assign new_new_n16817__ = ~new_new_n164__ & ~new_new_n990__;
  assign new_new_n16818__ = ~new_new_n473__ & ~new_new_n749__;
  assign new_new_n16819__ = ~new_new_n1398__ & ~new_new_n1515__;
  assign new_new_n16820__ = new_new_n16818__ & new_new_n16819__;
  assign new_new_n16821__ = ~new_new_n189__ & new_new_n1309__;
  assign new_new_n16822__ = new_new_n2426__ & new_new_n5413__;
  assign new_new_n16823__ = new_new_n6321__ & new_new_n16817__;
  assign new_new_n16824__ = new_new_n16822__ & new_new_n16823__;
  assign new_new_n16825__ = new_new_n16820__ & new_new_n16821__;
  assign new_new_n16826__ = new_new_n592__ & new_new_n962__;
  assign new_new_n16827__ = new_new_n1295__ & new_new_n1450__;
  assign new_new_n16828__ = new_new_n16812__ & new_new_n16827__;
  assign new_new_n16829__ = new_new_n16825__ & new_new_n16826__;
  assign new_new_n16830__ = new_new_n2089__ & new_new_n16824__;
  assign new_new_n16831__ = new_new_n16829__ & new_new_n16830__;
  assign new_new_n16832__ = new_new_n669__ & new_new_n16828__;
  assign new_new_n16833__ = new_new_n16816__ & new_new_n16832__;
  assign new_new_n16834__ = new_new_n6164__ & new_new_n16831__;
  assign new_new_n16835__ = new_new_n16833__ & new_new_n16834__;
  assign new_new_n16836__ = new_new_n3384__ & new_new_n16835__;
  assign new_new_n16837__ = new_new_n4436__ & new_new_n16836__;
  assign new_new_n16838__ = new_new_n16811__ & ~new_new_n16837__;
  assign new_new_n16839__ = new_new_n16765__ & ~new_new_n16838__;
  assign new_new_n16840__ = new_new_n16810__ & new_new_n16837__;
  assign new_new_n16841__ = ~new_new_n16781__ & new_new_n16840__;
  assign new_new_n16842__ = ~new_new_n16765__ & ~new_new_n16841__;
  assign new_new_n16843__ = ~pi14 & ~new_new_n6989__;
  assign new_new_n16844__ = ~new_new_n6987__ & ~new_new_n16843__;
  assign new_new_n16845__ = ~new_new_n388__ & ~new_new_n510__;
  assign new_new_n16846__ = ~new_new_n1212__ & new_new_n16845__;
  assign new_new_n16847__ = ~new_new_n1073__ & new_new_n1859__;
  assign new_new_n16848__ = new_new_n2116__ & new_new_n16847__;
  assign new_new_n16849__ = new_new_n16846__ & new_new_n16848__;
  assign new_new_n16850__ = new_new_n67__ & ~new_new_n15853__;
  assign new_new_n16851__ = new_new_n100__ & new_new_n16850__;
  assign new_new_n16852__ = ~new_new_n1070__ & new_new_n1366__;
  assign new_new_n16853__ = ~new_new_n379__ & ~new_new_n2170__;
  assign new_new_n16854__ = ~new_new_n192__ & new_new_n16853__;
  assign new_new_n16855__ = ~new_new_n280__ & ~new_new_n781__;
  assign new_new_n16856__ = new_new_n1368__ & ~new_new_n16851__;
  assign new_new_n16857__ = new_new_n16855__ & new_new_n16856__;
  assign new_new_n16858__ = new_new_n2771__ & new_new_n16854__;
  assign new_new_n16859__ = new_new_n5365__ & new_new_n5415__;
  assign new_new_n16860__ = new_new_n16852__ & new_new_n16859__;
  assign new_new_n16861__ = new_new_n16857__ & new_new_n16858__;
  assign new_new_n16862__ = new_new_n2990__ & new_new_n3586__;
  assign new_new_n16863__ = new_new_n16861__ & new_new_n16862__;
  assign new_new_n16864__ = new_new_n1229__ & new_new_n16860__;
  assign new_new_n16865__ = new_new_n16849__ & new_new_n16864__;
  assign new_new_n16866__ = new_new_n2243__ & new_new_n16863__;
  assign new_new_n16867__ = new_new_n16865__ & new_new_n16866__;
  assign new_new_n16868__ = new_new_n2286__ & new_new_n16867__;
  assign new_new_n16869__ = new_new_n7743__ & new_new_n16868__;
  assign new_new_n16870__ = new_new_n16844__ & ~new_new_n16869__;
  assign new_new_n16871__ = ~new_new_n16844__ & new_new_n16869__;
  assign new_new_n16872__ = ~new_new_n247__ & ~new_new_n298__;
  assign new_new_n16873__ = ~new_new_n939__ & new_new_n16872__;
  assign new_new_n16874__ = new_new_n6323__ & new_new_n16873__;
  assign new_new_n16875__ = new_new_n6319__ & new_new_n16874__;
  assign new_new_n16876__ = ~new_new_n283__ & ~new_new_n671__;
  assign new_new_n16877__ = ~new_new_n249__ & ~new_new_n253__;
  assign new_new_n16878__ = ~new_new_n701__ & ~new_new_n896__;
  assign new_new_n16879__ = ~new_new_n1212__ & new_new_n16878__;
  assign new_new_n16880__ = new_new_n3625__ & new_new_n16877__;
  assign new_new_n16881__ = new_new_n16876__ & new_new_n16880__;
  assign new_new_n16882__ = ~new_new_n607__ & new_new_n16879__;
  assign new_new_n16883__ = new_new_n743__ & new_new_n2991__;
  assign new_new_n16884__ = new_new_n3931__ & new_new_n16883__;
  assign new_new_n16885__ = new_new_n16881__ & new_new_n16882__;
  assign new_new_n16886__ = new_new_n16884__ & new_new_n16885__;
  assign new_new_n16887__ = new_new_n1857__ & new_new_n16886__;
  assign new_new_n16888__ = new_new_n3036__ & new_new_n16887__;
  assign new_new_n16889__ = new_new_n1192__ & new_new_n16888__;
  assign new_new_n16890__ = new_new_n16875__ & new_new_n16889__;
  assign new_new_n16891__ = ~new_new_n16871__ & ~new_new_n16890__;
  assign new_new_n16892__ = ~new_new_n16870__ & ~new_new_n16891__;
  assign new_new_n16893__ = ~new_new_n16842__ & new_new_n16892__;
  assign new_new_n16894__ = ~new_new_n306__ & new_new_n2158__;
  assign new_new_n16895__ = ~new_new_n150__ & ~new_new_n715__;
  assign new_new_n16896__ = new_new_n2644__ & new_new_n16895__;
  assign new_new_n16897__ = ~new_new_n322__ & new_new_n474__;
  assign new_new_n16898__ = new_new_n672__ & ~new_new_n959__;
  assign new_new_n16899__ = ~new_new_n1003__ & new_new_n16898__;
  assign new_new_n16900__ = ~new_new_n115__ & new_new_n16897__;
  assign new_new_n16901__ = new_new_n542__ & new_new_n743__;
  assign new_new_n16902__ = new_new_n1905__ & new_new_n2909__;
  assign new_new_n16903__ = new_new_n4981__ & new_new_n7724__;
  assign new_new_n16904__ = new_new_n16894__ & new_new_n16903__;
  assign new_new_n16905__ = new_new_n16901__ & new_new_n16902__;
  assign new_new_n16906__ = new_new_n16899__ & new_new_n16900__;
  assign new_new_n16907__ = new_new_n16896__ & new_new_n16906__;
  assign new_new_n16908__ = new_new_n16904__ & new_new_n16905__;
  assign new_new_n16909__ = new_new_n16907__ & new_new_n16908__;
  assign new_new_n16910__ = new_new_n3221__ & new_new_n16139__;
  assign new_new_n16911__ = new_new_n16909__ & new_new_n16910__;
  assign new_new_n16912__ = new_new_n3787__ & new_new_n16911__;
  assign new_new_n16913__ = new_new_n5607__ & new_new_n16912__;
  assign new_new_n16914__ = ~new_new_n10337__ & ~new_new_n16913__;
  assign new_new_n16915__ = ~new_new_n10340__ & new_new_n16913__;
  assign new_new_n16916__ = ~new_new_n6958__ & ~new_new_n16914__;
  assign new_new_n16917__ = ~new_new_n16915__ & new_new_n16916__;
  assign new_new_n16918__ = ~pi17 & ~new_new_n16913__;
  assign new_new_n16919__ = pi17 & new_new_n16913__;
  assign new_new_n16920__ = pi17 & ~new_new_n10340__;
  assign new_new_n16921__ = ~new_new_n10337__ & new_new_n16913__;
  assign new_new_n16922__ = ~new_new_n6958__ & ~new_new_n16920__;
  assign new_new_n16923__ = ~new_new_n16921__ & new_new_n16922__;
  assign new_new_n16924__ = ~new_new_n16918__ & ~new_new_n16919__;
  assign new_new_n16925__ = ~new_new_n16923__ & new_new_n16924__;
  assign new_new_n16926__ = ~new_new_n16917__ & ~new_new_n16925__;
  assign new_new_n16927__ = ~new_new_n16839__ & ~new_new_n16926__;
  assign new_new_n16928__ = ~new_new_n16893__ & new_new_n16927__;
  assign new_new_n16929__ = new_new_n16837__ & new_new_n16926__;
  assign new_new_n16930__ = ~new_new_n16765__ & new_new_n16811__;
  assign new_new_n16931__ = ~new_new_n16929__ & ~new_new_n16930__;
  assign new_new_n16932__ = ~new_new_n16781__ & new_new_n16810__;
  assign new_new_n16933__ = new_new_n16765__ & new_new_n16932__;
  assign new_new_n16934__ = new_new_n16929__ & ~new_new_n16933__;
  assign new_new_n16935__ = new_new_n16892__ & ~new_new_n16934__;
  assign new_new_n16936__ = ~new_new_n16931__ & ~new_new_n16935__;
  assign new_new_n16937__ = ~new_new_n16928__ & ~new_new_n16936__;
  assign new_new_n16938__ = new_new_n4212__ & ~new_new_n15273__;
  assign new_new_n16939__ = ~new_new_n4818__ & ~new_new_n15321__;
  assign new_new_n16940__ = new_new_n4815__ & new_new_n15285__;
  assign new_new_n16941__ = ~new_new_n16938__ & ~new_new_n16939__;
  assign new_new_n16942__ = ~new_new_n16940__ & new_new_n16941__;
  assign new_new_n16943__ = new_new_n4214__ & new_new_n16078__;
  assign new_new_n16944__ = pi29 & ~new_new_n16943__;
  assign new_new_n16945__ = new_new_n4825__ & new_new_n16078__;
  assign new_new_n16946__ = ~new_new_n16944__ & ~new_new_n16945__;
  assign new_new_n16947__ = new_new_n16942__ & ~new_new_n16946__;
  assign new_new_n16948__ = ~pi29 & ~new_new_n16942__;
  assign new_new_n16949__ = ~new_new_n16947__ & ~new_new_n16948__;
  assign new_new_n16950__ = new_new_n16937__ & new_new_n16949__;
  assign new_new_n16951__ = new_new_n16913__ & ~new_new_n16926__;
  assign new_new_n16952__ = ~new_new_n16929__ & ~new_new_n16951__;
  assign new_new_n16953__ = new_new_n5021__ & ~new_new_n15349__;
  assign new_new_n16954__ = new_new_n15390__ & ~new_new_n15826__;
  assign new_new_n16955__ = ~new_new_n15390__ & ~new_new_n15828__;
  assign new_new_n16956__ = ~new_new_n16954__ & ~new_new_n16955__;
  assign new_new_n16957__ = new_new_n15349__ & new_new_n16956__;
  assign new_new_n16958__ = new_new_n16451__ & new_new_n16954__;
  assign new_new_n16959__ = ~new_new_n16957__ & ~new_new_n16958__;
  assign new_new_n16960__ = ~new_new_n15853__ & ~new_new_n16959__;
  assign new_new_n16961__ = ~new_new_n16451__ & ~new_new_n16956__;
  assign new_new_n16962__ = ~new_new_n161__ & ~new_new_n16961__;
  assign new_new_n16963__ = ~new_new_n71__ & ~new_new_n15390__;
  assign new_new_n16964__ = ~new_new_n16962__ & new_new_n16963__;
  assign new_new_n16965__ = ~new_new_n16960__ & ~new_new_n16964__;
  assign new_new_n16966__ = new_new_n4147__ & new_new_n16965__;
  assign new_new_n16967__ = pi31 & ~new_new_n16965__;
  assign new_new_n16968__ = ~new_new_n5052__ & ~new_new_n15398__;
  assign new_new_n16969__ = ~new_new_n16967__ & new_new_n16968__;
  assign new_new_n16970__ = ~new_new_n16953__ & ~new_new_n16966__;
  assign new_new_n16971__ = ~new_new_n16969__ & new_new_n16970__;
  assign new_new_n16972__ = new_new_n16952__ & ~new_new_n16971__;
  assign new_new_n16973__ = ~new_new_n16952__ & new_new_n16971__;
  assign new_new_n16974__ = new_new_n16181__ & ~new_new_n16973__;
  assign new_new_n16975__ = ~new_new_n16972__ & ~new_new_n16974__;
  assign new_new_n16976__ = ~new_new_n16950__ & ~new_new_n16975__;
  assign new_new_n16977__ = new_new_n16506__ & ~new_new_n16512__;
  assign new_new_n16978__ = ~new_new_n16506__ & new_new_n16514__;
  assign new_new_n16979__ = ~new_new_n16977__ & ~new_new_n16978__;
  assign new_new_n16980__ = ~new_new_n16976__ & new_new_n16979__;
  assign new_new_n16981__ = ~new_new_n16972__ & new_new_n16979__;
  assign new_new_n16982__ = new_new_n16181__ & ~new_new_n16981__;
  assign new_new_n16983__ = ~new_new_n16937__ & ~new_new_n16949__;
  assign new_new_n16984__ = ~new_new_n16973__ & ~new_new_n16979__;
  assign new_new_n16985__ = ~new_new_n16982__ & ~new_new_n16984__;
  assign new_new_n16986__ = ~new_new_n16983__ & new_new_n16985__;
  assign new_new_n16987__ = new_new_n16950__ & new_new_n16975__;
  assign new_new_n16988__ = ~new_new_n16980__ & ~new_new_n16987__;
  assign new_new_n16989__ = ~new_new_n16986__ & new_new_n16988__;
  assign new_new_n16990__ = ~new_new_n16732__ & new_new_n16989__;
  assign new_new_n16991__ = new_new_n16732__ & ~new_new_n16989__;
  assign new_new_n16992__ = ~new_new_n16537__ & ~new_new_n16991__;
  assign new_new_n16993__ = ~new_new_n16990__ & ~new_new_n16992__;
  assign new_new_n16994__ = ~new_new_n16696__ & ~new_new_n16993__;
  assign new_new_n16995__ = ~new_new_n16695__ & ~new_new_n16994__;
  assign new_new_n16996__ = ~new_new_n16671__ & new_new_n16995__;
  assign new_new_n16997__ = new_new_n16671__ & ~new_new_n16995__;
  assign new_new_n16998__ = ~pi23 & ~new_new_n5186__;
  assign new_new_n16999__ = ~new_new_n5189__ & ~new_new_n16998__;
  assign new_new_n17000__ = ~new_new_n16997__ & new_new_n16999__;
  assign new_new_n17001__ = ~new_new_n16996__ & ~new_new_n17000__;
  assign new_new_n17002__ = new_new_n16667__ & ~new_new_n17001__;
  assign new_new_n17003__ = ~new_new_n16667__ & new_new_n17001__;
  assign new_new_n17004__ = new_new_n5215__ & new_new_n16025__;
  assign new_new_n17005__ = new_new_n5191__ & new_new_n15237__;
  assign new_new_n17006__ = new_new_n5183__ & new_new_n15905__;
  assign new_new_n17007__ = ~new_new_n17005__ & ~new_new_n17006__;
  assign new_new_n17008__ = ~new_new_n17004__ & new_new_n17007__;
  assign new_new_n17009__ = new_new_n5195__ & ~new_new_n15998__;
  assign new_new_n17010__ = pi23 & ~new_new_n17009__;
  assign new_new_n17011__ = new_new_n5974__ & ~new_new_n15998__;
  assign new_new_n17012__ = ~new_new_n17010__ & ~new_new_n17011__;
  assign new_new_n17013__ = new_new_n17008__ & ~new_new_n17012__;
  assign new_new_n17014__ = ~pi23 & ~new_new_n17008__;
  assign new_new_n17015__ = ~new_new_n17013__ & ~new_new_n17014__;
  assign new_new_n17016__ = new_new_n3311__ & new_new_n15244__;
  assign new_new_n17017__ = new_new_n873__ & ~new_new_n15248__;
  assign new_new_n17018__ = ~new_new_n333__ & ~new_new_n15314__;
  assign new_new_n17019__ = ~new_new_n4900__ & new_new_n16378__;
  assign new_new_n17020__ = ~new_new_n17017__ & ~new_new_n17018__;
  assign new_new_n17021__ = ~new_new_n17016__ & new_new_n17020__;
  assign new_new_n17022__ = ~new_new_n17019__ & new_new_n17021__;
  assign new_new_n17023__ = pi26 & ~new_new_n17022__;
  assign new_new_n17024__ = ~pi26 & new_new_n17022__;
  assign new_new_n17025__ = ~new_new_n17023__ & ~new_new_n17024__;
  assign new_new_n17026__ = ~new_new_n16972__ & ~new_new_n16973__;
  assign new_new_n17027__ = ~new_new_n16950__ & ~new_new_n16983__;
  assign new_new_n17028__ = ~new_new_n16181__ & new_new_n17027__;
  assign new_new_n17029__ = new_new_n16181__ & ~new_new_n17027__;
  assign new_new_n17030__ = ~new_new_n17028__ & ~new_new_n17029__;
  assign new_new_n17031__ = new_new_n17026__ & ~new_new_n17030__;
  assign new_new_n17032__ = ~new_new_n17026__ & new_new_n17030__;
  assign new_new_n17033__ = ~new_new_n17031__ & ~new_new_n17032__;
  assign new_new_n17034__ = new_new_n17025__ & new_new_n17033__;
  assign new_new_n17035__ = ~new_new_n17025__ & ~new_new_n17033__;
  assign new_new_n17036__ = ~new_new_n17034__ & ~new_new_n17035__;
  assign new_new_n17037__ = new_new_n16765__ & ~new_new_n16926__;
  assign new_new_n17038__ = ~new_new_n16765__ & new_new_n16926__;
  assign new_new_n17039__ = ~new_new_n17037__ & ~new_new_n17038__;
  assign new_new_n17040__ = new_new_n16837__ & new_new_n17039__;
  assign new_new_n17041__ = ~new_new_n16837__ & ~new_new_n17039__;
  assign new_new_n17042__ = ~new_new_n17040__ & ~new_new_n17041__;
  assign new_new_n17043__ = new_new_n4212__ & ~new_new_n15349__;
  assign new_new_n17044__ = ~new_new_n4818__ & ~new_new_n15398__;
  assign new_new_n17045__ = new_new_n4815__ & ~new_new_n15321__;
  assign new_new_n17046__ = ~new_new_n17043__ & ~new_new_n17044__;
  assign new_new_n17047__ = ~new_new_n17045__ & new_new_n17046__;
  assign new_new_n17048__ = new_new_n4214__ & new_new_n16458__;
  assign new_new_n17049__ = ~pi29 & ~new_new_n17048__;
  assign new_new_n17050__ = new_new_n5732__ & new_new_n16458__;
  assign new_new_n17051__ = ~new_new_n17049__ & ~new_new_n17050__;
  assign new_new_n17052__ = new_new_n17047__ & ~new_new_n17051__;
  assign new_new_n17053__ = pi29 & ~new_new_n17047__;
  assign new_new_n17054__ = ~new_new_n17052__ & ~new_new_n17053__;
  assign new_new_n17055__ = new_new_n5059__ & ~new_new_n15432__;
  assign new_new_n17056__ = new_new_n5053__ & ~new_new_n15362__;
  assign new_new_n17057__ = pi31 & new_new_n15829__;
  assign new_new_n17058__ = ~new_new_n15390__ & ~new_new_n17057__;
  assign new_new_n17059__ = new_new_n15390__ & new_new_n17057__;
  assign new_new_n17060__ = new_new_n765__ & ~new_new_n17058__;
  assign new_new_n17061__ = ~new_new_n17059__ & new_new_n17060__;
  assign new_new_n17062__ = ~new_new_n17055__ & ~new_new_n17056__;
  assign new_new_n17063__ = ~new_new_n17061__ & new_new_n17062__;
  assign new_new_n17064__ = ~new_new_n17054__ & new_new_n17063__;
  assign new_new_n17065__ = new_new_n16811__ & ~new_new_n16892__;
  assign new_new_n17066__ = ~new_new_n16837__ & ~new_new_n17065__;
  assign new_new_n17067__ = new_new_n16810__ & ~new_new_n16892__;
  assign new_new_n17068__ = new_new_n16932__ & ~new_new_n17067__;
  assign new_new_n17069__ = ~new_new_n17066__ & ~new_new_n17068__;
  assign new_new_n17070__ = new_new_n17064__ & new_new_n17069__;
  assign new_new_n17071__ = ~new_new_n17065__ & ~new_new_n17068__;
  assign new_new_n17072__ = ~new_new_n16810__ & ~new_new_n16837__;
  assign new_new_n17073__ = ~new_new_n16840__ & ~new_new_n17072__;
  assign new_new_n17074__ = ~new_new_n17071__ & new_new_n17073__;
  assign new_new_n17075__ = new_new_n17054__ & ~new_new_n17063__;
  assign new_new_n17076__ = ~new_new_n17064__ & ~new_new_n17075__;
  assign new_new_n17077__ = ~new_new_n17074__ & new_new_n17076__;
  assign new_new_n17078__ = ~new_new_n17069__ & new_new_n17075__;
  assign new_new_n17079__ = ~new_new_n17070__ & ~new_new_n17078__;
  assign new_new_n17080__ = ~new_new_n17077__ & new_new_n17079__;
  assign new_new_n17081__ = ~new_new_n17042__ & ~new_new_n17080__;
  assign new_new_n17082__ = new_new_n17065__ & new_new_n17075__;
  assign new_new_n17083__ = ~new_new_n16810__ & new_new_n16892__;
  assign new_new_n17084__ = new_new_n16781__ & ~new_new_n17083__;
  assign new_new_n17085__ = ~new_new_n17067__ & ~new_new_n17084__;
  assign new_new_n17086__ = ~new_new_n17064__ & ~new_new_n17085__;
  assign new_new_n17087__ = ~new_new_n17075__ & ~new_new_n17086__;
  assign new_new_n17088__ = new_new_n16810__ & new_new_n17087__;
  assign new_new_n17089__ = new_new_n17064__ & new_new_n17085__;
  assign new_new_n17090__ = ~new_new_n17088__ & ~new_new_n17089__;
  assign new_new_n17091__ = ~new_new_n16837__ & ~new_new_n17090__;
  assign new_new_n17092__ = ~new_new_n16810__ & ~new_new_n17087__;
  assign new_new_n17093__ = new_new_n17075__ & ~new_new_n17085__;
  assign new_new_n17094__ = ~new_new_n17092__ & ~new_new_n17093__;
  assign new_new_n17095__ = new_new_n16837__ & ~new_new_n17094__;
  assign new_new_n17096__ = new_new_n17064__ & new_new_n17068__;
  assign new_new_n17097__ = ~new_new_n17082__ & ~new_new_n17096__;
  assign new_new_n17098__ = ~new_new_n17091__ & new_new_n17097__;
  assign new_new_n17099__ = ~new_new_n17095__ & new_new_n17098__;
  assign new_new_n17100__ = new_new_n17042__ & ~new_new_n17099__;
  assign new_new_n17101__ = ~new_new_n17081__ & ~new_new_n17100__;
  assign new_new_n17102__ = ~new_new_n15321__ & ~new_new_n16516__;
  assign new_new_n17103__ = ~new_new_n16517__ & ~new_new_n17102__;
  assign new_new_n17104__ = new_new_n4813__ & ~new_new_n17103__;
  assign new_new_n17105__ = ~new_new_n4818__ & ~new_new_n15349__;
  assign new_new_n17106__ = new_new_n4212__ & ~new_new_n15321__;
  assign new_new_n17107__ = ~new_new_n17105__ & ~new_new_n17106__;
  assign new_new_n17108__ = ~new_new_n17104__ & new_new_n17107__;
  assign new_new_n17109__ = new_new_n4214__ & ~new_new_n15273__;
  assign new_new_n17110__ = pi29 & ~new_new_n17109__;
  assign new_new_n17111__ = new_new_n5732__ & ~new_new_n15273__;
  assign new_new_n17112__ = ~new_new_n17110__ & ~new_new_n17111__;
  assign new_new_n17113__ = new_new_n17108__ & ~new_new_n17112__;
  assign new_new_n17114__ = ~pi29 & ~new_new_n17108__;
  assign new_new_n17115__ = ~new_new_n17113__ & ~new_new_n17114__;
  assign new_new_n17116__ = new_new_n17101__ & new_new_n17115__;
  assign new_new_n17117__ = ~new_new_n17069__ & new_new_n17100__;
  assign new_new_n17118__ = new_new_n17069__ & new_new_n17081__;
  assign new_new_n17119__ = ~new_new_n17117__ & ~new_new_n17118__;
  assign new_new_n17120__ = ~new_new_n17116__ & new_new_n17119__;
  assign new_new_n17121__ = new_new_n17036__ & ~new_new_n17120__;
  assign new_new_n17122__ = ~new_new_n17036__ & new_new_n17120__;
  assign new_new_n17123__ = ~new_new_n17121__ & ~new_new_n17122__;
  assign new_new_n17124__ = new_new_n17015__ & new_new_n17123__;
  assign new_new_n17125__ = ~new_new_n17015__ & ~new_new_n17123__;
  assign new_new_n17126__ = ~new_new_n17124__ & ~new_new_n17125__;
  assign new_new_n17127__ = new_new_n873__ & ~new_new_n15314__;
  assign new_new_n17128__ = ~new_new_n333__ & new_new_n15285__;
  assign new_new_n17129__ = new_new_n3311__ & ~new_new_n15248__;
  assign new_new_n17130__ = ~new_new_n17127__ & ~new_new_n17128__;
  assign new_new_n17131__ = ~new_new_n17129__ & new_new_n17130__;
  assign new_new_n17132__ = ~pi26 & ~new_new_n17131__;
  assign new_new_n17133__ = new_new_n512__ & new_new_n16725__;
  assign new_new_n17134__ = new_new_n801__ & new_new_n16725__;
  assign new_new_n17135__ = pi26 & ~new_new_n17134__;
  assign new_new_n17136__ = ~new_new_n17133__ & ~new_new_n17135__;
  assign new_new_n17137__ = new_new_n17131__ & ~new_new_n17136__;
  assign new_new_n17138__ = ~new_new_n17132__ & ~new_new_n17137__;
  assign new_new_n17139__ = ~new_new_n15314__ & new_new_n16082__;
  assign new_new_n17140__ = ~new_new_n16091__ & ~new_new_n17139__;
  assign new_new_n17141__ = ~new_new_n4900__ & new_new_n17140__;
  assign new_new_n17142__ = ~new_new_n333__ & ~new_new_n15273__;
  assign new_new_n17143__ = new_new_n873__ & new_new_n15285__;
  assign new_new_n17144__ = ~new_new_n17142__ & ~new_new_n17143__;
  assign new_new_n17145__ = ~new_new_n17141__ & new_new_n17144__;
  assign new_new_n17146__ = ~pi26 & ~new_new_n17145__;
  assign new_new_n17147__ = new_new_n4898__ & ~new_new_n15314__;
  assign new_new_n17148__ = new_new_n801__ & ~new_new_n15314__;
  assign new_new_n17149__ = pi26 & ~new_new_n17148__;
  assign new_new_n17150__ = ~new_new_n17147__ & ~new_new_n17149__;
  assign new_new_n17151__ = new_new_n17145__ & ~new_new_n17150__;
  assign new_new_n17152__ = ~new_new_n17146__ & ~new_new_n17151__;
  assign new_new_n17153__ = new_new_n68__ & new_new_n15390__;
  assign new_new_n17154__ = pi29 & ~new_new_n17153__;
  assign new_new_n17155__ = pi28 & new_new_n15390__;
  assign new_new_n17156__ = new_new_n3889__ & new_new_n17155__;
  assign new_new_n17157__ = ~new_new_n17154__ & ~new_new_n17156__;
  assign new_new_n17158__ = new_new_n4815__ & ~new_new_n15349__;
  assign new_new_n17159__ = new_new_n4212__ & ~new_new_n15398__;
  assign new_new_n17160__ = ~new_new_n15349__ & new_new_n16448__;
  assign new_new_n17161__ = new_new_n15362__ & new_new_n16443__;
  assign new_new_n17162__ = new_new_n15349__ & new_new_n16441__;
  assign new_new_n17163__ = ~new_new_n15824__ & new_new_n17162__;
  assign new_new_n17164__ = ~new_new_n17161__ & ~new_new_n17163__;
  assign new_new_n17165__ = new_new_n15432__ & ~new_new_n17164__;
  assign new_new_n17166__ = ~new_new_n15824__ & new_new_n16443__;
  assign new_new_n17167__ = ~new_new_n17162__ & ~new_new_n17166__;
  assign new_new_n17168__ = new_new_n15362__ & ~new_new_n17167__;
  assign new_new_n17169__ = new_new_n15349__ & new_new_n16447__;
  assign new_new_n17170__ = new_new_n15824__ & new_new_n17169__;
  assign new_new_n17171__ = ~new_new_n15362__ & new_new_n16450__;
  assign new_new_n17172__ = ~new_new_n17170__ & ~new_new_n17171__;
  assign new_new_n17173__ = ~new_new_n15432__ & ~new_new_n17172__;
  assign new_new_n17174__ = new_new_n15824__ & new_new_n16450__;
  assign new_new_n17175__ = ~new_new_n17169__ & ~new_new_n17174__;
  assign new_new_n17176__ = ~new_new_n15362__ & ~new_new_n17175__;
  assign new_new_n17177__ = ~new_new_n17165__ & ~new_new_n17168__;
  assign new_new_n17178__ = ~new_new_n17173__ & ~new_new_n17176__;
  assign new_new_n17179__ = new_new_n17177__ & new_new_n17178__;
  assign new_new_n17180__ = ~new_new_n17160__ & new_new_n17179__;
  assign new_new_n17181__ = new_new_n4813__ & ~new_new_n17180__;
  assign new_new_n17182__ = ~new_new_n17158__ & ~new_new_n17159__;
  assign new_new_n17183__ = ~new_new_n17181__ & new_new_n17182__;
  assign new_new_n17184__ = ~new_new_n17157__ & new_new_n17183__;
  assign new_new_n17185__ = ~pi29 & ~new_new_n17183__;
  assign new_new_n17186__ = ~new_new_n17184__ & ~new_new_n17185__;
  assign new_new_n17187__ = new_new_n5021__ & ~new_new_n15432__;
  assign new_new_n17188__ = ~new_new_n15440__ & ~new_new_n15475__;
  assign new_new_n17189__ = new_new_n15820__ & new_new_n17188__;
  assign new_new_n17190__ = new_new_n15440__ & ~new_new_n15464__;
  assign new_new_n17191__ = new_new_n15471__ & new_new_n15475__;
  assign new_new_n17192__ = ~new_new_n17190__ & ~new_new_n17191__;
  assign new_new_n17193__ = ~new_new_n15811__ & ~new_new_n17192__;
  assign new_new_n17194__ = new_new_n15439__ & ~new_new_n15464__;
  assign new_new_n17195__ = ~new_new_n15439__ & new_new_n15471__;
  assign new_new_n17196__ = ~new_new_n17194__ & ~new_new_n17195__;
  assign new_new_n17197__ = ~new_new_n15819__ & new_new_n17196__;
  assign new_new_n17198__ = new_new_n17188__ & new_new_n17197__;
  assign new_new_n17199__ = ~new_new_n15439__ & ~new_new_n15819__;
  assign new_new_n17200__ = ~new_new_n15464__ & ~new_new_n17188__;
  assign new_new_n17201__ = ~new_new_n17199__ & new_new_n17200__;
  assign new_new_n17202__ = ~new_new_n17189__ & ~new_new_n17198__;
  assign new_new_n17203__ = ~new_new_n17193__ & new_new_n17202__;
  assign new_new_n17204__ = ~new_new_n17201__ & new_new_n17203__;
  assign new_new_n17205__ = ~new_new_n161__ & new_new_n17204__;
  assign new_new_n17206__ = new_new_n161__ & new_new_n15464__;
  assign new_new_n17207__ = ~new_new_n71__ & ~new_new_n17206__;
  assign new_new_n17208__ = ~new_new_n17205__ & new_new_n17207__;
  assign new_new_n17209__ = new_new_n4147__ & ~new_new_n17208__;
  assign new_new_n17210__ = pi31 & new_new_n17208__;
  assign new_new_n17211__ = ~new_new_n5052__ & ~new_new_n15439__;
  assign new_new_n17212__ = ~new_new_n17210__ & new_new_n17211__;
  assign new_new_n17213__ = ~new_new_n17187__ & ~new_new_n17209__;
  assign new_new_n17214__ = ~new_new_n17212__ & new_new_n17213__;
  assign new_new_n17215__ = new_new_n765__ & ~new_new_n15439__;
  assign new_new_n17216__ = ~new_new_n17206__ & ~new_new_n17215__;
  assign new_new_n17217__ = ~pi31 & ~new_new_n17216__;
  assign new_new_n17218__ = new_new_n71__ & new_new_n15464__;
  assign new_new_n17219__ = new_new_n161__ & ~new_new_n15471__;
  assign new_new_n17220__ = ~new_new_n15439__ & new_new_n15816__;
  assign new_new_n17221__ = new_new_n15472__ & new_new_n15809__;
  assign new_new_n17222__ = new_new_n15439__ & new_new_n15814__;
  assign new_new_n17223__ = new_new_n15779__ & new_new_n17222__;
  assign new_new_n17224__ = ~new_new_n17221__ & ~new_new_n17223__;
  assign new_new_n17225__ = new_new_n15487__ & ~new_new_n17224__;
  assign new_new_n17226__ = ~new_new_n15809__ & new_new_n17195__;
  assign new_new_n17227__ = new_new_n15439__ & new_new_n15815__;
  assign new_new_n17228__ = ~new_new_n15779__ & new_new_n17227__;
  assign new_new_n17229__ = ~new_new_n17226__ & ~new_new_n17228__;
  assign new_new_n17230__ = ~new_new_n15487__ & ~new_new_n17229__;
  assign new_new_n17231__ = ~new_new_n15779__ & new_new_n17195__;
  assign new_new_n17232__ = ~new_new_n17227__ & ~new_new_n17231__;
  assign new_new_n17233__ = ~new_new_n15809__ & ~new_new_n17232__;
  assign new_new_n17234__ = new_new_n15472__ & new_new_n15779__;
  assign new_new_n17235__ = ~new_new_n17222__ & ~new_new_n17234__;
  assign new_new_n17236__ = new_new_n15809__ & ~new_new_n17235__;
  assign new_new_n17237__ = ~new_new_n17233__ & ~new_new_n17236__;
  assign new_new_n17238__ = ~new_new_n17225__ & new_new_n17237__;
  assign new_new_n17239__ = ~new_new_n17230__ & new_new_n17238__;
  assign new_new_n17240__ = ~new_new_n17220__ & new_new_n17239__;
  assign new_new_n17241__ = new_new_n765__ & ~new_new_n17240__;
  assign new_new_n17242__ = ~new_new_n17218__ & ~new_new_n17219__;
  assign new_new_n17243__ = ~new_new_n17241__ & new_new_n17242__;
  assign new_new_n17244__ = pi31 & ~new_new_n17243__;
  assign new_new_n17245__ = ~new_new_n17217__ & ~new_new_n17244__;
  assign new_new_n17246__ = new_new_n2290__ & new_new_n4314__;
  assign new_new_n17247__ = ~new_new_n242__ & ~new_new_n425__;
  assign new_new_n17248__ = ~new_new_n632__ & new_new_n17247__;
  assign new_new_n17249__ = ~new_new_n1073__ & new_new_n17248__;
  assign new_new_n17250__ = ~new_new_n508__ & ~new_new_n809__;
  assign new_new_n17251__ = new_new_n1564__ & new_new_n3635__;
  assign new_new_n17252__ = new_new_n17250__ & new_new_n17251__;
  assign new_new_n17253__ = new_new_n2896__ & new_new_n17249__;
  assign new_new_n17254__ = new_new_n17246__ & new_new_n17253__;
  assign new_new_n17255__ = new_new_n17252__ & new_new_n17254__;
  assign new_new_n17256__ = ~new_new_n274__ & ~new_new_n336__;
  assign new_new_n17257__ = ~new_new_n106__ & ~new_new_n138__;
  assign new_new_n17258__ = new_new_n660__ & ~new_new_n829__;
  assign new_new_n17259__ = ~new_new_n427__ & new_new_n7517__;
  assign new_new_n17260__ = new_new_n17258__ & new_new_n17259__;
  assign new_new_n17261__ = ~new_new_n637__ & ~new_new_n942__;
  assign new_new_n17262__ = ~new_new_n166__ & new_new_n17261__;
  assign new_new_n17263__ = ~new_new_n1064__ & new_new_n1368__;
  assign new_new_n17264__ = new_new_n1628__ & ~new_new_n2697__;
  assign new_new_n17265__ = new_new_n3957__ & new_new_n17257__;
  assign new_new_n17266__ = new_new_n17264__ & new_new_n17265__;
  assign new_new_n17267__ = new_new_n17262__ & new_new_n17263__;
  assign new_new_n17268__ = new_new_n1825__ & new_new_n4389__;
  assign new_new_n17269__ = new_new_n17267__ & new_new_n17268__;
  assign new_new_n17270__ = new_new_n378__ & new_new_n17266__;
  assign new_new_n17271__ = new_new_n1704__ & new_new_n17260__;
  assign new_new_n17272__ = new_new_n17270__ & new_new_n17271__;
  assign new_new_n17273__ = new_new_n1144__ & new_new_n17269__;
  assign new_new_n17274__ = new_new_n17272__ & new_new_n17273__;
  assign new_new_n17275__ = new_new_n121__ & ~new_new_n489__;
  assign new_new_n17276__ = ~new_new_n939__ & new_new_n1709__;
  assign new_new_n17277__ = new_new_n2033__ & new_new_n16282__;
  assign new_new_n17278__ = new_new_n17276__ & new_new_n17277__;
  assign new_new_n17279__ = new_new_n1216__ & new_new_n17275__;
  assign new_new_n17280__ = new_new_n1226__ & new_new_n3386__;
  assign new_new_n17281__ = new_new_n3387__ & new_new_n5566__;
  assign new_new_n17282__ = new_new_n17256__ & new_new_n17281__;
  assign new_new_n17283__ = new_new_n17279__ & new_new_n17280__;
  assign new_new_n17284__ = new_new_n2588__ & new_new_n17278__;
  assign new_new_n17285__ = new_new_n17283__ & new_new_n17284__;
  assign new_new_n17286__ = new_new_n17282__ & new_new_n17285__;
  assign new_new_n17287__ = new_new_n4503__ & new_new_n17286__;
  assign new_new_n17288__ = new_new_n17255__ & new_new_n17274__;
  assign new_new_n17289__ = new_new_n17287__ & new_new_n17288__;
  assign new_new_n17290__ = new_new_n2671__ & new_new_n17289__;
  assign new_new_n17291__ = ~new_new_n17245__ & ~new_new_n17290__;
  assign new_new_n17292__ = new_new_n17245__ & new_new_n17290__;
  assign new_new_n17293__ = ~new_new_n16870__ & ~new_new_n16871__;
  assign new_new_n17294__ = new_new_n17292__ & ~new_new_n17293__;
  assign new_new_n17295__ = new_new_n16890__ & ~new_new_n17294__;
  assign new_new_n17296__ = ~new_new_n17291__ & ~new_new_n17295__;
  assign new_new_n17297__ = ~new_new_n17214__ & ~new_new_n17296__;
  assign new_new_n17298__ = ~new_new_n17292__ & new_new_n17293__;
  assign new_new_n17299__ = new_new_n17295__ & new_new_n17298__;
  assign new_new_n17300__ = new_new_n17214__ & ~new_new_n17291__;
  assign new_new_n17301__ = ~new_new_n16890__ & ~new_new_n17293__;
  assign new_new_n17302__ = ~new_new_n17300__ & new_new_n17301__;
  assign new_new_n17303__ = ~new_new_n17299__ & ~new_new_n17302__;
  assign new_new_n17304__ = ~new_new_n17297__ & new_new_n17303__;
  assign new_new_n17305__ = ~new_new_n17186__ & ~new_new_n17304__;
  assign new_new_n17306__ = new_new_n17186__ & new_new_n17304__;
  assign new_new_n17307__ = ~new_new_n17067__ & ~new_new_n17083__;
  assign new_new_n17308__ = new_new_n16781__ & new_new_n17307__;
  assign new_new_n17309__ = ~new_new_n16781__ & ~new_new_n17307__;
  assign new_new_n17310__ = ~new_new_n17308__ & ~new_new_n17309__;
  assign new_new_n17311__ = ~new_new_n17306__ & new_new_n17310__;
  assign new_new_n17312__ = ~new_new_n17305__ & ~new_new_n17311__;
  assign new_new_n17313__ = new_new_n17152__ & new_new_n17312__;
  assign new_new_n17314__ = ~new_new_n17152__ & ~new_new_n17312__;
  assign new_new_n17315__ = new_new_n17073__ & ~new_new_n17085__;
  assign new_new_n17316__ = ~new_new_n17073__ & new_new_n17085__;
  assign new_new_n17317__ = ~new_new_n17315__ & ~new_new_n17316__;
  assign new_new_n17318__ = ~new_new_n17076__ & new_new_n17317__;
  assign new_new_n17319__ = new_new_n17076__ & ~new_new_n17317__;
  assign new_new_n17320__ = ~new_new_n17318__ & ~new_new_n17319__;
  assign new_new_n17321__ = ~new_new_n17314__ & ~new_new_n17320__;
  assign new_new_n17322__ = ~new_new_n17313__ & ~new_new_n17321__;
  assign new_new_n17323__ = new_new_n17138__ & ~new_new_n17322__;
  assign new_new_n17324__ = ~new_new_n17138__ & new_new_n17322__;
  assign new_new_n17325__ = ~new_new_n17101__ & ~new_new_n17115__;
  assign new_new_n17326__ = ~new_new_n17116__ & ~new_new_n17325__;
  assign new_new_n17327__ = ~new_new_n17324__ & new_new_n17326__;
  assign new_new_n17328__ = ~new_new_n17323__ & ~new_new_n17327__;
  assign new_new_n17329__ = new_new_n17126__ & ~new_new_n17328__;
  assign new_new_n17330__ = ~new_new_n17126__ & new_new_n17328__;
  assign new_new_n17331__ = ~new_new_n17329__ & ~new_new_n17330__;
  assign new_new_n17332__ = ~pi20 & new_new_n6631__;
  assign new_new_n17333__ = ~pi19 & ~new_new_n16056__;
  assign new_new_n17334__ = ~pi18 & ~new_new_n6633__;
  assign new_new_n17335__ = ~new_new_n7015__ & new_new_n17334__;
  assign new_new_n17336__ = ~new_new_n17333__ & new_new_n17335__;
  assign new_new_n17337__ = new_new_n6620__ & new_new_n16056__;
  assign new_new_n17338__ = pi18 & ~new_new_n6632__;
  assign new_new_n17339__ = ~new_new_n6640__ & new_new_n17338__;
  assign new_new_n17340__ = ~new_new_n17337__ & new_new_n17339__;
  assign new_new_n17341__ = ~new_new_n17332__ & ~new_new_n17336__;
  assign new_new_n17342__ = ~new_new_n17340__ & new_new_n17341__;
  assign new_new_n17343__ = ~new_new_n17331__ & ~new_new_n17342__;
  assign new_new_n17344__ = new_new_n17331__ & new_new_n17342__;
  assign new_new_n17345__ = new_new_n873__ & ~new_new_n15273__;
  assign new_new_n17346__ = ~new_new_n333__ & ~new_new_n15321__;
  assign new_new_n17347__ = new_new_n3311__ & new_new_n15285__;
  assign new_new_n17348__ = ~new_new_n17345__ & ~new_new_n17346__;
  assign new_new_n17349__ = ~new_new_n17347__ & new_new_n17348__;
  assign new_new_n17350__ = ~pi26 & ~new_new_n17349__;
  assign new_new_n17351__ = new_new_n512__ & new_new_n16078__;
  assign new_new_n17352__ = new_new_n801__ & new_new_n16078__;
  assign new_new_n17353__ = pi26 & ~new_new_n17352__;
  assign new_new_n17354__ = ~new_new_n17351__ & ~new_new_n17353__;
  assign new_new_n17355__ = new_new_n17349__ & ~new_new_n17354__;
  assign new_new_n17356__ = ~new_new_n17350__ & ~new_new_n17355__;
  assign new_new_n17357__ = new_new_n4212__ & new_new_n15390__;
  assign new_new_n17358__ = ~new_new_n4818__ & ~new_new_n15362__;
  assign new_new_n17359__ = ~new_new_n17357__ & ~new_new_n17358__;
  assign new_new_n17360__ = ~new_new_n15398__ & ~new_new_n16956__;
  assign new_new_n17361__ = new_new_n4214__ & new_new_n17360__;
  assign new_new_n17362__ = new_new_n17359__ & ~new_new_n17361__;
  assign new_new_n17363__ = pi29 & ~new_new_n17362__;
  assign new_new_n17364__ = new_new_n15398__ & ~new_new_n16956__;
  assign new_new_n17365__ = new_new_n4214__ & ~new_new_n17364__;
  assign new_new_n17366__ = ~pi29 & ~new_new_n17365__;
  assign new_new_n17367__ = ~pi28 & ~new_new_n15398__;
  assign new_new_n17368__ = pi28 & new_new_n15398__;
  assign new_new_n17369__ = new_new_n4214__ & ~new_new_n17367__;
  assign new_new_n17370__ = ~new_new_n17368__ & new_new_n17369__;
  assign new_new_n17371__ = new_new_n16956__ & new_new_n17370__;
  assign new_new_n17372__ = ~new_new_n17366__ & ~new_new_n17371__;
  assign new_new_n17373__ = new_new_n17359__ & ~new_new_n17372__;
  assign new_new_n17374__ = ~new_new_n17363__ & ~new_new_n17373__;
  assign new_new_n17375__ = new_new_n765__ & new_new_n15464__;
  assign new_new_n17376__ = ~new_new_n17219__ & ~new_new_n17375__;
  assign new_new_n17377__ = ~pi31 & ~new_new_n17376__;
  assign new_new_n17378__ = new_new_n71__ & ~new_new_n15471__;
  assign new_new_n17379__ = new_new_n161__ & ~new_new_n15809__;
  assign new_new_n17380__ = new_new_n765__ & new_new_n15819__;
  assign new_new_n17381__ = ~new_new_n17378__ & ~new_new_n17379__;
  assign new_new_n17382__ = ~new_new_n17380__ & new_new_n17381__;
  assign new_new_n17383__ = pi31 & ~new_new_n17382__;
  assign new_new_n17384__ = ~new_new_n17377__ & ~new_new_n17383__;
  assign new_new_n17385__ = new_new_n167__ & new_new_n936__;
  assign new_new_n17386__ = ~new_new_n476__ & ~new_new_n700__;
  assign new_new_n17387__ = ~new_new_n947__ & ~new_new_n1080__;
  assign new_new_n17388__ = new_new_n17386__ & new_new_n17387__;
  assign new_new_n17389__ = ~new_new_n945__ & new_new_n17388__;
  assign new_new_n17390__ = ~new_new_n254__ & new_new_n17389__;
  assign new_new_n17391__ = new_new_n91__ & ~new_new_n1107__;
  assign new_new_n17392__ = ~new_new_n213__ & ~new_new_n701__;
  assign new_new_n17393__ = ~new_new_n1008__ & new_new_n17392__;
  assign new_new_n17394__ = new_new_n1383__ & ~new_new_n1506__;
  assign new_new_n17395__ = new_new_n2606__ & new_new_n6186__;
  assign new_new_n17396__ = ~new_new_n17391__ & new_new_n17395__;
  assign new_new_n17397__ = new_new_n17393__ & new_new_n17394__;
  assign new_new_n17398__ = new_new_n782__ & new_new_n1114__;
  assign new_new_n17399__ = new_new_n17397__ & new_new_n17398__;
  assign new_new_n17400__ = new_new_n17396__ & new_new_n17399__;
  assign new_new_n17401__ = ~new_new_n179__ & ~new_new_n240__;
  assign new_new_n17402__ = ~new_new_n441__ & ~new_new_n600__;
  assign new_new_n17403__ = ~new_new_n942__ & new_new_n17402__;
  assign new_new_n17404__ = ~new_new_n828__ & new_new_n17401__;
  assign new_new_n17405__ = ~new_new_n1512__ & new_new_n1740__;
  assign new_new_n17406__ = new_new_n2607__ & new_new_n17257__;
  assign new_new_n17407__ = new_new_n17405__ & new_new_n17406__;
  assign new_new_n17408__ = new_new_n17403__ & new_new_n17404__;
  assign new_new_n17409__ = ~new_new_n115__ & new_new_n1846__;
  assign new_new_n17410__ = new_new_n2066__ & new_new_n3363__;
  assign new_new_n17411__ = new_new_n6122__ & new_new_n17410__;
  assign new_new_n17412__ = new_new_n17408__ & new_new_n17409__;
  assign new_new_n17413__ = new_new_n17407__ & new_new_n17412__;
  assign new_new_n17414__ = new_new_n669__ & new_new_n17411__;
  assign new_new_n17415__ = new_new_n17385__ & new_new_n17390__;
  assign new_new_n17416__ = new_new_n17414__ & new_new_n17415__;
  assign new_new_n17417__ = new_new_n17400__ & new_new_n17413__;
  assign new_new_n17418__ = new_new_n17416__ & new_new_n17417__;
  assign new_new_n17419__ = new_new_n3310__ & new_new_n17418__;
  assign new_new_n17420__ = new_new_n7124__ & new_new_n17419__;
  assign new_new_n17421__ = ~new_new_n282__ & ~new_new_n715__;
  assign new_new_n17422__ = ~new_new_n211__ & ~new_new_n224__;
  assign new_new_n17423__ = new_new_n241__ & ~new_new_n17422__;
  assign new_new_n17424__ = ~new_new_n200__ & ~new_new_n591__;
  assign new_new_n17425__ = ~new_new_n496__ & ~new_new_n724__;
  assign new_new_n17426__ = new_new_n1740__ & new_new_n17425__;
  assign new_new_n17427__ = ~new_new_n17423__ & new_new_n17426__;
  assign new_new_n17428__ = new_new_n17424__ & new_new_n17427__;
  assign new_new_n17429__ = ~new_new_n154__ & ~new_new_n208__;
  assign new_new_n17430__ = ~new_new_n383__ & new_new_n17429__;
  assign new_new_n17431__ = new_new_n16876__ & new_new_n17421__;
  assign new_new_n17432__ = new_new_n17430__ & new_new_n17431__;
  assign new_new_n17433__ = new_new_n964__ & new_new_n1705__;
  assign new_new_n17434__ = new_new_n3513__ & new_new_n4989__;
  assign new_new_n17435__ = new_new_n17433__ & new_new_n17434__;
  assign new_new_n17436__ = new_new_n1160__ & new_new_n17432__;
  assign new_new_n17437__ = new_new_n5412__ & new_new_n17436__;
  assign new_new_n17438__ = new_new_n17428__ & new_new_n17435__;
  assign new_new_n17439__ = new_new_n17437__ & new_new_n17438__;
  assign new_new_n17440__ = new_new_n1839__ & new_new_n17439__;
  assign new_new_n17441__ = new_new_n3580__ & new_new_n6772__;
  assign new_new_n17442__ = new_new_n17440__ & new_new_n17441__;
  assign new_new_n17443__ = new_new_n3662__ & new_new_n17442__;
  assign new_new_n17444__ = new_new_n17420__ & new_new_n17443__;
  assign new_new_n17445__ = ~new_new_n17420__ & ~new_new_n17443__;
  assign new_new_n17446__ = ~pi11 & ~new_new_n8477__;
  assign new_new_n17447__ = ~new_new_n8855__ & ~new_new_n17446__;
  assign new_new_n17448__ = ~new_new_n17445__ & ~new_new_n17447__;
  assign new_new_n17449__ = ~new_new_n17444__ & ~new_new_n17448__;
  assign new_new_n17450__ = ~new_new_n17384__ & new_new_n17449__;
  assign new_new_n17451__ = new_new_n4212__ & ~new_new_n15432__;
  assign new_new_n17452__ = ~new_new_n4215__ & ~new_new_n16771__;
  assign new_new_n17453__ = new_new_n4215__ & new_new_n15362__;
  assign new_new_n17454__ = new_new_n4214__ & ~new_new_n17453__;
  assign new_new_n17455__ = ~new_new_n17452__ & new_new_n17454__;
  assign new_new_n17456__ = ~new_new_n17451__ & ~new_new_n17455__;
  assign new_new_n17457__ = ~pi29 & ~new_new_n17456__;
  assign new_new_n17458__ = new_new_n4221__ & ~new_new_n15439__;
  assign new_new_n17459__ = pi29 & ~new_new_n17458__;
  assign new_new_n17460__ = new_new_n66__ & ~new_new_n15439__;
  assign new_new_n17461__ = ~new_new_n17459__ & ~new_new_n17460__;
  assign new_new_n17462__ = new_new_n17456__ & ~new_new_n17461__;
  assign new_new_n17463__ = ~new_new_n17457__ & ~new_new_n17462__;
  assign new_new_n17464__ = ~new_new_n15487__ & ~new_new_n15809__;
  assign new_new_n17465__ = new_new_n15779__ & ~new_new_n15809__;
  assign new_new_n17466__ = ~new_new_n15780__ & ~new_new_n15853__;
  assign new_new_n17467__ = ~new_new_n17465__ & new_new_n17466__;
  assign new_new_n17468__ = ~new_new_n17464__ & ~new_new_n17467__;
  assign new_new_n17469__ = ~new_new_n15471__ & ~new_new_n17468__;
  assign new_new_n17470__ = new_new_n15471__ & new_new_n15809__;
  assign new_new_n17471__ = ~new_new_n15779__ & new_new_n17470__;
  assign new_new_n17472__ = ~new_new_n161__ & ~new_new_n17471__;
  assign new_new_n17473__ = ~new_new_n71__ & ~new_new_n15487__;
  assign new_new_n17474__ = ~new_new_n17472__ & new_new_n17473__;
  assign new_new_n17475__ = ~new_new_n71__ & ~new_new_n15776__;
  assign new_new_n17476__ = ~new_new_n161__ & ~new_new_n15809__;
  assign new_new_n17477__ = ~new_new_n17475__ & new_new_n17476__;
  assign new_new_n17478__ = ~new_new_n17474__ & ~new_new_n17477__;
  assign new_new_n17479__ = ~new_new_n17469__ & new_new_n17478__;
  assign new_new_n17480__ = pi31 & ~new_new_n17479__;
  assign new_new_n17481__ = new_new_n765__ & ~new_new_n15471__;
  assign new_new_n17482__ = ~new_new_n17379__ & ~new_new_n17481__;
  assign new_new_n17483__ = ~pi31 & ~new_new_n17482__;
  assign new_new_n17484__ = ~new_new_n17480__ & ~new_new_n17483__;
  assign new_new_n17485__ = ~new_new_n17444__ & ~new_new_n17445__;
  assign new_new_n17486__ = new_new_n17447__ & ~new_new_n17485__;
  assign new_new_n17487__ = ~new_new_n17444__ & new_new_n17448__;
  assign new_new_n17488__ = ~new_new_n17486__ & ~new_new_n17487__;
  assign new_new_n17489__ = new_new_n17484__ & new_new_n17488__;
  assign new_new_n17490__ = ~new_new_n17484__ & ~new_new_n17488__;
  assign new_new_n17491__ = ~new_new_n282__ & ~new_new_n510__;
  assign new_new_n17492__ = ~new_new_n632__ & new_new_n17491__;
  assign new_new_n17493__ = ~new_new_n226__ & ~new_new_n483__;
  assign new_new_n17494__ = ~new_new_n939__ & new_new_n17493__;
  assign new_new_n17495__ = new_new_n1341__ & new_new_n17492__;
  assign new_new_n17496__ = new_new_n2161__ & new_new_n7725__;
  assign new_new_n17497__ = new_new_n17495__ & new_new_n17496__;
  assign new_new_n17498__ = new_new_n2580__ & new_new_n17494__;
  assign new_new_n17499__ = new_new_n17497__ & new_new_n17498__;
  assign new_new_n17500__ = ~new_new_n1033__ & ~new_new_n2170__;
  assign new_new_n17501__ = ~new_new_n189__ & ~new_new_n945__;
  assign new_new_n17502__ = ~new_new_n270__ & ~new_new_n445__;
  assign new_new_n17503__ = ~new_new_n382__ & new_new_n17500__;
  assign new_new_n17504__ = new_new_n17502__ & new_new_n17503__;
  assign new_new_n17505__ = new_new_n17501__ & new_new_n17504__;
  assign new_new_n17506__ = ~new_new_n240__ & ~new_new_n472__;
  assign new_new_n17507__ = ~new_new_n584__ & ~new_new_n603__;
  assign new_new_n17508__ = ~new_new_n933__ & ~new_new_n1113__;
  assign new_new_n17509__ = ~new_new_n1291__ & new_new_n17508__;
  assign new_new_n17510__ = new_new_n17506__ & new_new_n17507__;
  assign new_new_n17511__ = ~new_new_n255__ & new_new_n16794__;
  assign new_new_n17512__ = new_new_n17510__ & new_new_n17511__;
  assign new_new_n17513__ = ~new_new_n519__ & new_new_n17509__;
  assign new_new_n17514__ = new_new_n1225__ & new_new_n1252__;
  assign new_new_n17515__ = new_new_n2706__ & new_new_n2763__;
  assign new_new_n17516__ = new_new_n2994__ & new_new_n7401__;
  assign new_new_n17517__ = new_new_n17515__ & new_new_n17516__;
  assign new_new_n17518__ = new_new_n17513__ & new_new_n17514__;
  assign new_new_n17519__ = new_new_n17512__ & new_new_n17518__;
  assign new_new_n17520__ = new_new_n17505__ & new_new_n17517__;
  assign new_new_n17521__ = new_new_n17519__ & new_new_n17520__;
  assign new_new_n17522__ = new_new_n17499__ & new_new_n17521__;
  assign new_new_n17523__ = new_new_n1874__ & new_new_n17522__;
  assign new_new_n17524__ = new_new_n3927__ & new_new_n17523__;
  assign new_new_n17525__ = ~new_new_n235__ & ~new_new_n1007__;
  assign new_new_n17526__ = ~new_new_n198__ & ~new_new_n282__;
  assign new_new_n17527__ = ~new_new_n258__ & ~new_new_n816__;
  assign new_new_n17528__ = ~new_new_n1217__ & new_new_n1423__;
  assign new_new_n17529__ = new_new_n2506__ & new_new_n17525__;
  assign new_new_n17530__ = new_new_n17528__ & new_new_n17529__;
  assign new_new_n17531__ = new_new_n17526__ & new_new_n17527__;
  assign new_new_n17532__ = ~new_new_n935__ & new_new_n1216__;
  assign new_new_n17533__ = new_new_n5698__ & new_new_n17532__;
  assign new_new_n17534__ = new_new_n17530__ & new_new_n17531__;
  assign new_new_n17535__ = new_new_n5791__ & new_new_n17534__;
  assign new_new_n17536__ = new_new_n17533__ & new_new_n17535__;
  assign new_new_n17537__ = ~new_new_n212__ & ~new_new_n425__;
  assign new_new_n17538__ = ~new_new_n1109__ & new_new_n17537__;
  assign new_new_n17539__ = ~new_new_n346__ & ~new_new_n732__;
  assign new_new_n17540__ = new_new_n3056__ & new_new_n17539__;
  assign new_new_n17541__ = new_new_n1153__ & new_new_n17538__;
  assign new_new_n17542__ = new_new_n3203__ & new_new_n17541__;
  assign new_new_n17543__ = new_new_n985__ & new_new_n17540__;
  assign new_new_n17544__ = new_new_n17542__ & new_new_n17543__;
  assign new_new_n17545__ = ~new_new_n890__ & ~new_new_n995__;
  assign new_new_n17546__ = ~new_new_n143__ & ~new_new_n317__;
  assign new_new_n17547__ = ~new_new_n353__ & ~new_new_n489__;
  assign new_new_n17548__ = ~new_new_n1073__ & new_new_n17545__;
  assign new_new_n17549__ = ~new_new_n2697__ & new_new_n3485__;
  assign new_new_n17550__ = new_new_n17548__ & new_new_n17549__;
  assign new_new_n17551__ = new_new_n17546__ & new_new_n17547__;
  assign new_new_n17552__ = ~new_new_n115__ & new_new_n1268__;
  assign new_new_n17553__ = new_new_n1448__ & new_new_n2911__;
  assign new_new_n17554__ = new_new_n4729__ & new_new_n17553__;
  assign new_new_n17555__ = new_new_n17551__ & new_new_n17552__;
  assign new_new_n17556__ = new_new_n256__ & new_new_n17550__;
  assign new_new_n17557__ = new_new_n4398__ & new_new_n17556__;
  assign new_new_n17558__ = new_new_n17554__ & new_new_n17555__;
  assign new_new_n17559__ = new_new_n17557__ & new_new_n17558__;
  assign new_new_n17560__ = new_new_n17544__ & new_new_n17559__;
  assign new_new_n17561__ = new_new_n16294__ & new_new_n17536__;
  assign new_new_n17562__ = new_new_n17560__ & new_new_n17561__;
  assign new_new_n17563__ = new_new_n3413__ & new_new_n17562__;
  assign new_new_n17564__ = ~new_new_n17524__ & ~new_new_n17563__;
  assign new_new_n17565__ = new_new_n17524__ & new_new_n17563__;
  assign new_new_n17566__ = pi05 & new_new_n10712__;
  assign new_new_n17567__ = ~pi05 & new_new_n10709__;
  assign new_new_n17568__ = ~pi08 & ~new_new_n17567__;
  assign new_new_n17569__ = ~new_new_n17566__ & ~new_new_n17568__;
  assign new_new_n17570__ = ~new_new_n17565__ & new_new_n17569__;
  assign new_new_n17571__ = ~new_new_n17564__ & ~new_new_n17570__;
  assign new_new_n17572__ = new_new_n161__ & new_new_n15524__;
  assign new_new_n17573__ = new_new_n765__ & ~new_new_n15487__;
  assign new_new_n17574__ = ~new_new_n17572__ & ~new_new_n17573__;
  assign new_new_n17575__ = ~pi31 & ~new_new_n17574__;
  assign new_new_n17576__ = new_new_n15487__ & ~new_new_n15524__;
  assign new_new_n17577__ = new_new_n15533__ & ~new_new_n15779__;
  assign new_new_n17578__ = ~new_new_n17576__ & ~new_new_n17577__;
  assign new_new_n17579__ = ~new_new_n15520__ & ~new_new_n17578__;
  assign new_new_n17580__ = new_new_n15533__ & new_new_n17576__;
  assign new_new_n17581__ = ~new_new_n15520__ & ~new_new_n15774__;
  assign new_new_n17582__ = ~new_new_n17580__ & ~new_new_n17581__;
  assign new_new_n17583__ = new_new_n15771__ & ~new_new_n17582__;
  assign new_new_n17584__ = ~new_new_n15487__ & new_new_n15524__;
  assign new_new_n17585__ = ~new_new_n15779__ & ~new_new_n17584__;
  assign new_new_n17586__ = ~new_new_n17583__ & ~new_new_n17585__;
  assign new_new_n17587__ = ~new_new_n17579__ & new_new_n17586__;
  assign new_new_n17588__ = new_new_n765__ & ~new_new_n17587__;
  assign new_new_n17589__ = new_new_n161__ & ~new_new_n15520__;
  assign new_new_n17590__ = new_new_n71__ & ~new_new_n15524__;
  assign new_new_n17591__ = pi31 & ~new_new_n17590__;
  assign new_new_n17592__ = ~new_new_n17589__ & new_new_n17591__;
  assign new_new_n17593__ = ~new_new_n17588__ & new_new_n17592__;
  assign new_new_n17594__ = ~new_new_n17575__ & ~new_new_n17593__;
  assign new_new_n17595__ = new_new_n17571__ & new_new_n17594__;
  assign new_new_n17596__ = new_new_n17420__ & ~new_new_n17595__;
  assign new_new_n17597__ = ~new_new_n76__ & ~new_new_n346__;
  assign new_new_n17598__ = new_new_n6124__ & new_new_n17597__;
  assign new_new_n17599__ = ~new_new_n826__ & ~new_new_n869__;
  assign new_new_n17600__ = ~new_new_n952__ & new_new_n17599__;
  assign new_new_n17601__ = new_new_n1569__ & new_new_n17600__;
  assign new_new_n17602__ = ~new_new_n657__ & ~new_new_n2170__;
  assign new_new_n17603__ = new_new_n779__ & new_new_n17602__;
  assign new_new_n17604__ = ~new_new_n1167__ & new_new_n5817__;
  assign new_new_n17605__ = new_new_n17603__ & new_new_n17604__;
  assign new_new_n17606__ = ~new_new_n630__ & new_new_n1114__;
  assign new_new_n17607__ = new_new_n1905__ & new_new_n4979__;
  assign new_new_n17608__ = new_new_n17424__ & new_new_n17607__;
  assign new_new_n17609__ = new_new_n17605__ & new_new_n17606__;
  assign new_new_n17610__ = new_new_n709__ & new_new_n3180__;
  assign new_new_n17611__ = new_new_n3321__ & new_new_n17598__;
  assign new_new_n17612__ = new_new_n17610__ & new_new_n17611__;
  assign new_new_n17613__ = new_new_n17608__ & new_new_n17609__;
  assign new_new_n17614__ = new_new_n728__ & new_new_n17613__;
  assign new_new_n17615__ = new_new_n17601__ & new_new_n17612__;
  assign new_new_n17616__ = new_new_n17614__ & new_new_n17615__;
  assign new_new_n17617__ = new_new_n2437__ & new_new_n17616__;
  assign new_new_n17618__ = ~new_new_n312__ & ~new_new_n320__;
  assign new_new_n17619__ = ~new_new_n875__ & ~new_new_n1398__;
  assign new_new_n17620__ = new_new_n17618__ & new_new_n17619__;
  assign new_new_n17621__ = ~new_new_n329__ & ~new_new_n635__;
  assign new_new_n17622__ = ~new_new_n1009__ & new_new_n1570__;
  assign new_new_n17623__ = new_new_n3439__ & new_new_n17622__;
  assign new_new_n17624__ = new_new_n17620__ & new_new_n17621__;
  assign new_new_n17625__ = ~new_new_n316__ & new_new_n17624__;
  assign new_new_n17626__ = new_new_n17623__ & new_new_n17625__;
  assign new_new_n17627__ = ~new_new_n438__ & ~new_new_n445__;
  assign new_new_n17628__ = ~new_new_n600__ & ~new_new_n658__;
  assign new_new_n17629__ = ~new_new_n776__ & ~new_new_n1080__;
  assign new_new_n17630__ = ~new_new_n1343__ & new_new_n17629__;
  assign new_new_n17631__ = new_new_n17627__ & new_new_n17628__;
  assign new_new_n17632__ = ~new_new_n816__ & new_new_n1370__;
  assign new_new_n17633__ = new_new_n1629__ & new_new_n3283__;
  assign new_new_n17634__ = new_new_n4948__ & new_new_n17633__;
  assign new_new_n17635__ = new_new_n17631__ & new_new_n17632__;
  assign new_new_n17636__ = new_new_n751__ & new_new_n17630__;
  assign new_new_n17637__ = new_new_n1078__ & new_new_n2889__;
  assign new_new_n17638__ = new_new_n17636__ & new_new_n17637__;
  assign new_new_n17639__ = new_new_n17634__ & new_new_n17635__;
  assign new_new_n17640__ = ~new_new_n1539__ & new_new_n17639__;
  assign new_new_n17641__ = new_new_n17638__ & new_new_n17640__;
  assign new_new_n17642__ = new_new_n17626__ & new_new_n17641__;
  assign new_new_n17643__ = new_new_n5472__ & new_new_n17642__;
  assign new_new_n17644__ = new_new_n17617__ & new_new_n17643__;
  assign new_new_n17645__ = ~new_new_n17596__ & new_new_n17644__;
  assign new_new_n17646__ = ~new_new_n17571__ & ~new_new_n17594__;
  assign new_new_n17647__ = ~new_new_n17420__ & ~new_new_n17646__;
  assign new_new_n17648__ = ~new_new_n17645__ & ~new_new_n17647__;
  assign new_new_n17649__ = ~new_new_n17490__ & ~new_new_n17648__;
  assign new_new_n17650__ = ~new_new_n17489__ & ~new_new_n17649__;
  assign new_new_n17651__ = new_new_n17463__ & ~new_new_n17650__;
  assign new_new_n17652__ = ~new_new_n17463__ & new_new_n17650__;
  assign new_new_n17653__ = new_new_n17384__ & ~new_new_n17449__;
  assign new_new_n17654__ = ~new_new_n17450__ & ~new_new_n17653__;
  assign new_new_n17655__ = new_new_n16890__ & new_new_n17654__;
  assign new_new_n17656__ = ~new_new_n16890__ & ~new_new_n17654__;
  assign new_new_n17657__ = ~new_new_n17655__ & ~new_new_n17656__;
  assign new_new_n17658__ = ~new_new_n17652__ & ~new_new_n17657__;
  assign new_new_n17659__ = ~new_new_n17651__ & ~new_new_n17658__;
  assign new_new_n17660__ = new_new_n17450__ & new_new_n17659__;
  assign new_new_n17661__ = ~new_new_n17291__ & ~new_new_n17292__;
  assign new_new_n17662__ = ~new_new_n16890__ & new_new_n17450__;
  assign new_new_n17663__ = ~new_new_n17659__ & ~new_new_n17662__;
  assign new_new_n17664__ = new_new_n16890__ & new_new_n17653__;
  assign new_new_n17665__ = new_new_n17661__ & ~new_new_n17664__;
  assign new_new_n17666__ = ~new_new_n17663__ & new_new_n17665__;
  assign new_new_n17667__ = new_new_n17653__ & ~new_new_n17659__;
  assign new_new_n17668__ = new_new_n16890__ & ~new_new_n17661__;
  assign new_new_n17669__ = ~new_new_n17667__ & new_new_n17668__;
  assign new_new_n17670__ = ~new_new_n17660__ & ~new_new_n17666__;
  assign new_new_n17671__ = ~new_new_n17669__ & new_new_n17670__;
  assign new_new_n17672__ = new_new_n17374__ & ~new_new_n17671__;
  assign new_new_n17673__ = ~new_new_n17374__ & new_new_n17671__;
  assign new_new_n17674__ = new_new_n16890__ & ~new_new_n17292__;
  assign new_new_n17675__ = ~new_new_n16890__ & ~new_new_n17291__;
  assign new_new_n17676__ = ~new_new_n17674__ & ~new_new_n17675__;
  assign new_new_n17677__ = ~new_new_n17214__ & new_new_n17293__;
  assign new_new_n17678__ = new_new_n17214__ & ~new_new_n17293__;
  assign new_new_n17679__ = ~new_new_n17677__ & ~new_new_n17678__;
  assign new_new_n17680__ = new_new_n17676__ & new_new_n17679__;
  assign new_new_n17681__ = ~new_new_n17676__ & ~new_new_n17679__;
  assign new_new_n17682__ = ~new_new_n17680__ & ~new_new_n17681__;
  assign new_new_n17683__ = ~new_new_n17673__ & ~new_new_n17682__;
  assign new_new_n17684__ = ~new_new_n17672__ & ~new_new_n17683__;
  assign new_new_n17685__ = new_new_n17356__ & new_new_n17684__;
  assign new_new_n17686__ = ~new_new_n17356__ & ~new_new_n17684__;
  assign new_new_n17687__ = ~new_new_n17305__ & ~new_new_n17306__;
  assign new_new_n17688__ = new_new_n17310__ & new_new_n17687__;
  assign new_new_n17689__ = ~new_new_n17310__ & ~new_new_n17687__;
  assign new_new_n17690__ = ~new_new_n17688__ & ~new_new_n17689__;
  assign new_new_n17691__ = ~new_new_n17686__ & ~new_new_n17690__;
  assign new_new_n17692__ = ~new_new_n17685__ & ~new_new_n17691__;
  assign new_new_n17693__ = ~new_new_n17313__ & ~new_new_n17314__;
  assign new_new_n17694__ = ~new_new_n17320__ & new_new_n17693__;
  assign new_new_n17695__ = new_new_n17320__ & ~new_new_n17693__;
  assign new_new_n17696__ = ~new_new_n17694__ & ~new_new_n17695__;
  assign new_new_n17697__ = new_new_n17692__ & ~new_new_n17696__;
  assign new_new_n17698__ = ~new_new_n17692__ & new_new_n17696__;
  assign new_new_n17699__ = new_new_n5213__ & new_new_n15237__;
  assign new_new_n17700__ = new_new_n5183__ & new_new_n15244__;
  assign new_new_n17701__ = new_new_n5191__ & ~new_new_n15248__;
  assign new_new_n17702__ = new_new_n5215__ & ~new_new_n16603__;
  assign new_new_n17703__ = ~new_new_n17700__ & ~new_new_n17701__;
  assign new_new_n17704__ = ~new_new_n17699__ & new_new_n17703__;
  assign new_new_n17705__ = ~new_new_n17702__ & new_new_n17704__;
  assign new_new_n17706__ = ~new_new_n17697__ & ~new_new_n17698__;
  assign new_new_n17707__ = pi23 & ~new_new_n17706__;
  assign new_new_n17708__ = ~pi23 & new_new_n17706__;
  assign new_new_n17709__ = ~new_new_n17707__ & ~new_new_n17708__;
  assign new_new_n17710__ = new_new_n17705__ & new_new_n17709__;
  assign new_new_n17711__ = ~new_new_n17705__ & ~new_new_n17709__;
  assign new_new_n17712__ = ~new_new_n17710__ & ~new_new_n17711__;
  assign new_new_n17713__ = ~new_new_n17698__ & ~new_new_n17712__;
  assign new_new_n17714__ = ~new_new_n17697__ & ~new_new_n17713__;
  assign new_new_n17715__ = ~new_new_n17323__ & ~new_new_n17324__;
  assign new_new_n17716__ = ~new_new_n17326__ & ~new_new_n17715__;
  assign new_new_n17717__ = new_new_n17326__ & new_new_n17715__;
  assign new_new_n17718__ = ~new_new_n17716__ & ~new_new_n17717__;
  assign new_new_n17719__ = new_new_n17714__ & new_new_n17718__;
  assign new_new_n17720__ = ~new_new_n17714__ & ~new_new_n17718__;
  assign new_new_n17721__ = new_new_n5191__ & new_new_n15244__;
  assign new_new_n17722__ = new_new_n5183__ & new_new_n15237__;
  assign new_new_n17723__ = ~new_new_n5212__ & ~new_new_n15905__;
  assign new_new_n17724__ = new_new_n5212__ & new_new_n15917__;
  assign new_new_n17725__ = new_new_n5195__ & ~new_new_n17723__;
  assign new_new_n17726__ = ~new_new_n17724__ & new_new_n17725__;
  assign new_new_n17727__ = ~new_new_n17722__ & ~new_new_n17726__;
  assign new_new_n17728__ = ~new_new_n17721__ & new_new_n17727__;
  assign new_new_n17729__ = pi23 & ~new_new_n17728__;
  assign new_new_n17730__ = new_new_n9374__ & ~new_new_n15244__;
  assign new_new_n17731__ = ~new_new_n5190__ & ~new_new_n17730__;
  assign new_new_n17732__ = ~pi23 & ~new_new_n17731__;
  assign new_new_n17733__ = new_new_n17727__ & new_new_n17732__;
  assign new_new_n17734__ = ~new_new_n17729__ & ~new_new_n17733__;
  assign new_new_n17735__ = ~new_new_n17720__ & ~new_new_n17734__;
  assign new_new_n17736__ = ~new_new_n17719__ & ~new_new_n17735__;
  assign new_new_n17737__ = ~new_new_n17344__ & new_new_n17736__;
  assign new_new_n17738__ = ~new_new_n17343__ & ~new_new_n17737__;
  assign new_new_n17739__ = new_new_n5183__ & ~new_new_n15998__;
  assign new_new_n17740__ = new_new_n5212__ & new_new_n16051__;
  assign new_new_n17741__ = new_new_n5195__ & ~new_new_n16056__;
  assign new_new_n17742__ = ~new_new_n17740__ & new_new_n17741__;
  assign new_new_n17743__ = ~new_new_n17739__ & ~new_new_n17742__;
  assign new_new_n17744__ = new_new_n5185__ & new_new_n15905__;
  assign new_new_n17745__ = pi23 & ~new_new_n17744__;
  assign new_new_n17746__ = new_new_n5188__ & new_new_n15905__;
  assign new_new_n17747__ = ~pi23 & ~new_new_n17746__;
  assign new_new_n17748__ = pi20 & ~new_new_n17747__;
  assign new_new_n17749__ = ~new_new_n17745__ & ~new_new_n17748__;
  assign new_new_n17750__ = new_new_n17743__ & ~new_new_n17749__;
  assign new_new_n17751__ = ~pi23 & ~new_new_n17743__;
  assign new_new_n17752__ = ~new_new_n17750__ & ~new_new_n17751__;
  assign new_new_n17753__ = ~new_new_n17034__ & ~new_new_n17120__;
  assign new_new_n17754__ = ~new_new_n17035__ & ~new_new_n17753__;
  assign new_new_n17755__ = ~new_new_n17752__ & new_new_n17754__;
  assign new_new_n17756__ = new_new_n17752__ & ~new_new_n17754__;
  assign new_new_n17757__ = ~new_new_n17755__ & ~new_new_n17756__;
  assign new_new_n17758__ = new_new_n4212__ & new_new_n15285__;
  assign new_new_n17759__ = ~new_new_n4818__ & ~new_new_n15273__;
  assign new_new_n17760__ = ~new_new_n17758__ & ~new_new_n17759__;
  assign new_new_n17761__ = new_new_n4214__ & ~new_new_n16091__;
  assign new_new_n17762__ = ~new_new_n15314__ & ~new_new_n16082__;
  assign new_new_n17763__ = new_new_n17761__ & new_new_n17762__;
  assign new_new_n17764__ = new_new_n17760__ & ~new_new_n17763__;
  assign new_new_n17765__ = ~pi29 & ~new_new_n17764__;
  assign new_new_n17766__ = ~pi29 & ~new_new_n17761__;
  assign new_new_n17767__ = pi28 & new_new_n15314__;
  assign new_new_n17768__ = ~pi28 & ~new_new_n17140__;
  assign new_new_n17769__ = new_new_n17761__ & ~new_new_n17767__;
  assign new_new_n17770__ = ~new_new_n17768__ & new_new_n17769__;
  assign new_new_n17771__ = new_new_n17760__ & ~new_new_n17766__;
  assign new_new_n17772__ = ~new_new_n17770__ & new_new_n17771__;
  assign new_new_n17773__ = ~new_new_n17765__ & ~new_new_n17772__;
  assign new_new_n17774__ = ~new_new_n4900__ & ~new_new_n16603__;
  assign new_new_n17775__ = ~new_new_n333__ & ~new_new_n15248__;
  assign new_new_n17776__ = new_new_n873__ & new_new_n15244__;
  assign new_new_n17777__ = ~new_new_n17775__ & ~new_new_n17776__;
  assign new_new_n17778__ = ~new_new_n17774__ & new_new_n17777__;
  assign new_new_n17779__ = pi26 & ~new_new_n17778__;
  assign new_new_n17780__ = new_new_n512__ & new_new_n15237__;
  assign new_new_n17781__ = new_new_n801__ & new_new_n15237__;
  assign new_new_n17782__ = ~pi26 & ~new_new_n17781__;
  assign new_new_n17783__ = ~new_new_n17780__ & ~new_new_n17782__;
  assign new_new_n17784__ = new_new_n17778__ & ~new_new_n17783__;
  assign new_new_n17785__ = ~new_new_n17779__ & ~new_new_n17784__;
  assign new_new_n17786__ = new_new_n16975__ & ~new_new_n16983__;
  assign new_new_n17787__ = ~new_new_n16976__ & ~new_new_n17786__;
  assign new_new_n17788__ = new_new_n16181__ & new_new_n16972__;
  assign new_new_n17789__ = ~new_new_n16181__ & new_new_n16973__;
  assign new_new_n17790__ = ~new_new_n17788__ & ~new_new_n17789__;
  assign new_new_n17791__ = new_new_n17027__ & new_new_n17790__;
  assign new_new_n17792__ = ~new_new_n17787__ & ~new_new_n17791__;
  assign new_new_n17793__ = ~new_new_n16979__ & ~new_new_n17792__;
  assign new_new_n17794__ = new_new_n16950__ & new_new_n16973__;
  assign new_new_n17795__ = new_new_n16950__ & new_new_n16971__;
  assign new_new_n17796__ = ~new_new_n16950__ & ~new_new_n16971__;
  assign new_new_n17797__ = ~new_new_n16952__ & ~new_new_n16983__;
  assign new_new_n17798__ = ~new_new_n17796__ & new_new_n17797__;
  assign new_new_n17799__ = ~new_new_n17795__ & ~new_new_n17798__;
  assign new_new_n17800__ = ~new_new_n16181__ & ~new_new_n17799__;
  assign new_new_n17801__ = ~new_new_n16973__ & new_new_n16983__;
  assign new_new_n17802__ = new_new_n16952__ & new_new_n17796__;
  assign new_new_n17803__ = ~new_new_n17801__ & ~new_new_n17802__;
  assign new_new_n17804__ = new_new_n16181__ & ~new_new_n17803__;
  assign new_new_n17805__ = new_new_n16972__ & new_new_n16983__;
  assign new_new_n17806__ = ~new_new_n17794__ & ~new_new_n17805__;
  assign new_new_n17807__ = ~new_new_n17800__ & new_new_n17806__;
  assign new_new_n17808__ = ~new_new_n17804__ & new_new_n17807__;
  assign new_new_n17809__ = new_new_n16979__ & ~new_new_n17808__;
  assign new_new_n17810__ = ~new_new_n17793__ & ~new_new_n17809__;
  assign new_new_n17811__ = ~new_new_n17785__ & new_new_n17810__;
  assign new_new_n17812__ = new_new_n17785__ & ~new_new_n17810__;
  assign new_new_n17813__ = ~new_new_n17811__ & ~new_new_n17812__;
  assign new_new_n17814__ = new_new_n17773__ & new_new_n17813__;
  assign new_new_n17815__ = ~new_new_n17773__ & ~new_new_n17813__;
  assign new_new_n17816__ = ~new_new_n17814__ & ~new_new_n17815__;
  assign new_new_n17817__ = new_new_n17757__ & new_new_n17816__;
  assign new_new_n17818__ = ~new_new_n17757__ & ~new_new_n17816__;
  assign new_new_n17819__ = ~new_new_n17817__ & ~new_new_n17818__;
  assign new_new_n17820__ = ~new_new_n17738__ & new_new_n17819__;
  assign new_new_n17821__ = ~new_new_n17756__ & ~new_new_n17814__;
  assign new_new_n17822__ = ~new_new_n17815__ & new_new_n17821__;
  assign new_new_n17823__ = ~new_new_n17755__ & ~new_new_n17822__;
  assign new_new_n17824__ = ~new_new_n4900__ & ~new_new_n15917__;
  assign new_new_n17825__ = ~new_new_n333__ & new_new_n15244__;
  assign new_new_n17826__ = new_new_n873__ & new_new_n15237__;
  assign new_new_n17827__ = ~new_new_n17825__ & ~new_new_n17826__;
  assign new_new_n17828__ = ~new_new_n17824__ & new_new_n17827__;
  assign new_new_n17829__ = pi26 & ~new_new_n17828__;
  assign new_new_n17830__ = new_new_n512__ & new_new_n15905__;
  assign new_new_n17831__ = new_new_n801__ & new_new_n15905__;
  assign new_new_n17832__ = ~pi26 & ~new_new_n17831__;
  assign new_new_n17833__ = ~new_new_n17830__ & ~new_new_n17832__;
  assign new_new_n17834__ = new_new_n17828__ & ~new_new_n17833__;
  assign new_new_n17835__ = ~new_new_n17829__ & ~new_new_n17834__;
  assign new_new_n17836__ = new_new_n17773__ & ~new_new_n17785__;
  assign new_new_n17837__ = ~new_new_n17773__ & new_new_n17785__;
  assign new_new_n17838__ = ~new_new_n17810__ & ~new_new_n17837__;
  assign new_new_n17839__ = ~new_new_n17836__ & ~new_new_n17838__;
  assign new_new_n17840__ = new_new_n17835__ & new_new_n17839__;
  assign new_new_n17841__ = ~new_new_n17835__ & ~new_new_n17839__;
  assign new_new_n17842__ = ~new_new_n17840__ & ~new_new_n17841__;
  assign new_new_n17843__ = ~new_new_n16990__ & ~new_new_n16991__;
  assign new_new_n17844__ = ~new_new_n16537__ & new_new_n17843__;
  assign new_new_n17845__ = new_new_n16537__ & ~new_new_n17843__;
  assign new_new_n17846__ = ~new_new_n17844__ & ~new_new_n17845__;
  assign new_new_n17847__ = new_new_n17842__ & ~new_new_n17846__;
  assign new_new_n17848__ = ~new_new_n17842__ & new_new_n17846__;
  assign new_new_n17849__ = ~new_new_n17847__ & ~new_new_n17848__;
  assign new_new_n17850__ = new_new_n17823__ & new_new_n17849__;
  assign new_new_n17851__ = ~new_new_n17823__ & ~new_new_n17849__;
  assign new_new_n17852__ = ~new_new_n17850__ & ~new_new_n17851__;
  assign new_new_n17853__ = new_new_n5191__ & ~new_new_n15998__;
  assign new_new_n17854__ = new_new_n5212__ & ~new_new_n16630__;
  assign new_new_n17855__ = new_new_n5195__ & ~new_new_n17854__;
  assign new_new_n17856__ = new_new_n5183__ & ~new_new_n16056__;
  assign new_new_n17857__ = ~new_new_n17853__ & ~new_new_n17856__;
  assign new_new_n17858__ = ~new_new_n17855__ & new_new_n17857__;
  assign new_new_n17859__ = pi23 & ~new_new_n17858__;
  assign new_new_n17860__ = ~pi23 & new_new_n17858__;
  assign new_new_n17861__ = ~new_new_n17859__ & ~new_new_n17860__;
  assign new_new_n17862__ = new_new_n17852__ & new_new_n17861__;
  assign new_new_n17863__ = ~new_new_n17852__ & ~new_new_n17861__;
  assign new_new_n17864__ = ~new_new_n17862__ & ~new_new_n17863__;
  assign new_new_n17865__ = new_new_n17820__ & new_new_n17864__;
  assign new_new_n17866__ = new_new_n17738__ & ~new_new_n17819__;
  assign new_new_n17867__ = ~new_new_n17124__ & new_new_n17328__;
  assign new_new_n17868__ = ~new_new_n17125__ & ~new_new_n17867__;
  assign new_new_n17869__ = new_new_n5191__ & ~new_new_n15314__;
  assign new_new_n17870__ = new_new_n5183__ & ~new_new_n15248__;
  assign new_new_n17871__ = new_new_n5213__ & new_new_n15244__;
  assign new_new_n17872__ = ~new_new_n17869__ & ~new_new_n17870__;
  assign new_new_n17873__ = ~new_new_n17871__ & new_new_n17872__;
  assign new_new_n17874__ = new_new_n5195__ & new_new_n16378__;
  assign new_new_n17875__ = pi23 & ~new_new_n17874__;
  assign new_new_n17876__ = new_new_n7878__ & new_new_n16378__;
  assign new_new_n17877__ = ~new_new_n17875__ & ~new_new_n17876__;
  assign new_new_n17878__ = new_new_n17873__ & ~new_new_n17877__;
  assign new_new_n17879__ = ~pi23 & ~new_new_n17873__;
  assign new_new_n17880__ = ~new_new_n17878__ & ~new_new_n17879__;
  assign new_new_n17881__ = new_new_n3311__ & ~new_new_n15273__;
  assign new_new_n17882__ = ~new_new_n333__ & ~new_new_n15349__;
  assign new_new_n17883__ = new_new_n873__ & ~new_new_n15321__;
  assign new_new_n17884__ = ~new_new_n17882__ & ~new_new_n17883__;
  assign new_new_n17885__ = ~new_new_n17881__ & new_new_n17884__;
  assign new_new_n17886__ = pi26 & ~new_new_n17885__;
  assign new_new_n17887__ = new_new_n4898__ & ~new_new_n17103__;
  assign new_new_n17888__ = new_new_n801__ & ~new_new_n17103__;
  assign new_new_n17889__ = ~pi26 & ~new_new_n17888__;
  assign new_new_n17890__ = ~new_new_n17887__ & ~new_new_n17889__;
  assign new_new_n17891__ = new_new_n17885__ & ~new_new_n17890__;
  assign new_new_n17892__ = ~new_new_n17886__ & ~new_new_n17891__;
  assign new_new_n17893__ = ~new_new_n17672__ & ~new_new_n17673__;
  assign new_new_n17894__ = new_new_n17682__ & ~new_new_n17893__;
  assign new_new_n17895__ = ~new_new_n17682__ & new_new_n17893__;
  assign new_new_n17896__ = ~new_new_n17894__ & ~new_new_n17895__;
  assign new_new_n17897__ = new_new_n17892__ & new_new_n17896__;
  assign new_new_n17898__ = ~new_new_n17892__ & ~new_new_n17896__;
  assign new_new_n17899__ = new_new_n873__ & ~new_new_n15349__;
  assign new_new_n17900__ = ~new_new_n333__ & ~new_new_n15398__;
  assign new_new_n17901__ = new_new_n3311__ & ~new_new_n15321__;
  assign new_new_n17902__ = ~new_new_n17899__ & ~new_new_n17900__;
  assign new_new_n17903__ = ~new_new_n17901__ & new_new_n17902__;
  assign new_new_n17904__ = pi26 & ~new_new_n17903__;
  assign new_new_n17905__ = new_new_n4898__ & new_new_n16458__;
  assign new_new_n17906__ = new_new_n801__ & new_new_n16458__;
  assign new_new_n17907__ = ~pi26 & ~new_new_n17906__;
  assign new_new_n17908__ = ~new_new_n17905__ & ~new_new_n17907__;
  assign new_new_n17909__ = new_new_n17903__ & ~new_new_n17908__;
  assign new_new_n17910__ = ~new_new_n17904__ & ~new_new_n17909__;
  assign new_new_n17911__ = ~new_new_n4818__ & ~new_new_n15432__;
  assign new_new_n17912__ = new_new_n4212__ & ~new_new_n15362__;
  assign new_new_n17913__ = ~new_new_n17911__ & ~new_new_n17912__;
  assign new_new_n17914__ = new_new_n15390__ & ~new_new_n15829__;
  assign new_new_n17915__ = new_new_n4214__ & new_new_n17914__;
  assign new_new_n17916__ = new_new_n17913__ & ~new_new_n17915__;
  assign new_new_n17917__ = pi29 & ~new_new_n17916__;
  assign new_new_n17918__ = ~new_new_n15390__ & ~new_new_n15829__;
  assign new_new_n17919__ = new_new_n4214__ & ~new_new_n17918__;
  assign new_new_n17920__ = ~pi29 & ~new_new_n17919__;
  assign new_new_n17921__ = ~pi28 & ~new_new_n15390__;
  assign new_new_n17922__ = ~new_new_n17155__ & ~new_new_n17921__;
  assign new_new_n17923__ = new_new_n4214__ & new_new_n15829__;
  assign new_new_n17924__ = ~new_new_n17922__ & new_new_n17923__;
  assign new_new_n17925__ = ~new_new_n17920__ & ~new_new_n17924__;
  assign new_new_n17926__ = new_new_n17913__ & ~new_new_n17925__;
  assign new_new_n17927__ = ~new_new_n17917__ & ~new_new_n17926__;
  assign new_new_n17928__ = new_new_n17910__ & new_new_n17927__;
  assign new_new_n17929__ = ~new_new_n17910__ & ~new_new_n17927__;
  assign new_new_n17930__ = ~new_new_n17928__ & ~new_new_n17929__;
  assign new_new_n17931__ = ~new_new_n17662__ & ~new_new_n17664__;
  assign new_new_n17932__ = new_new_n17245__ & ~new_new_n17931__;
  assign new_new_n17933__ = ~new_new_n17245__ & new_new_n17931__;
  assign new_new_n17934__ = ~new_new_n17932__ & ~new_new_n17933__;
  assign new_new_n17935__ = new_new_n17290__ & ~new_new_n17659__;
  assign new_new_n17936__ = ~new_new_n17290__ & new_new_n17659__;
  assign new_new_n17937__ = ~new_new_n17935__ & ~new_new_n17936__;
  assign new_new_n17938__ = new_new_n17934__ & new_new_n17937__;
  assign new_new_n17939__ = ~new_new_n17934__ & ~new_new_n17937__;
  assign new_new_n17940__ = ~new_new_n17938__ & ~new_new_n17939__;
  assign new_new_n17941__ = new_new_n17930__ & ~new_new_n17940__;
  assign new_new_n17942__ = ~new_new_n17928__ & ~new_new_n17941__;
  assign new_new_n17943__ = ~new_new_n17898__ & ~new_new_n17942__;
  assign new_new_n17944__ = ~new_new_n17897__ & ~new_new_n17943__;
  assign new_new_n17945__ = ~new_new_n17880__ & ~new_new_n17944__;
  assign new_new_n17946__ = new_new_n17880__ & new_new_n17944__;
  assign new_new_n17947__ = ~new_new_n17685__ & ~new_new_n17686__;
  assign new_new_n17948__ = ~new_new_n17690__ & new_new_n17947__;
  assign new_new_n17949__ = new_new_n17690__ & ~new_new_n17947__;
  assign new_new_n17950__ = ~new_new_n17948__ & ~new_new_n17949__;
  assign new_new_n17951__ = ~new_new_n17946__ & ~new_new_n17950__;
  assign new_new_n17952__ = ~new_new_n17945__ & ~new_new_n17951__;
  assign new_new_n17953__ = ~new_new_n17712__ & new_new_n17952__;
  assign new_new_n17954__ = new_new_n17712__ & ~new_new_n17952__;
  assign new_new_n17955__ = new_new_n6631__ & ~new_new_n16056__;
  assign new_new_n17956__ = pi20 & ~new_new_n16051__;
  assign new_new_n17957__ = new_new_n6629__ & ~new_new_n15998__;
  assign new_new_n17958__ = ~new_new_n6625__ & new_new_n15905__;
  assign new_new_n17959__ = ~new_new_n17957__ & ~new_new_n17958__;
  assign new_new_n17960__ = pi19 & new_new_n16051__;
  assign new_new_n17961__ = new_new_n17959__ & new_new_n17960__;
  assign new_new_n17962__ = ~new_new_n17956__ & ~new_new_n17961__;
  assign new_new_n17963__ = new_new_n17955__ & ~new_new_n17962__;
  assign new_new_n17964__ = pi20 & ~new_new_n17959__;
  assign new_new_n17965__ = ~pi20 & ~new_new_n17955__;
  assign new_new_n17966__ = new_new_n17959__ & new_new_n17965__;
  assign new_new_n17967__ = ~new_new_n17964__ & ~new_new_n17966__;
  assign new_new_n17968__ = ~new_new_n17963__ & new_new_n17967__;
  assign new_new_n17969__ = ~new_new_n17954__ & ~new_new_n17968__;
  assign new_new_n17970__ = ~new_new_n17953__ & ~new_new_n17969__;
  assign new_new_n17971__ = new_new_n6629__ & new_new_n15237__;
  assign new_new_n17972__ = ~new_new_n6625__ & new_new_n15244__;
  assign new_new_n17973__ = ~new_new_n17971__ & ~new_new_n17972__;
  assign new_new_n17974__ = new_new_n15905__ & ~new_new_n15917__;
  assign new_new_n17975__ = new_new_n6631__ & new_new_n17974__;
  assign new_new_n17976__ = new_new_n17973__ & ~new_new_n17975__;
  assign new_new_n17977__ = pi20 & ~new_new_n17976__;
  assign new_new_n17978__ = ~new_new_n15905__ & new_new_n15917__;
  assign new_new_n17979__ = new_new_n6631__ & ~new_new_n17978__;
  assign new_new_n17980__ = ~pi20 & ~new_new_n17979__;
  assign new_new_n17981__ = ~new_new_n15905__ & ~new_new_n15917__;
  assign new_new_n17982__ = ~pi19 & ~new_new_n17981__;
  assign new_new_n17983__ = new_new_n15905__ & new_new_n15917__;
  assign new_new_n17984__ = pi19 & ~new_new_n17983__;
  assign new_new_n17985__ = new_new_n6631__ & ~new_new_n17982__;
  assign new_new_n17986__ = ~new_new_n17984__ & new_new_n17985__;
  assign new_new_n17987__ = ~new_new_n17980__ & ~new_new_n17986__;
  assign new_new_n17988__ = new_new_n17973__ & ~new_new_n17987__;
  assign new_new_n17989__ = ~new_new_n17977__ & ~new_new_n17988__;
  assign new_new_n17990__ = new_new_n5183__ & ~new_new_n15314__;
  assign new_new_n17991__ = new_new_n5191__ & new_new_n15285__;
  assign new_new_n17992__ = new_new_n5213__ & ~new_new_n15248__;
  assign new_new_n17993__ = new_new_n5215__ & new_new_n16725__;
  assign new_new_n17994__ = ~new_new_n17990__ & ~new_new_n17991__;
  assign new_new_n17995__ = ~new_new_n17992__ & new_new_n17994__;
  assign new_new_n17996__ = ~new_new_n17993__ & new_new_n17995__;
  assign new_new_n17997__ = pi23 & ~new_new_n17996__;
  assign new_new_n17998__ = ~pi23 & new_new_n17996__;
  assign new_new_n17999__ = ~new_new_n17997__ & ~new_new_n17998__;
  assign new_new_n18000__ = ~new_new_n17897__ & ~new_new_n17898__;
  assign new_new_n18001__ = ~new_new_n17942__ & new_new_n18000__;
  assign new_new_n18002__ = new_new_n17942__ & ~new_new_n18000__;
  assign new_new_n18003__ = ~new_new_n18001__ & ~new_new_n18002__;
  assign new_new_n18004__ = ~new_new_n17651__ & ~new_new_n17652__;
  assign new_new_n18005__ = new_new_n17657__ & ~new_new_n18004__;
  assign new_new_n18006__ = ~new_new_n17657__ & new_new_n18004__;
  assign new_new_n18007__ = ~new_new_n18005__ & ~new_new_n18006__;
  assign new_new_n18008__ = ~new_new_n17489__ & ~new_new_n17490__;
  assign new_new_n18009__ = ~new_new_n17648__ & new_new_n18008__;
  assign new_new_n18010__ = new_new_n17648__ & ~new_new_n18008__;
  assign new_new_n18011__ = ~new_new_n18009__ & ~new_new_n18010__;
  assign new_new_n18012__ = new_new_n161__ & ~new_new_n15487__;
  assign new_new_n18013__ = new_new_n765__ & ~new_new_n15809__;
  assign new_new_n18014__ = ~new_new_n18012__ & ~new_new_n18013__;
  assign new_new_n18015__ = ~pi31 & ~new_new_n18014__;
  assign new_new_n18016__ = new_new_n71__ & ~new_new_n15487__;
  assign new_new_n18017__ = ~new_new_n15775__ & ~new_new_n15780__;
  assign new_new_n18018__ = ~new_new_n15809__ & new_new_n18017__;
  assign new_new_n18019__ = new_new_n15809__ & ~new_new_n18017__;
  assign new_new_n18020__ = ~new_new_n18018__ & ~new_new_n18019__;
  assign new_new_n18021__ = new_new_n765__ & new_new_n18020__;
  assign new_new_n18022__ = ~new_new_n17572__ & ~new_new_n18016__;
  assign new_new_n18023__ = ~new_new_n18021__ & new_new_n18022__;
  assign new_new_n18024__ = pi31 & ~new_new_n18023__;
  assign new_new_n18025__ = ~new_new_n18015__ & ~new_new_n18024__;
  assign new_new_n18026__ = new_new_n4813__ & ~new_new_n17240__;
  assign new_new_n18027__ = ~new_new_n4818__ & ~new_new_n15471__;
  assign new_new_n18028__ = new_new_n4212__ & new_new_n15464__;
  assign new_new_n18029__ = ~new_new_n18027__ & ~new_new_n18028__;
  assign new_new_n18030__ = ~new_new_n18026__ & new_new_n18029__;
  assign new_new_n18031__ = new_new_n4214__ & ~new_new_n15439__;
  assign new_new_n18032__ = ~pi29 & ~new_new_n18031__;
  assign new_new_n18033__ = new_new_n4825__ & ~new_new_n15439__;
  assign new_new_n18034__ = ~new_new_n18032__ & ~new_new_n18033__;
  assign new_new_n18035__ = new_new_n18030__ & ~new_new_n18034__;
  assign new_new_n18036__ = pi29 & ~new_new_n18030__;
  assign new_new_n18037__ = ~new_new_n18035__ & ~new_new_n18036__;
  assign new_new_n18038__ = new_new_n18025__ & ~new_new_n18037__;
  assign new_new_n18039__ = ~new_new_n18025__ & new_new_n18037__;
  assign new_new_n18040__ = ~new_new_n17596__ & ~new_new_n17647__;
  assign new_new_n18041__ = new_new_n17644__ & ~new_new_n18040__;
  assign new_new_n18042__ = ~new_new_n17644__ & new_new_n18040__;
  assign new_new_n18043__ = ~new_new_n18041__ & ~new_new_n18042__;
  assign new_new_n18044__ = ~new_new_n18039__ & ~new_new_n18043__;
  assign new_new_n18045__ = ~new_new_n18038__ & ~new_new_n18044__;
  assign new_new_n18046__ = new_new_n18011__ & ~new_new_n18045__;
  assign new_new_n18047__ = ~new_new_n18011__ & new_new_n18045__;
  assign new_new_n18048__ = new_new_n4815__ & ~new_new_n15432__;
  assign new_new_n18049__ = new_new_n4212__ & ~new_new_n15439__;
  assign new_new_n18050__ = ~new_new_n4818__ & new_new_n15464__;
  assign new_new_n18051__ = new_new_n4813__ & new_new_n17204__;
  assign new_new_n18052__ = ~new_new_n18049__ & ~new_new_n18050__;
  assign new_new_n18053__ = ~new_new_n18048__ & new_new_n18052__;
  assign new_new_n18054__ = ~new_new_n18051__ & new_new_n18053__;
  assign new_new_n18055__ = pi29 & ~new_new_n18054__;
  assign new_new_n18056__ = ~pi29 & new_new_n18054__;
  assign new_new_n18057__ = ~new_new_n18055__ & ~new_new_n18056__;
  assign new_new_n18058__ = ~new_new_n18047__ & ~new_new_n18057__;
  assign new_new_n18059__ = ~new_new_n18046__ & ~new_new_n18058__;
  assign new_new_n18060__ = ~new_new_n18007__ & new_new_n18059__;
  assign new_new_n18061__ = new_new_n18007__ & ~new_new_n18059__;
  assign new_new_n18062__ = new_new_n3311__ & ~new_new_n15349__;
  assign new_new_n18063__ = new_new_n873__ & ~new_new_n15398__;
  assign new_new_n18064__ = ~new_new_n333__ & new_new_n15390__;
  assign new_new_n18065__ = ~new_new_n4900__ & ~new_new_n17180__;
  assign new_new_n18066__ = ~new_new_n18063__ & ~new_new_n18064__;
  assign new_new_n18067__ = ~new_new_n18062__ & new_new_n18066__;
  assign new_new_n18068__ = ~new_new_n18065__ & new_new_n18067__;
  assign new_new_n18069__ = pi26 & ~new_new_n18068__;
  assign new_new_n18070__ = ~pi26 & new_new_n18068__;
  assign new_new_n18071__ = ~new_new_n18069__ & ~new_new_n18070__;
  assign new_new_n18072__ = ~new_new_n18061__ & new_new_n18071__;
  assign new_new_n18073__ = ~new_new_n18060__ & ~new_new_n18072__;
  assign new_new_n18074__ = ~new_new_n17930__ & new_new_n17940__;
  assign new_new_n18075__ = ~new_new_n17941__ & ~new_new_n18074__;
  assign new_new_n18076__ = new_new_n5213__ & ~new_new_n15314__;
  assign new_new_n18077__ = new_new_n5191__ & ~new_new_n15273__;
  assign new_new_n18078__ = new_new_n5183__ & new_new_n15285__;
  assign new_new_n18079__ = ~new_new_n18077__ & ~new_new_n18078__;
  assign new_new_n18080__ = ~new_new_n18076__ & new_new_n18079__;
  assign new_new_n18081__ = new_new_n5195__ & new_new_n17140__;
  assign new_new_n18082__ = pi23 & ~new_new_n18081__;
  assign new_new_n18083__ = new_new_n7878__ & new_new_n17140__;
  assign new_new_n18084__ = ~new_new_n18082__ & ~new_new_n18083__;
  assign new_new_n18085__ = new_new_n18080__ & ~new_new_n18084__;
  assign new_new_n18086__ = ~pi23 & ~new_new_n18080__;
  assign new_new_n18087__ = ~new_new_n18085__ & ~new_new_n18086__;
  assign new_new_n18088__ = new_new_n18075__ & ~new_new_n18087__;
  assign new_new_n18089__ = new_new_n18073__ & ~new_new_n18088__;
  assign new_new_n18090__ = ~new_new_n18075__ & new_new_n18087__;
  assign new_new_n18091__ = ~new_new_n18089__ & ~new_new_n18090__;
  assign new_new_n18092__ = new_new_n18003__ & new_new_n18091__;
  assign new_new_n18093__ = ~new_new_n18003__ & ~new_new_n18091__;
  assign new_new_n18094__ = ~new_new_n18092__ & ~new_new_n18093__;
  assign new_new_n18095__ = new_new_n17999__ & ~new_new_n18094__;
  assign new_new_n18096__ = ~new_new_n17999__ & new_new_n18094__;
  assign new_new_n18097__ = ~new_new_n18095__ & ~new_new_n18096__;
  assign new_new_n18098__ = new_new_n17989__ & ~new_new_n18097__;
  assign new_new_n18099__ = ~new_new_n17989__ & new_new_n18097__;
  assign new_new_n18100__ = ~new_new_n333__ & ~new_new_n15362__;
  assign new_new_n18101__ = new_new_n873__ & new_new_n15390__;
  assign new_new_n18102__ = ~new_new_n18100__ & ~new_new_n18101__;
  assign new_new_n18103__ = new_new_n801__ & new_new_n17360__;
  assign new_new_n18104__ = new_new_n18102__ & ~new_new_n18103__;
  assign new_new_n18105__ = pi26 & ~new_new_n18104__;
  assign new_new_n18106__ = new_new_n801__ & ~new_new_n17364__;
  assign new_new_n18107__ = ~pi26 & ~new_new_n18106__;
  assign new_new_n18108__ = pi25 & new_new_n15398__;
  assign new_new_n18109__ = ~pi25 & ~new_new_n15398__;
  assign new_new_n18110__ = ~new_new_n110__ & ~new_new_n18108__;
  assign new_new_n18111__ = ~new_new_n18109__ & new_new_n18110__;
  assign new_new_n18112__ = new_new_n16956__ & new_new_n18111__;
  assign new_new_n18113__ = ~new_new_n18107__ & ~new_new_n18112__;
  assign new_new_n18114__ = new_new_n18102__ & ~new_new_n18113__;
  assign new_new_n18115__ = ~new_new_n18105__ & ~new_new_n18114__;
  assign new_new_n18116__ = ~new_new_n18038__ & ~new_new_n18039__;
  assign new_new_n18117__ = ~new_new_n18043__ & new_new_n18116__;
  assign new_new_n18118__ = new_new_n18043__ & ~new_new_n18116__;
  assign new_new_n18119__ = ~new_new_n18117__ & ~new_new_n18118__;
  assign new_new_n18120__ = ~new_new_n17564__ & ~new_new_n17565__;
  assign new_new_n18121__ = ~new_new_n17569__ & new_new_n18120__;
  assign new_new_n18122__ = new_new_n17569__ & ~new_new_n18120__;
  assign new_new_n18123__ = ~new_new_n18121__ & ~new_new_n18122__;
  assign new_new_n18124__ = ~new_new_n15520__ & new_new_n15533__;
  assign new_new_n18125__ = ~new_new_n15533__ & new_new_n15771__;
  assign new_new_n18126__ = ~new_new_n15777__ & ~new_new_n18125__;
  assign new_new_n18127__ = new_new_n765__ & ~new_new_n18126__;
  assign new_new_n18128__ = ~new_new_n18124__ & ~new_new_n18127__;
  assign new_new_n18129__ = ~new_new_n15524__ & ~new_new_n18128__;
  assign new_new_n18130__ = ~new_new_n161__ & ~new_new_n15520__;
  assign new_new_n18131__ = ~new_new_n71__ & ~new_new_n15773__;
  assign new_new_n18132__ = new_new_n18130__ & ~new_new_n18131__;
  assign new_new_n18133__ = new_new_n15525__ & new_new_n15771__;
  assign new_new_n18134__ = ~new_new_n161__ & ~new_new_n18133__;
  assign new_new_n18135__ = ~new_new_n71__ & new_new_n15533__;
  assign new_new_n18136__ = ~new_new_n18134__ & new_new_n18135__;
  assign new_new_n18137__ = pi31 & ~new_new_n18132__;
  assign new_new_n18138__ = ~new_new_n18136__ & new_new_n18137__;
  assign new_new_n18139__ = ~new_new_n18129__ & new_new_n18138__;
  assign new_new_n18140__ = ~new_new_n161__ & ~new_new_n15524__;
  assign new_new_n18141__ = new_new_n4876__ & ~new_new_n18140__;
  assign new_new_n18142__ = ~new_new_n17589__ & new_new_n18141__;
  assign new_new_n18143__ = ~new_new_n18139__ & ~new_new_n18142__;
  assign new_new_n18144__ = ~new_new_n18123__ & ~new_new_n18143__;
  assign new_new_n18145__ = new_new_n18123__ & new_new_n18143__;
  assign new_new_n18146__ = ~pi02 & ~new_new_n14393__;
  assign new_new_n18147__ = ~pi05 & ~new_new_n11466__;
  assign new_new_n18148__ = new_new_n18146__ & new_new_n18147__;
  assign new_new_n18149__ = ~new_new_n120__ & new_new_n1263__;
  assign new_new_n18150__ = ~new_new_n383__ & ~new_new_n657__;
  assign new_new_n18151__ = new_new_n596__ & new_new_n18150__;
  assign new_new_n18152__ = new_new_n2119__ & new_new_n18151__;
  assign new_new_n18153__ = new_new_n984__ & new_new_n1230__;
  assign new_new_n18154__ = new_new_n1307__ & new_new_n2168__;
  assign new_new_n18155__ = new_new_n3129__ & new_new_n18154__;
  assign new_new_n18156__ = new_new_n18152__ & new_new_n18153__;
  assign new_new_n18157__ = new_new_n789__ & new_new_n18156__;
  assign new_new_n18158__ = new_new_n18155__ & new_new_n18157__;
  assign new_new_n18159__ = new_new_n1145__ & ~new_new_n1539__;
  assign new_new_n18160__ = ~new_new_n698__ & new_new_n17598__;
  assign new_new_n18161__ = new_new_n18159__ & new_new_n18160__;
  assign new_new_n18162__ = ~new_new_n874__ & ~new_new_n937__;
  assign new_new_n18163__ = ~new_new_n130__ & ~new_new_n250__;
  assign new_new_n18164__ = ~new_new_n284__ & ~new_new_n1162__;
  assign new_new_n18165__ = new_new_n18163__ & new_new_n18164__;
  assign new_new_n18166__ = new_new_n1563__ & new_new_n18165__;
  assign new_new_n18167__ = new_new_n3277__ & new_new_n16852__;
  assign new_new_n18168__ = new_new_n18162__ & new_new_n18167__;
  assign new_new_n18169__ = new_new_n3320__ & new_new_n18166__;
  assign new_new_n18170__ = new_new_n18168__ & new_new_n18169__;
  assign new_new_n18171__ = new_new_n3201__ & new_new_n4719__;
  assign new_new_n18172__ = new_new_n17385__ & new_new_n18171__;
  assign new_new_n18173__ = new_new_n18161__ & new_new_n18170__;
  assign new_new_n18174__ = new_new_n18172__ & new_new_n18173__;
  assign new_new_n18175__ = new_new_n18158__ & new_new_n18174__;
  assign new_new_n18176__ = ~new_new_n379__ & ~new_new_n634__;
  assign new_new_n18177__ = ~new_new_n990__ & ~new_new_n1343__;
  assign new_new_n18178__ = new_new_n18176__ & new_new_n18177__;
  assign new_new_n18179__ = new_new_n4465__ & new_new_n18178__;
  assign new_new_n18180__ = ~new_new_n124__ & new_new_n1428__;
  assign new_new_n18181__ = new_new_n1961__ & new_new_n18149__;
  assign new_new_n18182__ = new_new_n18180__ & new_new_n18181__;
  assign new_new_n18183__ = ~new_new_n652__ & new_new_n18179__;
  assign new_new_n18184__ = new_new_n7522__ & new_new_n18183__;
  assign new_new_n18185__ = new_new_n4572__ & new_new_n18182__;
  assign new_new_n18186__ = new_new_n7130__ & new_new_n18185__;
  assign new_new_n18187__ = new_new_n17400__ & new_new_n18184__;
  assign new_new_n18188__ = new_new_n18186__ & new_new_n18187__;
  assign new_new_n18189__ = new_new_n18175__ & new_new_n18188__;
  assign new_new_n18190__ = pi02 & pi04;
  assign new_new_n18191__ = pi05 & ~new_new_n18190__;
  assign new_new_n18192__ = pi03 & ~new_new_n18191__;
  assign new_new_n18193__ = ~pi02 & ~pi04;
  assign new_new_n18194__ = ~pi05 & ~new_new_n18193__;
  assign new_new_n18195__ = ~new_new_n18146__ & ~new_new_n18194__;
  assign new_new_n18196__ = ~new_new_n18192__ & new_new_n18195__;
  assign new_new_n18197__ = new_new_n18189__ & ~new_new_n18196__;
  assign new_new_n18198__ = ~new_new_n18148__ & ~new_new_n18197__;
  assign new_new_n18199__ = ~new_new_n15560__ & ~new_new_n15767__;
  assign new_new_n18200__ = ~new_new_n15761__ & new_new_n15767__;
  assign new_new_n18201__ = new_new_n15560__ & new_new_n15761__;
  assign new_new_n18202__ = ~new_new_n18200__ & ~new_new_n18201__;
  assign new_new_n18203__ = new_new_n765__ & ~new_new_n18202__;
  assign new_new_n18204__ = ~new_new_n18199__ & ~new_new_n18203__;
  assign new_new_n18205__ = new_new_n15533__ & ~new_new_n18204__;
  assign new_new_n18206__ = ~new_new_n71__ & ~new_new_n15763__;
  assign new_new_n18207__ = ~new_new_n161__ & ~new_new_n15767__;
  assign new_new_n18208__ = ~new_new_n18206__ & new_new_n18207__;
  assign new_new_n18209__ = ~new_new_n15533__ & new_new_n15767__;
  assign new_new_n18210__ = new_new_n15761__ & new_new_n18209__;
  assign new_new_n18211__ = ~new_new_n161__ & ~new_new_n18210__;
  assign new_new_n18212__ = ~new_new_n71__ & ~new_new_n15560__;
  assign new_new_n18213__ = ~new_new_n18211__ & new_new_n18212__;
  assign new_new_n18214__ = ~new_new_n18208__ & ~new_new_n18213__;
  assign new_new_n18215__ = ~new_new_n18205__ & new_new_n18214__;
  assign new_new_n18216__ = pi31 & ~new_new_n18215__;
  assign new_new_n18217__ = new_new_n765__ & ~new_new_n15533__;
  assign new_new_n18218__ = new_new_n161__ & new_new_n15767__;
  assign new_new_n18219__ = ~pi31 & ~new_new_n18218__;
  assign new_new_n18220__ = ~new_new_n18217__ & new_new_n18219__;
  assign new_new_n18221__ = ~new_new_n18216__ & ~new_new_n18220__;
  assign new_new_n18222__ = ~new_new_n277__ & ~new_new_n1372__;
  assign new_new_n18223__ = new_new_n81__ & ~new_new_n5390__;
  assign new_new_n18224__ = ~new_new_n168__ & ~new_new_n213__;
  assign new_new_n18225__ = ~new_new_n1113__ & new_new_n18224__;
  assign new_new_n18226__ = ~new_new_n189__ & ~new_new_n961__;
  assign new_new_n18227__ = ~new_new_n1008__ & new_new_n1740__;
  assign new_new_n18228__ = new_new_n3958__ & new_new_n17500__;
  assign new_new_n18229__ = ~new_new_n18223__ & new_new_n18228__;
  assign new_new_n18230__ = new_new_n18226__ & new_new_n18227__;
  assign new_new_n18231__ = new_new_n3564__ & new_new_n18225__;
  assign new_new_n18232__ = new_new_n4963__ & new_new_n18222__;
  assign new_new_n18233__ = new_new_n18231__ & new_new_n18232__;
  assign new_new_n18234__ = new_new_n18229__ & new_new_n18230__;
  assign new_new_n18235__ = new_new_n116__ & ~new_new_n1539__;
  assign new_new_n18236__ = new_new_n18234__ & new_new_n18235__;
  assign new_new_n18237__ = new_new_n834__ & new_new_n18233__;
  assign new_new_n18238__ = new_new_n18236__ & new_new_n18237__;
  assign new_new_n18239__ = new_new_n742__ & new_new_n18238__;
  assign new_new_n18240__ = new_new_n2255__ & new_new_n18239__;
  assign new_new_n18241__ = new_new_n2452__ & new_new_n18240__;
  assign new_new_n18242__ = new_new_n18221__ & ~new_new_n18241__;
  assign new_new_n18243__ = ~new_new_n17563__ & ~new_new_n18242__;
  assign new_new_n18244__ = new_new_n18198__ & ~new_new_n18243__;
  assign new_new_n18245__ = ~new_new_n18221__ & new_new_n18241__;
  assign new_new_n18246__ = new_new_n17563__ & ~new_new_n18245__;
  assign new_new_n18247__ = ~new_new_n18244__ & ~new_new_n18246__;
  assign new_new_n18248__ = ~new_new_n18145__ & ~new_new_n18247__;
  assign new_new_n18249__ = ~new_new_n18144__ & ~new_new_n18248__;
  assign new_new_n18250__ = new_new_n4815__ & new_new_n15464__;
  assign new_new_n18251__ = new_new_n4212__ & ~new_new_n15471__;
  assign new_new_n18252__ = new_new_n4813__ & new_new_n15819__;
  assign new_new_n18253__ = ~new_new_n18250__ & ~new_new_n18251__;
  assign new_new_n18254__ = ~new_new_n18252__ & new_new_n18253__;
  assign new_new_n18255__ = ~pi29 & ~new_new_n18254__;
  assign new_new_n18256__ = new_new_n4221__ & ~new_new_n15809__;
  assign new_new_n18257__ = pi29 & ~new_new_n18256__;
  assign new_new_n18258__ = new_new_n66__ & ~new_new_n15809__;
  assign new_new_n18259__ = ~new_new_n18257__ & ~new_new_n18258__;
  assign new_new_n18260__ = new_new_n18254__ & ~new_new_n18259__;
  assign new_new_n18261__ = ~new_new_n18255__ & ~new_new_n18260__;
  assign new_new_n18262__ = new_new_n18249__ & new_new_n18261__;
  assign new_new_n18263__ = ~new_new_n18249__ & ~new_new_n18261__;
  assign new_new_n18264__ = ~new_new_n17595__ & ~new_new_n17646__;
  assign new_new_n18265__ = new_new_n17420__ & ~new_new_n18264__;
  assign new_new_n18266__ = ~new_new_n17420__ & new_new_n18264__;
  assign new_new_n18267__ = ~new_new_n18265__ & ~new_new_n18266__;
  assign new_new_n18268__ = ~new_new_n18263__ & new_new_n18267__;
  assign new_new_n18269__ = ~new_new_n18262__ & ~new_new_n18268__;
  assign new_new_n18270__ = ~new_new_n18119__ & new_new_n18269__;
  assign new_new_n18271__ = new_new_n18119__ & ~new_new_n18269__;
  assign new_new_n18272__ = ~new_new_n333__ & ~new_new_n15432__;
  assign new_new_n18273__ = new_new_n873__ & ~new_new_n15362__;
  assign new_new_n18274__ = ~new_new_n18272__ & ~new_new_n18273__;
  assign new_new_n18275__ = new_new_n801__ & ~new_new_n17918__;
  assign new_new_n18276__ = pi26 & ~new_new_n18275__;
  assign new_new_n18277__ = pi25 & new_new_n15390__;
  assign new_new_n18278__ = ~pi25 & ~new_new_n15390__;
  assign new_new_n18279__ = ~new_new_n110__ & new_new_n15829__;
  assign new_new_n18280__ = ~new_new_n18277__ & ~new_new_n18278__;
  assign new_new_n18281__ = new_new_n18279__ & new_new_n18280__;
  assign new_new_n18282__ = ~new_new_n18276__ & ~new_new_n18281__;
  assign new_new_n18283__ = new_new_n18274__ & ~new_new_n18282__;
  assign new_new_n18284__ = new_new_n801__ & new_new_n17914__;
  assign new_new_n18285__ = new_new_n18274__ & ~new_new_n18284__;
  assign new_new_n18286__ = ~pi26 & ~new_new_n18285__;
  assign new_new_n18287__ = ~new_new_n18283__ & ~new_new_n18286__;
  assign new_new_n18288__ = ~new_new_n18271__ & ~new_new_n18287__;
  assign new_new_n18289__ = ~new_new_n18270__ & ~new_new_n18288__;
  assign new_new_n18290__ = new_new_n18115__ & ~new_new_n18289__;
  assign new_new_n18291__ = ~new_new_n18115__ & new_new_n18289__;
  assign new_new_n18292__ = ~new_new_n18290__ & ~new_new_n18291__;
  assign new_new_n18293__ = ~new_new_n18046__ & ~new_new_n18047__;
  assign new_new_n18294__ = ~new_new_n18057__ & new_new_n18293__;
  assign new_new_n18295__ = new_new_n18057__ & ~new_new_n18293__;
  assign new_new_n18296__ = ~new_new_n18294__ & ~new_new_n18295__;
  assign new_new_n18297__ = new_new_n18292__ & ~new_new_n18296__;
  assign new_new_n18298__ = ~new_new_n18290__ & ~new_new_n18297__;
  assign new_new_n18299__ = ~new_new_n18060__ & ~new_new_n18061__;
  assign new_new_n18300__ = ~new_new_n18071__ & ~new_new_n18299__;
  assign new_new_n18301__ = new_new_n18071__ & new_new_n18299__;
  assign new_new_n18302__ = ~new_new_n18300__ & ~new_new_n18301__;
  assign new_new_n18303__ = ~new_new_n18298__ & new_new_n18302__;
  assign new_new_n18304__ = new_new_n18298__ & ~new_new_n18302__;
  assign new_new_n18305__ = new_new_n5213__ & new_new_n15285__;
  assign new_new_n18306__ = new_new_n5191__ & ~new_new_n15321__;
  assign new_new_n18307__ = new_new_n5183__ & ~new_new_n15273__;
  assign new_new_n18308__ = new_new_n5215__ & new_new_n16078__;
  assign new_new_n18309__ = ~new_new_n18306__ & ~new_new_n18307__;
  assign new_new_n18310__ = ~new_new_n18305__ & new_new_n18309__;
  assign new_new_n18311__ = ~new_new_n18308__ & new_new_n18310__;
  assign new_new_n18312__ = ~pi23 & ~new_new_n18311__;
  assign new_new_n18313__ = pi23 & new_new_n18311__;
  assign new_new_n18314__ = ~new_new_n18312__ & ~new_new_n18313__;
  assign new_new_n18315__ = ~new_new_n18304__ & ~new_new_n18314__;
  assign new_new_n18316__ = ~new_new_n18303__ & ~new_new_n18315__;
  assign new_new_n18317__ = new_new_n6936__ & ~new_new_n16603__;
  assign new_new_n18318__ = new_new_n6629__ & new_new_n15244__;
  assign new_new_n18319__ = new_new_n6634__ & new_new_n15237__;
  assign new_new_n18320__ = ~new_new_n18318__ & ~new_new_n18319__;
  assign new_new_n18321__ = ~new_new_n18317__ & new_new_n18320__;
  assign new_new_n18322__ = ~pi20 & ~new_new_n18321__;
  assign new_new_n18323__ = new_new_n6623__ & ~new_new_n15248__;
  assign new_new_n18324__ = pi20 & ~new_new_n18323__;
  assign new_new_n18325__ = new_new_n9920__ & ~new_new_n15248__;
  assign new_new_n18326__ = ~new_new_n18324__ & ~new_new_n18325__;
  assign new_new_n18327__ = new_new_n18321__ & ~new_new_n18326__;
  assign new_new_n18328__ = ~new_new_n18322__ & ~new_new_n18327__;
  assign new_new_n18329__ = new_new_n18073__ & ~new_new_n18328__;
  assign new_new_n18330__ = ~new_new_n18073__ & new_new_n18328__;
  assign new_new_n18331__ = ~new_new_n18329__ & ~new_new_n18330__;
  assign new_new_n18332__ = ~new_new_n18088__ & ~new_new_n18090__;
  assign new_new_n18333__ = new_new_n18331__ & new_new_n18332__;
  assign new_new_n18334__ = ~new_new_n18331__ & ~new_new_n18332__;
  assign new_new_n18335__ = ~new_new_n18333__ & ~new_new_n18334__;
  assign new_new_n18336__ = ~new_new_n18316__ & ~new_new_n18335__;
  assign new_new_n18337__ = ~new_new_n18328__ & new_new_n18335__;
  assign new_new_n18338__ = ~new_new_n18336__ & ~new_new_n18337__;
  assign new_new_n18339__ = ~new_new_n18099__ & ~new_new_n18338__;
  assign new_new_n18340__ = ~new_new_n18098__ & ~new_new_n18339__;
  assign new_new_n18341__ = ~new_new_n18098__ & ~new_new_n18099__;
  assign new_new_n18342__ = new_new_n18338__ & new_new_n18341__;
  assign new_new_n18343__ = ~new_new_n18338__ & ~new_new_n18341__;
  assign new_new_n18344__ = ~new_new_n18342__ & ~new_new_n18343__;
  assign new_new_n18345__ = new_new_n6968__ & ~new_new_n15998__;
  assign new_new_n18346__ = new_new_n6955__ & new_new_n16051__;
  assign new_new_n18347__ = new_new_n6958__ & ~new_new_n16056__;
  assign new_new_n18348__ = ~new_new_n18346__ & new_new_n18347__;
  assign new_new_n18349__ = ~new_new_n18345__ & ~new_new_n18348__;
  assign new_new_n18350__ = new_new_n10337__ & new_new_n15905__;
  assign new_new_n18351__ = pi17 & ~new_new_n18350__;
  assign new_new_n18352__ = new_new_n10340__ & new_new_n15905__;
  assign new_new_n18353__ = ~pi17 & ~new_new_n18352__;
  assign new_new_n18354__ = pi14 & ~new_new_n18353__;
  assign new_new_n18355__ = ~new_new_n18351__ & ~new_new_n18354__;
  assign new_new_n18356__ = new_new_n18349__ & ~new_new_n18355__;
  assign new_new_n18357__ = ~pi17 & ~new_new_n18349__;
  assign new_new_n18358__ = ~new_new_n18356__ & ~new_new_n18357__;
  assign new_new_n18359__ = new_new_n18316__ & new_new_n18335__;
  assign new_new_n18360__ = ~new_new_n18336__ & ~new_new_n18359__;
  assign new_new_n18361__ = new_new_n6634__ & new_new_n15244__;
  assign new_new_n18362__ = new_new_n6629__ & ~new_new_n15248__;
  assign new_new_n18363__ = ~new_new_n6625__ & ~new_new_n15314__;
  assign new_new_n18364__ = ~new_new_n18362__ & ~new_new_n18363__;
  assign new_new_n18365__ = ~new_new_n18361__ & new_new_n18364__;
  assign new_new_n18366__ = new_new_n6631__ & new_new_n16378__;
  assign new_new_n18367__ = ~pi20 & ~new_new_n18366__;
  assign new_new_n18368__ = new_new_n7015__ & new_new_n16378__;
  assign new_new_n18369__ = ~new_new_n18367__ & ~new_new_n18368__;
  assign new_new_n18370__ = new_new_n18365__ & ~new_new_n18369__;
  assign new_new_n18371__ = pi20 & ~new_new_n18365__;
  assign new_new_n18372__ = ~new_new_n18370__ & ~new_new_n18371__;
  assign new_new_n18373__ = ~new_new_n18303__ & ~new_new_n18304__;
  assign new_new_n18374__ = ~new_new_n18314__ & new_new_n18373__;
  assign new_new_n18375__ = new_new_n18314__ & ~new_new_n18373__;
  assign new_new_n18376__ = ~new_new_n18374__ & ~new_new_n18375__;
  assign new_new_n18377__ = ~new_new_n18372__ & ~new_new_n18376__;
  assign new_new_n18378__ = new_new_n18372__ & new_new_n18376__;
  assign new_new_n18379__ = new_new_n5213__ & ~new_new_n15273__;
  assign new_new_n18380__ = new_new_n5191__ & ~new_new_n15349__;
  assign new_new_n18381__ = new_new_n5183__ & ~new_new_n15321__;
  assign new_new_n18382__ = ~new_new_n18380__ & ~new_new_n18381__;
  assign new_new_n18383__ = ~new_new_n18379__ & new_new_n18382__;
  assign new_new_n18384__ = new_new_n5195__ & ~new_new_n17103__;
  assign new_new_n18385__ = pi23 & ~new_new_n18384__;
  assign new_new_n18386__ = new_new_n7878__ & ~new_new_n17103__;
  assign new_new_n18387__ = ~new_new_n18385__ & ~new_new_n18386__;
  assign new_new_n18388__ = new_new_n18383__ & ~new_new_n18387__;
  assign new_new_n18389__ = ~pi23 & ~new_new_n18383__;
  assign new_new_n18390__ = ~new_new_n18388__ & ~new_new_n18389__;
  assign new_new_n18391__ = ~new_new_n18292__ & new_new_n18296__;
  assign new_new_n18392__ = ~new_new_n18297__ & ~new_new_n18391__;
  assign new_new_n18393__ = new_new_n5183__ & ~new_new_n15349__;
  assign new_new_n18394__ = new_new_n5191__ & ~new_new_n15398__;
  assign new_new_n18395__ = new_new_n5213__ & ~new_new_n15321__;
  assign new_new_n18396__ = ~new_new_n18393__ & ~new_new_n18394__;
  assign new_new_n18397__ = ~new_new_n18395__ & new_new_n18396__;
  assign new_new_n18398__ = new_new_n5195__ & new_new_n16458__;
  assign new_new_n18399__ = pi23 & ~new_new_n18398__;
  assign new_new_n18400__ = new_new_n7878__ & new_new_n16458__;
  assign new_new_n18401__ = ~new_new_n18399__ & ~new_new_n18400__;
  assign new_new_n18402__ = new_new_n18397__ & ~new_new_n18401__;
  assign new_new_n18403__ = ~pi23 & ~new_new_n18397__;
  assign new_new_n18404__ = ~new_new_n18402__ & ~new_new_n18403__;
  assign new_new_n18405__ = ~new_new_n18270__ & ~new_new_n18271__;
  assign new_new_n18406__ = new_new_n18287__ & new_new_n18405__;
  assign new_new_n18407__ = ~new_new_n18287__ & ~new_new_n18405__;
  assign new_new_n18408__ = ~new_new_n18406__ & ~new_new_n18407__;
  assign new_new_n18409__ = new_new_n18404__ & new_new_n18408__;
  assign new_new_n18410__ = ~new_new_n18404__ & ~new_new_n18408__;
  assign new_new_n18411__ = new_new_n3311__ & ~new_new_n15362__;
  assign new_new_n18412__ = new_new_n873__ & ~new_new_n15432__;
  assign new_new_n18413__ = ~new_new_n4900__ & new_new_n16771__;
  assign new_new_n18414__ = ~new_new_n18411__ & ~new_new_n18412__;
  assign new_new_n18415__ = ~new_new_n18413__ & new_new_n18414__;
  assign new_new_n18416__ = new_new_n303__ & ~new_new_n15439__;
  assign new_new_n18417__ = pi26 & ~new_new_n18416__;
  assign new_new_n18418__ = new_new_n145__ & ~new_new_n15439__;
  assign new_new_n18419__ = ~pi26 & ~new_new_n18418__;
  assign new_new_n18420__ = pi23 & ~new_new_n18419__;
  assign new_new_n18421__ = ~new_new_n18417__ & ~new_new_n18420__;
  assign new_new_n18422__ = new_new_n18415__ & ~new_new_n18421__;
  assign new_new_n18423__ = ~pi26 & ~new_new_n18415__;
  assign new_new_n18424__ = ~new_new_n18422__ & ~new_new_n18423__;
  assign new_new_n18425__ = new_new_n71__ & new_new_n15533__;
  assign new_new_n18426__ = ~new_new_n71__ & new_new_n15520__;
  assign new_new_n18427__ = new_new_n18125__ & new_new_n18426__;
  assign new_new_n18428__ = ~new_new_n161__ & ~new_new_n18427__;
  assign new_new_n18429__ = ~new_new_n15767__ & ~new_new_n18428__;
  assign new_new_n18430__ = new_new_n15533__ & new_new_n15770__;
  assign new_new_n18431__ = ~new_new_n15520__ & ~new_new_n18125__;
  assign new_new_n18432__ = ~new_new_n18430__ & new_new_n18431__;
  assign new_new_n18433__ = new_new_n18430__ & ~new_new_n18431__;
  assign new_new_n18434__ = ~new_new_n18432__ & ~new_new_n18433__;
  assign new_new_n18435__ = new_new_n765__ & ~new_new_n18434__;
  assign new_new_n18436__ = ~new_new_n18429__ & ~new_new_n18435__;
  assign new_new_n18437__ = pi31 & ~new_new_n18436__;
  assign new_new_n18438__ = pi29 & ~new_new_n15533__;
  assign new_new_n18439__ = new_new_n15853__ & ~new_new_n18438__;
  assign new_new_n18440__ = ~new_new_n18130__ & ~new_new_n18439__;
  assign new_new_n18441__ = ~pi31 & ~new_new_n18440__;
  assign new_new_n18442__ = ~new_new_n18425__ & ~new_new_n18441__;
  assign new_new_n18443__ = ~new_new_n18437__ & new_new_n18442__;
  assign new_new_n18444__ = new_new_n161__ & new_new_n15560__;
  assign new_new_n18445__ = new_new_n765__ & new_new_n15767__;
  assign new_new_n18446__ = ~new_new_n18444__ & ~new_new_n18445__;
  assign new_new_n18447__ = ~pi31 & ~new_new_n18446__;
  assign new_new_n18448__ = new_new_n71__ & new_new_n15560__;
  assign new_new_n18449__ = new_new_n161__ & new_new_n15572__;
  assign new_new_n18450__ = new_new_n15761__ & ~new_new_n15767__;
  assign new_new_n18451__ = ~new_new_n18200__ & ~new_new_n18450__;
  assign new_new_n18452__ = ~new_new_n15560__ & new_new_n18451__;
  assign new_new_n18453__ = new_new_n15560__ & ~new_new_n18451__;
  assign new_new_n18454__ = ~new_new_n18452__ & ~new_new_n18453__;
  assign new_new_n18455__ = new_new_n765__ & ~new_new_n18454__;
  assign new_new_n18456__ = ~new_new_n18448__ & ~new_new_n18449__;
  assign new_new_n18457__ = ~new_new_n18455__ & new_new_n18456__;
  assign new_new_n18458__ = pi31 & ~new_new_n18457__;
  assign new_new_n18459__ = ~new_new_n18447__ & ~new_new_n18458__;
  assign new_new_n18460__ = new_new_n11466__ & ~new_new_n14393__;
  assign new_new_n18461__ = ~new_new_n14393__ & new_new_n18189__;
  assign new_new_n18462__ = ~new_new_n11466__ & ~new_new_n18461__;
  assign new_new_n18463__ = ~pi02 & ~new_new_n18460__;
  assign new_new_n18464__ = ~new_new_n18462__ & new_new_n18463__;
  assign new_new_n18465__ = new_new_n18189__ & ~new_new_n18464__;
  assign new_new_n18466__ = new_new_n18146__ & new_new_n18462__;
  assign new_new_n18467__ = ~new_new_n18465__ & ~new_new_n18466__;
  assign new_new_n18468__ = ~pi05 & ~new_new_n18467__;
  assign new_new_n18469__ = new_new_n6811__ & ~new_new_n11467__;
  assign new_new_n18470__ = ~pi02 & new_new_n14393__;
  assign new_new_n18471__ = ~new_new_n18147__ & new_new_n18470__;
  assign new_new_n18472__ = ~new_new_n18469__ & ~new_new_n18471__;
  assign new_new_n18473__ = ~new_new_n18189__ & ~new_new_n18472__;
  assign new_new_n18474__ = ~new_new_n12828__ & ~new_new_n18146__;
  assign new_new_n18475__ = ~new_new_n12829__ & ~new_new_n18474__;
  assign new_new_n18476__ = new_new_n18189__ & new_new_n18475__;
  assign new_new_n18477__ = ~new_new_n18473__ & ~new_new_n18476__;
  assign new_new_n18478__ = ~new_new_n18468__ & new_new_n18477__;
  assign new_new_n18479__ = ~new_new_n18459__ & ~new_new_n18478__;
  assign new_new_n18480__ = new_new_n18459__ & new_new_n18478__;
  assign new_new_n18481__ = ~new_new_n747__ & ~new_new_n1080__;
  assign new_new_n18482__ = ~new_new_n385__ & ~new_new_n624__;
  assign new_new_n18483__ = ~new_new_n724__ & new_new_n18482__;
  assign new_new_n18484__ = new_new_n6296__ & new_new_n18483__;
  assign new_new_n18485__ = new_new_n227__ & new_new_n743__;
  assign new_new_n18486__ = new_new_n1037__ & new_new_n2331__;
  assign new_new_n18487__ = new_new_n2453__ & new_new_n3904__;
  assign new_new_n18488__ = new_new_n5566__ & new_new_n18222__;
  assign new_new_n18489__ = new_new_n18481__ & new_new_n18488__;
  assign new_new_n18490__ = new_new_n18486__ & new_new_n18487__;
  assign new_new_n18491__ = new_new_n18484__ & new_new_n18485__;
  assign new_new_n18492__ = new_new_n2478__ & new_new_n4235__;
  assign new_new_n18493__ = new_new_n18491__ & new_new_n18492__;
  assign new_new_n18494__ = new_new_n18489__ & new_new_n18490__;
  assign new_new_n18495__ = new_new_n1290__ & new_new_n16263__;
  assign new_new_n18496__ = new_new_n18494__ & new_new_n18495__;
  assign new_new_n18497__ = new_new_n1407__ & new_new_n18493__;
  assign new_new_n18498__ = new_new_n18496__ & new_new_n18497__;
  assign new_new_n18499__ = new_new_n18175__ & new_new_n18498__;
  assign new_new_n18500__ = new_new_n71__ & new_new_n15615__;
  assign new_new_n18501__ = pi31 & ~new_new_n18500__;
  assign new_new_n18502__ = new_new_n161__ & new_new_n15615__;
  assign new_new_n18503__ = ~new_new_n161__ & ~new_new_n15564__;
  assign new_new_n18504__ = ~new_new_n71__ & ~new_new_n18502__;
  assign new_new_n18505__ = ~new_new_n18503__ & new_new_n18504__;
  assign new_new_n18506__ = ~new_new_n18501__ & ~new_new_n18505__;
  assign new_new_n18507__ = new_new_n15564__ & new_new_n15755__;
  assign new_new_n18508__ = ~new_new_n15564__ & ~new_new_n15755__;
  assign new_new_n18509__ = ~new_new_n18507__ & ~new_new_n18508__;
  assign new_new_n18510__ = ~new_new_n15615__ & ~new_new_n18509__;
  assign new_new_n18511__ = new_new_n15615__ & new_new_n18509__;
  assign new_new_n18512__ = ~new_new_n18510__ & ~new_new_n18511__;
  assign new_new_n18513__ = ~new_new_n71__ & ~new_new_n18512__;
  assign new_new_n18514__ = ~new_new_n161__ & ~new_new_n18513__;
  assign new_new_n18515__ = new_new_n161__ & new_new_n15743__;
  assign new_new_n18516__ = pi31 & ~new_new_n18515__;
  assign new_new_n18517__ = ~new_new_n18514__ & new_new_n18516__;
  assign new_new_n18518__ = ~new_new_n18506__ & ~new_new_n18517__;
  assign new_new_n18519__ = new_new_n2077__ & new_new_n6240__;
  assign new_new_n18520__ = new_new_n16223__ & new_new_n18519__;
  assign new_new_n18521__ = new_new_n697__ & new_new_n18520__;
  assign new_new_n18522__ = ~new_new_n895__ & new_new_n18521__;
  assign new_new_n18523__ = ~new_new_n482__ & ~new_new_n510__;
  assign new_new_n18524__ = ~new_new_n693__ & ~new_new_n890__;
  assign new_new_n18525__ = new_new_n18523__ & new_new_n18524__;
  assign new_new_n18526__ = new_new_n1942__ & new_new_n2166__;
  assign new_new_n18527__ = new_new_n2333__ & new_new_n2708__;
  assign new_new_n18528__ = ~new_new_n7417__ & new_new_n18527__;
  assign new_new_n18529__ = new_new_n18525__ & new_new_n18526__;
  assign new_new_n18530__ = ~new_new_n607__ & new_new_n18529__;
  assign new_new_n18531__ = new_new_n440__ & new_new_n18528__;
  assign new_new_n18532__ = new_new_n3791__ & new_new_n18531__;
  assign new_new_n18533__ = new_new_n18530__ & new_new_n18532__;
  assign new_new_n18534__ = new_new_n2321__ & new_new_n18522__;
  assign new_new_n18535__ = new_new_n18533__ & new_new_n18534__;
  assign new_new_n18536__ = ~new_new_n671__ & ~new_new_n781__;
  assign new_new_n18537__ = ~new_new_n88__ & ~new_new_n383__;
  assign new_new_n18538__ = ~new_new_n634__ & new_new_n18537__;
  assign new_new_n18539__ = new_new_n2424__ & new_new_n18538__;
  assign new_new_n18540__ = new_new_n18536__ & new_new_n18539__;
  assign new_new_n18541__ = new_new_n18535__ & new_new_n18540__;
  assign new_new_n18542__ = ~new_new_n106__ & ~new_new_n248__;
  assign new_new_n18543__ = ~new_new_n480__ & ~new_new_n838__;
  assign new_new_n18544__ = ~new_new_n1212__ & new_new_n18543__;
  assign new_new_n18545__ = ~new_new_n123__ & new_new_n18542__;
  assign new_new_n18546__ = ~new_new_n828__ & new_new_n18545__;
  assign new_new_n18547__ = new_new_n720__ & new_new_n18544__;
  assign new_new_n18548__ = new_new_n18546__ & new_new_n18547__;
  assign new_new_n18549__ = ~new_new_n379__ & ~new_new_n509__;
  assign new_new_n18550__ = ~new_new_n937__ & new_new_n18549__;
  assign new_new_n18551__ = ~new_new_n17391__ & new_new_n18550__;
  assign new_new_n18552__ = new_new_n1215__ & new_new_n2540__;
  assign new_new_n18553__ = new_new_n6322__ & new_new_n18552__;
  assign new_new_n18554__ = new_new_n1969__ & new_new_n18551__;
  assign new_new_n18555__ = new_new_n2028__ & new_new_n17598__;
  assign new_new_n18556__ = new_new_n18554__ & new_new_n18555__;
  assign new_new_n18557__ = new_new_n2327__ & new_new_n18553__;
  assign new_new_n18558__ = new_new_n18548__ & new_new_n18557__;
  assign new_new_n18559__ = new_new_n18556__ & new_new_n18558__;
  assign new_new_n18560__ = new_new_n16486__ & new_new_n18559__;
  assign new_new_n18561__ = new_new_n18541__ & new_new_n18560__;
  assign new_new_n18562__ = new_new_n18518__ & ~new_new_n18561__;
  assign new_new_n18563__ = ~new_new_n18499__ & new_new_n18562__;
  assign new_new_n18564__ = ~new_new_n18146__ & ~new_new_n18563__;
  assign new_new_n18565__ = ~new_new_n18518__ & new_new_n18561__;
  assign new_new_n18566__ = new_new_n18499__ & new_new_n18565__;
  assign new_new_n18567__ = ~new_new_n18564__ & ~new_new_n18566__;
  assign new_new_n18568__ = ~new_new_n701__ & ~new_new_n851__;
  assign new_new_n18569__ = ~new_new_n192__ & ~new_new_n322__;
  assign new_new_n18570__ = ~new_new_n835__ & ~new_new_n921__;
  assign new_new_n18571__ = ~new_new_n959__ & new_new_n4980__;
  assign new_new_n18572__ = new_new_n18568__ & new_new_n18571__;
  assign new_new_n18573__ = new_new_n18569__ & new_new_n18570__;
  assign new_new_n18574__ = new_new_n2515__ & new_new_n3687__;
  assign new_new_n18575__ = new_new_n6142__ & new_new_n18574__;
  assign new_new_n18576__ = new_new_n18572__ & new_new_n18573__;
  assign new_new_n18577__ = new_new_n7147__ & new_new_n18576__;
  assign new_new_n18578__ = new_new_n1776__ & new_new_n18575__;
  assign new_new_n18579__ = new_new_n3316__ & new_new_n18578__;
  assign new_new_n18580__ = new_new_n3966__ & new_new_n18577__;
  assign new_new_n18581__ = new_new_n18579__ & new_new_n18580__;
  assign new_new_n18582__ = new_new_n297__ & new_new_n18581__;
  assign new_new_n18583__ = new_new_n4497__ & new_new_n18582__;
  assign new_new_n18584__ = ~new_new_n18567__ & new_new_n18583__;
  assign new_new_n18585__ = new_new_n18146__ & ~new_new_n18584__;
  assign new_new_n18586__ = new_new_n18563__ & ~new_new_n18583__;
  assign new_new_n18587__ = ~new_new_n18585__ & ~new_new_n18586__;
  assign new_new_n18588__ = ~new_new_n18480__ & ~new_new_n18587__;
  assign new_new_n18589__ = ~new_new_n18479__ & ~new_new_n18588__;
  assign new_new_n18590__ = ~new_new_n4818__ & new_new_n15520__;
  assign new_new_n18591__ = new_new_n4212__ & new_new_n15524__;
  assign new_new_n18592__ = new_new_n4815__ & ~new_new_n15487__;
  assign new_new_n18593__ = ~new_new_n18590__ & ~new_new_n18591__;
  assign new_new_n18594__ = ~new_new_n18592__ & new_new_n18593__;
  assign new_new_n18595__ = new_new_n4214__ & new_new_n17587__;
  assign new_new_n18596__ = ~pi29 & ~new_new_n18595__;
  assign new_new_n18597__ = new_new_n5732__ & new_new_n17587__;
  assign new_new_n18598__ = ~new_new_n18596__ & ~new_new_n18597__;
  assign new_new_n18599__ = new_new_n18594__ & ~new_new_n18598__;
  assign new_new_n18600__ = pi29 & ~new_new_n18594__;
  assign new_new_n18601__ = ~new_new_n18599__ & ~new_new_n18600__;
  assign new_new_n18602__ = new_new_n18589__ & ~new_new_n18601__;
  assign new_new_n18603__ = ~new_new_n18589__ & new_new_n18601__;
  assign new_new_n18604__ = ~new_new_n18198__ & new_new_n18221__;
  assign new_new_n18605__ = new_new_n18198__ & ~new_new_n18221__;
  assign new_new_n18606__ = ~new_new_n18604__ & ~new_new_n18605__;
  assign new_new_n18607__ = new_new_n17563__ & new_new_n18606__;
  assign new_new_n18608__ = ~new_new_n17563__ & ~new_new_n18606__;
  assign new_new_n18609__ = ~new_new_n18607__ & ~new_new_n18608__;
  assign new_new_n18610__ = ~new_new_n18603__ & new_new_n18609__;
  assign new_new_n18611__ = ~new_new_n18602__ & ~new_new_n18610__;
  assign new_new_n18612__ = new_new_n18443__ & new_new_n18611__;
  assign new_new_n18613__ = ~new_new_n18443__ & ~new_new_n18611__;
  assign new_new_n18614__ = ~new_new_n18242__ & ~new_new_n18245__;
  assign new_new_n18615__ = ~new_new_n17563__ & ~new_new_n18604__;
  assign new_new_n18616__ = ~new_new_n18605__ & ~new_new_n18615__;
  assign new_new_n18617__ = new_new_n18614__ & new_new_n18616__;
  assign new_new_n18618__ = ~new_new_n18614__ & ~new_new_n18616__;
  assign new_new_n18619__ = ~new_new_n18617__ & ~new_new_n18618__;
  assign new_new_n18620__ = ~new_new_n18613__ & new_new_n18619__;
  assign new_new_n18621__ = ~new_new_n18612__ & ~new_new_n18620__;
  assign new_new_n18622__ = ~new_new_n18144__ & ~new_new_n18145__;
  assign new_new_n18623__ = new_new_n18247__ & ~new_new_n18622__;
  assign new_new_n18624__ = ~new_new_n18247__ & new_new_n18622__;
  assign new_new_n18625__ = ~new_new_n18623__ & ~new_new_n18624__;
  assign new_new_n18626__ = ~new_new_n18621__ & new_new_n18625__;
  assign new_new_n18627__ = new_new_n18621__ & ~new_new_n18625__;
  assign new_new_n18628__ = new_new_n15487__ & new_new_n15809__;
  assign new_new_n18629__ = ~new_new_n17464__ & ~new_new_n18628__;
  assign new_new_n18630__ = ~new_new_n18017__ & new_new_n18629__;
  assign new_new_n18631__ = ~new_new_n15471__ & ~new_new_n18630__;
  assign new_new_n18632__ = new_new_n15471__ & new_new_n18630__;
  assign new_new_n18633__ = ~new_new_n18631__ & ~new_new_n18632__;
  assign new_new_n18634__ = new_new_n4813__ & ~new_new_n18633__;
  assign new_new_n18635__ = ~new_new_n4818__ & ~new_new_n15487__;
  assign new_new_n18636__ = new_new_n4212__ & ~new_new_n15809__;
  assign new_new_n18637__ = new_new_n4815__ & ~new_new_n15471__;
  assign new_new_n18638__ = ~new_new_n18635__ & ~new_new_n18636__;
  assign new_new_n18639__ = ~new_new_n18637__ & new_new_n18638__;
  assign new_new_n18640__ = ~new_new_n18634__ & new_new_n18639__;
  assign new_new_n18641__ = pi29 & ~new_new_n18640__;
  assign new_new_n18642__ = ~pi29 & new_new_n18640__;
  assign new_new_n18643__ = ~new_new_n18641__ & ~new_new_n18642__;
  assign new_new_n18644__ = ~new_new_n18627__ & new_new_n18643__;
  assign new_new_n18645__ = ~new_new_n18626__ & ~new_new_n18644__;
  assign new_new_n18646__ = new_new_n18424__ & new_new_n18645__;
  assign new_new_n18647__ = ~new_new_n18424__ & ~new_new_n18645__;
  assign new_new_n18648__ = ~new_new_n18262__ & ~new_new_n18263__;
  assign new_new_n18649__ = ~new_new_n18267__ & new_new_n18648__;
  assign new_new_n18650__ = new_new_n18267__ & ~new_new_n18648__;
  assign new_new_n18651__ = ~new_new_n18649__ & ~new_new_n18650__;
  assign new_new_n18652__ = ~new_new_n18647__ & ~new_new_n18651__;
  assign new_new_n18653__ = ~new_new_n18646__ & ~new_new_n18652__;
  assign new_new_n18654__ = ~new_new_n18410__ & ~new_new_n18653__;
  assign new_new_n18655__ = ~new_new_n18409__ & ~new_new_n18654__;
  assign new_new_n18656__ = new_new_n18392__ & new_new_n18655__;
  assign new_new_n18657__ = new_new_n18390__ & ~new_new_n18656__;
  assign new_new_n18658__ = ~new_new_n18392__ & ~new_new_n18655__;
  assign new_new_n18659__ = ~new_new_n18657__ & ~new_new_n18658__;
  assign new_new_n18660__ = ~new_new_n18378__ & ~new_new_n18659__;
  assign new_new_n18661__ = ~new_new_n18377__ & ~new_new_n18660__;
  assign new_new_n18662__ = new_new_n18360__ & new_new_n18661__;
  assign new_new_n18663__ = new_new_n18358__ & ~new_new_n18662__;
  assign new_new_n18664__ = ~new_new_n18360__ & ~new_new_n18661__;
  assign new_new_n18665__ = ~new_new_n18663__ & ~new_new_n18664__;
  assign new_new_n18666__ = new_new_n18344__ & ~new_new_n18665__;
  assign new_new_n18667__ = ~new_new_n18344__ & new_new_n18665__;
  assign new_new_n18668__ = new_new_n6964__ & ~new_new_n15998__;
  assign new_new_n18669__ = new_new_n6959__ & new_new_n16630__;
  assign new_new_n18670__ = new_new_n6968__ & ~new_new_n16056__;
  assign new_new_n18671__ = ~new_new_n7935__ & ~new_new_n18670__;
  assign new_new_n18672__ = ~new_new_n18668__ & new_new_n18671__;
  assign new_new_n18673__ = ~new_new_n18669__ & new_new_n18672__;
  assign new_new_n18674__ = pi17 & ~new_new_n18673__;
  assign new_new_n18675__ = ~pi17 & new_new_n18673__;
  assign new_new_n18676__ = ~new_new_n18674__ & ~new_new_n18675__;
  assign new_new_n18677__ = ~new_new_n18667__ & ~new_new_n18676__;
  assign new_new_n18678__ = ~new_new_n18666__ & ~new_new_n18677__;
  assign new_new_n18679__ = new_new_n18340__ & ~new_new_n18678__;
  assign new_new_n18680__ = new_new_n6634__ & ~new_new_n15998__;
  assign new_new_n18681__ = ~new_new_n6625__ & new_new_n15237__;
  assign new_new_n18682__ = new_new_n6629__ & new_new_n15905__;
  assign new_new_n18683__ = new_new_n6936__ & new_new_n16025__;
  assign new_new_n18684__ = ~new_new_n18681__ & ~new_new_n18682__;
  assign new_new_n18685__ = ~new_new_n18680__ & new_new_n18684__;
  assign new_new_n18686__ = ~new_new_n18683__ & new_new_n18685__;
  assign new_new_n18687__ = pi20 & ~new_new_n18686__;
  assign new_new_n18688__ = ~pi20 & new_new_n18686__;
  assign new_new_n18689__ = ~new_new_n18687__ & ~new_new_n18688__;
  assign new_new_n18690__ = ~new_new_n17999__ & ~new_new_n18092__;
  assign new_new_n18691__ = ~new_new_n18093__ & ~new_new_n18690__;
  assign new_new_n18692__ = ~new_new_n18689__ & ~new_new_n18691__;
  assign new_new_n18693__ = new_new_n18689__ & new_new_n18691__;
  assign new_new_n18694__ = ~new_new_n17945__ & ~new_new_n17946__;
  assign new_new_n18695__ = ~new_new_n17950__ & new_new_n18694__;
  assign new_new_n18696__ = new_new_n17950__ & ~new_new_n18694__;
  assign new_new_n18697__ = ~new_new_n18695__ & ~new_new_n18696__;
  assign new_new_n18698__ = ~new_new_n18693__ & ~new_new_n18697__;
  assign new_new_n18699__ = ~new_new_n18692__ & ~new_new_n18698__;
  assign new_new_n18700__ = pi17 & ~new_new_n6962__;
  assign new_new_n18701__ = ~new_new_n6961__ & ~new_new_n18700__;
  assign new_new_n18702__ = new_new_n18699__ & new_new_n18701__;
  assign new_new_n18703__ = ~new_new_n18699__ & ~new_new_n18701__;
  assign new_new_n18704__ = ~new_new_n18702__ & ~new_new_n18703__;
  assign new_new_n18705__ = ~new_new_n17954__ & new_new_n17970__;
  assign new_new_n18706__ = ~new_new_n17953__ & new_new_n17969__;
  assign new_new_n18707__ = ~new_new_n17968__ & ~new_new_n18706__;
  assign new_new_n18708__ = ~new_new_n18705__ & ~new_new_n18707__;
  assign new_new_n18709__ = new_new_n18704__ & ~new_new_n18708__;
  assign new_new_n18710__ = ~new_new_n18704__ & new_new_n18708__;
  assign new_new_n18711__ = ~new_new_n18709__ & ~new_new_n18710__;
  assign new_new_n18712__ = new_new_n18679__ & new_new_n18711__;
  assign new_new_n18713__ = ~new_new_n18692__ & ~new_new_n18693__;
  assign new_new_n18714__ = new_new_n18697__ & ~new_new_n18713__;
  assign new_new_n18715__ = ~new_new_n18697__ & new_new_n18713__;
  assign new_new_n18716__ = ~new_new_n18714__ & ~new_new_n18715__;
  assign new_new_n18717__ = ~pi14 & new_new_n6994__;
  assign new_new_n18718__ = pi13 & ~new_new_n16056__;
  assign new_new_n18719__ = new_new_n10772__ & ~new_new_n18718__;
  assign new_new_n18720__ = pi12 & ~new_new_n8820__;
  assign new_new_n18721__ = ~new_new_n18719__ & new_new_n18720__;
  assign new_new_n18722__ = pi14 & ~new_new_n6994__;
  assign new_new_n18723__ = new_new_n16056__ & new_new_n18722__;
  assign new_new_n18724__ = ~pi13 & ~new_new_n18723__;
  assign new_new_n18725__ = ~pi12 & ~new_new_n10771__;
  assign new_new_n18726__ = ~new_new_n18724__ & new_new_n18725__;
  assign new_new_n18727__ = ~new_new_n18717__ & ~new_new_n18721__;
  assign new_new_n18728__ = ~new_new_n18726__ & new_new_n18727__;
  assign new_new_n18729__ = new_new_n6959__ & new_new_n16025__;
  assign new_new_n18730__ = new_new_n6964__ & new_new_n15237__;
  assign new_new_n18731__ = new_new_n6968__ & new_new_n15905__;
  assign new_new_n18732__ = ~new_new_n18730__ & ~new_new_n18731__;
  assign new_new_n18733__ = ~new_new_n18729__ & new_new_n18732__;
  assign new_new_n18734__ = new_new_n6958__ & ~new_new_n15998__;
  assign new_new_n18735__ = ~pi17 & ~new_new_n18734__;
  assign new_new_n18736__ = new_new_n7942__ & ~new_new_n15998__;
  assign new_new_n18737__ = ~new_new_n18735__ & ~new_new_n18736__;
  assign new_new_n18738__ = new_new_n18733__ & ~new_new_n18737__;
  assign new_new_n18739__ = pi17 & ~new_new_n18733__;
  assign new_new_n18740__ = ~new_new_n18738__ & ~new_new_n18739__;
  assign new_new_n18741__ = new_new_n18392__ & ~new_new_n18655__;
  assign new_new_n18742__ = ~new_new_n18392__ & new_new_n18655__;
  assign new_new_n18743__ = ~new_new_n18741__ & ~new_new_n18742__;
  assign new_new_n18744__ = new_new_n18390__ & new_new_n18743__;
  assign new_new_n18745__ = ~new_new_n18390__ & ~new_new_n18743__;
  assign new_new_n18746__ = ~new_new_n18744__ & ~new_new_n18745__;
  assign new_new_n18747__ = new_new_n6629__ & new_new_n15285__;
  assign new_new_n18748__ = ~new_new_n6625__ & ~new_new_n15273__;
  assign new_new_n18749__ = new_new_n6936__ & new_new_n17140__;
  assign new_new_n18750__ = ~new_new_n18747__ & ~new_new_n18748__;
  assign new_new_n18751__ = ~new_new_n18749__ & new_new_n18750__;
  assign new_new_n18752__ = new_new_n6631__ & ~new_new_n15314__;
  assign new_new_n18753__ = ~pi20 & ~new_new_n18752__;
  assign new_new_n18754__ = new_new_n6640__ & ~new_new_n15314__;
  assign new_new_n18755__ = ~new_new_n18753__ & ~new_new_n18754__;
  assign new_new_n18756__ = new_new_n18751__ & ~new_new_n18755__;
  assign new_new_n18757__ = pi20 & ~new_new_n18751__;
  assign new_new_n18758__ = ~new_new_n18756__ & ~new_new_n18757__;
  assign new_new_n18759__ = ~new_new_n18409__ & ~new_new_n18410__;
  assign new_new_n18760__ = ~new_new_n18653__ & new_new_n18759__;
  assign new_new_n18761__ = new_new_n18653__ & ~new_new_n18759__;
  assign new_new_n18762__ = ~new_new_n18760__ & ~new_new_n18761__;
  assign new_new_n18763__ = ~new_new_n18758__ & new_new_n18762__;
  assign new_new_n18764__ = new_new_n18758__ & ~new_new_n18762__;
  assign new_new_n18765__ = ~new_new_n18646__ & ~new_new_n18647__;
  assign new_new_n18766__ = ~new_new_n18651__ & new_new_n18765__;
  assign new_new_n18767__ = new_new_n18651__ & ~new_new_n18765__;
  assign new_new_n18768__ = ~new_new_n18766__ & ~new_new_n18767__;
  assign new_new_n18769__ = new_new_n4815__ & ~new_new_n15809__;
  assign new_new_n18770__ = new_new_n4212__ & ~new_new_n15487__;
  assign new_new_n18771__ = new_new_n4813__ & new_new_n18020__;
  assign new_new_n18772__ = ~new_new_n18769__ & ~new_new_n18770__;
  assign new_new_n18773__ = ~new_new_n18771__ & new_new_n18772__;
  assign new_new_n18774__ = ~pi29 & ~new_new_n18773__;
  assign new_new_n18775__ = new_new_n66__ & new_new_n15524__;
  assign new_new_n18776__ = ~pi28 & new_new_n15524__;
  assign new_new_n18777__ = new_new_n4209__ & new_new_n18776__;
  assign new_new_n18778__ = pi29 & ~new_new_n18777__;
  assign new_new_n18779__ = ~new_new_n18775__ & ~new_new_n18778__;
  assign new_new_n18780__ = new_new_n18773__ & ~new_new_n18779__;
  assign new_new_n18781__ = ~new_new_n18774__ & ~new_new_n18780__;
  assign new_new_n18782__ = ~new_new_n18612__ & ~new_new_n18613__;
  assign new_new_n18783__ = new_new_n18619__ & new_new_n18782__;
  assign new_new_n18784__ = ~new_new_n18619__ & ~new_new_n18782__;
  assign new_new_n18785__ = ~new_new_n18783__ & ~new_new_n18784__;
  assign new_new_n18786__ = new_new_n18781__ & ~new_new_n18785__;
  assign new_new_n18787__ = ~new_new_n18781__ & new_new_n18785__;
  assign new_new_n18788__ = ~new_new_n4900__ & ~new_new_n17240__;
  assign new_new_n18789__ = ~new_new_n333__ & ~new_new_n15471__;
  assign new_new_n18790__ = new_new_n873__ & new_new_n15464__;
  assign new_new_n18791__ = ~new_new_n18789__ & ~new_new_n18790__;
  assign new_new_n18792__ = ~new_new_n18788__ & new_new_n18791__;
  assign new_new_n18793__ = pi26 & ~new_new_n18792__;
  assign new_new_n18794__ = new_new_n512__ & ~new_new_n15439__;
  assign new_new_n18795__ = new_new_n801__ & ~new_new_n15439__;
  assign new_new_n18796__ = ~pi26 & ~new_new_n18795__;
  assign new_new_n18797__ = ~new_new_n18794__ & ~new_new_n18796__;
  assign new_new_n18798__ = new_new_n18792__ & ~new_new_n18797__;
  assign new_new_n18799__ = ~new_new_n18793__ & ~new_new_n18798__;
  assign new_new_n18800__ = ~new_new_n18787__ & ~new_new_n18799__;
  assign new_new_n18801__ = ~new_new_n18786__ & ~new_new_n18800__;
  assign new_new_n18802__ = ~new_new_n18626__ & ~new_new_n18627__;
  assign new_new_n18803__ = new_new_n18643__ & new_new_n18802__;
  assign new_new_n18804__ = ~new_new_n18643__ & ~new_new_n18802__;
  assign new_new_n18805__ = ~new_new_n18803__ & ~new_new_n18804__;
  assign new_new_n18806__ = ~new_new_n18801__ & ~new_new_n18805__;
  assign new_new_n18807__ = new_new_n18801__ & new_new_n18805__;
  assign new_new_n18808__ = new_new_n3311__ & ~new_new_n15432__;
  assign new_new_n18809__ = new_new_n873__ & ~new_new_n15439__;
  assign new_new_n18810__ = ~new_new_n333__ & new_new_n15464__;
  assign new_new_n18811__ = ~new_new_n4900__ & new_new_n17204__;
  assign new_new_n18812__ = ~new_new_n18809__ & ~new_new_n18810__;
  assign new_new_n18813__ = ~new_new_n18808__ & new_new_n18812__;
  assign new_new_n18814__ = ~new_new_n18811__ & new_new_n18813__;
  assign new_new_n18815__ = pi26 & ~new_new_n18814__;
  assign new_new_n18816__ = ~pi26 & new_new_n18814__;
  assign new_new_n18817__ = ~new_new_n18815__ & ~new_new_n18816__;
  assign new_new_n18818__ = ~new_new_n18807__ & ~new_new_n18817__;
  assign new_new_n18819__ = ~new_new_n18806__ & ~new_new_n18818__;
  assign new_new_n18820__ = new_new_n18768__ & ~new_new_n18819__;
  assign new_new_n18821__ = ~new_new_n18768__ & new_new_n18819__;
  assign new_new_n18822__ = new_new_n5213__ & ~new_new_n15349__;
  assign new_new_n18823__ = new_new_n5183__ & ~new_new_n15398__;
  assign new_new_n18824__ = new_new_n5191__ & new_new_n15390__;
  assign new_new_n18825__ = new_new_n5215__ & ~new_new_n17180__;
  assign new_new_n18826__ = ~new_new_n18823__ & ~new_new_n18824__;
  assign new_new_n18827__ = ~new_new_n18822__ & new_new_n18826__;
  assign new_new_n18828__ = ~new_new_n18825__ & new_new_n18827__;
  assign new_new_n18829__ = pi23 & ~new_new_n18828__;
  assign new_new_n18830__ = ~pi23 & new_new_n18828__;
  assign new_new_n18831__ = ~new_new_n18829__ & ~new_new_n18830__;
  assign new_new_n18832__ = ~new_new_n18821__ & ~new_new_n18831__;
  assign new_new_n18833__ = ~new_new_n18820__ & ~new_new_n18832__;
  assign new_new_n18834__ = ~new_new_n18764__ & ~new_new_n18833__;
  assign new_new_n18835__ = ~new_new_n18763__ & ~new_new_n18834__;
  assign new_new_n18836__ = ~new_new_n18746__ & ~new_new_n18835__;
  assign new_new_n18837__ = new_new_n18746__ & new_new_n18835__;
  assign new_new_n18838__ = new_new_n6629__ & ~new_new_n15314__;
  assign new_new_n18839__ = new_new_n6634__ & ~new_new_n15248__;
  assign new_new_n18840__ = ~new_new_n6625__ & new_new_n15285__;
  assign new_new_n18841__ = new_new_n6936__ & new_new_n16725__;
  assign new_new_n18842__ = ~new_new_n18838__ & ~new_new_n18840__;
  assign new_new_n18843__ = ~new_new_n18839__ & new_new_n18842__;
  assign new_new_n18844__ = ~new_new_n18841__ & new_new_n18843__;
  assign new_new_n18845__ = ~pi20 & ~new_new_n18844__;
  assign new_new_n18846__ = pi20 & new_new_n18844__;
  assign new_new_n18847__ = ~new_new_n18845__ & ~new_new_n18846__;
  assign new_new_n18848__ = ~new_new_n18837__ & new_new_n18847__;
  assign new_new_n18849__ = ~new_new_n18836__ & ~new_new_n18848__;
  assign new_new_n18850__ = ~new_new_n18740__ & ~new_new_n18849__;
  assign new_new_n18851__ = new_new_n18740__ & new_new_n18849__;
  assign new_new_n18852__ = ~new_new_n18850__ & ~new_new_n18851__;
  assign new_new_n18853__ = ~new_new_n18377__ & ~new_new_n18378__;
  assign new_new_n18854__ = ~new_new_n18659__ & new_new_n18853__;
  assign new_new_n18855__ = new_new_n18659__ & ~new_new_n18853__;
  assign new_new_n18856__ = ~new_new_n18854__ & ~new_new_n18855__;
  assign new_new_n18857__ = new_new_n18852__ & ~new_new_n18856__;
  assign new_new_n18858__ = ~new_new_n18852__ & new_new_n18856__;
  assign new_new_n18859__ = ~new_new_n18857__ & ~new_new_n18858__;
  assign new_new_n18860__ = new_new_n18728__ & ~new_new_n18859__;
  assign new_new_n18861__ = ~new_new_n18728__ & new_new_n18859__;
  assign new_new_n18862__ = new_new_n6959__ & ~new_new_n15917__;
  assign new_new_n18863__ = new_new_n6964__ & new_new_n15244__;
  assign new_new_n18864__ = new_new_n6968__ & new_new_n15237__;
  assign new_new_n18865__ = ~new_new_n18863__ & ~new_new_n18864__;
  assign new_new_n18866__ = ~new_new_n18862__ & new_new_n18865__;
  assign new_new_n18867__ = new_new_n6958__ & new_new_n15905__;
  assign new_new_n18868__ = pi17 & ~new_new_n18867__;
  assign new_new_n18869__ = new_new_n8160__ & new_new_n15905__;
  assign new_new_n18870__ = ~new_new_n18868__ & ~new_new_n18869__;
  assign new_new_n18871__ = new_new_n18866__ & ~new_new_n18870__;
  assign new_new_n18872__ = ~pi17 & ~new_new_n18866__;
  assign new_new_n18873__ = ~new_new_n18871__ & ~new_new_n18872__;
  assign new_new_n18874__ = new_new_n6629__ & ~new_new_n15273__;
  assign new_new_n18875__ = ~new_new_n6625__ & ~new_new_n15321__;
  assign new_new_n18876__ = new_new_n6634__ & new_new_n15285__;
  assign new_new_n18877__ = ~new_new_n18874__ & ~new_new_n18875__;
  assign new_new_n18878__ = ~new_new_n18876__ & new_new_n18877__;
  assign new_new_n18879__ = new_new_n6631__ & new_new_n16078__;
  assign new_new_n18880__ = pi20 & ~new_new_n18879__;
  assign new_new_n18881__ = new_new_n6640__ & new_new_n16078__;
  assign new_new_n18882__ = ~new_new_n18880__ & ~new_new_n18881__;
  assign new_new_n18883__ = new_new_n18878__ & ~new_new_n18882__;
  assign new_new_n18884__ = ~pi20 & ~new_new_n18878__;
  assign new_new_n18885__ = ~new_new_n18883__ & ~new_new_n18884__;
  assign new_new_n18886__ = ~new_new_n18820__ & ~new_new_n18821__;
  assign new_new_n18887__ = ~new_new_n18831__ & new_new_n18886__;
  assign new_new_n18888__ = new_new_n18831__ & ~new_new_n18886__;
  assign new_new_n18889__ = ~new_new_n18887__ & ~new_new_n18888__;
  assign new_new_n18890__ = new_new_n18885__ & new_new_n18889__;
  assign new_new_n18891__ = ~new_new_n18885__ & ~new_new_n18889__;
  assign new_new_n18892__ = ~new_new_n18806__ & ~new_new_n18807__;
  assign new_new_n18893__ = ~new_new_n18817__ & new_new_n18892__;
  assign new_new_n18894__ = new_new_n18817__ & ~new_new_n18892__;
  assign new_new_n18895__ = ~new_new_n18893__ & ~new_new_n18894__;
  assign new_new_n18896__ = new_new_n3311__ & new_new_n15464__;
  assign new_new_n18897__ = ~new_new_n333__ & ~new_new_n15809__;
  assign new_new_n18898__ = new_new_n873__ & ~new_new_n15471__;
  assign new_new_n18899__ = ~new_new_n18897__ & ~new_new_n18898__;
  assign new_new_n18900__ = ~new_new_n18896__ & new_new_n18899__;
  assign new_new_n18901__ = pi26 & ~new_new_n18900__;
  assign new_new_n18902__ = new_new_n4898__ & new_new_n15819__;
  assign new_new_n18903__ = new_new_n801__ & new_new_n15819__;
  assign new_new_n18904__ = ~pi26 & ~new_new_n18903__;
  assign new_new_n18905__ = ~new_new_n18902__ & ~new_new_n18904__;
  assign new_new_n18906__ = new_new_n18900__ & ~new_new_n18905__;
  assign new_new_n18907__ = ~new_new_n18901__ & ~new_new_n18906__;
  assign new_new_n18908__ = ~new_new_n4818__ & ~new_new_n15533__;
  assign new_new_n18909__ = new_new_n4212__ & new_new_n15520__;
  assign new_new_n18910__ = ~new_new_n18908__ & ~new_new_n18909__;
  assign new_new_n18911__ = ~new_new_n15767__ & new_new_n18125__;
  assign new_new_n18912__ = ~new_new_n15777__ & ~new_new_n18124__;
  assign new_new_n18913__ = ~new_new_n18911__ & new_new_n18912__;
  assign new_new_n18914__ = ~new_new_n15524__ & ~new_new_n18913__;
  assign new_new_n18915__ = new_new_n4214__ & ~new_new_n18914__;
  assign new_new_n18916__ = pi29 & ~new_new_n18915__;
  assign new_new_n18917__ = pi28 & ~new_new_n15524__;
  assign new_new_n18918__ = ~new_new_n18776__ & ~new_new_n18917__;
  assign new_new_n18919__ = new_new_n4214__ & ~new_new_n18918__;
  assign new_new_n18920__ = new_new_n18913__ & new_new_n18919__;
  assign new_new_n18921__ = ~new_new_n18916__ & ~new_new_n18920__;
  assign new_new_n18922__ = new_new_n18910__ & ~new_new_n18921__;
  assign new_new_n18923__ = new_new_n15524__ & ~new_new_n18913__;
  assign new_new_n18924__ = new_new_n4214__ & new_new_n18923__;
  assign new_new_n18925__ = new_new_n18910__ & ~new_new_n18924__;
  assign new_new_n18926__ = ~pi29 & ~new_new_n18925__;
  assign new_new_n18927__ = ~new_new_n18922__ & ~new_new_n18926__;
  assign new_new_n18928__ = new_new_n765__ & new_new_n15560__;
  assign new_new_n18929__ = ~new_new_n18449__ & ~new_new_n18928__;
  assign new_new_n18930__ = ~pi31 & ~new_new_n18929__;
  assign new_new_n18931__ = ~new_new_n15615__ & ~new_new_n15755__;
  assign new_new_n18932__ = ~new_new_n15564__ & ~new_new_n18931__;
  assign new_new_n18933__ = new_new_n15572__ & ~new_new_n18932__;
  assign new_new_n18934__ = ~new_new_n15560__ & new_new_n18933__;
  assign new_new_n18935__ = new_new_n15615__ & new_new_n18507__;
  assign new_new_n18936__ = new_new_n15564__ & ~new_new_n18935__;
  assign new_new_n18937__ = ~new_new_n15572__ & ~new_new_n18936__;
  assign new_new_n18938__ = ~new_new_n15560__ & new_new_n18937__;
  assign new_new_n18939__ = ~new_new_n18934__ & ~new_new_n18938__;
  assign new_new_n18940__ = ~new_new_n15564__ & ~new_new_n15572__;
  assign new_new_n18941__ = ~new_new_n18933__ & ~new_new_n18935__;
  assign new_new_n18942__ = ~new_new_n18940__ & new_new_n18941__;
  assign new_new_n18943__ = new_new_n15560__ & new_new_n18942__;
  assign new_new_n18944__ = new_new_n18939__ & ~new_new_n18943__;
  assign new_new_n18945__ = new_new_n765__ & ~new_new_n18944__;
  assign new_new_n18946__ = new_new_n71__ & ~new_new_n15572__;
  assign new_new_n18947__ = new_new_n161__ & ~new_new_n15564__;
  assign new_new_n18948__ = pi31 & ~new_new_n18947__;
  assign new_new_n18949__ = ~new_new_n18946__ & new_new_n18948__;
  assign new_new_n18950__ = ~new_new_n18945__ & new_new_n18949__;
  assign new_new_n18951__ = ~new_new_n18930__ & ~new_new_n18950__;
  assign new_new_n18952__ = ~new_new_n18562__ & ~new_new_n18565__;
  assign new_new_n18953__ = new_new_n18518__ & ~new_new_n18535__;
  assign new_new_n18954__ = new_new_n18952__ & ~new_new_n18953__;
  assign new_new_n18955__ = ~new_new_n18499__ & new_new_n18954__;
  assign new_new_n18956__ = ~new_new_n18499__ & new_new_n18518__;
  assign new_new_n18957__ = ~new_new_n18566__ & ~new_new_n18956__;
  assign new_new_n18958__ = new_new_n18146__ & ~new_new_n18957__;
  assign new_new_n18959__ = new_new_n18499__ & ~new_new_n18562__;
  assign new_new_n18960__ = ~new_new_n18146__ & ~new_new_n18956__;
  assign new_new_n18961__ = ~new_new_n18959__ & new_new_n18960__;
  assign new_new_n18962__ = ~new_new_n18955__ & ~new_new_n18961__;
  assign new_new_n18963__ = ~new_new_n18958__ & new_new_n18962__;
  assign new_new_n18964__ = new_new_n4212__ & new_new_n15560__;
  assign new_new_n18965__ = ~new_new_n4215__ & new_new_n18454__;
  assign new_new_n18966__ = new_new_n4215__ & ~new_new_n15767__;
  assign new_new_n18967__ = new_new_n4214__ & ~new_new_n18966__;
  assign new_new_n18968__ = ~new_new_n18965__ & new_new_n18967__;
  assign new_new_n18969__ = ~new_new_n18964__ & ~new_new_n18968__;
  assign new_new_n18970__ = new_new_n67__ & new_new_n15572__;
  assign new_new_n18971__ = pi29 & ~new_new_n18970__;
  assign new_new_n18972__ = new_new_n65__ & new_new_n15572__;
  assign new_new_n18973__ = ~pi29 & ~new_new_n18972__;
  assign new_new_n18974__ = pi26 & ~new_new_n18973__;
  assign new_new_n18975__ = ~new_new_n18971__ & ~new_new_n18974__;
  assign new_new_n18976__ = new_new_n18969__ & ~new_new_n18975__;
  assign new_new_n18977__ = ~pi29 & ~new_new_n18969__;
  assign new_new_n18978__ = ~new_new_n18976__ & ~new_new_n18977__;
  assign new_new_n18979__ = new_new_n18146__ & ~new_new_n18952__;
  assign new_new_n18980__ = ~new_new_n18146__ & new_new_n18954__;
  assign new_new_n18981__ = ~new_new_n18979__ & ~new_new_n18980__;
  assign new_new_n18982__ = ~new_new_n18978__ & ~new_new_n18981__;
  assign new_new_n18983__ = new_new_n18978__ & new_new_n18981__;
  assign new_new_n18984__ = new_new_n765__ & ~new_new_n15615__;
  assign new_new_n18985__ = ~new_new_n18515__ & ~new_new_n18984__;
  assign new_new_n18986__ = ~pi31 & ~new_new_n18985__;
  assign new_new_n18987__ = new_new_n15615__ & ~new_new_n15743__;
  assign new_new_n18988__ = new_new_n15582__ & new_new_n18987__;
  assign new_new_n18989__ = new_new_n15638__ & new_new_n15743__;
  assign new_new_n18990__ = ~new_new_n15615__ & new_new_n18989__;
  assign new_new_n18991__ = ~new_new_n15736__ & new_new_n18990__;
  assign new_new_n18992__ = ~new_new_n18988__ & ~new_new_n18991__;
  assign new_new_n18993__ = new_new_n15647__ & ~new_new_n18992__;
  assign new_new_n18994__ = ~new_new_n15736__ & new_new_n18987__;
  assign new_new_n18995__ = ~new_new_n18990__ & ~new_new_n18994__;
  assign new_new_n18996__ = new_new_n15582__ & ~new_new_n18995__;
  assign new_new_n18997__ = ~new_new_n15615__ & new_new_n15743__;
  assign new_new_n18998__ = ~new_new_n15638__ & ~new_new_n15743__;
  assign new_new_n18999__ = ~new_new_n18989__ & ~new_new_n18998__;
  assign new_new_n19000__ = new_new_n15615__ & new_new_n18999__;
  assign new_new_n19001__ = ~new_new_n15746__ & ~new_new_n19000__;
  assign new_new_n19002__ = ~new_new_n15751__ & new_new_n19001__;
  assign new_new_n19003__ = ~new_new_n18997__ & ~new_new_n19002__;
  assign new_new_n19004__ = ~new_new_n18993__ & ~new_new_n18996__;
  assign new_new_n19005__ = ~new_new_n19003__ & new_new_n19004__;
  assign new_new_n19006__ = new_new_n765__ & ~new_new_n19005__;
  assign new_new_n19007__ = new_new_n71__ & ~new_new_n15743__;
  assign new_new_n19008__ = new_new_n161__ & new_new_n15638__;
  assign new_new_n19009__ = pi31 & ~new_new_n19008__;
  assign new_new_n19010__ = ~new_new_n19007__ & new_new_n19009__;
  assign new_new_n19011__ = ~new_new_n19006__ & new_new_n19010__;
  assign new_new_n19012__ = ~new_new_n18986__ & ~new_new_n19011__;
  assign new_new_n19013__ = ~new_new_n313__ & ~new_new_n1167__;
  assign new_new_n19014__ = ~new_new_n235__ & ~new_new_n783__;
  assign new_new_n19015__ = new_new_n1036__ & new_new_n19014__;
  assign new_new_n19016__ = new_new_n2026__ & new_new_n19015__;
  assign new_new_n19017__ = ~new_new_n119__ & ~new_new_n168__;
  assign new_new_n19018__ = ~new_new_n302__ & new_new_n7131__;
  assign new_new_n19019__ = new_new_n210__ & new_new_n19017__;
  assign new_new_n19020__ = ~new_new_n232__ & new_new_n1154__;
  assign new_new_n19021__ = ~new_new_n2697__ & new_new_n3058__;
  assign new_new_n19022__ = new_new_n19020__ & new_new_n19021__;
  assign new_new_n19023__ = new_new_n19018__ & new_new_n19019__;
  assign new_new_n19024__ = ~new_new_n124__ & new_new_n830__;
  assign new_new_n19025__ = new_new_n1065__ & new_new_n19013__;
  assign new_new_n19026__ = new_new_n19024__ & new_new_n19025__;
  assign new_new_n19027__ = new_new_n19022__ & new_new_n19023__;
  assign new_new_n19028__ = new_new_n3585__ & new_new_n19027__;
  assign new_new_n19029__ = new_new_n17390__ & new_new_n19026__;
  assign new_new_n19030__ = new_new_n19016__ & new_new_n19029__;
  assign new_new_n19031__ = new_new_n2767__ & new_new_n19028__;
  assign new_new_n19032__ = new_new_n19030__ & new_new_n19031__;
  assign new_new_n19033__ = new_new_n1538__ & new_new_n19032__;
  assign new_new_n19034__ = new_new_n5608__ & new_new_n19033__;
  assign new_new_n19035__ = ~new_new_n19012__ & ~new_new_n19034__;
  assign new_new_n19036__ = ~new_new_n242__ & ~new_new_n473__;
  assign new_new_n19037__ = ~new_new_n657__ & ~new_new_n768__;
  assign new_new_n19038__ = new_new_n19036__ & new_new_n19037__;
  assign new_new_n19039__ = ~new_new_n483__ & ~new_new_n1632__;
  assign new_new_n19040__ = new_new_n5378__ & new_new_n16487__;
  assign new_new_n19041__ = new_new_n19039__ & new_new_n19040__;
  assign new_new_n19042__ = new_new_n2003__ & new_new_n19038__;
  assign new_new_n19043__ = new_new_n2769__ & new_new_n19042__;
  assign new_new_n19044__ = new_new_n810__ & new_new_n19041__;
  assign new_new_n19045__ = new_new_n3982__ & new_new_n19044__;
  assign new_new_n19046__ = new_new_n16160__ & new_new_n19043__;
  assign new_new_n19047__ = new_new_n19045__ & new_new_n19046__;
  assign new_new_n19048__ = new_new_n3150__ & new_new_n19047__;
  assign new_new_n19049__ = new_new_n2402__ & new_new_n19048__;
  assign new_new_n19050__ = new_new_n18541__ & new_new_n19049__;
  assign new_new_n19051__ = new_new_n15647__ & ~new_new_n15736__;
  assign new_new_n19052__ = new_new_n15582__ & new_new_n15736__;
  assign new_new_n19053__ = ~new_new_n15853__ & ~new_new_n19051__;
  assign new_new_n19054__ = ~new_new_n19052__ & new_new_n19053__;
  assign new_new_n19055__ = ~new_new_n15711__ & ~new_new_n19054__;
  assign new_new_n19056__ = new_new_n15638__ & ~new_new_n19055__;
  assign new_new_n19057__ = ~new_new_n71__ & new_new_n15647__;
  assign new_new_n19058__ = ~new_new_n15582__ & ~new_new_n15736__;
  assign new_new_n19059__ = ~new_new_n15638__ & new_new_n19058__;
  assign new_new_n19060__ = ~new_new_n161__ & ~new_new_n19059__;
  assign new_new_n19061__ = new_new_n19057__ & ~new_new_n19060__;
  assign new_new_n19062__ = ~new_new_n71__ & ~new_new_n15748__;
  assign new_new_n19063__ = ~new_new_n161__ & ~new_new_n19057__;
  assign new_new_n19064__ = new_new_n15582__ & new_new_n19063__;
  assign new_new_n19065__ = ~new_new_n19062__ & new_new_n19064__;
  assign new_new_n19066__ = ~new_new_n19061__ & ~new_new_n19065__;
  assign new_new_n19067__ = ~new_new_n19056__ & new_new_n19066__;
  assign new_new_n19068__ = pi31 & ~new_new_n19067__;
  assign new_new_n19069__ = new_new_n161__ & ~new_new_n15582__;
  assign new_new_n19070__ = new_new_n765__ & ~new_new_n15638__;
  assign new_new_n19071__ = ~pi31 & ~new_new_n19069__;
  assign new_new_n19072__ = ~new_new_n19070__ & new_new_n19071__;
  assign new_new_n19073__ = ~new_new_n19068__ & ~new_new_n19072__;
  assign new_new_n19074__ = new_new_n19050__ & ~new_new_n19073__;
  assign new_new_n19075__ = ~new_new_n19050__ & new_new_n19073__;
  assign new_new_n19076__ = new_new_n161__ & ~new_new_n15647__;
  assign new_new_n19077__ = new_new_n765__ & ~new_new_n15582__;
  assign new_new_n19078__ = ~new_new_n19076__ & ~new_new_n19077__;
  assign new_new_n19079__ = ~pi31 & ~new_new_n19078__;
  assign new_new_n19080__ = new_new_n765__ & new_new_n15736__;
  assign new_new_n19081__ = new_new_n161__ & new_new_n15710__;
  assign new_new_n19082__ = new_new_n71__ & new_new_n15647__;
  assign new_new_n19083__ = pi31 & ~new_new_n19081__;
  assign new_new_n19084__ = ~new_new_n19082__ & new_new_n19083__;
  assign new_new_n19085__ = ~new_new_n19080__ & new_new_n19084__;
  assign new_new_n19086__ = ~new_new_n19079__ & ~new_new_n19085__;
  assign new_new_n19087__ = new_new_n161__ & ~new_new_n15710__;
  assign new_new_n19088__ = new_new_n765__ & ~new_new_n15647__;
  assign new_new_n19089__ = ~new_new_n19087__ & ~new_new_n19088__;
  assign new_new_n19090__ = ~pi31 & ~new_new_n19089__;
  assign new_new_n19091__ = new_new_n71__ & ~new_new_n15710__;
  assign new_new_n19092__ = new_new_n161__ & new_new_n15656__;
  assign new_new_n19093__ = new_new_n15656__ & ~new_new_n15710__;
  assign new_new_n19094__ = ~new_new_n15656__ & new_new_n15710__;
  assign new_new_n19095__ = ~new_new_n19093__ & ~new_new_n19094__;
  assign new_new_n19096__ = ~new_new_n15647__ & ~new_new_n19095__;
  assign new_new_n19097__ = new_new_n15643__ & new_new_n15722__;
  assign new_new_n19098__ = new_new_n15656__ & new_new_n15723__;
  assign new_new_n19099__ = new_new_n15680__ & new_new_n19098__;
  assign new_new_n19100__ = ~new_new_n19097__ & ~new_new_n19099__;
  assign new_new_n19101__ = ~new_new_n15661__ & ~new_new_n19100__;
  assign new_new_n19102__ = ~new_new_n15647__ & new_new_n15710__;
  assign new_new_n19103__ = ~new_new_n15643__ & new_new_n19102__;
  assign new_new_n19104__ = ~new_new_n15656__ & ~new_new_n15710__;
  assign new_new_n19105__ = new_new_n15647__ & new_new_n19104__;
  assign new_new_n19106__ = ~new_new_n15680__ & new_new_n19105__;
  assign new_new_n19107__ = ~new_new_n19103__ & ~new_new_n19106__;
  assign new_new_n19108__ = new_new_n15661__ & ~new_new_n19107__;
  assign new_new_n19109__ = ~new_new_n15680__ & new_new_n19102__;
  assign new_new_n19110__ = ~new_new_n19105__ & ~new_new_n19109__;
  assign new_new_n19111__ = ~new_new_n15643__ & ~new_new_n19110__;
  assign new_new_n19112__ = new_new_n15680__ & new_new_n15722__;
  assign new_new_n19113__ = ~new_new_n19098__ & ~new_new_n19112__;
  assign new_new_n19114__ = new_new_n15643__ & ~new_new_n19113__;
  assign new_new_n19115__ = ~new_new_n19111__ & ~new_new_n19114__;
  assign new_new_n19116__ = ~new_new_n19101__ & new_new_n19115__;
  assign new_new_n19117__ = ~new_new_n19108__ & new_new_n19116__;
  assign new_new_n19118__ = ~new_new_n19096__ & new_new_n19117__;
  assign new_new_n19119__ = new_new_n765__ & ~new_new_n19118__;
  assign new_new_n19120__ = ~new_new_n19091__ & ~new_new_n19092__;
  assign new_new_n19121__ = ~new_new_n19119__ & new_new_n19120__;
  assign new_new_n19122__ = pi31 & ~new_new_n19121__;
  assign new_new_n19123__ = ~new_new_n19090__ & ~new_new_n19122__;
  assign new_new_n19124__ = ~new_new_n140__ & ~new_new_n3746__;
  assign new_new_n19125__ = new_new_n225__ & new_new_n19124__;
  assign new_new_n19126__ = ~new_new_n379__ & ~new_new_n586__;
  assign new_new_n19127__ = ~new_new_n671__ & ~new_new_n723__;
  assign new_new_n19128__ = new_new_n19126__ & new_new_n19127__;
  assign new_new_n19129__ = ~new_new_n696__ & ~new_new_n732__;
  assign new_new_n19130__ = ~new_new_n871__ & ~new_new_n1166__;
  assign new_new_n19131__ = new_new_n1709__ & new_new_n2698__;
  assign new_new_n19132__ = new_new_n3179__ & new_new_n4414__;
  assign new_new_n19133__ = ~new_new_n19125__ & new_new_n19132__;
  assign new_new_n19134__ = new_new_n19130__ & new_new_n19131__;
  assign new_new_n19135__ = new_new_n19128__ & new_new_n19129__;
  assign new_new_n19136__ = ~new_new_n316__ & new_new_n19135__;
  assign new_new_n19137__ = new_new_n19133__ & new_new_n19134__;
  assign new_new_n19138__ = new_new_n562__ & ~new_new_n895__;
  assign new_new_n19139__ = new_new_n985__ & new_new_n7630__;
  assign new_new_n19140__ = new_new_n19138__ & new_new_n19139__;
  assign new_new_n19141__ = new_new_n19136__ & new_new_n19137__;
  assign new_new_n19142__ = new_new_n19140__ & new_new_n19141__;
  assign new_new_n19143__ = ~new_new_n300__ & ~new_new_n935__;
  assign new_new_n19144__ = ~new_new_n119__ & ~new_new_n336__;
  assign new_new_n19145__ = ~new_new_n482__ & ~new_new_n995__;
  assign new_new_n19146__ = new_new_n19144__ & new_new_n19145__;
  assign new_new_n19147__ = new_new_n2575__ & new_new_n3967__;
  assign new_new_n19148__ = new_new_n19146__ & new_new_n19147__;
  assign new_new_n19149__ = ~new_new_n344__ & ~new_new_n630__;
  assign new_new_n19150__ = new_new_n1283__ & new_new_n1806__;
  assign new_new_n19151__ = new_new_n4391__ & new_new_n5566__;
  assign new_new_n19152__ = new_new_n19150__ & new_new_n19151__;
  assign new_new_n19153__ = new_new_n19148__ & new_new_n19149__;
  assign new_new_n19154__ = new_new_n19143__ & new_new_n19153__;
  assign new_new_n19155__ = new_new_n4321__ & new_new_n19152__;
  assign new_new_n19156__ = new_new_n19154__ & new_new_n19155__;
  assign new_new_n19157__ = new_new_n7500__ & new_new_n19156__;
  assign new_new_n19158__ = ~new_new_n384__ & ~new_new_n388__;
  assign new_new_n19159__ = ~new_new_n511__ & ~new_new_n1070__;
  assign new_new_n19160__ = new_new_n19158__ & new_new_n19159__;
  assign new_new_n19161__ = ~new_new_n348__ & new_new_n1741__;
  assign new_new_n19162__ = new_new_n19160__ & new_new_n19161__;
  assign new_new_n19163__ = new_new_n743__ & new_new_n944__;
  assign new_new_n19164__ = new_new_n2159__ & new_new_n2501__;
  assign new_new_n19165__ = new_new_n4229__ & new_new_n19164__;
  assign new_new_n19166__ = new_new_n19162__ & new_new_n19163__;
  assign new_new_n19167__ = new_new_n1400__ & new_new_n2478__;
  assign new_new_n19168__ = new_new_n3019__ & new_new_n3024__;
  assign new_new_n19169__ = new_new_n7727__ & new_new_n19168__;
  assign new_new_n19170__ = new_new_n19166__ & new_new_n19167__;
  assign new_new_n19171__ = new_new_n669__ & new_new_n19165__;
  assign new_new_n19172__ = new_new_n19170__ & new_new_n19171__;
  assign new_new_n19173__ = new_new_n19169__ & new_new_n19172__;
  assign new_new_n19174__ = new_new_n17255__ & new_new_n19142__;
  assign new_new_n19175__ = new_new_n19173__ & new_new_n19174__;
  assign new_new_n19176__ = new_new_n19157__ & new_new_n19175__;
  assign new_new_n19177__ = ~new_new_n19123__ & ~new_new_n19176__;
  assign new_new_n19178__ = new_new_n19123__ & new_new_n19176__;
  assign new_new_n19179__ = new_new_n15678__ & new_new_n15710__;
  assign new_new_n19180__ = ~new_new_n161__ & ~new_new_n19093__;
  assign new_new_n19181__ = ~new_new_n19179__ & new_new_n19180__;
  assign new_new_n19182__ = new_new_n15643__ & ~new_new_n19181__;
  assign new_new_n19183__ = ~new_new_n15643__ & new_new_n15656__;
  assign new_new_n19184__ = new_new_n15710__ & new_new_n19183__;
  assign new_new_n19185__ = ~new_new_n19104__ & ~new_new_n19184__;
  assign new_new_n19186__ = new_new_n15687__ & ~new_new_n19185__;
  assign new_new_n19187__ = ~new_new_n15643__ & ~new_new_n15687__;
  assign new_new_n19188__ = ~new_new_n15710__ & new_new_n19187__;
  assign new_new_n19189__ = ~new_new_n19186__ & ~new_new_n19188__;
  assign new_new_n19190__ = ~new_new_n161__ & ~new_new_n19189__;
  assign new_new_n19191__ = new_new_n4147__ & ~new_new_n19182__;
  assign new_new_n19192__ = ~new_new_n19190__ & new_new_n19191__;
  assign new_new_n19193__ = ~new_new_n71__ & new_new_n19092__;
  assign new_new_n19194__ = new_new_n71__ & ~new_new_n15656__;
  assign new_new_n19195__ = pi31 & ~new_new_n19194__;
  assign new_new_n19196__ = ~new_new_n15710__ & ~new_new_n15853__;
  assign new_new_n19197__ = ~new_new_n19193__ & ~new_new_n19195__;
  assign new_new_n19198__ = ~new_new_n19196__ & new_new_n19197__;
  assign new_new_n19199__ = ~new_new_n19192__ & ~new_new_n19198__;
  assign new_new_n19200__ = ~new_new_n15643__ & new_new_n15673__;
  assign new_new_n19201__ = ~new_new_n15675__ & ~new_new_n19200__;
  assign new_new_n19202__ = ~new_new_n161__ & ~new_new_n19201__;
  assign new_new_n19203__ = ~new_new_n15643__ & ~new_new_n15668__;
  assign new_new_n19204__ = ~new_new_n71__ & ~new_new_n19203__;
  assign new_new_n19205__ = ~new_new_n19202__ & new_new_n19204__;
  assign new_new_n19206__ = new_new_n15661__ & ~new_new_n19205__;
  assign new_new_n19207__ = new_new_n161__ & ~new_new_n15668__;
  assign new_new_n19208__ = ~new_new_n161__ & ~new_new_n15643__;
  assign new_new_n19209__ = new_new_n15668__ & ~new_new_n19208__;
  assign new_new_n19210__ = ~new_new_n15661__ & new_new_n19204__;
  assign new_new_n19211__ = ~new_new_n19209__ & new_new_n19210__;
  assign new_new_n19212__ = pi31 & ~new_new_n19207__;
  assign new_new_n19213__ = ~new_new_n19211__ & new_new_n19212__;
  assign new_new_n19214__ = ~new_new_n19206__ & new_new_n19213__;
  assign new_new_n19215__ = new_new_n161__ & ~new_new_n15661__;
  assign new_new_n19216__ = new_new_n765__ & new_new_n15643__;
  assign new_new_n19217__ = ~new_new_n19215__ & ~new_new_n19216__;
  assign new_new_n19218__ = ~pi31 & ~new_new_n19217__;
  assign new_new_n19219__ = ~new_new_n19214__ & ~new_new_n19218__;
  assign new_new_n19220__ = ~new_new_n98__ & new_new_n110__;
  assign new_new_n19221__ = new_new_n95__ & ~new_new_n4898__;
  assign new_new_n19222__ = ~new_new_n19220__ & new_new_n19221__;
  assign new_new_n19223__ = ~new_new_n260__ & ~new_new_n783__;
  assign new_new_n19224__ = ~new_new_n382__ & new_new_n19223__;
  assign new_new_n19225__ = new_new_n3194__ & new_new_n19224__;
  assign new_new_n19226__ = new_new_n3420__ & new_new_n4365__;
  assign new_new_n19227__ = ~new_new_n19222__ & new_new_n19226__;
  assign new_new_n19228__ = new_new_n2641__ & new_new_n19225__;
  assign new_new_n19229__ = new_new_n7421__ & new_new_n16235__;
  assign new_new_n19230__ = new_new_n19228__ & new_new_n19229__;
  assign new_new_n19231__ = new_new_n3171__ & new_new_n19227__;
  assign new_new_n19232__ = new_new_n19230__ & new_new_n19231__;
  assign new_new_n19233__ = new_new_n3785__ & new_new_n6148__;
  assign new_new_n19234__ = new_new_n19232__ & new_new_n19233__;
  assign new_new_n19235__ = new_new_n4089__ & new_new_n19234__;
  assign new_new_n19236__ = new_new_n4364__ & new_new_n19235__;
  assign new_new_n19237__ = ~new_new_n19219__ & ~new_new_n19236__;
  assign new_new_n19238__ = new_new_n19219__ & new_new_n19236__;
  assign new_new_n19239__ = new_new_n765__ & new_new_n15669__;
  assign new_new_n19240__ = ~new_new_n161__ & new_new_n15661__;
  assign new_new_n19241__ = new_new_n15673__ & ~new_new_n19240__;
  assign new_new_n19242__ = ~new_new_n15682__ & ~new_new_n19241__;
  assign new_new_n19243__ = ~new_new_n71__ & ~new_new_n19242__;
  assign new_new_n19244__ = pi31 & ~new_new_n19243__;
  assign new_new_n19245__ = new_new_n4876__ & ~new_new_n19240__;
  assign new_new_n19246__ = ~new_new_n19244__ & ~new_new_n19245__;
  assign new_new_n19247__ = new_new_n15668__ & ~new_new_n19246__;
  assign new_new_n19248__ = new_new_n5059__ & ~new_new_n15673__;
  assign new_new_n19249__ = ~new_new_n19239__ & ~new_new_n19248__;
  assign new_new_n19250__ = ~new_new_n19247__ & new_new_n19249__;
  assign new_new_n19251__ = ~new_new_n238__ & ~new_new_n308__;
  assign new_new_n19252__ = ~new_new_n701__ & new_new_n19251__;
  assign new_new_n19253__ = ~new_new_n945__ & ~new_new_n1073__;
  assign new_new_n19254__ = new_new_n1154__ & new_new_n1558__;
  assign new_new_n19255__ = new_new_n19253__ & new_new_n19254__;
  assign new_new_n19256__ = new_new_n542__ & new_new_n19252__;
  assign new_new_n19257__ = new_new_n1919__ & new_new_n2549__;
  assign new_new_n19258__ = new_new_n3294__ & new_new_n19257__;
  assign new_new_n19259__ = new_new_n4712__ & new_new_n19256__;
  assign new_new_n19260__ = new_new_n3100__ & new_new_n19255__;
  assign new_new_n19261__ = new_new_n3791__ & new_new_n4504__;
  assign new_new_n19262__ = new_new_n19260__ & new_new_n19261__;
  assign new_new_n19263__ = new_new_n19258__ & new_new_n19259__;
  assign new_new_n19264__ = new_new_n18548__ & new_new_n19263__;
  assign new_new_n19265__ = new_new_n19262__ & new_new_n19264__;
  assign new_new_n19266__ = new_new_n16318__ & new_new_n19265__;
  assign new_new_n19267__ = new_new_n17617__ & new_new_n19266__;
  assign new_new_n19268__ = ~new_new_n19250__ & ~new_new_n19267__;
  assign new_new_n19269__ = new_new_n19250__ & new_new_n19267__;
  assign new_new_n19270__ = ~new_new_n267__ & ~new_new_n768__;
  assign new_new_n19271__ = ~new_new_n472__ & ~new_new_n476__;
  assign new_new_n19272__ = ~new_new_n692__ & new_new_n19271__;
  assign new_new_n19273__ = ~new_new_n1507__ & new_new_n1711__;
  assign new_new_n19274__ = new_new_n19272__ & new_new_n19273__;
  assign new_new_n19275__ = new_new_n743__ & new_new_n19274__;
  assign new_new_n19276__ = ~new_new_n327__ & ~new_new_n637__;
  assign new_new_n19277__ = new_new_n2822__ & new_new_n19276__;
  assign new_new_n19278__ = new_new_n5397__ & new_new_n19277__;
  assign new_new_n19279__ = new_new_n16148__ & new_new_n19278__;
  assign new_new_n19280__ = new_new_n2547__ & new_new_n19279__;
  assign new_new_n19281__ = ~new_new_n384__ & ~new_new_n937__;
  assign new_new_n19282__ = ~new_new_n232__ & new_new_n19281__;
  assign new_new_n19283__ = ~new_new_n606__ & new_new_n702__;
  assign new_new_n19284__ = new_new_n19270__ & new_new_n19283__;
  assign new_new_n19285__ = ~new_new_n519__ & new_new_n19282__;
  assign new_new_n19286__ = new_new_n1645__ & new_new_n19285__;
  assign new_new_n19287__ = new_new_n627__ & new_new_n19284__;
  assign new_new_n19288__ = new_new_n3933__ & new_new_n16265__;
  assign new_new_n19289__ = new_new_n19287__ & new_new_n19288__;
  assign new_new_n19290__ = new_new_n19275__ & new_new_n19286__;
  assign new_new_n19291__ = new_new_n19289__ & new_new_n19290__;
  assign new_new_n19292__ = new_new_n19280__ & new_new_n19291__;
  assign new_new_n19293__ = ~new_new_n108__ & ~new_new_n238__;
  assign new_new_n19294__ = ~new_new_n950__ & ~new_new_n1176__;
  assign new_new_n19295__ = new_new_n19293__ & new_new_n19294__;
  assign new_new_n19296__ = ~new_new_n781__ & new_new_n1571__;
  assign new_new_n19297__ = new_new_n2079__ & new_new_n19296__;
  assign new_new_n19298__ = ~new_new_n373__ & new_new_n19295__;
  assign new_new_n19299__ = new_new_n953__ & new_new_n19298__;
  assign new_new_n19300__ = new_new_n216__ & new_new_n19297__;
  assign new_new_n19301__ = new_new_n440__ & new_new_n1400__;
  assign new_new_n19302__ = new_new_n19300__ & new_new_n19301__;
  assign new_new_n19303__ = new_new_n2657__ & new_new_n19299__;
  assign new_new_n19304__ = new_new_n2678__ & new_new_n19303__;
  assign new_new_n19305__ = new_new_n7534__ & new_new_n19302__;
  assign new_new_n19306__ = new_new_n19304__ & new_new_n19305__;
  assign new_new_n19307__ = new_new_n19292__ & new_new_n19306__;
  assign new_new_n19308__ = new_new_n2941__ & new_new_n19307__;
  assign new_new_n19309__ = new_new_n8646__ & ~new_new_n15673__;
  assign new_new_n19310__ = new_new_n15668__ & ~new_new_n15853__;
  assign new_new_n19311__ = new_new_n19309__ & new_new_n19310__;
  assign new_new_n19312__ = ~new_new_n19309__ & ~new_new_n19310__;
  assign new_new_n19313__ = ~new_new_n19308__ & ~new_new_n19311__;
  assign new_new_n19314__ = ~new_new_n19312__ & new_new_n19313__;
  assign new_new_n19315__ = ~new_new_n19269__ & new_new_n19314__;
  assign new_new_n19316__ = ~new_new_n19268__ & ~new_new_n19315__;
  assign new_new_n19317__ = ~new_new_n19238__ & ~new_new_n19316__;
  assign new_new_n19318__ = ~new_new_n19237__ & ~new_new_n19317__;
  assign new_new_n19319__ = ~new_new_n249__ & ~new_new_n383__;
  assign new_new_n19320__ = ~new_new_n258__ & new_new_n19319__;
  assign new_new_n19321__ = new_new_n3639__ & new_new_n19320__;
  assign new_new_n19322__ = new_new_n4390__ & new_new_n19321__;
  assign new_new_n19323__ = ~new_new_n652__ & new_new_n19322__;
  assign new_new_n19324__ = new_new_n91__ & ~new_new_n7416__;
  assign new_new_n19325__ = ~new_new_n1162__ & new_new_n16817__;
  assign new_new_n19326__ = ~new_new_n19324__ & new_new_n19325__;
  assign new_new_n19327__ = ~new_new_n106__ & ~new_new_n222__;
  assign new_new_n19328__ = ~new_new_n302__ & ~new_new_n335__;
  assign new_new_n19329__ = new_new_n19327__ & new_new_n19328__;
  assign new_new_n19330__ = new_new_n131__ & ~new_new_n155__;
  assign new_new_n19331__ = ~new_new_n280__ & ~new_new_n606__;
  assign new_new_n19332__ = ~new_new_n894__ & ~new_new_n1035__;
  assign new_new_n19333__ = new_new_n4595__ & new_new_n19332__;
  assign new_new_n19334__ = new_new_n19330__ & new_new_n19331__;
  assign new_new_n19335__ = new_new_n2911__ & new_new_n19329__;
  assign new_new_n19336__ = new_new_n19334__ & new_new_n19335__;
  assign new_new_n19337__ = new_new_n19326__ & new_new_n19333__;
  assign new_new_n19338__ = new_new_n19336__ & new_new_n19337__;
  assign new_new_n19339__ = new_new_n17626__ & new_new_n19338__;
  assign new_new_n19340__ = new_new_n19323__ & new_new_n19339__;
  assign new_new_n19341__ = ~new_new_n242__ & ~new_new_n282__;
  assign new_new_n19342__ = ~new_new_n480__ & new_new_n19341__;
  assign new_new_n19343__ = ~new_new_n696__ & new_new_n19342__;
  assign new_new_n19344__ = new_new_n543__ & new_new_n1428__;
  assign new_new_n19345__ = new_new_n1677__ & new_new_n3280__;
  assign new_new_n19346__ = new_new_n5698__ & new_new_n19345__;
  assign new_new_n19347__ = new_new_n19343__ & new_new_n19344__;
  assign new_new_n19348__ = new_new_n6256__ & new_new_n19347__;
  assign new_new_n19349__ = new_new_n1222__ & new_new_n19346__;
  assign new_new_n19350__ = new_new_n5612__ & new_new_n19349__;
  assign new_new_n19351__ = new_new_n3429__ & new_new_n19348__;
  assign new_new_n19352__ = new_new_n19350__ & new_new_n19351__;
  assign new_new_n19353__ = new_new_n1992__ & new_new_n19352__;
  assign new_new_n19354__ = new_new_n19340__ & new_new_n19353__;
  assign new_new_n19355__ = new_new_n19318__ & new_new_n19354__;
  assign new_new_n19356__ = ~new_new_n19318__ & ~new_new_n19354__;
  assign new_new_n19357__ = ~new_new_n19355__ & ~new_new_n19356__;
  assign new_new_n19358__ = new_new_n161__ & new_new_n15643__;
  assign new_new_n19359__ = new_new_n765__ & new_new_n15656__;
  assign new_new_n19360__ = ~new_new_n19358__ & ~new_new_n19359__;
  assign new_new_n19361__ = ~pi31 & ~new_new_n19360__;
  assign new_new_n19362__ = new_new_n71__ & ~new_new_n15643__;
  assign new_new_n19363__ = ~new_new_n15656__ & ~new_new_n15680__;
  assign new_new_n19364__ = new_new_n15656__ & ~new_new_n15681__;
  assign new_new_n19365__ = ~new_new_n19363__ & ~new_new_n19364__;
  assign new_new_n19366__ = new_new_n19240__ & ~new_new_n19365__;
  assign new_new_n19367__ = new_new_n15680__ & new_new_n19183__;
  assign new_new_n19368__ = new_new_n15643__ & ~new_new_n15656__;
  assign new_new_n19369__ = ~new_new_n15661__ & ~new_new_n19368__;
  assign new_new_n19370__ = ~new_new_n19367__ & new_new_n19369__;
  assign new_new_n19371__ = ~new_new_n19366__ & ~new_new_n19370__;
  assign new_new_n19372__ = ~new_new_n15643__ & new_new_n19363__;
  assign new_new_n19373__ = ~new_new_n19371__ & ~new_new_n19372__;
  assign new_new_n19374__ = ~new_new_n71__ & ~new_new_n19215__;
  assign new_new_n19375__ = ~new_new_n19373__ & new_new_n19374__;
  assign new_new_n19376__ = pi31 & ~new_new_n19362__;
  assign new_new_n19377__ = ~new_new_n19375__ & new_new_n19376__;
  assign new_new_n19378__ = ~new_new_n19361__ & ~new_new_n19377__;
  assign new_new_n19379__ = new_new_n19357__ & new_new_n19378__;
  assign new_new_n19380__ = ~new_new_n19355__ & ~new_new_n19379__;
  assign new_new_n19381__ = new_new_n19199__ & new_new_n19380__;
  assign new_new_n19382__ = ~new_new_n19199__ & ~new_new_n19380__;
  assign new_new_n19383__ = new_new_n628__ & ~new_new_n1064__;
  assign new_new_n19384__ = ~new_new_n252__ & ~new_new_n656__;
  assign new_new_n19385__ = ~new_new_n586__ & ~new_new_n729__;
  assign new_new_n19386__ = ~new_new_n829__ & ~new_new_n846__;
  assign new_new_n19387__ = new_new_n19385__ & new_new_n19386__;
  assign new_new_n19388__ = new_new_n2868__ & new_new_n4730__;
  assign new_new_n19389__ = new_new_n19384__ & new_new_n19388__;
  assign new_new_n19390__ = new_new_n167__ & new_new_n19387__;
  assign new_new_n19391__ = new_new_n844__ & new_new_n1037__;
  assign new_new_n19392__ = new_new_n1840__ & new_new_n2453__;
  assign new_new_n19393__ = new_new_n2508__ & new_new_n19392__;
  assign new_new_n19394__ = new_new_n19390__ & new_new_n19391__;
  assign new_new_n19395__ = new_new_n3700__ & new_new_n19389__;
  assign new_new_n19396__ = new_new_n19394__ & new_new_n19395__;
  assign new_new_n19397__ = new_new_n19393__ & new_new_n19396__;
  assign new_new_n19398__ = new_new_n3496__ & new_new_n17499__;
  assign new_new_n19399__ = new_new_n19397__ & new_new_n19398__;
  assign new_new_n19400__ = ~new_new_n130__ & ~new_new_n351__;
  assign new_new_n19401__ = ~new_new_n724__ & ~new_new_n768__;
  assign new_new_n19402__ = new_new_n4261__ & new_new_n19401__;
  assign new_new_n19403__ = ~new_new_n270__ & new_new_n19400__;
  assign new_new_n19404__ = ~new_new_n427__ & new_new_n1424__;
  assign new_new_n19405__ = new_new_n1713__ & new_new_n2078__;
  assign new_new_n19406__ = new_new_n19404__ & new_new_n19405__;
  assign new_new_n19407__ = new_new_n19402__ & new_new_n19403__;
  assign new_new_n19408__ = new_new_n144__ & ~new_new_n344__;
  assign new_new_n19409__ = new_new_n1703__ & new_new_n2467__;
  assign new_new_n19410__ = new_new_n2894__ & new_new_n19409__;
  assign new_new_n19411__ = new_new_n19407__ & new_new_n19408__;
  assign new_new_n19412__ = new_new_n2271__ & new_new_n19406__;
  assign new_new_n19413__ = new_new_n5815__ & new_new_n7658__;
  assign new_new_n19414__ = new_new_n19383__ & new_new_n19413__;
  assign new_new_n19415__ = new_new_n19411__ & new_new_n19412__;
  assign new_new_n19416__ = new_new_n19410__ & new_new_n19415__;
  assign new_new_n19417__ = new_new_n19414__ & new_new_n19416__;
  assign new_new_n19418__ = new_new_n4742__ & new_new_n19417__;
  assign new_new_n19419__ = new_new_n19399__ & new_new_n19418__;
  assign new_new_n19420__ = ~new_new_n19382__ & ~new_new_n19419__;
  assign new_new_n19421__ = ~new_new_n19381__ & ~new_new_n19420__;
  assign new_new_n19422__ = ~new_new_n19178__ & ~new_new_n19421__;
  assign new_new_n19423__ = ~new_new_n19177__ & ~new_new_n19422__;
  assign new_new_n19424__ = ~new_new_n19086__ & ~new_new_n19423__;
  assign new_new_n19425__ = new_new_n19086__ & new_new_n19423__;
  assign new_new_n19426__ = ~new_new_n168__ & ~new_new_n853__;
  assign new_new_n19427__ = ~new_new_n990__ & new_new_n19426__;
  assign new_new_n19428__ = ~new_new_n382__ & ~new_new_n489__;
  assign new_new_n19429__ = ~new_new_n993__ & new_new_n19428__;
  assign new_new_n19430__ = new_new_n1097__ & new_new_n19427__;
  assign new_new_n19431__ = new_new_n2003__ & new_new_n4001__;
  assign new_new_n19432__ = new_new_n16790__ & new_new_n19431__;
  assign new_new_n19433__ = new_new_n19429__ & new_new_n19430__;
  assign new_new_n19434__ = new_new_n7630__ & new_new_n19143__;
  assign new_new_n19435__ = new_new_n19433__ & new_new_n19434__;
  assign new_new_n19436__ = new_new_n3668__ & new_new_n19432__;
  assign new_new_n19437__ = new_new_n19275__ & new_new_n19436__;
  assign new_new_n19438__ = new_new_n19435__ & new_new_n19437__;
  assign new_new_n19439__ = new_new_n4313__ & new_new_n19438__;
  assign new_new_n19440__ = new_new_n4617__ & new_new_n19439__;
  assign new_new_n19441__ = ~new_new_n19425__ & ~new_new_n19440__;
  assign new_new_n19442__ = ~new_new_n19424__ & ~new_new_n19441__;
  assign new_new_n19443__ = ~new_new_n19075__ & new_new_n19442__;
  assign new_new_n19444__ = ~new_new_n19074__ & ~new_new_n19443__;
  assign new_new_n19445__ = new_new_n71__ & ~new_new_n15638__;
  assign new_new_n19446__ = new_new_n15582__ & new_new_n15638__;
  assign new_new_n19447__ = ~new_new_n15582__ & new_new_n15638__;
  assign new_new_n19448__ = ~new_new_n15710__ & new_new_n19447__;
  assign new_new_n19449__ = ~new_new_n15673__ & ~new_new_n19184__;
  assign new_new_n19450__ = new_new_n15661__ & ~new_new_n19449__;
  assign new_new_n19451__ = new_new_n15668__ & ~new_new_n19450__;
  assign new_new_n19452__ = new_new_n15661__ & new_new_n19104__;
  assign new_new_n19453__ = ~new_new_n19184__ & ~new_new_n19452__;
  assign new_new_n19454__ = ~new_new_n19451__ & ~new_new_n19453__;
  assign new_new_n19455__ = ~new_new_n15661__ & new_new_n19093__;
  assign new_new_n19456__ = ~new_new_n15673__ & new_new_n19368__;
  assign new_new_n19457__ = new_new_n15710__ & new_new_n19456__;
  assign new_new_n19458__ = ~new_new_n19455__ & ~new_new_n19457__;
  assign new_new_n19459__ = new_new_n15668__ & ~new_new_n19458__;
  assign new_new_n19460__ = new_new_n15643__ & new_new_n19095__;
  assign new_new_n19461__ = ~new_new_n15656__ & new_new_n15661__;
  assign new_new_n19462__ = new_new_n15643__ & ~new_new_n19461__;
  assign new_new_n19463__ = ~new_new_n19104__ & ~new_new_n19462__;
  assign new_new_n19464__ = ~new_new_n19460__ & ~new_new_n19463__;
  assign new_new_n19465__ = ~new_new_n19459__ & ~new_new_n19464__;
  assign new_new_n19466__ = ~new_new_n19454__ & new_new_n19465__;
  assign new_new_n19467__ = ~new_new_n15638__ & new_new_n15718__;
  assign new_new_n19468__ = new_new_n19466__ & new_new_n19467__;
  assign new_new_n19469__ = ~new_new_n19448__ & ~new_new_n19468__;
  assign new_new_n19470__ = new_new_n15656__ & ~new_new_n19469__;
  assign new_new_n19471__ = new_new_n19447__ & new_new_n19466__;
  assign new_new_n19472__ = ~new_new_n19467__ & ~new_new_n19471__;
  assign new_new_n19473__ = ~new_new_n15710__ & ~new_new_n19472__;
  assign new_new_n19474__ = ~new_new_n15638__ & new_new_n15716__;
  assign new_new_n19475__ = new_new_n19446__ & ~new_new_n19466__;
  assign new_new_n19476__ = ~new_new_n19474__ & ~new_new_n19475__;
  assign new_new_n19477__ = new_new_n15710__ & ~new_new_n19476__;
  assign new_new_n19478__ = new_new_n15710__ & new_new_n19446__;
  assign new_new_n19479__ = ~new_new_n19466__ & new_new_n19474__;
  assign new_new_n19480__ = ~new_new_n19478__ & ~new_new_n19479__;
  assign new_new_n19481__ = ~new_new_n15656__ & ~new_new_n19480__;
  assign new_new_n19482__ = ~new_new_n15716__ & ~new_new_n15718__;
  assign new_new_n19483__ = new_new_n15638__ & new_new_n19482__;
  assign new_new_n19484__ = ~new_new_n19470__ & ~new_new_n19483__;
  assign new_new_n19485__ = ~new_new_n19473__ & ~new_new_n19477__;
  assign new_new_n19486__ = ~new_new_n19481__ & new_new_n19485__;
  assign new_new_n19487__ = new_new_n19484__ & new_new_n19486__;
  assign new_new_n19488__ = new_new_n15638__ & ~new_new_n19487__;
  assign new_new_n19489__ = new_new_n15582__ & new_new_n19487__;
  assign new_new_n19490__ = ~new_new_n19488__ & ~new_new_n19489__;
  assign new_new_n19491__ = ~new_new_n19446__ & ~new_new_n19490__;
  assign new_new_n19492__ = ~new_new_n15743__ & ~new_new_n19491__;
  assign new_new_n19493__ = new_new_n15743__ & new_new_n19491__;
  assign new_new_n19494__ = ~new_new_n19492__ & ~new_new_n19493__;
  assign new_new_n19495__ = new_new_n765__ & new_new_n19494__;
  assign new_new_n19496__ = ~new_new_n19069__ & ~new_new_n19445__;
  assign new_new_n19497__ = ~new_new_n19495__ & new_new_n19496__;
  assign new_new_n19498__ = pi31 & ~new_new_n19497__;
  assign new_new_n19499__ = ~new_new_n161__ & ~new_new_n15743__;
  assign new_new_n19500__ = new_new_n4876__ & ~new_new_n19008__;
  assign new_new_n19501__ = ~new_new_n19499__ & new_new_n19500__;
  assign new_new_n19502__ = ~new_new_n19498__ & ~new_new_n19501__;
  assign new_new_n19503__ = new_new_n19444__ & ~new_new_n19502__;
  assign new_new_n19504__ = ~new_new_n851__ & ~new_new_n1176__;
  assign new_new_n19505__ = ~new_new_n143__ & ~new_new_n1515__;
  assign new_new_n19506__ = ~new_new_n348__ & ~new_new_n945__;
  assign new_new_n19507__ = new_new_n15877__ & new_new_n19504__;
  assign new_new_n19508__ = new_new_n19506__ & new_new_n19507__;
  assign new_new_n19509__ = ~new_new_n479__ & new_new_n19505__;
  assign new_new_n19510__ = new_new_n2336__ & new_new_n3370__;
  assign new_new_n19511__ = new_new_n16147__ & new_new_n19510__;
  assign new_new_n19512__ = new_new_n19508__ & new_new_n19509__;
  assign new_new_n19513__ = new_new_n985__ & ~new_new_n1539__;
  assign new_new_n19514__ = new_new_n19512__ & new_new_n19513__;
  assign new_new_n19515__ = new_new_n2918__ & new_new_n19511__;
  assign new_new_n19516__ = new_new_n19514__ & new_new_n19515__;
  assign new_new_n19517__ = new_new_n4072__ & new_new_n7154__;
  assign new_new_n19518__ = new_new_n19516__ & new_new_n19517__;
  assign new_new_n19519__ = new_new_n1282__ & new_new_n19518__;
  assign new_new_n19520__ = new_new_n1626__ & new_new_n19519__;
  assign new_new_n19521__ = ~new_new_n19503__ & new_new_n19520__;
  assign new_new_n19522__ = new_new_n19012__ & new_new_n19034__;
  assign new_new_n19523__ = ~new_new_n19444__ & new_new_n19502__;
  assign new_new_n19524__ = ~new_new_n19522__ & ~new_new_n19523__;
  assign new_new_n19525__ = ~new_new_n19521__ & new_new_n19524__;
  assign new_new_n19526__ = ~new_new_n19035__ & ~new_new_n19525__;
  assign new_new_n19527__ = ~new_new_n18983__ & ~new_new_n19526__;
  assign new_new_n19528__ = ~new_new_n18982__ & ~new_new_n19527__;
  assign new_new_n19529__ = ~new_new_n18963__ & ~new_new_n19528__;
  assign new_new_n19530__ = new_new_n18963__ & new_new_n19528__;
  assign new_new_n19531__ = new_new_n5059__ & ~new_new_n15615__;
  assign new_new_n19532__ = new_new_n5053__ & new_new_n15564__;
  assign new_new_n19533__ = ~new_new_n18931__ & ~new_new_n18935__;
  assign new_new_n19534__ = ~new_new_n18936__ & ~new_new_n19533__;
  assign new_new_n19535__ = pi31 & new_new_n19534__;
  assign new_new_n19536__ = ~new_new_n15572__ & ~new_new_n19535__;
  assign new_new_n19537__ = new_new_n15572__ & new_new_n19535__;
  assign new_new_n19538__ = new_new_n765__ & ~new_new_n19536__;
  assign new_new_n19539__ = ~new_new_n19537__ & new_new_n19538__;
  assign new_new_n19540__ = ~new_new_n19531__ & ~new_new_n19532__;
  assign new_new_n19541__ = ~new_new_n19539__ & new_new_n19540__;
  assign new_new_n19542__ = ~new_new_n19530__ & ~new_new_n19541__;
  assign new_new_n19543__ = ~new_new_n19529__ & ~new_new_n19542__;
  assign new_new_n19544__ = new_new_n18951__ & new_new_n19543__;
  assign new_new_n19545__ = ~new_new_n18951__ & ~new_new_n19543__;
  assign new_new_n19546__ = new_new_n18567__ & ~new_new_n18583__;
  assign new_new_n19547__ = ~new_new_n18584__ & ~new_new_n19546__;
  assign new_new_n19548__ = ~new_new_n18146__ & ~new_new_n19547__;
  assign new_new_n19549__ = new_new_n18146__ & new_new_n19547__;
  assign new_new_n19550__ = ~new_new_n19548__ & ~new_new_n19549__;
  assign new_new_n19551__ = ~new_new_n19545__ & ~new_new_n19550__;
  assign new_new_n19552__ = ~new_new_n19544__ & ~new_new_n19551__;
  assign new_new_n19553__ = ~new_new_n18927__ & new_new_n19552__;
  assign new_new_n19554__ = new_new_n18927__ & ~new_new_n19552__;
  assign new_new_n19555__ = ~new_new_n18479__ & ~new_new_n18480__;
  assign new_new_n19556__ = ~new_new_n18585__ & ~new_new_n19546__;
  assign new_new_n19557__ = new_new_n19555__ & ~new_new_n19556__;
  assign new_new_n19558__ = ~new_new_n19555__ & new_new_n19556__;
  assign new_new_n19559__ = ~new_new_n19557__ & ~new_new_n19558__;
  assign new_new_n19560__ = ~new_new_n19554__ & new_new_n19559__;
  assign new_new_n19561__ = ~new_new_n19553__ & ~new_new_n19560__;
  assign new_new_n19562__ = ~new_new_n18907__ & new_new_n19561__;
  assign new_new_n19563__ = new_new_n18907__ & ~new_new_n19561__;
  assign new_new_n19564__ = ~new_new_n18602__ & ~new_new_n18603__;
  assign new_new_n19565__ = ~new_new_n17563__ & new_new_n18606__;
  assign new_new_n19566__ = new_new_n17563__ & ~new_new_n18606__;
  assign new_new_n19567__ = ~new_new_n19565__ & ~new_new_n19566__;
  assign new_new_n19568__ = new_new_n19564__ & new_new_n19567__;
  assign new_new_n19569__ = ~new_new_n19564__ & ~new_new_n19567__;
  assign new_new_n19570__ = ~new_new_n19568__ & ~new_new_n19569__;
  assign new_new_n19571__ = ~new_new_n19563__ & ~new_new_n19570__;
  assign new_new_n19572__ = ~new_new_n19562__ & ~new_new_n19571__;
  assign new_new_n19573__ = new_new_n5191__ & ~new_new_n15432__;
  assign new_new_n19574__ = new_new_n5183__ & ~new_new_n15362__;
  assign new_new_n19575__ = ~new_new_n19573__ & ~new_new_n19574__;
  assign new_new_n19576__ = new_new_n5195__ & new_new_n17914__;
  assign new_new_n19577__ = new_new_n19575__ & ~new_new_n19576__;
  assign new_new_n19578__ = pi23 & ~new_new_n19577__;
  assign new_new_n19579__ = new_new_n5195__ & ~new_new_n17918__;
  assign new_new_n19580__ = ~pi23 & ~new_new_n19579__;
  assign new_new_n19581__ = ~pi22 & new_new_n15390__;
  assign new_new_n19582__ = pi22 & ~new_new_n15390__;
  assign new_new_n19583__ = new_new_n5195__ & new_new_n15829__;
  assign new_new_n19584__ = ~new_new_n19581__ & ~new_new_n19582__;
  assign new_new_n19585__ = new_new_n19583__ & new_new_n19584__;
  assign new_new_n19586__ = ~new_new_n19580__ & ~new_new_n19585__;
  assign new_new_n19587__ = new_new_n19575__ & ~new_new_n19586__;
  assign new_new_n19588__ = ~new_new_n19578__ & ~new_new_n19587__;
  assign new_new_n19589__ = ~new_new_n18786__ & ~new_new_n18787__;
  assign new_new_n19590__ = new_new_n18799__ & new_new_n19589__;
  assign new_new_n19591__ = ~new_new_n18799__ & ~new_new_n19589__;
  assign new_new_n19592__ = ~new_new_n19590__ & ~new_new_n19591__;
  assign new_new_n19593__ = new_new_n19588__ & new_new_n19592__;
  assign new_new_n19594__ = ~new_new_n19572__ & ~new_new_n19593__;
  assign new_new_n19595__ = ~new_new_n19588__ & ~new_new_n19592__;
  assign new_new_n19596__ = ~new_new_n19594__ & ~new_new_n19595__;
  assign new_new_n19597__ = new_new_n18895__ & ~new_new_n19596__;
  assign new_new_n19598__ = ~new_new_n18895__ & new_new_n19596__;
  assign new_new_n19599__ = new_new_n5183__ & new_new_n15390__;
  assign new_new_n19600__ = new_new_n5191__ & ~new_new_n15362__;
  assign new_new_n19601__ = ~new_new_n19599__ & ~new_new_n19600__;
  assign new_new_n19602__ = new_new_n5195__ & ~new_new_n17364__;
  assign new_new_n19603__ = pi23 & ~new_new_n19602__;
  assign new_new_n19604__ = ~pi22 & new_new_n15398__;
  assign new_new_n19605__ = pi22 & ~new_new_n15398__;
  assign new_new_n19606__ = new_new_n5195__ & ~new_new_n19604__;
  assign new_new_n19607__ = ~new_new_n19605__ & new_new_n19606__;
  assign new_new_n19608__ = new_new_n16956__ & new_new_n19607__;
  assign new_new_n19609__ = ~new_new_n19603__ & ~new_new_n19608__;
  assign new_new_n19610__ = new_new_n19601__ & ~new_new_n19609__;
  assign new_new_n19611__ = new_new_n5195__ & new_new_n17360__;
  assign new_new_n19612__ = new_new_n19601__ & ~new_new_n19611__;
  assign new_new_n19613__ = ~pi23 & ~new_new_n19612__;
  assign new_new_n19614__ = ~new_new_n19610__ & ~new_new_n19613__;
  assign new_new_n19615__ = ~new_new_n19598__ & new_new_n19614__;
  assign new_new_n19616__ = ~new_new_n19597__ & ~new_new_n19615__;
  assign new_new_n19617__ = ~new_new_n18891__ & ~new_new_n19616__;
  assign new_new_n19618__ = ~new_new_n18890__ & ~new_new_n19617__;
  assign new_new_n19619__ = ~new_new_n18763__ & ~new_new_n18764__;
  assign new_new_n19620__ = ~new_new_n18833__ & new_new_n19619__;
  assign new_new_n19621__ = new_new_n18833__ & ~new_new_n19619__;
  assign new_new_n19622__ = ~new_new_n19620__ & ~new_new_n19621__;
  assign new_new_n19623__ = new_new_n19618__ & ~new_new_n19622__;
  assign new_new_n19624__ = ~new_new_n19618__ & new_new_n19622__;
  assign new_new_n19625__ = new_new_n7935__ & new_new_n15237__;
  assign new_new_n19626__ = new_new_n6968__ & new_new_n15244__;
  assign new_new_n19627__ = new_new_n6964__ & ~new_new_n15248__;
  assign new_new_n19628__ = new_new_n6959__ & ~new_new_n16603__;
  assign new_new_n19629__ = ~new_new_n19626__ & ~new_new_n19627__;
  assign new_new_n19630__ = ~new_new_n19625__ & new_new_n19629__;
  assign new_new_n19631__ = ~new_new_n19628__ & new_new_n19630__;
  assign new_new_n19632__ = ~pi17 & ~new_new_n19631__;
  assign new_new_n19633__ = pi17 & new_new_n19631__;
  assign new_new_n19634__ = ~new_new_n19632__ & ~new_new_n19633__;
  assign new_new_n19635__ = ~new_new_n19624__ & ~new_new_n19634__;
  assign new_new_n19636__ = ~new_new_n19623__ & ~new_new_n19635__;
  assign new_new_n19637__ = new_new_n18873__ & new_new_n19636__;
  assign new_new_n19638__ = ~new_new_n18873__ & ~new_new_n19636__;
  assign new_new_n19639__ = ~pi20 & new_new_n18835__;
  assign new_new_n19640__ = pi20 & ~new_new_n18835__;
  assign new_new_n19641__ = ~new_new_n19639__ & ~new_new_n19640__;
  assign new_new_n19642__ = ~new_new_n18844__ & new_new_n19641__;
  assign new_new_n19643__ = new_new_n18844__ & ~new_new_n19641__;
  assign new_new_n19644__ = ~new_new_n19642__ & ~new_new_n19643__;
  assign new_new_n19645__ = new_new_n18746__ & new_new_n19644__;
  assign new_new_n19646__ = ~new_new_n18746__ & ~new_new_n19644__;
  assign new_new_n19647__ = ~new_new_n19645__ & ~new_new_n19646__;
  assign new_new_n19648__ = ~new_new_n19638__ & new_new_n19647__;
  assign new_new_n19649__ = ~new_new_n19637__ & ~new_new_n19648__;
  assign new_new_n19650__ = ~new_new_n18861__ & ~new_new_n19649__;
  assign new_new_n19651__ = ~new_new_n18860__ & ~new_new_n19650__;
  assign new_new_n19652__ = pi14 & new_new_n16630__;
  assign new_new_n19653__ = pi13 & ~new_new_n16630__;
  assign new_new_n19654__ = new_new_n6994__ & ~new_new_n19652__;
  assign new_new_n19655__ = ~new_new_n19653__ & new_new_n19654__;
  assign new_new_n19656__ = new_new_n6991__ & ~new_new_n15998__;
  assign new_new_n19657__ = new_new_n6985__ & ~new_new_n16056__;
  assign new_new_n19658__ = ~new_new_n19656__ & ~new_new_n19657__;
  assign new_new_n19659__ = ~pi14 & ~new_new_n19658__;
  assign new_new_n19660__ = new_new_n18722__ & new_new_n19658__;
  assign new_new_n19661__ = ~new_new_n19659__ & ~new_new_n19660__;
  assign new_new_n19662__ = ~new_new_n19655__ & new_new_n19661__;
  assign new_new_n19663__ = ~new_new_n19623__ & ~new_new_n19624__;
  assign new_new_n19664__ = new_new_n19634__ & new_new_n19663__;
  assign new_new_n19665__ = ~new_new_n19634__ & ~new_new_n19663__;
  assign new_new_n19666__ = ~new_new_n19664__ & ~new_new_n19665__;
  assign new_new_n19667__ = new_new_n6634__ & ~new_new_n15273__;
  assign new_new_n19668__ = new_new_n6629__ & ~new_new_n15321__;
  assign new_new_n19669__ = ~new_new_n6625__ & ~new_new_n15349__;
  assign new_new_n19670__ = new_new_n6936__ & ~new_new_n17103__;
  assign new_new_n19671__ = ~new_new_n19668__ & ~new_new_n19669__;
  assign new_new_n19672__ = ~new_new_n19667__ & new_new_n19671__;
  assign new_new_n19673__ = ~new_new_n19670__ & new_new_n19672__;
  assign new_new_n19674__ = ~pi20 & ~new_new_n19673__;
  assign new_new_n19675__ = pi20 & new_new_n19673__;
  assign new_new_n19676__ = ~new_new_n19674__ & ~new_new_n19675__;
  assign new_new_n19677__ = ~pi19 & ~new_new_n15398__;
  assign new_new_n19678__ = new_new_n6622__ & new_new_n19677__;
  assign new_new_n19679__ = pi20 & ~new_new_n19678__;
  assign new_new_n19680__ = ~new_new_n15398__ & new_new_n16182__;
  assign new_new_n19681__ = ~new_new_n19679__ & ~new_new_n19680__;
  assign new_new_n19682__ = new_new_n6936__ & new_new_n16458__;
  assign new_new_n19683__ = new_new_n6629__ & ~new_new_n15349__;
  assign new_new_n19684__ = new_new_n6634__ & ~new_new_n15321__;
  assign new_new_n19685__ = ~new_new_n19683__ & ~new_new_n19684__;
  assign new_new_n19686__ = ~new_new_n19682__ & new_new_n19685__;
  assign new_new_n19687__ = ~new_new_n19681__ & new_new_n19686__;
  assign new_new_n19688__ = ~pi20 & ~new_new_n19686__;
  assign new_new_n19689__ = ~new_new_n19687__ & ~new_new_n19688__;
  assign new_new_n19690__ = ~new_new_n19562__ & ~new_new_n19563__;
  assign new_new_n19691__ = ~new_new_n19570__ & new_new_n19690__;
  assign new_new_n19692__ = new_new_n19570__ & ~new_new_n19690__;
  assign new_new_n19693__ = ~new_new_n19691__ & ~new_new_n19692__;
  assign new_new_n19694__ = ~new_new_n4900__ & ~new_new_n18633__;
  assign new_new_n19695__ = ~new_new_n333__ & ~new_new_n15487__;
  assign new_new_n19696__ = new_new_n873__ & ~new_new_n15809__;
  assign new_new_n19697__ = ~new_new_n19695__ & ~new_new_n19696__;
  assign new_new_n19698__ = ~new_new_n19694__ & new_new_n19697__;
  assign new_new_n19699__ = pi26 & ~new_new_n19698__;
  assign new_new_n19700__ = new_new_n512__ & ~new_new_n15471__;
  assign new_new_n19701__ = new_new_n801__ & ~new_new_n15471__;
  assign new_new_n19702__ = ~pi26 & ~new_new_n19701__;
  assign new_new_n19703__ = ~new_new_n19700__ & ~new_new_n19702__;
  assign new_new_n19704__ = new_new_n19698__ & ~new_new_n19703__;
  assign new_new_n19705__ = ~new_new_n19699__ & ~new_new_n19704__;
  assign new_new_n19706__ = ~new_new_n4900__ & new_new_n18020__;
  assign new_new_n19707__ = ~new_new_n333__ & new_new_n15524__;
  assign new_new_n19708__ = new_new_n873__ & ~new_new_n15487__;
  assign new_new_n19709__ = ~new_new_n19707__ & ~new_new_n19708__;
  assign new_new_n19710__ = ~new_new_n19706__ & new_new_n19709__;
  assign new_new_n19711__ = pi26 & ~new_new_n19710__;
  assign new_new_n19712__ = new_new_n512__ & ~new_new_n15809__;
  assign new_new_n19713__ = new_new_n801__ & ~new_new_n15809__;
  assign new_new_n19714__ = ~pi26 & ~new_new_n19713__;
  assign new_new_n19715__ = ~new_new_n19712__ & ~new_new_n19714__;
  assign new_new_n19716__ = new_new_n19710__ & ~new_new_n19715__;
  assign new_new_n19717__ = ~new_new_n19711__ & ~new_new_n19716__;
  assign new_new_n19718__ = ~new_new_n19544__ & ~new_new_n19545__;
  assign new_new_n19719__ = ~new_new_n19550__ & new_new_n19718__;
  assign new_new_n19720__ = new_new_n19550__ & ~new_new_n19718__;
  assign new_new_n19721__ = ~new_new_n19719__ & ~new_new_n19720__;
  assign new_new_n19722__ = new_new_n19717__ & ~new_new_n19721__;
  assign new_new_n19723__ = ~new_new_n19717__ & new_new_n19721__;
  assign new_new_n19724__ = new_new_n4815__ & new_new_n15520__;
  assign new_new_n19725__ = ~new_new_n4818__ & new_new_n15767__;
  assign new_new_n19726__ = new_new_n4212__ & ~new_new_n15533__;
  assign new_new_n19727__ = ~new_new_n19725__ & ~new_new_n19726__;
  assign new_new_n19728__ = ~new_new_n19724__ & new_new_n19727__;
  assign new_new_n19729__ = ~new_new_n18430__ & ~new_new_n18911__;
  assign new_new_n19730__ = new_new_n15520__ & ~new_new_n19729__;
  assign new_new_n19731__ = ~new_new_n18432__ & ~new_new_n19730__;
  assign new_new_n19732__ = new_new_n4214__ & new_new_n19731__;
  assign new_new_n19733__ = pi29 & ~new_new_n19732__;
  assign new_new_n19734__ = new_new_n4825__ & new_new_n19731__;
  assign new_new_n19735__ = ~new_new_n19733__ & ~new_new_n19734__;
  assign new_new_n19736__ = new_new_n19728__ & ~new_new_n19735__;
  assign new_new_n19737__ = ~pi29 & ~new_new_n19728__;
  assign new_new_n19738__ = ~new_new_n19736__ & ~new_new_n19737__;
  assign new_new_n19739__ = ~new_new_n19723__ & ~new_new_n19738__;
  assign new_new_n19740__ = ~new_new_n19722__ & ~new_new_n19739__;
  assign new_new_n19741__ = new_new_n19705__ & ~new_new_n19740__;
  assign new_new_n19742__ = ~new_new_n19705__ & new_new_n19740__;
  assign new_new_n19743__ = ~new_new_n19553__ & ~new_new_n19554__;
  assign new_new_n19744__ = new_new_n19559__ & new_new_n19743__;
  assign new_new_n19745__ = ~new_new_n19559__ & ~new_new_n19743__;
  assign new_new_n19746__ = ~new_new_n19744__ & ~new_new_n19745__;
  assign new_new_n19747__ = ~new_new_n19742__ & new_new_n19746__;
  assign new_new_n19748__ = ~new_new_n19741__ & ~new_new_n19747__;
  assign new_new_n19749__ = ~new_new_n19693__ & ~new_new_n19748__;
  assign new_new_n19750__ = new_new_n19693__ & new_new_n19748__;
  assign new_new_n19751__ = new_new_n5183__ & ~new_new_n15432__;
  assign new_new_n19752__ = new_new_n5191__ & ~new_new_n15439__;
  assign new_new_n19753__ = new_new_n5212__ & ~new_new_n16771__;
  assign new_new_n19754__ = ~new_new_n5212__ & new_new_n15362__;
  assign new_new_n19755__ = new_new_n5195__ & ~new_new_n19754__;
  assign new_new_n19756__ = ~new_new_n19753__ & new_new_n19755__;
  assign new_new_n19757__ = ~new_new_n19751__ & ~new_new_n19752__;
  assign new_new_n19758__ = ~new_new_n19756__ & new_new_n19757__;
  assign new_new_n19759__ = ~pi23 & ~new_new_n19758__;
  assign new_new_n19760__ = pi23 & new_new_n19758__;
  assign new_new_n19761__ = ~new_new_n19759__ & ~new_new_n19760__;
  assign new_new_n19762__ = ~new_new_n19750__ & ~new_new_n19761__;
  assign new_new_n19763__ = ~new_new_n19749__ & ~new_new_n19762__;
  assign new_new_n19764__ = ~new_new_n19588__ & new_new_n19763__;
  assign new_new_n19765__ = new_new_n19588__ & ~new_new_n19763__;
  assign new_new_n19766__ = ~new_new_n19764__ & ~new_new_n19765__;
  assign new_new_n19767__ = ~new_new_n19572__ & new_new_n19766__;
  assign new_new_n19768__ = new_new_n19572__ & ~new_new_n19766__;
  assign new_new_n19769__ = ~new_new_n19767__ & ~new_new_n19768__;
  assign new_new_n19770__ = new_new_n19592__ & new_new_n19769__;
  assign new_new_n19771__ = ~new_new_n19592__ & ~new_new_n19769__;
  assign new_new_n19772__ = ~new_new_n19770__ & ~new_new_n19771__;
  assign new_new_n19773__ = new_new_n19689__ & ~new_new_n19772__;
  assign new_new_n19774__ = new_new_n19763__ & new_new_n19772__;
  assign new_new_n19775__ = ~new_new_n19773__ & ~new_new_n19774__;
  assign new_new_n19776__ = new_new_n19676__ & ~new_new_n19775__;
  assign new_new_n19777__ = ~new_new_n19676__ & new_new_n19775__;
  assign new_new_n19778__ = ~new_new_n19597__ & ~new_new_n19598__;
  assign new_new_n19779__ = ~new_new_n19614__ & ~new_new_n19778__;
  assign new_new_n19780__ = new_new_n19614__ & new_new_n19778__;
  assign new_new_n19781__ = ~new_new_n19779__ & ~new_new_n19780__;
  assign new_new_n19782__ = ~new_new_n19777__ & new_new_n19781__;
  assign new_new_n19783__ = ~new_new_n19776__ & ~new_new_n19782__;
  assign new_new_n19784__ = ~new_new_n18890__ & ~new_new_n18891__;
  assign new_new_n19785__ = ~new_new_n19616__ & new_new_n19784__;
  assign new_new_n19786__ = new_new_n19616__ & ~new_new_n19784__;
  assign new_new_n19787__ = ~new_new_n19785__ & ~new_new_n19786__;
  assign new_new_n19788__ = new_new_n19783__ & ~new_new_n19787__;
  assign new_new_n19789__ = ~new_new_n19783__ & new_new_n19787__;
  assign new_new_n19790__ = new_new_n6964__ & ~new_new_n15314__;
  assign new_new_n19791__ = new_new_n6968__ & ~new_new_n15248__;
  assign new_new_n19792__ = new_new_n7935__ & new_new_n15244__;
  assign new_new_n19793__ = ~new_new_n19790__ & ~new_new_n19791__;
  assign new_new_n19794__ = ~new_new_n19792__ & new_new_n19793__;
  assign new_new_n19795__ = new_new_n6958__ & new_new_n16378__;
  assign new_new_n19796__ = pi17 & ~new_new_n19795__;
  assign new_new_n19797__ = new_new_n7942__ & new_new_n16378__;
  assign new_new_n19798__ = ~new_new_n19796__ & ~new_new_n19797__;
  assign new_new_n19799__ = new_new_n19794__ & ~new_new_n19798__;
  assign new_new_n19800__ = ~pi17 & ~new_new_n19794__;
  assign new_new_n19801__ = ~new_new_n19799__ & ~new_new_n19800__;
  assign new_new_n19802__ = ~new_new_n19789__ & ~new_new_n19801__;
  assign new_new_n19803__ = ~new_new_n19788__ & ~new_new_n19802__;
  assign new_new_n19804__ = ~pi14 & ~new_new_n16051__;
  assign new_new_n19805__ = ~pi13 & new_new_n16051__;
  assign new_new_n19806__ = new_new_n6994__ & ~new_new_n16056__;
  assign new_new_n19807__ = ~new_new_n19804__ & new_new_n19806__;
  assign new_new_n19808__ = ~new_new_n19805__ & new_new_n19807__;
  assign new_new_n19809__ = new_new_n6985__ & ~new_new_n15998__;
  assign new_new_n19810__ = new_new_n6991__ & new_new_n15905__;
  assign new_new_n19811__ = ~new_new_n19809__ & ~new_new_n19810__;
  assign new_new_n19812__ = pi14 & ~new_new_n19811__;
  assign new_new_n19813__ = ~pi14 & ~new_new_n19806__;
  assign new_new_n19814__ = new_new_n19811__ & new_new_n19813__;
  assign new_new_n19815__ = ~new_new_n19812__ & ~new_new_n19814__;
  assign new_new_n19816__ = ~new_new_n19808__ & new_new_n19815__;
  assign new_new_n19817__ = new_new_n19803__ & ~new_new_n19816__;
  assign new_new_n19818__ = ~new_new_n19803__ & new_new_n19816__;
  assign new_new_n19819__ = ~new_new_n19817__ & ~new_new_n19818__;
  assign new_new_n19820__ = new_new_n19666__ & new_new_n19819__;
  assign new_new_n19821__ = ~new_new_n19666__ & ~new_new_n19819__;
  assign new_new_n19822__ = ~new_new_n19820__ & ~new_new_n19821__;
  assign new_new_n19823__ = pi12 & pi13;
  assign new_new_n19824__ = ~pi12 & ~pi13;
  assign new_new_n19825__ = ~new_new_n19823__ & ~new_new_n19824__;
  assign new_new_n19826__ = new_new_n15905__ & new_new_n19825__;
  assign new_new_n19827__ = pi14 & ~new_new_n19824__;
  assign new_new_n19828__ = ~pi14 & ~new_new_n19823__;
  assign new_new_n19829__ = ~new_new_n19827__ & ~new_new_n19828__;
  assign new_new_n19830__ = new_new_n15237__ & new_new_n19829__;
  assign new_new_n19831__ = ~new_new_n19826__ & ~new_new_n19830__;
  assign new_new_n19832__ = ~new_new_n6994__ & ~new_new_n19831__;
  assign new_new_n19833__ = new_new_n6994__ & ~new_new_n15998__;
  assign new_new_n19834__ = new_new_n16025__ & new_new_n19833__;
  assign new_new_n19835__ = ~new_new_n19832__ & ~new_new_n19834__;
  assign new_new_n19836__ = ~pi14 & ~new_new_n19835__;
  assign new_new_n19837__ = ~pi13 & ~new_new_n16684__;
  assign new_new_n19838__ = pi13 & ~new_new_n16682__;
  assign new_new_n19839__ = new_new_n6994__ & ~new_new_n19837__;
  assign new_new_n19840__ = ~new_new_n19838__ & new_new_n19839__;
  assign new_new_n19841__ = new_new_n6994__ & ~new_new_n16679__;
  assign new_new_n19842__ = pi14 & ~new_new_n19832__;
  assign new_new_n19843__ = ~new_new_n19841__ & new_new_n19842__;
  assign new_new_n19844__ = ~new_new_n19836__ & ~new_new_n19840__;
  assign new_new_n19845__ = ~new_new_n19843__ & new_new_n19844__;
  assign new_new_n19846__ = new_new_n7935__ & ~new_new_n15314__;
  assign new_new_n19847__ = new_new_n6964__ & ~new_new_n15273__;
  assign new_new_n19848__ = new_new_n6968__ & new_new_n15285__;
  assign new_new_n19849__ = ~new_new_n19847__ & ~new_new_n19848__;
  assign new_new_n19850__ = ~new_new_n19846__ & new_new_n19849__;
  assign new_new_n19851__ = new_new_n6958__ & new_new_n17140__;
  assign new_new_n19852__ = pi17 & ~new_new_n19851__;
  assign new_new_n19853__ = new_new_n7942__ & new_new_n17140__;
  assign new_new_n19854__ = ~new_new_n19852__ & ~new_new_n19853__;
  assign new_new_n19855__ = new_new_n19850__ & ~new_new_n19854__;
  assign new_new_n19856__ = ~pi17 & ~new_new_n19850__;
  assign new_new_n19857__ = ~new_new_n19855__ & ~new_new_n19856__;
  assign new_new_n19858__ = ~new_new_n19749__ & ~new_new_n19750__;
  assign new_new_n19859__ = ~new_new_n19761__ & new_new_n19858__;
  assign new_new_n19860__ = new_new_n19761__ & ~new_new_n19858__;
  assign new_new_n19861__ = ~new_new_n19859__ & ~new_new_n19860__;
  assign new_new_n19862__ = new_new_n5213__ & ~new_new_n15439__;
  assign new_new_n19863__ = new_new_n5191__ & ~new_new_n15471__;
  assign new_new_n19864__ = new_new_n5183__ & new_new_n15464__;
  assign new_new_n19865__ = new_new_n5215__ & ~new_new_n17240__;
  assign new_new_n19866__ = ~new_new_n19862__ & ~new_new_n19863__;
  assign new_new_n19867__ = ~new_new_n19864__ & new_new_n19866__;
  assign new_new_n19868__ = ~new_new_n19865__ & new_new_n19867__;
  assign new_new_n19869__ = pi23 & ~new_new_n19868__;
  assign new_new_n19870__ = ~pi23 & new_new_n19868__;
  assign new_new_n19871__ = ~new_new_n19869__ & ~new_new_n19870__;
  assign new_new_n19872__ = ~new_new_n333__ & new_new_n15520__;
  assign new_new_n19873__ = new_new_n873__ & new_new_n15524__;
  assign new_new_n19874__ = new_new_n3311__ & ~new_new_n15487__;
  assign new_new_n19875__ = ~new_new_n19872__ & ~new_new_n19873__;
  assign new_new_n19876__ = ~new_new_n19874__ & new_new_n19875__;
  assign new_new_n19877__ = ~pi26 & ~new_new_n19876__;
  assign new_new_n19878__ = new_new_n512__ & new_new_n17587__;
  assign new_new_n19879__ = new_new_n801__ & new_new_n17587__;
  assign new_new_n19880__ = pi26 & ~new_new_n19879__;
  assign new_new_n19881__ = ~new_new_n19878__ & ~new_new_n19880__;
  assign new_new_n19882__ = new_new_n19876__ & ~new_new_n19881__;
  assign new_new_n19883__ = ~new_new_n19877__ & ~new_new_n19882__;
  assign new_new_n19884__ = ~new_new_n4818__ & new_new_n15560__;
  assign new_new_n19885__ = new_new_n4212__ & new_new_n15767__;
  assign new_new_n19886__ = new_new_n4815__ & ~new_new_n15533__;
  assign new_new_n19887__ = ~new_new_n19884__ & ~new_new_n19885__;
  assign new_new_n19888__ = ~new_new_n19886__ & new_new_n19887__;
  assign new_new_n19889__ = ~new_new_n18201__ & ~new_new_n18934__;
  assign new_new_n19890__ = new_new_n18451__ & new_new_n19889__;
  assign new_new_n19891__ = ~new_new_n15533__ & new_new_n19890__;
  assign new_new_n19892__ = new_new_n15533__ & ~new_new_n19890__;
  assign new_new_n19893__ = ~new_new_n19891__ & ~new_new_n19892__;
  assign new_new_n19894__ = new_new_n4214__ & new_new_n19893__;
  assign new_new_n19895__ = pi29 & ~new_new_n19894__;
  assign new_new_n19896__ = new_new_n4825__ & new_new_n19893__;
  assign new_new_n19897__ = ~new_new_n19895__ & ~new_new_n19896__;
  assign new_new_n19898__ = new_new_n19888__ & ~new_new_n19897__;
  assign new_new_n19899__ = ~pi29 & ~new_new_n19888__;
  assign new_new_n19900__ = ~new_new_n19898__ & ~new_new_n19899__;
  assign new_new_n19901__ = new_new_n19883__ & new_new_n19900__;
  assign new_new_n19902__ = ~new_new_n19883__ & ~new_new_n19900__;
  assign new_new_n19903__ = ~new_new_n19529__ & ~new_new_n19530__;
  assign new_new_n19904__ = new_new_n19541__ & ~new_new_n19903__;
  assign new_new_n19905__ = ~new_new_n19541__ & new_new_n19903__;
  assign new_new_n19906__ = ~new_new_n19904__ & ~new_new_n19905__;
  assign new_new_n19907__ = ~new_new_n19902__ & ~new_new_n19906__;
  assign new_new_n19908__ = ~new_new_n19901__ & ~new_new_n19907__;
  assign new_new_n19909__ = ~new_new_n19871__ & ~new_new_n19908__;
  assign new_new_n19910__ = new_new_n19871__ & new_new_n19908__;
  assign new_new_n19911__ = ~new_new_n19722__ & ~new_new_n19723__;
  assign new_new_n19912__ = ~new_new_n19738__ & new_new_n19911__;
  assign new_new_n19913__ = new_new_n19738__ & ~new_new_n19911__;
  assign new_new_n19914__ = ~new_new_n19912__ & ~new_new_n19913__;
  assign new_new_n19915__ = ~new_new_n19910__ & ~new_new_n19914__;
  assign new_new_n19916__ = ~new_new_n19909__ & ~new_new_n19915__;
  assign new_new_n19917__ = ~new_new_n19741__ & ~new_new_n19742__;
  assign new_new_n19918__ = new_new_n19746__ & new_new_n19917__;
  assign new_new_n19919__ = ~new_new_n19746__ & ~new_new_n19917__;
  assign new_new_n19920__ = ~new_new_n19918__ & ~new_new_n19919__;
  assign new_new_n19921__ = ~new_new_n19916__ & ~new_new_n19920__;
  assign new_new_n19922__ = new_new_n19916__ & new_new_n19920__;
  assign new_new_n19923__ = new_new_n5213__ & ~new_new_n15432__;
  assign new_new_n19924__ = new_new_n5183__ & ~new_new_n15439__;
  assign new_new_n19925__ = new_new_n5191__ & new_new_n15464__;
  assign new_new_n19926__ = new_new_n5215__ & new_new_n17204__;
  assign new_new_n19927__ = ~new_new_n19924__ & ~new_new_n19925__;
  assign new_new_n19928__ = ~new_new_n19923__ & new_new_n19927__;
  assign new_new_n19929__ = ~new_new_n19926__ & new_new_n19928__;
  assign new_new_n19930__ = pi23 & ~new_new_n19929__;
  assign new_new_n19931__ = ~pi23 & new_new_n19929__;
  assign new_new_n19932__ = ~new_new_n19930__ & ~new_new_n19931__;
  assign new_new_n19933__ = ~new_new_n19922__ & ~new_new_n19932__;
  assign new_new_n19934__ = ~new_new_n19921__ & ~new_new_n19933__;
  assign new_new_n19935__ = ~new_new_n19861__ & ~new_new_n19934__;
  assign new_new_n19936__ = new_new_n19861__ & new_new_n19934__;
  assign new_new_n19937__ = new_new_n6634__ & ~new_new_n15349__;
  assign new_new_n19938__ = ~new_new_n6625__ & new_new_n15390__;
  assign new_new_n19939__ = new_new_n6629__ & ~new_new_n15398__;
  assign new_new_n19940__ = new_new_n6936__ & ~new_new_n17180__;
  assign new_new_n19941__ = ~new_new_n19938__ & ~new_new_n19939__;
  assign new_new_n19942__ = ~new_new_n19937__ & new_new_n19941__;
  assign new_new_n19943__ = ~new_new_n19940__ & new_new_n19942__;
  assign new_new_n19944__ = pi20 & ~new_new_n19943__;
  assign new_new_n19945__ = ~pi20 & new_new_n19943__;
  assign new_new_n19946__ = ~new_new_n19944__ & ~new_new_n19945__;
  assign new_new_n19947__ = ~new_new_n19936__ & ~new_new_n19946__;
  assign new_new_n19948__ = ~new_new_n19935__ & ~new_new_n19947__;
  assign new_new_n19949__ = new_new_n19857__ & ~new_new_n19948__;
  assign new_new_n19950__ = ~new_new_n19857__ & new_new_n19948__;
  assign new_new_n19951__ = ~new_new_n19689__ & new_new_n19772__;
  assign new_new_n19952__ = ~new_new_n19773__ & ~new_new_n19951__;
  assign new_new_n19953__ = ~new_new_n19950__ & new_new_n19952__;
  assign new_new_n19954__ = ~new_new_n19949__ & ~new_new_n19953__;
  assign new_new_n19955__ = ~new_new_n19776__ & ~new_new_n19777__;
  assign new_new_n19956__ = new_new_n19781__ & new_new_n19955__;
  assign new_new_n19957__ = ~new_new_n19781__ & ~new_new_n19955__;
  assign new_new_n19958__ = ~new_new_n19956__ & ~new_new_n19957__;
  assign new_new_n19959__ = ~new_new_n19954__ & new_new_n19958__;
  assign new_new_n19960__ = new_new_n19954__ & ~new_new_n19958__;
  assign new_new_n19961__ = new_new_n6968__ & ~new_new_n15314__;
  assign new_new_n19962__ = new_new_n7935__ & ~new_new_n15248__;
  assign new_new_n19963__ = new_new_n6964__ & new_new_n15285__;
  assign new_new_n19964__ = new_new_n6959__ & new_new_n16725__;
  assign new_new_n19965__ = ~new_new_n19961__ & ~new_new_n19963__;
  assign new_new_n19966__ = ~new_new_n19962__ & new_new_n19965__;
  assign new_new_n19967__ = ~new_new_n19964__ & new_new_n19966__;
  assign new_new_n19968__ = pi17 & ~new_new_n19967__;
  assign new_new_n19969__ = ~pi17 & new_new_n19967__;
  assign new_new_n19970__ = ~new_new_n19968__ & ~new_new_n19969__;
  assign new_new_n19971__ = ~new_new_n19960__ & ~new_new_n19970__;
  assign new_new_n19972__ = ~new_new_n19959__ & ~new_new_n19971__;
  assign new_new_n19973__ = ~new_new_n19845__ & new_new_n19972__;
  assign new_new_n19974__ = new_new_n19845__ & ~new_new_n19972__;
  assign new_new_n19975__ = ~new_new_n19788__ & ~new_new_n19789__;
  assign new_new_n19976__ = ~new_new_n19801__ & new_new_n19975__;
  assign new_new_n19977__ = new_new_n19801__ & ~new_new_n19975__;
  assign new_new_n19978__ = ~new_new_n19976__ & ~new_new_n19977__;
  assign new_new_n19979__ = ~new_new_n19974__ & new_new_n19978__;
  assign new_new_n19980__ = ~new_new_n19973__ & ~new_new_n19979__;
  assign new_new_n19981__ = ~new_new_n19822__ & ~new_new_n19980__;
  assign new_new_n19982__ = new_new_n19822__ & new_new_n19980__;
  assign new_new_n19983__ = ~new_new_n17447__ & ~new_new_n19982__;
  assign new_new_n19984__ = ~new_new_n19981__ & ~new_new_n19983__;
  assign new_new_n19985__ = ~new_new_n19637__ & ~new_new_n19638__;
  assign new_new_n19986__ = new_new_n19647__ & new_new_n19985__;
  assign new_new_n19987__ = ~new_new_n19647__ & ~new_new_n19985__;
  assign new_new_n19988__ = ~new_new_n19986__ & ~new_new_n19987__;
  assign new_new_n19989__ = new_new_n19984__ & new_new_n19988__;
  assign new_new_n19990__ = ~new_new_n19973__ & ~new_new_n19974__;
  assign new_new_n19991__ = ~new_new_n19978__ & new_new_n19990__;
  assign new_new_n19992__ = new_new_n19978__ & ~new_new_n19990__;
  assign new_new_n19993__ = ~new_new_n19991__ & ~new_new_n19992__;
  assign new_new_n19994__ = ~pi10 & new_new_n16056__;
  assign new_new_n19995__ = pi11 & ~new_new_n19994__;
  assign new_new_n19996__ = ~pi08 & new_new_n8302__;
  assign new_new_n19997__ = ~new_new_n19995__ & ~new_new_n19996__;
  assign new_new_n19998__ = ~pi09 & ~new_new_n19997__;
  assign new_new_n19999__ = new_new_n8467__ & ~new_new_n8469__;
  assign new_new_n20000__ = new_new_n16056__ & new_new_n19999__;
  assign new_new_n20001__ = ~new_new_n8466__ & ~new_new_n20000__;
  assign new_new_n20002__ = pi09 & ~new_new_n20001__;
  assign new_new_n20003__ = pi11 & new_new_n8469__;
  assign new_new_n20004__ = ~new_new_n20002__ & ~new_new_n20003__;
  assign new_new_n20005__ = ~new_new_n19998__ & new_new_n20004__;
  assign new_new_n20006__ = ~new_new_n19993__ & new_new_n20005__;
  assign new_new_n20007__ = new_new_n19993__ & ~new_new_n20005__;
  assign new_new_n20008__ = ~new_new_n19959__ & ~new_new_n19960__;
  assign new_new_n20009__ = ~new_new_n19970__ & new_new_n20008__;
  assign new_new_n20010__ = new_new_n19970__ & ~new_new_n20008__;
  assign new_new_n20011__ = ~new_new_n20009__ & ~new_new_n20010__;
  assign new_new_n20012__ = new_new_n6994__ & new_new_n15852__;
  assign new_new_n20013__ = new_new_n6985__ & ~new_new_n15244__;
  assign new_new_n20014__ = ~new_new_n10998__ & new_new_n15248__;
  assign new_new_n20015__ = ~new_new_n10772__ & ~new_new_n10998__;
  assign new_new_n20016__ = ~new_new_n20014__ & ~new_new_n20015__;
  assign new_new_n20017__ = ~new_new_n20013__ & new_new_n20016__;
  assign new_new_n20018__ = ~new_new_n20012__ & new_new_n20017__;
  assign new_new_n20019__ = pi14 & ~new_new_n20018__;
  assign new_new_n20020__ = pi13 & new_new_n16602__;
  assign new_new_n20021__ = ~pi13 & ~new_new_n15850__;
  assign new_new_n20022__ = new_new_n15912__ & new_new_n20021__;
  assign new_new_n20023__ = ~new_new_n20020__ & ~new_new_n20022__;
  assign new_new_n20024__ = new_new_n6994__ & ~new_new_n20023__;
  assign new_new_n20025__ = new_new_n6994__ & ~new_new_n16601__;
  assign new_new_n20026__ = ~pi14 & new_new_n20017__;
  assign new_new_n20027__ = ~new_new_n20025__ & new_new_n20026__;
  assign new_new_n20028__ = ~new_new_n20019__ & ~new_new_n20027__;
  assign new_new_n20029__ = ~new_new_n20024__ & new_new_n20028__;
  assign new_new_n20030__ = ~new_new_n19935__ & ~new_new_n19936__;
  assign new_new_n20031__ = ~new_new_n19946__ & new_new_n20030__;
  assign new_new_n20032__ = new_new_n19946__ & ~new_new_n20030__;
  assign new_new_n20033__ = ~new_new_n20031__ & ~new_new_n20032__;
  assign new_new_n20034__ = new_new_n6629__ & new_new_n15390__;
  assign new_new_n20035__ = ~new_new_n6625__ & ~new_new_n15362__;
  assign new_new_n20036__ = ~new_new_n20034__ & ~new_new_n20035__;
  assign new_new_n20037__ = new_new_n6631__ & ~new_new_n17364__;
  assign new_new_n20038__ = pi20 & ~new_new_n20037__;
  assign new_new_n20039__ = pi19 & new_new_n15398__;
  assign new_new_n20040__ = ~new_new_n19677__ & ~new_new_n20039__;
  assign new_new_n20041__ = new_new_n6631__ & new_new_n16956__;
  assign new_new_n20042__ = ~new_new_n20040__ & new_new_n20041__;
  assign new_new_n20043__ = ~new_new_n20038__ & ~new_new_n20042__;
  assign new_new_n20044__ = new_new_n20036__ & ~new_new_n20043__;
  assign new_new_n20045__ = new_new_n6631__ & new_new_n17360__;
  assign new_new_n20046__ = new_new_n20036__ & ~new_new_n20045__;
  assign new_new_n20047__ = ~pi20 & ~new_new_n20046__;
  assign new_new_n20048__ = ~new_new_n20044__ & ~new_new_n20047__;
  assign new_new_n20049__ = ~new_new_n19921__ & ~new_new_n19922__;
  assign new_new_n20050__ = new_new_n19932__ & ~new_new_n20049__;
  assign new_new_n20051__ = ~new_new_n19932__ & new_new_n20049__;
  assign new_new_n20052__ = ~new_new_n20050__ & ~new_new_n20051__;
  assign new_new_n20053__ = new_new_n20048__ & new_new_n20052__;
  assign new_new_n20054__ = ~new_new_n20048__ & ~new_new_n20052__;
  assign new_new_n20055__ = new_new_n6629__ & ~new_new_n15362__;
  assign new_new_n20056__ = ~new_new_n6633__ & new_new_n15829__;
  assign new_new_n20057__ = ~new_new_n15390__ & ~new_new_n20056__;
  assign new_new_n20058__ = new_new_n15390__ & new_new_n20056__;
  assign new_new_n20059__ = new_new_n6631__ & ~new_new_n20057__;
  assign new_new_n20060__ = ~new_new_n20058__ & new_new_n20059__;
  assign new_new_n20061__ = ~new_new_n20055__ & ~new_new_n20060__;
  assign new_new_n20062__ = ~pi20 & ~new_new_n20061__;
  assign new_new_n20063__ = new_new_n6623__ & ~new_new_n15432__;
  assign new_new_n20064__ = pi20 & ~new_new_n20063__;
  assign new_new_n20065__ = new_new_n9920__ & ~new_new_n15432__;
  assign new_new_n20066__ = ~new_new_n20064__ & ~new_new_n20065__;
  assign new_new_n20067__ = new_new_n20061__ & ~new_new_n20066__;
  assign new_new_n20068__ = ~new_new_n20062__ & ~new_new_n20067__;
  assign new_new_n20069__ = ~new_new_n19909__ & ~new_new_n19910__;
  assign new_new_n20070__ = ~new_new_n19914__ & new_new_n20069__;
  assign new_new_n20071__ = new_new_n19914__ & ~new_new_n20069__;
  assign new_new_n20072__ = ~new_new_n20070__ & ~new_new_n20071__;
  assign new_new_n20073__ = new_new_n20068__ & new_new_n20072__;
  assign new_new_n20074__ = ~new_new_n20068__ & ~new_new_n20072__;
  assign new_new_n20075__ = ~new_new_n19901__ & ~new_new_n19902__;
  assign new_new_n20076__ = new_new_n19906__ & ~new_new_n20075__;
  assign new_new_n20077__ = ~new_new_n19906__ & new_new_n20075__;
  assign new_new_n20078__ = ~new_new_n20076__ & ~new_new_n20077__;
  assign new_new_n20079__ = ~new_new_n333__ & ~new_new_n15533__;
  assign new_new_n20080__ = new_new_n873__ & new_new_n15520__;
  assign new_new_n20081__ = ~new_new_n20079__ & ~new_new_n20080__;
  assign new_new_n20082__ = pi25 & new_new_n15524__;
  assign new_new_n20083__ = ~pi25 & ~new_new_n15524__;
  assign new_new_n20084__ = ~new_new_n110__ & ~new_new_n20082__;
  assign new_new_n20085__ = ~new_new_n20083__ & new_new_n20084__;
  assign new_new_n20086__ = new_new_n18913__ & new_new_n20085__;
  assign new_new_n20087__ = new_new_n801__ & ~new_new_n18914__;
  assign new_new_n20088__ = pi26 & ~new_new_n20087__;
  assign new_new_n20089__ = ~new_new_n20086__ & ~new_new_n20088__;
  assign new_new_n20090__ = new_new_n20081__ & ~new_new_n20089__;
  assign new_new_n20091__ = new_new_n801__ & new_new_n18923__;
  assign new_new_n20092__ = new_new_n20081__ & ~new_new_n20091__;
  assign new_new_n20093__ = ~pi26 & ~new_new_n20092__;
  assign new_new_n20094__ = ~new_new_n20090__ & ~new_new_n20093__;
  assign new_new_n20095__ = ~new_new_n19503__ & ~new_new_n19523__;
  assign new_new_n20096__ = new_new_n19520__ & ~new_new_n20095__;
  assign new_new_n20097__ = ~new_new_n19520__ & new_new_n20095__;
  assign new_new_n20098__ = ~new_new_n20096__ & ~new_new_n20097__;
  assign new_new_n20099__ = ~new_new_n19035__ & new_new_n19525__;
  assign new_new_n20100__ = new_new_n19035__ & new_new_n19520__;
  assign new_new_n20101__ = new_new_n19502__ & new_new_n19522__;
  assign new_new_n20102__ = ~new_new_n20100__ & ~new_new_n20101__;
  assign new_new_n20103__ = ~new_new_n19444__ & ~new_new_n20102__;
  assign new_new_n20104__ = new_new_n19035__ & new_new_n19502__;
  assign new_new_n20105__ = new_new_n19520__ & new_new_n19522__;
  assign new_new_n20106__ = ~new_new_n20104__ & ~new_new_n20105__;
  assign new_new_n20107__ = new_new_n20098__ & ~new_new_n20106__;
  assign new_new_n20108__ = ~new_new_n20099__ & ~new_new_n20103__;
  assign new_new_n20109__ = ~new_new_n20107__ & new_new_n20108__;
  assign new_new_n20110__ = new_new_n4815__ & new_new_n15572__;
  assign new_new_n20111__ = new_new_n15572__ & ~new_new_n19534__;
  assign new_new_n20112__ = new_new_n4215__ & ~new_new_n20111__;
  assign new_new_n20113__ = ~new_new_n15572__ & new_new_n19534__;
  assign new_new_n20114__ = ~new_new_n20111__ & ~new_new_n20113__;
  assign new_new_n20115__ = new_new_n4214__ & ~new_new_n20112__;
  assign new_new_n20116__ = ~new_new_n20114__ & new_new_n20115__;
  assign new_new_n20117__ = ~new_new_n4818__ & ~new_new_n15615__;
  assign new_new_n20118__ = new_new_n4212__ & new_new_n15564__;
  assign new_new_n20119__ = ~new_new_n20117__ & ~new_new_n20118__;
  assign new_new_n20120__ = ~new_new_n20110__ & new_new_n20119__;
  assign new_new_n20121__ = ~new_new_n20116__ & new_new_n20120__;
  assign new_new_n20122__ = ~new_new_n20109__ & ~new_new_n20121__;
  assign new_new_n20123__ = ~pi29 & new_new_n20121__;
  assign new_new_n20124__ = ~new_new_n20122__ & ~new_new_n20123__;
  assign new_new_n20125__ = new_new_n4815__ & new_new_n15560__;
  assign new_new_n20126__ = new_new_n4212__ & new_new_n15572__;
  assign new_new_n20127__ = ~new_new_n4818__ & new_new_n15564__;
  assign new_new_n20128__ = new_new_n4813__ & new_new_n18944__;
  assign new_new_n20129__ = ~new_new_n20126__ & ~new_new_n20127__;
  assign new_new_n20130__ = ~new_new_n20125__ & new_new_n20129__;
  assign new_new_n20131__ = ~new_new_n20128__ & new_new_n20130__;
  assign new_new_n20132__ = ~new_new_n20124__ & new_new_n20131__;
  assign new_new_n20133__ = ~new_new_n20109__ & new_new_n20121__;
  assign new_new_n20134__ = new_new_n4815__ & ~new_new_n15615__;
  assign new_new_n20135__ = ~new_new_n4818__ & ~new_new_n15638__;
  assign new_new_n20136__ = new_new_n4212__ & new_new_n15743__;
  assign new_new_n20137__ = ~new_new_n20135__ & ~new_new_n20136__;
  assign new_new_n20138__ = ~new_new_n20134__ & new_new_n20137__;
  assign new_new_n20139__ = new_new_n4214__ & new_new_n19005__;
  assign new_new_n20140__ = pi29 & ~new_new_n20139__;
  assign new_new_n20141__ = new_new_n4825__ & new_new_n19005__;
  assign new_new_n20142__ = ~new_new_n20140__ & ~new_new_n20141__;
  assign new_new_n20143__ = new_new_n20138__ & ~new_new_n20142__;
  assign new_new_n20144__ = ~pi29 & ~new_new_n20138__;
  assign new_new_n20145__ = ~new_new_n20143__ & ~new_new_n20144__;
  assign new_new_n20146__ = new_new_n4815__ & ~new_new_n15638__;
  assign new_new_n20147__ = new_new_n4212__ & ~new_new_n15582__;
  assign new_new_n20148__ = ~new_new_n4818__ & ~new_new_n15647__;
  assign new_new_n20149__ = new_new_n4813__ & new_new_n19487__;
  assign new_new_n20150__ = ~new_new_n20147__ & ~new_new_n20148__;
  assign new_new_n20151__ = ~new_new_n20146__ & new_new_n20150__;
  assign new_new_n20152__ = ~new_new_n20149__ & new_new_n20151__;
  assign new_new_n20153__ = ~pi29 & ~new_new_n20152__;
  assign new_new_n20154__ = pi29 & new_new_n20152__;
  assign new_new_n20155__ = ~new_new_n20153__ & ~new_new_n20154__;
  assign new_new_n20156__ = new_new_n4815__ & ~new_new_n15582__;
  assign new_new_n20157__ = ~new_new_n4818__ & ~new_new_n15710__;
  assign new_new_n20158__ = new_new_n4212__ & ~new_new_n15647__;
  assign new_new_n20159__ = ~new_new_n20157__ & ~new_new_n20158__;
  assign new_new_n20160__ = ~new_new_n20156__ & new_new_n20159__;
  assign new_new_n20161__ = new_new_n4214__ & ~new_new_n15736__;
  assign new_new_n20162__ = ~pi29 & ~new_new_n20161__;
  assign new_new_n20163__ = new_new_n5732__ & ~new_new_n15736__;
  assign new_new_n20164__ = ~new_new_n20162__ & ~new_new_n20163__;
  assign new_new_n20165__ = new_new_n20160__ & ~new_new_n20164__;
  assign new_new_n20166__ = pi29 & ~new_new_n20160__;
  assign new_new_n20167__ = ~new_new_n20165__ & ~new_new_n20166__;
  assign new_new_n20168__ = ~new_new_n19237__ & ~new_new_n19238__;
  assign new_new_n20169__ = new_new_n19316__ & ~new_new_n20168__;
  assign new_new_n20170__ = ~new_new_n19316__ & new_new_n20168__;
  assign new_new_n20171__ = ~new_new_n20169__ & ~new_new_n20170__;
  assign new_new_n20172__ = new_new_n4212__ & ~new_new_n15661__;
  assign new_new_n20173__ = ~new_new_n4818__ & new_new_n15668__;
  assign new_new_n20174__ = ~new_new_n20172__ & ~new_new_n20173__;
  assign new_new_n20175__ = new_new_n15661__ & ~new_new_n15668__;
  assign new_new_n20176__ = ~new_new_n15683__ & ~new_new_n20175__;
  assign new_new_n20177__ = ~new_new_n15643__ & ~new_new_n20176__;
  assign new_new_n20178__ = new_new_n4214__ & ~new_new_n20177__;
  assign new_new_n20179__ = pi29 & ~new_new_n20178__;
  assign new_new_n20180__ = pi28 & ~new_new_n15643__;
  assign new_new_n20181__ = ~pi28 & new_new_n15643__;
  assign new_new_n20182__ = ~new_new_n20180__ & ~new_new_n20181__;
  assign new_new_n20183__ = new_new_n4214__ & new_new_n20176__;
  assign new_new_n20184__ = ~new_new_n20182__ & new_new_n20183__;
  assign new_new_n20185__ = ~new_new_n20179__ & ~new_new_n20184__;
  assign new_new_n20186__ = new_new_n20174__ & ~new_new_n20185__;
  assign new_new_n20187__ = new_new_n15643__ & ~new_new_n20176__;
  assign new_new_n20188__ = new_new_n4214__ & new_new_n20187__;
  assign new_new_n20189__ = new_new_n20174__ & ~new_new_n20188__;
  assign new_new_n20190__ = ~pi29 & ~new_new_n20189__;
  assign new_new_n20191__ = ~new_new_n20186__ & ~new_new_n20190__;
  assign new_new_n20192__ = ~new_new_n4818__ & ~new_new_n15673__;
  assign new_new_n20193__ = new_new_n4212__ & new_new_n15668__;
  assign new_new_n20194__ = ~new_new_n20192__ & ~new_new_n20193__;
  assign new_new_n20195__ = new_new_n15668__ & new_new_n15673__;
  assign new_new_n20196__ = new_new_n15661__ & ~new_new_n20195__;
  assign new_new_n20197__ = new_new_n4214__ & ~new_new_n20196__;
  assign new_new_n20198__ = pi29 & ~new_new_n20197__;
  assign new_new_n20199__ = ~pi28 & new_new_n15661__;
  assign new_new_n20200__ = pi28 & ~new_new_n15661__;
  assign new_new_n20201__ = new_new_n4214__ & new_new_n20195__;
  assign new_new_n20202__ = ~new_new_n20199__ & new_new_n20201__;
  assign new_new_n20203__ = ~new_new_n20200__ & new_new_n20202__;
  assign new_new_n20204__ = ~new_new_n20198__ & ~new_new_n20203__;
  assign new_new_n20205__ = new_new_n20194__ & ~new_new_n20204__;
  assign new_new_n20206__ = ~new_new_n15661__ & ~new_new_n20195__;
  assign new_new_n20207__ = new_new_n4214__ & new_new_n20206__;
  assign new_new_n20208__ = new_new_n20194__ & ~new_new_n20207__;
  assign new_new_n20209__ = ~pi29 & ~new_new_n20208__;
  assign new_new_n20210__ = ~new_new_n20205__ & ~new_new_n20209__;
  assign new_new_n20211__ = ~new_new_n4209__ & new_new_n15668__;
  assign new_new_n20212__ = new_new_n15673__ & ~new_new_n20211__;
  assign new_new_n20213__ = ~pi28 & ~new_new_n15673__;
  assign new_new_n20214__ = new_new_n3889__ & ~new_new_n20213__;
  assign new_new_n20215__ = ~new_new_n68__ & ~new_new_n20214__;
  assign new_new_n20216__ = ~new_new_n20212__ & new_new_n20215__;
  assign new_new_n20217__ = pi29 & ~new_new_n20216__;
  assign new_new_n20218__ = ~new_new_n20210__ & new_new_n20217__;
  assign new_new_n20219__ = new_new_n765__ & ~new_new_n15673__;
  assign new_new_n20220__ = ~new_new_n20218__ & ~new_new_n20219__;
  assign new_new_n20221__ = ~new_new_n20191__ & ~new_new_n20220__;
  assign new_new_n20222__ = new_new_n4813__ & new_new_n15687__;
  assign new_new_n20223__ = ~new_new_n4818__ & ~new_new_n15661__;
  assign new_new_n20224__ = new_new_n4212__ & new_new_n15643__;
  assign new_new_n20225__ = ~new_new_n20223__ & ~new_new_n20224__;
  assign new_new_n20226__ = ~new_new_n20222__ & new_new_n20225__;
  assign new_new_n20227__ = new_new_n4214__ & new_new_n15656__;
  assign new_new_n20228__ = pi29 & ~new_new_n20227__;
  assign new_new_n20229__ = new_new_n5732__ & new_new_n15656__;
  assign new_new_n20230__ = ~new_new_n20228__ & ~new_new_n20229__;
  assign new_new_n20231__ = new_new_n20226__ & ~new_new_n20230__;
  assign new_new_n20232__ = ~pi29 & ~new_new_n20226__;
  assign new_new_n20233__ = ~new_new_n20231__ & ~new_new_n20232__;
  assign new_new_n20234__ = ~new_new_n20221__ & new_new_n20233__;
  assign new_new_n20235__ = new_new_n20221__ & ~new_new_n20233__;
  assign new_new_n20236__ = new_new_n4147__ & new_new_n15674__;
  assign new_new_n20237__ = ~new_new_n19312__ & ~new_new_n20236__;
  assign new_new_n20238__ = new_new_n19308__ & ~new_new_n20237__;
  assign new_new_n20239__ = ~new_new_n19314__ & ~new_new_n20238__;
  assign new_new_n20240__ = ~new_new_n20235__ & ~new_new_n20239__;
  assign new_new_n20241__ = ~new_new_n20234__ & ~new_new_n20240__;
  assign new_new_n20242__ = new_new_n4815__ & ~new_new_n15710__;
  assign new_new_n20243__ = ~new_new_n4818__ & new_new_n15643__;
  assign new_new_n20244__ = new_new_n4212__ & new_new_n15656__;
  assign new_new_n20245__ = ~new_new_n20243__ & ~new_new_n20244__;
  assign new_new_n20246__ = ~new_new_n20242__ & new_new_n20245__;
  assign new_new_n20247__ = new_new_n4214__ & ~new_new_n19466__;
  assign new_new_n20248__ = ~pi29 & ~new_new_n20247__;
  assign new_new_n20249__ = new_new_n5732__ & ~new_new_n19466__;
  assign new_new_n20250__ = ~new_new_n20248__ & ~new_new_n20249__;
  assign new_new_n20251__ = new_new_n20246__ & ~new_new_n20250__;
  assign new_new_n20252__ = pi29 & ~new_new_n20246__;
  assign new_new_n20253__ = ~new_new_n20251__ & ~new_new_n20252__;
  assign new_new_n20254__ = ~new_new_n20241__ & ~new_new_n20253__;
  assign new_new_n20255__ = new_new_n20241__ & new_new_n20253__;
  assign new_new_n20256__ = ~new_new_n20254__ & ~new_new_n20255__;
  assign new_new_n20257__ = ~new_new_n19268__ & ~new_new_n19269__;
  assign new_new_n20258__ = new_new_n19314__ & ~new_new_n20257__;
  assign new_new_n20259__ = ~new_new_n19314__ & new_new_n20257__;
  assign new_new_n20260__ = ~new_new_n20258__ & ~new_new_n20259__;
  assign new_new_n20261__ = new_new_n20256__ & new_new_n20260__;
  assign new_new_n20262__ = ~new_new_n20254__ & ~new_new_n20261__;
  assign new_new_n20263__ = new_new_n20171__ & new_new_n20262__;
  assign new_new_n20264__ = ~new_new_n20171__ & ~new_new_n20262__;
  assign new_new_n20265__ = new_new_n4813__ & ~new_new_n19118__;
  assign new_new_n20266__ = ~new_new_n4818__ & new_new_n15656__;
  assign new_new_n20267__ = new_new_n4212__ & ~new_new_n15710__;
  assign new_new_n20268__ = new_new_n4815__ & ~new_new_n15647__;
  assign new_new_n20269__ = ~new_new_n20266__ & ~new_new_n20267__;
  assign new_new_n20270__ = ~new_new_n20268__ & new_new_n20269__;
  assign new_new_n20271__ = ~new_new_n20265__ & new_new_n20270__;
  assign new_new_n20272__ = pi29 & ~new_new_n20271__;
  assign new_new_n20273__ = ~pi29 & new_new_n20271__;
  assign new_new_n20274__ = ~new_new_n20272__ & ~new_new_n20273__;
  assign new_new_n20275__ = ~new_new_n20264__ & new_new_n20274__;
  assign new_new_n20276__ = ~new_new_n20263__ & ~new_new_n20275__;
  assign new_new_n20277__ = new_new_n20167__ & ~new_new_n20276__;
  assign new_new_n20278__ = ~new_new_n20167__ & new_new_n20276__;
  assign new_new_n20279__ = ~new_new_n19357__ & ~new_new_n19378__;
  assign new_new_n20280__ = ~new_new_n19379__ & ~new_new_n20279__;
  assign new_new_n20281__ = ~new_new_n20278__ & ~new_new_n20280__;
  assign new_new_n20282__ = ~new_new_n20277__ & ~new_new_n20281__;
  assign new_new_n20283__ = new_new_n20155__ & new_new_n20282__;
  assign new_new_n20284__ = ~new_new_n19381__ & ~new_new_n19382__;
  assign new_new_n20285__ = ~new_new_n17499__ & ~new_new_n20284__;
  assign new_new_n20286__ = ~new_new_n20155__ & ~new_new_n20282__;
  assign new_new_n20287__ = new_new_n19419__ & ~new_new_n20284__;
  assign new_new_n20288__ = ~new_new_n19419__ & new_new_n20284__;
  assign new_new_n20289__ = ~new_new_n20287__ & ~new_new_n20288__;
  assign new_new_n20290__ = ~new_new_n20285__ & ~new_new_n20289__;
  assign new_new_n20291__ = ~new_new_n20286__ & new_new_n20290__;
  assign new_new_n20292__ = ~new_new_n20283__ & ~new_new_n20291__;
  assign new_new_n20293__ = ~new_new_n19177__ & ~new_new_n19178__;
  assign new_new_n20294__ = ~new_new_n19421__ & new_new_n20293__;
  assign new_new_n20295__ = new_new_n19421__ & ~new_new_n20293__;
  assign new_new_n20296__ = ~new_new_n20294__ & ~new_new_n20295__;
  assign new_new_n20297__ = ~new_new_n20292__ & ~new_new_n20296__;
  assign new_new_n20298__ = new_new_n20292__ & new_new_n20296__;
  assign new_new_n20299__ = new_new_n4813__ & new_new_n19494__;
  assign new_new_n20300__ = ~new_new_n4818__ & ~new_new_n15582__;
  assign new_new_n20301__ = new_new_n4212__ & ~new_new_n15638__;
  assign new_new_n20302__ = new_new_n4815__ & new_new_n15743__;
  assign new_new_n20303__ = ~new_new_n20300__ & ~new_new_n20301__;
  assign new_new_n20304__ = ~new_new_n20302__ & new_new_n20303__;
  assign new_new_n20305__ = ~new_new_n20299__ & new_new_n20304__;
  assign new_new_n20306__ = pi29 & ~new_new_n20305__;
  assign new_new_n20307__ = ~pi29 & new_new_n20305__;
  assign new_new_n20308__ = ~new_new_n20306__ & ~new_new_n20307__;
  assign new_new_n20309__ = ~new_new_n20298__ & ~new_new_n20308__;
  assign new_new_n20310__ = ~new_new_n20297__ & ~new_new_n20309__;
  assign new_new_n20311__ = new_new_n20145__ & ~new_new_n20310__;
  assign new_new_n20312__ = ~new_new_n20145__ & new_new_n20310__;
  assign new_new_n20313__ = ~new_new_n19424__ & ~new_new_n19425__;
  assign new_new_n20314__ = new_new_n19440__ & ~new_new_n20313__;
  assign new_new_n20315__ = ~new_new_n19440__ & new_new_n20313__;
  assign new_new_n20316__ = ~new_new_n20314__ & ~new_new_n20315__;
  assign new_new_n20317__ = ~new_new_n20312__ & ~new_new_n20316__;
  assign new_new_n20318__ = ~new_new_n20311__ & ~new_new_n20317__;
  assign new_new_n20319__ = ~new_new_n19074__ & ~new_new_n19075__;
  assign new_new_n20320__ = new_new_n19442__ & new_new_n20319__;
  assign new_new_n20321__ = ~new_new_n19442__ & ~new_new_n20319__;
  assign new_new_n20322__ = ~new_new_n20320__ & ~new_new_n20321__;
  assign new_new_n20323__ = new_new_n20318__ & ~new_new_n20322__;
  assign new_new_n20324__ = ~new_new_n20318__ & new_new_n20322__;
  assign new_new_n20325__ = new_new_n4815__ & new_new_n15564__;
  assign new_new_n20326__ = new_new_n4212__ & ~new_new_n15615__;
  assign new_new_n20327__ = ~new_new_n4818__ & new_new_n15743__;
  assign new_new_n20328__ = new_new_n4813__ & new_new_n18512__;
  assign new_new_n20329__ = ~new_new_n20326__ & ~new_new_n20327__;
  assign new_new_n20330__ = ~new_new_n20325__ & new_new_n20329__;
  assign new_new_n20331__ = ~new_new_n20328__ & new_new_n20330__;
  assign new_new_n20332__ = pi29 & ~new_new_n20331__;
  assign new_new_n20333__ = ~pi29 & new_new_n20331__;
  assign new_new_n20334__ = ~new_new_n20332__ & ~new_new_n20333__;
  assign new_new_n20335__ = ~new_new_n20324__ & new_new_n20334__;
  assign new_new_n20336__ = ~new_new_n20323__ & ~new_new_n20335__;
  assign new_new_n20337__ = new_new_n20121__ & ~new_new_n20336__;
  assign new_new_n20338__ = pi29 & ~new_new_n20337__;
  assign new_new_n20339__ = ~new_new_n20133__ & ~new_new_n20338__;
  assign new_new_n20340__ = ~new_new_n20131__ & ~new_new_n20339__;
  assign new_new_n20341__ = ~pi29 & new_new_n20131__;
  assign new_new_n20342__ = new_new_n20109__ & ~new_new_n20341__;
  assign new_new_n20343__ = new_new_n20336__ & ~new_new_n20342__;
  assign new_new_n20344__ = ~new_new_n20132__ & ~new_new_n20343__;
  assign new_new_n20345__ = ~new_new_n20340__ & new_new_n20344__;
  assign new_new_n20346__ = ~new_new_n20098__ & ~new_new_n20345__;
  assign new_new_n20347__ = pi29 & ~new_new_n20109__;
  assign new_new_n20348__ = pi29 & ~new_new_n20121__;
  assign new_new_n20349__ = ~new_new_n20133__ & ~new_new_n20348__;
  assign new_new_n20350__ = new_new_n20336__ & ~new_new_n20349__;
  assign new_new_n20351__ = ~new_new_n20347__ & ~new_new_n20350__;
  assign new_new_n20352__ = ~new_new_n20131__ & ~new_new_n20351__;
  assign new_new_n20353__ = ~pi29 & ~new_new_n20109__;
  assign new_new_n20354__ = ~new_new_n20124__ & new_new_n20336__;
  assign new_new_n20355__ = ~new_new_n20353__ & ~new_new_n20354__;
  assign new_new_n20356__ = new_new_n20131__ & ~new_new_n20355__;
  assign new_new_n20357__ = ~new_new_n20352__ & ~new_new_n20356__;
  assign new_new_n20358__ = ~new_new_n20346__ & new_new_n20357__;
  assign new_new_n20359__ = new_new_n20094__ & ~new_new_n20358__;
  assign new_new_n20360__ = new_new_n18981__ & ~new_new_n19526__;
  assign new_new_n20361__ = ~new_new_n18981__ & new_new_n19526__;
  assign new_new_n20362__ = ~new_new_n20360__ & ~new_new_n20361__;
  assign new_new_n20363__ = ~new_new_n18978__ & new_new_n20362__;
  assign new_new_n20364__ = ~new_new_n20094__ & new_new_n20358__;
  assign new_new_n20365__ = new_new_n18978__ & ~new_new_n20362__;
  assign new_new_n20366__ = ~new_new_n20363__ & ~new_new_n20365__;
  assign new_new_n20367__ = ~new_new_n20364__ & new_new_n20366__;
  assign new_new_n20368__ = ~new_new_n20359__ & ~new_new_n20367__;
  assign new_new_n20369__ = new_new_n20078__ & ~new_new_n20368__;
  assign new_new_n20370__ = ~new_new_n20078__ & new_new_n20368__;
  assign new_new_n20371__ = new_new_n5213__ & new_new_n15464__;
  assign new_new_n20372__ = new_new_n5183__ & ~new_new_n15471__;
  assign new_new_n20373__ = new_new_n5191__ & ~new_new_n15809__;
  assign new_new_n20374__ = new_new_n5215__ & new_new_n15819__;
  assign new_new_n20375__ = ~new_new_n20372__ & ~new_new_n20373__;
  assign new_new_n20376__ = ~new_new_n20371__ & new_new_n20375__;
  assign new_new_n20377__ = ~new_new_n20374__ & new_new_n20376__;
  assign new_new_n20378__ = ~new_new_n20369__ & ~new_new_n20370__;
  assign new_new_n20379__ = pi23 & ~new_new_n20378__;
  assign new_new_n20380__ = ~pi23 & new_new_n20378__;
  assign new_new_n20381__ = ~new_new_n20379__ & ~new_new_n20380__;
  assign new_new_n20382__ = new_new_n20377__ & new_new_n20381__;
  assign new_new_n20383__ = ~new_new_n20377__ & ~new_new_n20381__;
  assign new_new_n20384__ = ~new_new_n20382__ & ~new_new_n20383__;
  assign new_new_n20385__ = ~new_new_n20370__ & new_new_n20384__;
  assign new_new_n20386__ = ~new_new_n20369__ & ~new_new_n20385__;
  assign new_new_n20387__ = ~new_new_n20074__ & ~new_new_n20386__;
  assign new_new_n20388__ = ~new_new_n20073__ & ~new_new_n20387__;
  assign new_new_n20389__ = ~new_new_n20054__ & ~new_new_n20388__;
  assign new_new_n20390__ = ~new_new_n20053__ & ~new_new_n20389__;
  assign new_new_n20391__ = new_new_n20033__ & ~new_new_n20390__;
  assign new_new_n20392__ = ~new_new_n20033__ & new_new_n20390__;
  assign new_new_n20393__ = new_new_n6959__ & new_new_n16078__;
  assign new_new_n20394__ = new_new_n6964__ & ~new_new_n15321__;
  assign new_new_n20395__ = new_new_n6968__ & ~new_new_n15273__;
  assign new_new_n20396__ = new_new_n7935__ & new_new_n15285__;
  assign new_new_n20397__ = ~new_new_n20394__ & ~new_new_n20395__;
  assign new_new_n20398__ = ~new_new_n20396__ & new_new_n20397__;
  assign new_new_n20399__ = ~new_new_n20393__ & new_new_n20398__;
  assign new_new_n20400__ = pi17 & ~new_new_n20399__;
  assign new_new_n20401__ = ~pi17 & new_new_n20399__;
  assign new_new_n20402__ = ~new_new_n20400__ & ~new_new_n20401__;
  assign new_new_n20403__ = ~new_new_n20392__ & ~new_new_n20402__;
  assign new_new_n20404__ = ~new_new_n20391__ & ~new_new_n20403__;
  assign new_new_n20405__ = ~new_new_n20029__ & new_new_n20404__;
  assign new_new_n20406__ = new_new_n20029__ & ~new_new_n20404__;
  assign new_new_n20407__ = ~new_new_n19949__ & ~new_new_n19950__;
  assign new_new_n20408__ = new_new_n19952__ & new_new_n20407__;
  assign new_new_n20409__ = ~new_new_n19952__ & ~new_new_n20407__;
  assign new_new_n20410__ = ~new_new_n20408__ & ~new_new_n20409__;
  assign new_new_n20411__ = ~new_new_n20406__ & ~new_new_n20410__;
  assign new_new_n20412__ = ~new_new_n20405__ & ~new_new_n20411__;
  assign new_new_n20413__ = ~new_new_n20011__ & ~new_new_n20412__;
  assign new_new_n20414__ = new_new_n20011__ & new_new_n20412__;
  assign new_new_n20415__ = new_new_n6985__ & new_new_n15237__;
  assign new_new_n20416__ = new_new_n6991__ & new_new_n15244__;
  assign new_new_n20417__ = ~new_new_n20415__ & ~new_new_n20416__;
  assign new_new_n20418__ = new_new_n6994__ & new_new_n17974__;
  assign new_new_n20419__ = new_new_n20417__ & ~new_new_n20418__;
  assign new_new_n20420__ = ~pi14 & ~new_new_n20419__;
  assign new_new_n20421__ = new_new_n6994__ & ~new_new_n17978__;
  assign new_new_n20422__ = pi14 & new_new_n20417__;
  assign new_new_n20423__ = ~new_new_n20421__ & new_new_n20422__;
  assign new_new_n20424__ = ~pi13 & ~new_new_n17983__;
  assign new_new_n20425__ = pi13 & ~new_new_n17981__;
  assign new_new_n20426__ = new_new_n6994__ & ~new_new_n20424__;
  assign new_new_n20427__ = ~new_new_n20425__ & new_new_n20426__;
  assign new_new_n20428__ = ~new_new_n20420__ & ~new_new_n20423__;
  assign new_new_n20429__ = ~new_new_n20427__ & new_new_n20428__;
  assign new_new_n20430__ = ~new_new_n20414__ & ~new_new_n20429__;
  assign new_new_n20431__ = ~new_new_n20413__ & ~new_new_n20430__;
  assign new_new_n20432__ = ~new_new_n20007__ & ~new_new_n20431__;
  assign new_new_n20433__ = ~new_new_n20006__ & ~new_new_n20432__;
  assign new_new_n20434__ = ~new_new_n20405__ & ~new_new_n20406__;
  assign new_new_n20435__ = ~new_new_n20410__ & new_new_n20434__;
  assign new_new_n20436__ = new_new_n20410__ & ~new_new_n20434__;
  assign new_new_n20437__ = ~new_new_n20435__ & ~new_new_n20436__;
  assign new_new_n20438__ = ~new_new_n8479__ & new_new_n15905__;
  assign new_new_n20439__ = new_new_n8474__ & ~new_new_n15998__;
  assign new_new_n20440__ = ~new_new_n8468__ & new_new_n16051__;
  assign new_new_n20441__ = new_new_n8469__ & ~new_new_n16056__;
  assign new_new_n20442__ = ~new_new_n20440__ & new_new_n20441__;
  assign new_new_n20443__ = ~new_new_n20438__ & ~new_new_n20439__;
  assign new_new_n20444__ = ~new_new_n20442__ & new_new_n20443__;
  assign new_new_n20445__ = new_new_n6985__ & ~new_new_n15248__;
  assign new_new_n20446__ = new_new_n6991__ & ~new_new_n15314__;
  assign new_new_n20447__ = ~new_new_n20445__ & ~new_new_n20446__;
  assign new_new_n20448__ = new_new_n6994__ & new_new_n15244__;
  assign new_new_n20449__ = new_new_n16378__ & new_new_n20448__;
  assign new_new_n20450__ = new_new_n20447__ & ~new_new_n20449__;
  assign new_new_n20451__ = pi14 & ~new_new_n20450__;
  assign new_new_n20452__ = ~pi13 & new_new_n15244__;
  assign new_new_n20453__ = ~new_new_n15244__ & ~new_new_n16378__;
  assign new_new_n20454__ = new_new_n6994__ & ~new_new_n20453__;
  assign new_new_n20455__ = pi13 & new_new_n16378__;
  assign new_new_n20456__ = ~new_new_n20452__ & ~new_new_n20455__;
  assign new_new_n20457__ = new_new_n20454__ & new_new_n20456__;
  assign new_new_n20458__ = ~pi14 & new_new_n20447__;
  assign new_new_n20459__ = ~new_new_n20454__ & new_new_n20458__;
  assign new_new_n20460__ = ~new_new_n20451__ & ~new_new_n20457__;
  assign new_new_n20461__ = ~new_new_n20459__ & new_new_n20460__;
  assign new_new_n20462__ = ~new_new_n20391__ & ~new_new_n20392__;
  assign new_new_n20463__ = ~new_new_n20402__ & new_new_n20462__;
  assign new_new_n20464__ = new_new_n20402__ & ~new_new_n20462__;
  assign new_new_n20465__ = ~new_new_n20463__ & ~new_new_n20464__;
  assign new_new_n20466__ = ~new_new_n20461__ & new_new_n20465__;
  assign new_new_n20467__ = new_new_n20461__ & ~new_new_n20465__;
  assign new_new_n20468__ = new_new_n6968__ & ~new_new_n15349__;
  assign new_new_n20469__ = new_new_n6964__ & ~new_new_n15398__;
  assign new_new_n20470__ = new_new_n7935__ & ~new_new_n15321__;
  assign new_new_n20471__ = ~new_new_n20468__ & ~new_new_n20469__;
  assign new_new_n20472__ = ~new_new_n20470__ & new_new_n20471__;
  assign new_new_n20473__ = new_new_n6958__ & new_new_n16458__;
  assign new_new_n20474__ = pi17 & ~new_new_n20473__;
  assign new_new_n20475__ = new_new_n7942__ & new_new_n16458__;
  assign new_new_n20476__ = ~new_new_n20474__ & ~new_new_n20475__;
  assign new_new_n20477__ = new_new_n20472__ & ~new_new_n20476__;
  assign new_new_n20478__ = ~pi17 & ~new_new_n20472__;
  assign new_new_n20479__ = ~new_new_n20477__ & ~new_new_n20478__;
  assign new_new_n20480__ = new_new_n6629__ & ~new_new_n15432__;
  assign new_new_n20481__ = ~new_new_n6625__ & ~new_new_n15439__;
  assign new_new_n20482__ = new_new_n6634__ & ~new_new_n15362__;
  assign new_new_n20483__ = ~new_new_n20480__ & ~new_new_n20481__;
  assign new_new_n20484__ = ~new_new_n20482__ & new_new_n20483__;
  assign new_new_n20485__ = new_new_n6631__ & new_new_n16771__;
  assign new_new_n20486__ = ~pi20 & ~new_new_n20485__;
  assign new_new_n20487__ = new_new_n7015__ & new_new_n16771__;
  assign new_new_n20488__ = ~new_new_n20486__ & ~new_new_n20487__;
  assign new_new_n20489__ = new_new_n20484__ & ~new_new_n20488__;
  assign new_new_n20490__ = pi20 & ~new_new_n20484__;
  assign new_new_n20491__ = ~new_new_n20489__ & ~new_new_n20490__;
  assign new_new_n20492__ = new_new_n20384__ & new_new_n20491__;
  assign new_new_n20493__ = ~new_new_n20384__ & ~new_new_n20491__;
  assign new_new_n20494__ = ~new_new_n20109__ & ~new_new_n20131__;
  assign new_new_n20495__ = new_new_n20109__ & new_new_n20131__;
  assign new_new_n20496__ = ~new_new_n20494__ & ~new_new_n20495__;
  assign new_new_n20497__ = new_new_n20098__ & ~new_new_n20336__;
  assign new_new_n20498__ = ~new_new_n20098__ & new_new_n20336__;
  assign new_new_n20499__ = ~new_new_n20497__ & ~new_new_n20498__;
  assign new_new_n20500__ = ~new_new_n20121__ & new_new_n20499__;
  assign new_new_n20501__ = ~pi29 & new_new_n20497__;
  assign new_new_n20502__ = pi29 & new_new_n20498__;
  assign new_new_n20503__ = ~new_new_n20496__ & ~new_new_n20501__;
  assign new_new_n20504__ = ~new_new_n20502__ & new_new_n20503__;
  assign new_new_n20505__ = ~new_new_n20500__ & new_new_n20504__;
  assign new_new_n20506__ = pi29 & new_new_n20497__;
  assign new_new_n20507__ = new_new_n20121__ & new_new_n20499__;
  assign new_new_n20508__ = ~pi29 & new_new_n20498__;
  assign new_new_n20509__ = new_new_n20496__ & ~new_new_n20506__;
  assign new_new_n20510__ = ~new_new_n20508__ & new_new_n20509__;
  assign new_new_n20511__ = ~new_new_n20507__ & new_new_n20510__;
  assign new_new_n20512__ = ~new_new_n20505__ & ~new_new_n20511__;
  assign new_new_n20513__ = ~new_new_n20123__ & ~new_new_n20348__;
  assign new_new_n20514__ = new_new_n20499__ & new_new_n20513__;
  assign new_new_n20515__ = ~new_new_n20499__ & ~new_new_n20513__;
  assign new_new_n20516__ = ~new_new_n20514__ & ~new_new_n20515__;
  assign new_new_n20517__ = ~new_new_n333__ & ~new_new_n15615__;
  assign new_new_n20518__ = new_new_n873__ & new_new_n15564__;
  assign new_new_n20519__ = ~new_new_n20517__ & ~new_new_n20518__;
  assign new_new_n20520__ = new_new_n801__ & new_new_n20111__;
  assign new_new_n20521__ = new_new_n20519__ & ~new_new_n20520__;
  assign new_new_n20522__ = pi26 & ~new_new_n20521__;
  assign new_new_n20523__ = ~pi25 & new_new_n15572__;
  assign new_new_n20524__ = pi25 & ~new_new_n15572__;
  assign new_new_n20525__ = ~new_new_n110__ & ~new_new_n20523__;
  assign new_new_n20526__ = ~new_new_n20524__ & new_new_n20525__;
  assign new_new_n20527__ = new_new_n19534__ & new_new_n20526__;
  assign new_new_n20528__ = ~new_new_n15572__ & ~new_new_n19534__;
  assign new_new_n20529__ = new_new_n801__ & ~new_new_n20528__;
  assign new_new_n20530__ = ~pi26 & ~new_new_n20529__;
  assign new_new_n20531__ = ~new_new_n20527__ & ~new_new_n20530__;
  assign new_new_n20532__ = new_new_n20519__ & ~new_new_n20531__;
  assign new_new_n20533__ = ~new_new_n20522__ & ~new_new_n20532__;
  assign new_new_n20534__ = ~new_new_n20297__ & ~new_new_n20298__;
  assign new_new_n20535__ = ~new_new_n20308__ & new_new_n20534__;
  assign new_new_n20536__ = new_new_n20308__ & ~new_new_n20534__;
  assign new_new_n20537__ = ~new_new_n20535__ & ~new_new_n20536__;
  assign new_new_n20538__ = new_new_n20533__ & ~new_new_n20537__;
  assign new_new_n20539__ = ~new_new_n20533__ & new_new_n20537__;
  assign new_new_n20540__ = ~new_new_n20283__ & new_new_n20291__;
  assign new_new_n20541__ = ~new_new_n20283__ & ~new_new_n20286__;
  assign new_new_n20542__ = new_new_n20289__ & ~new_new_n20541__;
  assign new_new_n20543__ = ~new_new_n20540__ & ~new_new_n20542__;
  assign new_new_n20544__ = new_new_n3311__ & ~new_new_n15615__;
  assign new_new_n20545__ = ~new_new_n333__ & ~new_new_n15638__;
  assign new_new_n20546__ = new_new_n873__ & new_new_n15743__;
  assign new_new_n20547__ = ~new_new_n20545__ & ~new_new_n20546__;
  assign new_new_n20548__ = ~new_new_n20544__ & new_new_n20547__;
  assign new_new_n20549__ = ~pi26 & ~new_new_n20548__;
  assign new_new_n20550__ = new_new_n512__ & new_new_n19005__;
  assign new_new_n20551__ = new_new_n801__ & new_new_n19005__;
  assign new_new_n20552__ = pi26 & ~new_new_n20551__;
  assign new_new_n20553__ = ~new_new_n20550__ & ~new_new_n20552__;
  assign new_new_n20554__ = new_new_n20548__ & ~new_new_n20553__;
  assign new_new_n20555__ = ~new_new_n20549__ & ~new_new_n20554__;
  assign new_new_n20556__ = ~new_new_n20263__ & ~new_new_n20264__;
  assign new_new_n20557__ = new_new_n20274__ & new_new_n20556__;
  assign new_new_n20558__ = ~new_new_n20274__ & ~new_new_n20556__;
  assign new_new_n20559__ = ~new_new_n20557__ & ~new_new_n20558__;
  assign new_new_n20560__ = new_new_n3311__ & ~new_new_n15638__;
  assign new_new_n20561__ = ~new_new_n333__ & ~new_new_n15647__;
  assign new_new_n20562__ = new_new_n873__ & ~new_new_n15582__;
  assign new_new_n20563__ = ~new_new_n20561__ & ~new_new_n20562__;
  assign new_new_n20564__ = ~new_new_n20560__ & new_new_n20563__;
  assign new_new_n20565__ = ~pi26 & ~new_new_n20564__;
  assign new_new_n20566__ = new_new_n512__ & new_new_n19487__;
  assign new_new_n20567__ = new_new_n801__ & new_new_n19487__;
  assign new_new_n20568__ = pi26 & ~new_new_n20567__;
  assign new_new_n20569__ = ~new_new_n20566__ & ~new_new_n20568__;
  assign new_new_n20570__ = new_new_n20564__ & ~new_new_n20569__;
  assign new_new_n20571__ = ~new_new_n20565__ & ~new_new_n20570__;
  assign new_new_n20572__ = ~new_new_n4900__ & ~new_new_n15736__;
  assign new_new_n20573__ = ~new_new_n333__ & ~new_new_n15710__;
  assign new_new_n20574__ = new_new_n873__ & ~new_new_n15647__;
  assign new_new_n20575__ = ~new_new_n20573__ & ~new_new_n20574__;
  assign new_new_n20576__ = ~new_new_n20572__ & new_new_n20575__;
  assign new_new_n20577__ = pi26 & ~new_new_n20576__;
  assign new_new_n20578__ = new_new_n512__ & ~new_new_n15582__;
  assign new_new_n20579__ = new_new_n801__ & ~new_new_n15582__;
  assign new_new_n20580__ = ~pi26 & ~new_new_n20579__;
  assign new_new_n20581__ = ~new_new_n20578__ & ~new_new_n20580__;
  assign new_new_n20582__ = new_new_n20576__ & ~new_new_n20581__;
  assign new_new_n20583__ = ~new_new_n20577__ & ~new_new_n20582__;
  assign new_new_n20584__ = ~new_new_n4900__ & ~new_new_n19118__;
  assign new_new_n20585__ = new_new_n873__ & ~new_new_n15710__;
  assign new_new_n20586__ = ~new_new_n333__ & new_new_n15656__;
  assign new_new_n20587__ = new_new_n3311__ & ~new_new_n15647__;
  assign new_new_n20588__ = ~new_new_n20585__ & ~new_new_n20586__;
  assign new_new_n20589__ = ~new_new_n20587__ & new_new_n20588__;
  assign new_new_n20590__ = ~new_new_n20584__ & new_new_n20589__;
  assign new_new_n20591__ = pi26 & ~new_new_n20590__;
  assign new_new_n20592__ = ~pi26 & new_new_n20590__;
  assign new_new_n20593__ = ~new_new_n20591__ & ~new_new_n20592__;
  assign new_new_n20594__ = new_new_n20191__ & new_new_n20220__;
  assign new_new_n20595__ = ~new_new_n20221__ & ~new_new_n20594__;
  assign new_new_n20596__ = ~pi30 & ~new_new_n15673__;
  assign new_new_n20597__ = new_new_n20218__ & new_new_n20596__;
  assign new_new_n20598__ = ~new_new_n20595__ & ~new_new_n20597__;
  assign new_new_n20599__ = new_new_n20593__ & ~new_new_n20598__;
  assign new_new_n20600__ = new_new_n3311__ & ~new_new_n15710__;
  assign new_new_n20601__ = ~new_new_n333__ & new_new_n15643__;
  assign new_new_n20602__ = new_new_n873__ & new_new_n15656__;
  assign new_new_n20603__ = ~new_new_n20601__ & ~new_new_n20602__;
  assign new_new_n20604__ = ~new_new_n20600__ & new_new_n20603__;
  assign new_new_n20605__ = pi26 & ~new_new_n20604__;
  assign new_new_n20606__ = new_new_n4898__ & ~new_new_n19466__;
  assign new_new_n20607__ = new_new_n801__ & ~new_new_n19466__;
  assign new_new_n20608__ = ~pi26 & ~new_new_n20607__;
  assign new_new_n20609__ = ~new_new_n20606__ & ~new_new_n20608__;
  assign new_new_n20610__ = new_new_n20604__ & ~new_new_n20609__;
  assign new_new_n20611__ = ~new_new_n20605__ & ~new_new_n20610__;
  assign new_new_n20612__ = new_new_n20210__ & new_new_n20595__;
  assign new_new_n20613__ = ~new_new_n20593__ & ~new_new_n20612__;
  assign new_new_n20614__ = ~new_new_n4900__ & new_new_n15687__;
  assign new_new_n20615__ = ~new_new_n333__ & ~new_new_n15661__;
  assign new_new_n20616__ = new_new_n873__ & new_new_n15643__;
  assign new_new_n20617__ = ~new_new_n20615__ & ~new_new_n20616__;
  assign new_new_n20618__ = ~new_new_n20614__ & new_new_n20617__;
  assign new_new_n20619__ = pi26 & ~new_new_n20618__;
  assign new_new_n20620__ = new_new_n512__ & new_new_n15656__;
  assign new_new_n20621__ = new_new_n801__ & new_new_n15656__;
  assign new_new_n20622__ = ~pi26 & ~new_new_n20621__;
  assign new_new_n20623__ = ~new_new_n20620__ & ~new_new_n20622__;
  assign new_new_n20624__ = new_new_n20618__ & ~new_new_n20623__;
  assign new_new_n20625__ = ~new_new_n20619__ & ~new_new_n20624__;
  assign new_new_n20626__ = new_new_n4214__ & ~new_new_n15673__;
  assign new_new_n20627__ = new_new_n873__ & ~new_new_n15673__;
  assign new_new_n20628__ = ~new_new_n15668__ & new_new_n15673__;
  assign new_new_n20629__ = new_new_n801__ & ~new_new_n20628__;
  assign new_new_n20630__ = ~new_new_n20627__ & ~new_new_n20629__;
  assign new_new_n20631__ = ~new_new_n333__ & ~new_new_n15673__;
  assign new_new_n20632__ = new_new_n873__ & new_new_n15668__;
  assign new_new_n20633__ = ~new_new_n447__ & new_new_n20195__;
  assign new_new_n20634__ = new_new_n15661__ & ~new_new_n20633__;
  assign new_new_n20635__ = ~new_new_n15661__ & new_new_n20633__;
  assign new_new_n20636__ = new_new_n801__ & ~new_new_n20634__;
  assign new_new_n20637__ = ~new_new_n20635__ & new_new_n20636__;
  assign new_new_n20638__ = ~new_new_n20631__ & ~new_new_n20632__;
  assign new_new_n20639__ = ~new_new_n20637__ & new_new_n20638__;
  assign new_new_n20640__ = pi26 & new_new_n20630__;
  assign new_new_n20641__ = new_new_n20639__ & new_new_n20640__;
  assign new_new_n20642__ = ~new_new_n20626__ & ~new_new_n20641__;
  assign new_new_n20643__ = new_new_n3311__ & new_new_n15643__;
  assign new_new_n20644__ = new_new_n15664__ & ~new_new_n15680__;
  assign new_new_n20645__ = ~new_new_n15664__ & new_new_n15680__;
  assign new_new_n20646__ = ~new_new_n20644__ & ~new_new_n20645__;
  assign new_new_n20647__ = ~new_new_n4900__ & new_new_n20646__;
  assign new_new_n20648__ = new_new_n873__ & ~new_new_n15661__;
  assign new_new_n20649__ = ~new_new_n20643__ & ~new_new_n20648__;
  assign new_new_n20650__ = ~new_new_n20647__ & new_new_n20649__;
  assign new_new_n20651__ = new_new_n303__ & new_new_n15668__;
  assign new_new_n20652__ = pi26 & ~new_new_n20651__;
  assign new_new_n20653__ = new_new_n145__ & new_new_n15668__;
  assign new_new_n20654__ = ~pi26 & ~new_new_n20653__;
  assign new_new_n20655__ = pi23 & ~new_new_n20654__;
  assign new_new_n20656__ = ~new_new_n20652__ & ~new_new_n20655__;
  assign new_new_n20657__ = new_new_n20650__ & ~new_new_n20656__;
  assign new_new_n20658__ = ~pi26 & ~new_new_n20650__;
  assign new_new_n20659__ = ~new_new_n20657__ & ~new_new_n20658__;
  assign new_new_n20660__ = ~new_new_n20642__ & ~new_new_n20659__;
  assign new_new_n20661__ = new_new_n4210__ & new_new_n15674__;
  assign new_new_n20662__ = ~new_new_n4214__ & new_new_n20195__;
  assign new_new_n20663__ = new_new_n4211__ & ~new_new_n20211__;
  assign new_new_n20664__ = ~new_new_n66__ & ~new_new_n20628__;
  assign new_new_n20665__ = ~new_new_n20661__ & new_new_n20664__;
  assign new_new_n20666__ = ~new_new_n20662__ & ~new_new_n20663__;
  assign new_new_n20667__ = new_new_n20665__ & new_new_n20666__;
  assign new_new_n20668__ = ~new_new_n20660__ & ~new_new_n20667__;
  assign new_new_n20669__ = new_new_n20625__ & ~new_new_n20668__;
  assign new_new_n20670__ = new_new_n20626__ & new_new_n20667__;
  assign new_new_n20671__ = ~new_new_n20659__ & new_new_n20670__;
  assign new_new_n20672__ = ~new_new_n20669__ & ~new_new_n20671__;
  assign new_new_n20673__ = new_new_n20611__ & ~new_new_n20672__;
  assign new_new_n20674__ = ~new_new_n20613__ & new_new_n20673__;
  assign new_new_n20675__ = ~new_new_n20593__ & new_new_n20598__;
  assign new_new_n20676__ = ~new_new_n20217__ & ~new_new_n20672__;
  assign new_new_n20677__ = ~new_new_n20611__ & ~new_new_n20676__;
  assign new_new_n20678__ = ~new_new_n20210__ & ~new_new_n20217__;
  assign new_new_n20679__ = new_new_n20210__ & new_new_n20217__;
  assign new_new_n20680__ = ~new_new_n20678__ & ~new_new_n20679__;
  assign new_new_n20681__ = ~new_new_n20677__ & ~new_new_n20680__;
  assign new_new_n20682__ = ~new_new_n20675__ & new_new_n20681__;
  assign new_new_n20683__ = ~new_new_n20599__ & ~new_new_n20674__;
  assign new_new_n20684__ = ~new_new_n20682__ & new_new_n20683__;
  assign new_new_n20685__ = new_new_n20583__ & ~new_new_n20684__;
  assign new_new_n20686__ = ~new_new_n20583__ & new_new_n20684__;
  assign new_new_n20687__ = ~new_new_n20234__ & ~new_new_n20235__;
  assign new_new_n20688__ = new_new_n20239__ & new_new_n20687__;
  assign new_new_n20689__ = ~new_new_n20239__ & ~new_new_n20687__;
  assign new_new_n20690__ = ~new_new_n20688__ & ~new_new_n20689__;
  assign new_new_n20691__ = ~new_new_n20686__ & new_new_n20690__;
  assign new_new_n20692__ = ~new_new_n20685__ & ~new_new_n20691__;
  assign new_new_n20693__ = ~new_new_n20571__ & ~new_new_n20692__;
  assign new_new_n20694__ = new_new_n20571__ & new_new_n20692__;
  assign new_new_n20695__ = ~new_new_n19314__ & new_new_n20256__;
  assign new_new_n20696__ = new_new_n19314__ & ~new_new_n20256__;
  assign new_new_n20697__ = ~new_new_n20695__ & ~new_new_n20696__;
  assign new_new_n20698__ = ~new_new_n17601__ & new_new_n19250__;
  assign new_new_n20699__ = ~new_new_n20257__ & ~new_new_n20698__;
  assign new_new_n20700__ = ~new_new_n20697__ & new_new_n20699__;
  assign new_new_n20701__ = new_new_n20257__ & new_new_n20697__;
  assign new_new_n20702__ = ~new_new_n20700__ & ~new_new_n20701__;
  assign new_new_n20703__ = ~new_new_n20694__ & ~new_new_n20702__;
  assign new_new_n20704__ = ~new_new_n20693__ & ~new_new_n20703__;
  assign new_new_n20705__ = ~new_new_n20559__ & new_new_n20704__;
  assign new_new_n20706__ = new_new_n20559__ & ~new_new_n20704__;
  assign new_new_n20707__ = ~new_new_n4900__ & new_new_n19494__;
  assign new_new_n20708__ = ~new_new_n333__ & ~new_new_n15582__;
  assign new_new_n20709__ = new_new_n873__ & ~new_new_n15638__;
  assign new_new_n20710__ = new_new_n3311__ & new_new_n15743__;
  assign new_new_n20711__ = ~new_new_n20708__ & ~new_new_n20709__;
  assign new_new_n20712__ = ~new_new_n20710__ & new_new_n20711__;
  assign new_new_n20713__ = ~new_new_n20707__ & new_new_n20712__;
  assign new_new_n20714__ = pi26 & ~new_new_n20713__;
  assign new_new_n20715__ = ~pi26 & new_new_n20713__;
  assign new_new_n20716__ = ~new_new_n20714__ & ~new_new_n20715__;
  assign new_new_n20717__ = ~new_new_n20706__ & ~new_new_n20716__;
  assign new_new_n20718__ = ~new_new_n20705__ & ~new_new_n20717__;
  assign new_new_n20719__ = new_new_n20555__ & ~new_new_n20718__;
  assign new_new_n20720__ = ~new_new_n20555__ & new_new_n20718__;
  assign new_new_n20721__ = new_new_n20167__ & ~new_new_n20280__;
  assign new_new_n20722__ = ~new_new_n20167__ & new_new_n20280__;
  assign new_new_n20723__ = ~new_new_n20721__ & ~new_new_n20722__;
  assign new_new_n20724__ = new_new_n20276__ & new_new_n20723__;
  assign new_new_n20725__ = ~new_new_n20276__ & ~new_new_n20723__;
  assign new_new_n20726__ = ~new_new_n20724__ & ~new_new_n20725__;
  assign new_new_n20727__ = ~new_new_n20720__ & new_new_n20726__;
  assign new_new_n20728__ = ~new_new_n20719__ & ~new_new_n20727__;
  assign new_new_n20729__ = new_new_n20543__ & ~new_new_n20728__;
  assign new_new_n20730__ = ~new_new_n20543__ & new_new_n20728__;
  assign new_new_n20731__ = ~new_new_n333__ & new_new_n15743__;
  assign new_new_n20732__ = new_new_n873__ & ~new_new_n15615__;
  assign new_new_n20733__ = ~new_new_n20731__ & ~new_new_n20732__;
  assign new_new_n20734__ = ~new_new_n110__ & new_new_n15564__;
  assign new_new_n20735__ = new_new_n18512__ & new_new_n20734__;
  assign new_new_n20736__ = new_new_n20733__ & ~new_new_n20735__;
  assign new_new_n20737__ = pi26 & ~new_new_n20736__;
  assign new_new_n20738__ = ~new_new_n15564__ & ~new_new_n18512__;
  assign new_new_n20739__ = new_new_n801__ & ~new_new_n20738__;
  assign new_new_n20740__ = ~pi26 & ~new_new_n20739__;
  assign new_new_n20741__ = ~new_new_n15564__ & new_new_n18512__;
  assign new_new_n20742__ = ~pi25 & ~new_new_n20741__;
  assign new_new_n20743__ = new_new_n15564__ & ~new_new_n18512__;
  assign new_new_n20744__ = pi25 & ~new_new_n20743__;
  assign new_new_n20745__ = ~new_new_n110__ & ~new_new_n20742__;
  assign new_new_n20746__ = ~new_new_n20744__ & new_new_n20745__;
  assign new_new_n20747__ = ~new_new_n20740__ & ~new_new_n20746__;
  assign new_new_n20748__ = new_new_n20733__ & ~new_new_n20747__;
  assign new_new_n20749__ = ~new_new_n20737__ & ~new_new_n20748__;
  assign new_new_n20750__ = ~new_new_n20730__ & ~new_new_n20749__;
  assign new_new_n20751__ = ~new_new_n20729__ & ~new_new_n20750__;
  assign new_new_n20752__ = ~new_new_n20539__ & new_new_n20751__;
  assign new_new_n20753__ = ~new_new_n20538__ & ~new_new_n20752__;
  assign new_new_n20754__ = ~new_new_n20311__ & ~new_new_n20312__;
  assign new_new_n20755__ = ~new_new_n20316__ & new_new_n20754__;
  assign new_new_n20756__ = new_new_n20316__ & ~new_new_n20754__;
  assign new_new_n20757__ = ~new_new_n20755__ & ~new_new_n20756__;
  assign new_new_n20758__ = ~new_new_n20753__ & ~new_new_n20757__;
  assign new_new_n20759__ = new_new_n20753__ & new_new_n20757__;
  assign new_new_n20760__ = new_new_n3311__ & new_new_n15560__;
  assign new_new_n20761__ = new_new_n873__ & new_new_n15572__;
  assign new_new_n20762__ = ~new_new_n333__ & new_new_n15564__;
  assign new_new_n20763__ = ~new_new_n4900__ & new_new_n18944__;
  assign new_new_n20764__ = ~new_new_n20761__ & ~new_new_n20762__;
  assign new_new_n20765__ = ~new_new_n20760__ & new_new_n20764__;
  assign new_new_n20766__ = ~new_new_n20763__ & new_new_n20765__;
  assign new_new_n20767__ = pi26 & ~new_new_n20766__;
  assign new_new_n20768__ = ~pi26 & new_new_n20766__;
  assign new_new_n20769__ = ~new_new_n20767__ & ~new_new_n20768__;
  assign new_new_n20770__ = ~new_new_n20759__ & new_new_n20769__;
  assign new_new_n20771__ = ~new_new_n20758__ & ~new_new_n20770__;
  assign new_new_n20772__ = ~new_new_n20323__ & ~new_new_n20324__;
  assign new_new_n20773__ = ~new_new_n20334__ & ~new_new_n20772__;
  assign new_new_n20774__ = new_new_n20334__ & new_new_n20772__;
  assign new_new_n20775__ = ~new_new_n20773__ & ~new_new_n20774__;
  assign new_new_n20776__ = ~new_new_n20771__ & new_new_n20775__;
  assign new_new_n20777__ = new_new_n20771__ & ~new_new_n20775__;
  assign new_new_n20778__ = new_new_n873__ & new_new_n15560__;
  assign new_new_n20779__ = new_new_n3311__ & new_new_n15767__;
  assign new_new_n20780__ = ~new_new_n333__ & new_new_n15572__;
  assign new_new_n20781__ = ~new_new_n4900__ & ~new_new_n18454__;
  assign new_new_n20782__ = ~new_new_n20779__ & ~new_new_n20780__;
  assign new_new_n20783__ = ~new_new_n20778__ & new_new_n20782__;
  assign new_new_n20784__ = ~new_new_n20781__ & new_new_n20783__;
  assign new_new_n20785__ = pi26 & ~new_new_n20784__;
  assign new_new_n20786__ = ~pi26 & new_new_n20784__;
  assign new_new_n20787__ = ~new_new_n20785__ & ~new_new_n20786__;
  assign new_new_n20788__ = ~new_new_n20777__ & new_new_n20787__;
  assign new_new_n20789__ = ~new_new_n20776__ & ~new_new_n20788__;
  assign new_new_n20790__ = ~new_new_n20516__ & new_new_n20789__;
  assign new_new_n20791__ = new_new_n20516__ & ~new_new_n20789__;
  assign new_new_n20792__ = new_new_n3311__ & ~new_new_n15533__;
  assign new_new_n20793__ = new_new_n873__ & new_new_n15767__;
  assign new_new_n20794__ = ~new_new_n333__ & new_new_n15560__;
  assign new_new_n20795__ = ~new_new_n4900__ & new_new_n19893__;
  assign new_new_n20796__ = ~new_new_n20793__ & ~new_new_n20794__;
  assign new_new_n20797__ = ~new_new_n20792__ & new_new_n20796__;
  assign new_new_n20798__ = ~new_new_n20795__ & new_new_n20797__;
  assign new_new_n20799__ = pi26 & ~new_new_n20798__;
  assign new_new_n20800__ = ~pi26 & new_new_n20798__;
  assign new_new_n20801__ = ~new_new_n20799__ & ~new_new_n20800__;
  assign new_new_n20802__ = ~new_new_n20791__ & ~new_new_n20801__;
  assign new_new_n20803__ = ~new_new_n20790__ & ~new_new_n20802__;
  assign new_new_n20804__ = new_new_n20512__ & ~new_new_n20803__;
  assign new_new_n20805__ = ~new_new_n20512__ & new_new_n20803__;
  assign new_new_n20806__ = new_new_n3311__ & new_new_n15520__;
  assign new_new_n20807__ = ~new_new_n333__ & new_new_n15767__;
  assign new_new_n20808__ = new_new_n873__ & ~new_new_n15533__;
  assign new_new_n20809__ = ~new_new_n20807__ & ~new_new_n20808__;
  assign new_new_n20810__ = ~new_new_n20806__ & new_new_n20809__;
  assign new_new_n20811__ = ~pi26 & ~new_new_n20810__;
  assign new_new_n20812__ = new_new_n512__ & new_new_n19731__;
  assign new_new_n20813__ = new_new_n801__ & new_new_n19731__;
  assign new_new_n20814__ = pi26 & ~new_new_n20813__;
  assign new_new_n20815__ = ~new_new_n20812__ & ~new_new_n20814__;
  assign new_new_n20816__ = new_new_n20810__ & ~new_new_n20815__;
  assign new_new_n20817__ = ~new_new_n20811__ & ~new_new_n20816__;
  assign new_new_n20818__ = ~new_new_n20805__ & new_new_n20817__;
  assign new_new_n20819__ = ~new_new_n20804__ & ~new_new_n20818__;
  assign new_new_n20820__ = ~new_new_n20359__ & ~new_new_n20364__;
  assign new_new_n20821__ = new_new_n20366__ & new_new_n20820__;
  assign new_new_n20822__ = ~new_new_n20366__ & ~new_new_n20820__;
  assign new_new_n20823__ = ~new_new_n20821__ & ~new_new_n20822__;
  assign new_new_n20824__ = new_new_n20819__ & ~new_new_n20823__;
  assign new_new_n20825__ = ~new_new_n20819__ & new_new_n20823__;
  assign new_new_n20826__ = new_new_n5183__ & ~new_new_n15809__;
  assign new_new_n20827__ = new_new_n5191__ & ~new_new_n15487__;
  assign new_new_n20828__ = new_new_n5213__ & ~new_new_n15471__;
  assign new_new_n20829__ = ~new_new_n20826__ & ~new_new_n20827__;
  assign new_new_n20830__ = ~new_new_n20828__ & new_new_n20829__;
  assign new_new_n20831__ = new_new_n5195__ & ~new_new_n18633__;
  assign new_new_n20832__ = pi23 & ~new_new_n20831__;
  assign new_new_n20833__ = new_new_n7878__ & ~new_new_n18633__;
  assign new_new_n20834__ = ~new_new_n20832__ & ~new_new_n20833__;
  assign new_new_n20835__ = new_new_n20830__ & ~new_new_n20834__;
  assign new_new_n20836__ = ~pi23 & ~new_new_n20830__;
  assign new_new_n20837__ = ~new_new_n20835__ & ~new_new_n20836__;
  assign new_new_n20838__ = ~new_new_n20825__ & ~new_new_n20837__;
  assign new_new_n20839__ = ~new_new_n20824__ & ~new_new_n20838__;
  assign new_new_n20840__ = ~new_new_n20493__ & ~new_new_n20839__;
  assign new_new_n20841__ = ~new_new_n20492__ & ~new_new_n20840__;
  assign new_new_n20842__ = new_new_n20479__ & new_new_n20841__;
  assign new_new_n20843__ = ~new_new_n20479__ & ~new_new_n20841__;
  assign new_new_n20844__ = ~new_new_n20073__ & ~new_new_n20074__;
  assign new_new_n20845__ = ~new_new_n20386__ & new_new_n20844__;
  assign new_new_n20846__ = new_new_n20386__ & ~new_new_n20844__;
  assign new_new_n20847__ = ~new_new_n20845__ & ~new_new_n20846__;
  assign new_new_n20848__ = ~new_new_n20843__ & new_new_n20847__;
  assign new_new_n20849__ = ~new_new_n20842__ & ~new_new_n20848__;
  assign new_new_n20850__ = new_new_n6959__ & ~new_new_n17103__;
  assign new_new_n20851__ = new_new_n6964__ & ~new_new_n15349__;
  assign new_new_n20852__ = new_new_n6968__ & ~new_new_n15321__;
  assign new_new_n20853__ = ~new_new_n20851__ & ~new_new_n20852__;
  assign new_new_n20854__ = ~new_new_n20850__ & new_new_n20853__;
  assign new_new_n20855__ = new_new_n6958__ & ~new_new_n15273__;
  assign new_new_n20856__ = ~pi17 & ~new_new_n20855__;
  assign new_new_n20857__ = new_new_n7942__ & ~new_new_n15273__;
  assign new_new_n20858__ = ~new_new_n20856__ & ~new_new_n20857__;
  assign new_new_n20859__ = new_new_n20854__ & ~new_new_n20858__;
  assign new_new_n20860__ = pi17 & ~new_new_n20854__;
  assign new_new_n20861__ = ~new_new_n20859__ & ~new_new_n20860__;
  assign new_new_n20862__ = ~new_new_n20849__ & ~new_new_n20861__;
  assign new_new_n20863__ = new_new_n20849__ & new_new_n20861__;
  assign new_new_n20864__ = ~new_new_n20053__ & ~new_new_n20054__;
  assign new_new_n20865__ = ~new_new_n20388__ & new_new_n20864__;
  assign new_new_n20866__ = new_new_n20388__ & ~new_new_n20864__;
  assign new_new_n20867__ = ~new_new_n20865__ & ~new_new_n20866__;
  assign new_new_n20868__ = ~new_new_n20863__ & new_new_n20867__;
  assign new_new_n20869__ = ~new_new_n20862__ & ~new_new_n20868__;
  assign new_new_n20870__ = ~new_new_n20467__ & ~new_new_n20869__;
  assign new_new_n20871__ = ~new_new_n20466__ & ~new_new_n20870__;
  assign new_new_n20872__ = pi11 & ~new_new_n20871__;
  assign new_new_n20873__ = ~pi11 & new_new_n20871__;
  assign new_new_n20874__ = ~new_new_n20872__ & ~new_new_n20873__;
  assign new_new_n20875__ = new_new_n20444__ & new_new_n20874__;
  assign new_new_n20876__ = ~new_new_n20444__ & ~new_new_n20874__;
  assign new_new_n20877__ = ~new_new_n20875__ & ~new_new_n20876__;
  assign new_new_n20878__ = ~new_new_n20437__ & new_new_n20877__;
  assign new_new_n20879__ = new_new_n20437__ & ~new_new_n20877__;
  assign new_new_n20880__ = ~new_new_n20878__ & ~new_new_n20879__;
  assign new_new_n20881__ = new_new_n17569__ & new_new_n20880__;
  assign new_new_n20882__ = ~new_new_n17569__ & ~new_new_n20880__;
  assign new_new_n20883__ = ~new_new_n20881__ & ~new_new_n20882__;
  assign new_new_n20884__ = ~pi13 & new_new_n15248__;
  assign new_new_n20885__ = pi14 & ~new_new_n15248__;
  assign new_new_n20886__ = ~new_new_n20884__ & ~new_new_n20885__;
  assign new_new_n20887__ = new_new_n16725__ & new_new_n20886__;
  assign new_new_n20888__ = ~pi14 & new_new_n15248__;
  assign new_new_n20889__ = pi13 & ~new_new_n15248__;
  assign new_new_n20890__ = ~new_new_n20888__ & ~new_new_n20889__;
  assign new_new_n20891__ = ~new_new_n16725__ & new_new_n20890__;
  assign new_new_n20892__ = ~new_new_n20887__ & ~new_new_n20891__;
  assign new_new_n20893__ = new_new_n6994__ & ~new_new_n20892__;
  assign new_new_n20894__ = ~pi14 & new_new_n19825__;
  assign new_new_n20895__ = ~new_new_n15314__ & new_new_n20894__;
  assign new_new_n20896__ = new_new_n15285__ & new_new_n19823__;
  assign new_new_n20897__ = ~new_new_n15314__ & new_new_n19825__;
  assign new_new_n20898__ = ~pi13 & new_new_n15285__;
  assign new_new_n20899__ = ~pi12 & new_new_n20898__;
  assign new_new_n20900__ = pi14 & ~new_new_n20899__;
  assign new_new_n20901__ = ~new_new_n20897__ & new_new_n20900__;
  assign new_new_n20902__ = ~new_new_n20895__ & ~new_new_n20896__;
  assign new_new_n20903__ = ~new_new_n20901__ & new_new_n20902__;
  assign new_new_n20904__ = ~new_new_n6994__ & ~new_new_n20903__;
  assign new_new_n20905__ = ~new_new_n20893__ & ~new_new_n20904__;
  assign new_new_n20906__ = ~pi13 & new_new_n16082__;
  assign new_new_n20907__ = ~pi14 & ~new_new_n16082__;
  assign new_new_n20908__ = ~new_new_n20906__ & ~new_new_n20907__;
  assign new_new_n20909__ = ~new_new_n15314__ & new_new_n20908__;
  assign new_new_n20910__ = new_new_n15314__ & ~new_new_n20908__;
  assign new_new_n20911__ = new_new_n6994__ & ~new_new_n20909__;
  assign new_new_n20912__ = ~new_new_n20910__ & new_new_n20911__;
  assign new_new_n20913__ = new_new_n15285__ & ~new_new_n19823__;
  assign new_new_n20914__ = new_new_n19827__ & new_new_n20913__;
  assign new_new_n20915__ = pi14 & new_new_n15273__;
  assign new_new_n20916__ = new_new_n19824__ & ~new_new_n20915__;
  assign new_new_n20917__ = ~new_new_n15273__ & new_new_n19823__;
  assign new_new_n20918__ = ~pi14 & ~new_new_n20917__;
  assign new_new_n20919__ = ~new_new_n20913__ & new_new_n20918__;
  assign new_new_n20920__ = ~new_new_n6994__ & ~new_new_n20916__;
  assign new_new_n20921__ = ~new_new_n20914__ & new_new_n20920__;
  assign new_new_n20922__ = ~new_new_n20919__ & new_new_n20921__;
  assign new_new_n20923__ = ~new_new_n20912__ & ~new_new_n20922__;
  assign new_new_n20924__ = ~new_new_n20842__ & ~new_new_n20843__;
  assign new_new_n20925__ = new_new_n20847__ & new_new_n20924__;
  assign new_new_n20926__ = ~new_new_n20847__ & ~new_new_n20924__;
  assign new_new_n20927__ = ~new_new_n20925__ & ~new_new_n20926__;
  assign new_new_n20928__ = ~new_new_n20923__ & ~new_new_n20927__;
  assign new_new_n20929__ = new_new_n20923__ & new_new_n20927__;
  assign new_new_n20930__ = ~new_new_n20492__ & ~new_new_n20493__;
  assign new_new_n20931__ = new_new_n20839__ & ~new_new_n20930__;
  assign new_new_n20932__ = ~new_new_n20839__ & new_new_n20930__;
  assign new_new_n20933__ = ~new_new_n20931__ & ~new_new_n20932__;
  assign new_new_n20934__ = new_new_n5183__ & ~new_new_n15487__;
  assign new_new_n20935__ = new_new_n5191__ & new_new_n15524__;
  assign new_new_n20936__ = ~new_new_n20934__ & ~new_new_n20935__;
  assign new_new_n20937__ = new_new_n5195__ & ~new_new_n15809__;
  assign new_new_n20938__ = new_new_n18020__ & new_new_n20937__;
  assign new_new_n20939__ = new_new_n20936__ & ~new_new_n20938__;
  assign new_new_n20940__ = pi23 & ~new_new_n20939__;
  assign new_new_n20941__ = new_new_n5195__ & ~new_new_n18019__;
  assign new_new_n20942__ = ~pi23 & ~new_new_n20941__;
  assign new_new_n20943__ = new_new_n15809__ & new_new_n18017__;
  assign new_new_n20944__ = ~pi22 & ~new_new_n20943__;
  assign new_new_n20945__ = pi22 & ~new_new_n18018__;
  assign new_new_n20946__ = new_new_n5195__ & ~new_new_n20944__;
  assign new_new_n20947__ = ~new_new_n20945__ & new_new_n20946__;
  assign new_new_n20948__ = ~new_new_n20942__ & ~new_new_n20947__;
  assign new_new_n20949__ = new_new_n20936__ & ~new_new_n20948__;
  assign new_new_n20950__ = ~new_new_n20940__ & ~new_new_n20949__;
  assign new_new_n20951__ = new_new_n5213__ & new_new_n15520__;
  assign new_new_n20952__ = new_new_n5191__ & new_new_n15767__;
  assign new_new_n20953__ = new_new_n5183__ & ~new_new_n15533__;
  assign new_new_n20954__ = ~new_new_n20952__ & ~new_new_n20953__;
  assign new_new_n20955__ = ~new_new_n20951__ & new_new_n20954__;
  assign new_new_n20956__ = new_new_n5195__ & new_new_n19731__;
  assign new_new_n20957__ = pi23 & ~new_new_n20956__;
  assign new_new_n20958__ = new_new_n7878__ & new_new_n19731__;
  assign new_new_n20959__ = ~new_new_n20957__ & ~new_new_n20958__;
  assign new_new_n20960__ = new_new_n20955__ & ~new_new_n20959__;
  assign new_new_n20961__ = ~pi23 & ~new_new_n20955__;
  assign new_new_n20962__ = ~new_new_n20960__ & ~new_new_n20961__;
  assign new_new_n20963__ = ~new_new_n20758__ & ~new_new_n20759__;
  assign new_new_n20964__ = new_new_n20769__ & new_new_n20963__;
  assign new_new_n20965__ = ~new_new_n20769__ & ~new_new_n20963__;
  assign new_new_n20966__ = ~new_new_n20964__ & ~new_new_n20965__;
  assign new_new_n20967__ = ~new_new_n20962__ & new_new_n20966__;
  assign new_new_n20968__ = new_new_n20962__ & ~new_new_n20966__;
  assign new_new_n20969__ = new_new_n5183__ & new_new_n15560__;
  assign new_new_n20970__ = new_new_n5191__ & new_new_n15572__;
  assign new_new_n20971__ = new_new_n5213__ & new_new_n15767__;
  assign new_new_n20972__ = ~new_new_n20970__ & ~new_new_n20971__;
  assign new_new_n20973__ = ~new_new_n20969__ & new_new_n20972__;
  assign new_new_n20974__ = new_new_n5195__ & ~new_new_n18454__;
  assign new_new_n20975__ = ~pi23 & ~new_new_n20974__;
  assign new_new_n20976__ = new_new_n5974__ & ~new_new_n18454__;
  assign new_new_n20977__ = ~new_new_n20975__ & ~new_new_n20976__;
  assign new_new_n20978__ = new_new_n20973__ & ~new_new_n20977__;
  assign new_new_n20979__ = pi23 & ~new_new_n20973__;
  assign new_new_n20980__ = ~new_new_n20978__ & ~new_new_n20979__;
  assign new_new_n20981__ = ~new_new_n20705__ & ~new_new_n20706__;
  assign new_new_n20982__ = ~new_new_n20716__ & new_new_n20981__;
  assign new_new_n20983__ = new_new_n20716__ & ~new_new_n20981__;
  assign new_new_n20984__ = ~new_new_n20982__ & ~new_new_n20983__;
  assign new_new_n20985__ = ~new_new_n20693__ & ~new_new_n20694__;
  assign new_new_n20986__ = new_new_n20257__ & ~new_new_n20697__;
  assign new_new_n20987__ = new_new_n20697__ & new_new_n20699__;
  assign new_new_n20988__ = ~new_new_n20986__ & ~new_new_n20987__;
  assign new_new_n20989__ = ~new_new_n20985__ & ~new_new_n20988__;
  assign new_new_n20990__ = ~new_new_n20702__ & new_new_n20985__;
  assign new_new_n20991__ = ~new_new_n20989__ & ~new_new_n20990__;
  assign new_new_n20992__ = ~new_new_n20599__ & ~new_new_n20675__;
  assign new_new_n20993__ = ~new_new_n20672__ & new_new_n20678__;
  assign new_new_n20994__ = ~new_new_n20611__ & ~new_new_n20993__;
  assign new_new_n20995__ = new_new_n20672__ & new_new_n20680__;
  assign new_new_n20996__ = ~new_new_n20994__ & ~new_new_n20995__;
  assign new_new_n20997__ = new_new_n20992__ & ~new_new_n20996__;
  assign new_new_n20998__ = ~new_new_n20992__ & new_new_n20996__;
  assign new_new_n20999__ = ~new_new_n20997__ & ~new_new_n20998__;
  assign new_new_n21000__ = new_new_n5215__ & new_new_n19487__;
  assign new_new_n21001__ = new_new_n5191__ & ~new_new_n15647__;
  assign new_new_n21002__ = new_new_n5183__ & ~new_new_n15582__;
  assign new_new_n21003__ = ~new_new_n21001__ & ~new_new_n21002__;
  assign new_new_n21004__ = ~new_new_n21000__ & new_new_n21003__;
  assign new_new_n21005__ = new_new_n5195__ & ~new_new_n15638__;
  assign new_new_n21006__ = pi23 & ~new_new_n21005__;
  assign new_new_n21007__ = new_new_n5974__ & ~new_new_n15638__;
  assign new_new_n21008__ = ~new_new_n21006__ & ~new_new_n21007__;
  assign new_new_n21009__ = new_new_n21004__ & ~new_new_n21008__;
  assign new_new_n21010__ = ~pi23 & ~new_new_n21004__;
  assign new_new_n21011__ = ~new_new_n21009__ & ~new_new_n21010__;
  assign new_new_n21012__ = new_new_n20625__ & ~new_new_n20667__;
  assign new_new_n21013__ = ~new_new_n20625__ & new_new_n20667__;
  assign new_new_n21014__ = ~new_new_n21012__ & ~new_new_n21013__;
  assign new_new_n21015__ = new_new_n20626__ & ~new_new_n21014__;
  assign new_new_n21016__ = new_new_n20641__ & new_new_n21012__;
  assign new_new_n21017__ = ~new_new_n21015__ & ~new_new_n21016__;
  assign new_new_n21018__ = ~new_new_n20659__ & ~new_new_n21017__;
  assign new_new_n21019__ = ~new_new_n20660__ & new_new_n21014__;
  assign new_new_n21020__ = ~new_new_n21018__ & ~new_new_n21019__;
  assign new_new_n21021__ = new_new_n5213__ & ~new_new_n15582__;
  assign new_new_n21022__ = new_new_n5191__ & ~new_new_n15710__;
  assign new_new_n21023__ = new_new_n5183__ & ~new_new_n15647__;
  assign new_new_n21024__ = ~new_new_n21022__ & ~new_new_n21023__;
  assign new_new_n21025__ = ~new_new_n21021__ & new_new_n21024__;
  assign new_new_n21026__ = new_new_n5195__ & ~new_new_n15736__;
  assign new_new_n21027__ = pi23 & ~new_new_n21026__;
  assign new_new_n21028__ = new_new_n7878__ & ~new_new_n15736__;
  assign new_new_n21029__ = ~new_new_n21027__ & ~new_new_n21028__;
  assign new_new_n21030__ = new_new_n21025__ & ~new_new_n21029__;
  assign new_new_n21031__ = ~pi23 & ~new_new_n21025__;
  assign new_new_n21032__ = ~new_new_n21030__ & ~new_new_n21031__;
  assign new_new_n21033__ = new_new_n21020__ & ~new_new_n21032__;
  assign new_new_n21034__ = ~new_new_n21020__ & new_new_n21032__;
  assign new_new_n21035__ = new_new_n5183__ & ~new_new_n15710__;
  assign new_new_n21036__ = new_new_n5191__ & new_new_n15656__;
  assign new_new_n21037__ = new_new_n5213__ & ~new_new_n15647__;
  assign new_new_n21038__ = ~new_new_n21035__ & ~new_new_n21036__;
  assign new_new_n21039__ = ~new_new_n21037__ & new_new_n21038__;
  assign new_new_n21040__ = new_new_n5195__ & ~new_new_n19118__;
  assign new_new_n21041__ = pi23 & ~new_new_n21040__;
  assign new_new_n21042__ = new_new_n7878__ & ~new_new_n19118__;
  assign new_new_n21043__ = ~new_new_n21041__ & ~new_new_n21042__;
  assign new_new_n21044__ = new_new_n21039__ & ~new_new_n21043__;
  assign new_new_n21045__ = ~pi23 & ~new_new_n21039__;
  assign new_new_n21046__ = ~new_new_n21044__ & ~new_new_n21045__;
  assign new_new_n21047__ = pi26 & ~new_new_n20630__;
  assign new_new_n21048__ = ~new_new_n20639__ & new_new_n21047__;
  assign new_new_n21049__ = new_new_n20639__ & ~new_new_n21047__;
  assign new_new_n21050__ = ~new_new_n21048__ & ~new_new_n21049__;
  assign new_new_n21051__ = new_new_n5213__ & new_new_n15656__;
  assign new_new_n21052__ = new_new_n5191__ & ~new_new_n15661__;
  assign new_new_n21053__ = new_new_n5183__ & new_new_n15643__;
  assign new_new_n21054__ = ~new_new_n21052__ & ~new_new_n21053__;
  assign new_new_n21055__ = ~new_new_n21051__ & new_new_n21054__;
  assign new_new_n21056__ = new_new_n5195__ & new_new_n15687__;
  assign new_new_n21057__ = pi23 & ~new_new_n21056__;
  assign new_new_n21058__ = new_new_n7878__ & new_new_n15687__;
  assign new_new_n21059__ = ~new_new_n21057__ & ~new_new_n21058__;
  assign new_new_n21060__ = new_new_n21055__ & ~new_new_n21059__;
  assign new_new_n21061__ = ~pi23 & ~new_new_n21055__;
  assign new_new_n21062__ = ~new_new_n21060__ & ~new_new_n21061__;
  assign new_new_n21063__ = ~new_new_n110__ & ~new_new_n15673__;
  assign new_new_n21064__ = ~new_new_n5185__ & ~new_new_n5188__;
  assign new_new_n21065__ = ~new_new_n15673__ & new_new_n21064__;
  assign new_new_n21066__ = new_new_n5195__ & ~new_new_n20628__;
  assign new_new_n21067__ = ~new_new_n21065__ & ~new_new_n21066__;
  assign new_new_n21068__ = new_new_n5191__ & ~new_new_n15673__;
  assign new_new_n21069__ = new_new_n5183__ & new_new_n15668__;
  assign new_new_n21070__ = new_new_n5212__ & new_new_n20195__;
  assign new_new_n21071__ = new_new_n15661__ & ~new_new_n21070__;
  assign new_new_n21072__ = ~new_new_n15661__ & new_new_n21070__;
  assign new_new_n21073__ = new_new_n5195__ & ~new_new_n21071__;
  assign new_new_n21074__ = ~new_new_n21072__ & new_new_n21073__;
  assign new_new_n21075__ = ~new_new_n21068__ & ~new_new_n21069__;
  assign new_new_n21076__ = ~new_new_n21074__ & new_new_n21075__;
  assign new_new_n21077__ = pi23 & new_new_n21067__;
  assign new_new_n21078__ = new_new_n21076__ & new_new_n21077__;
  assign new_new_n21079__ = ~new_new_n21063__ & ~new_new_n21078__;
  assign new_new_n21080__ = new_new_n5213__ & new_new_n15643__;
  assign new_new_n21081__ = new_new_n5191__ & new_new_n15668__;
  assign new_new_n21082__ = new_new_n5183__ & ~new_new_n15661__;
  assign new_new_n21083__ = ~new_new_n21081__ & ~new_new_n21082__;
  assign new_new_n21084__ = ~new_new_n21080__ & new_new_n21083__;
  assign new_new_n21085__ = new_new_n15643__ & new_new_n20176__;
  assign new_new_n21086__ = new_new_n5195__ & ~new_new_n20177__;
  assign new_new_n21087__ = ~new_new_n21085__ & new_new_n21086__;
  assign new_new_n21088__ = ~pi23 & ~new_new_n21087__;
  assign new_new_n21089__ = ~pi22 & new_new_n21087__;
  assign new_new_n21090__ = ~new_new_n21088__ & ~new_new_n21089__;
  assign new_new_n21091__ = new_new_n21084__ & ~new_new_n21090__;
  assign new_new_n21092__ = pi23 & ~new_new_n21084__;
  assign new_new_n21093__ = ~new_new_n21091__ & ~new_new_n21092__;
  assign new_new_n21094__ = ~new_new_n21079__ & new_new_n21093__;
  assign new_new_n21095__ = new_new_n419__ & new_new_n15674__;
  assign new_new_n21096__ = ~new_new_n104__ & new_new_n15668__;
  assign new_new_n21097__ = new_new_n389__ & ~new_new_n21096__;
  assign new_new_n21098__ = new_new_n110__ & new_new_n20195__;
  assign new_new_n21099__ = ~new_new_n146__ & ~new_new_n20628__;
  assign new_new_n21100__ = ~new_new_n21095__ & new_new_n21099__;
  assign new_new_n21101__ = ~new_new_n21097__ & ~new_new_n21098__;
  assign new_new_n21102__ = new_new_n21100__ & new_new_n21101__;
  assign new_new_n21103__ = ~new_new_n21094__ & ~new_new_n21102__;
  assign new_new_n21104__ = ~new_new_n21062__ & ~new_new_n21103__;
  assign new_new_n21105__ = new_new_n21063__ & new_new_n21102__;
  assign new_new_n21106__ = new_new_n21093__ & new_new_n21105__;
  assign new_new_n21107__ = ~new_new_n21104__ & ~new_new_n21106__;
  assign new_new_n21108__ = ~new_new_n21050__ & new_new_n21107__;
  assign new_new_n21109__ = new_new_n21050__ & ~new_new_n21107__;
  assign new_new_n21110__ = new_new_n5213__ & ~new_new_n15710__;
  assign new_new_n21111__ = new_new_n5183__ & new_new_n15656__;
  assign new_new_n21112__ = new_new_n5191__ & new_new_n15643__;
  assign new_new_n21113__ = new_new_n5215__ & ~new_new_n19466__;
  assign new_new_n21114__ = ~new_new_n21111__ & ~new_new_n21112__;
  assign new_new_n21115__ = ~new_new_n21110__ & new_new_n21114__;
  assign new_new_n21116__ = ~new_new_n21113__ & new_new_n21115__;
  assign new_new_n21117__ = pi23 & ~new_new_n21116__;
  assign new_new_n21118__ = ~pi23 & new_new_n21116__;
  assign new_new_n21119__ = ~new_new_n21117__ & ~new_new_n21118__;
  assign new_new_n21120__ = ~new_new_n21109__ & ~new_new_n21119__;
  assign new_new_n21121__ = ~new_new_n21108__ & ~new_new_n21120__;
  assign new_new_n21122__ = ~new_new_n21046__ & new_new_n21121__;
  assign new_new_n21123__ = new_new_n21046__ & ~new_new_n21121__;
  assign new_new_n21124__ = new_new_n20626__ & new_new_n20641__;
  assign new_new_n21125__ = ~new_new_n20659__ & ~new_new_n21124__;
  assign new_new_n21126__ = new_new_n20642__ & ~new_new_n21125__;
  assign new_new_n21127__ = ~new_new_n20642__ & new_new_n21125__;
  assign new_new_n21128__ = ~new_new_n21126__ & ~new_new_n21127__;
  assign new_new_n21129__ = ~new_new_n21123__ & new_new_n21128__;
  assign new_new_n21130__ = ~new_new_n21122__ & ~new_new_n21129__;
  assign new_new_n21131__ = ~new_new_n21034__ & ~new_new_n21130__;
  assign new_new_n21132__ = ~new_new_n21033__ & ~new_new_n21131__;
  assign new_new_n21133__ = ~new_new_n21011__ & ~new_new_n21132__;
  assign new_new_n21134__ = ~new_new_n20217__ & new_new_n20672__;
  assign new_new_n21135__ = new_new_n20217__ & ~new_new_n20672__;
  assign new_new_n21136__ = ~new_new_n21011__ & new_new_n21135__;
  assign new_new_n21137__ = ~new_new_n21134__ & ~new_new_n21136__;
  assign new_new_n21138__ = new_new_n21011__ & new_new_n21132__;
  assign new_new_n21139__ = new_new_n20210__ & ~new_new_n20611__;
  assign new_new_n21140__ = ~new_new_n20210__ & new_new_n20611__;
  assign new_new_n21141__ = ~new_new_n21139__ & ~new_new_n21140__;
  assign new_new_n21142__ = ~new_new_n21137__ & new_new_n21141__;
  assign new_new_n21143__ = ~new_new_n21138__ & new_new_n21142__;
  assign new_new_n21144__ = new_new_n20218__ & ~new_new_n20672__;
  assign new_new_n21145__ = ~new_new_n21134__ & ~new_new_n21144__;
  assign new_new_n21146__ = ~new_new_n21141__ & new_new_n21145__;
  assign new_new_n21147__ = ~new_new_n21138__ & new_new_n21146__;
  assign new_new_n21148__ = ~new_new_n21133__ & ~new_new_n21147__;
  assign new_new_n21149__ = ~new_new_n21143__ & new_new_n21148__;
  assign new_new_n21150__ = ~new_new_n20999__ & ~new_new_n21149__;
  assign new_new_n21151__ = new_new_n20999__ & new_new_n21149__;
  assign new_new_n21152__ = new_new_n5215__ & new_new_n19494__;
  assign new_new_n21153__ = new_new_n5191__ & ~new_new_n15582__;
  assign new_new_n21154__ = new_new_n5183__ & ~new_new_n15638__;
  assign new_new_n21155__ = new_new_n5213__ & new_new_n15743__;
  assign new_new_n21156__ = ~new_new_n21153__ & ~new_new_n21154__;
  assign new_new_n21157__ = ~new_new_n21155__ & new_new_n21156__;
  assign new_new_n21158__ = ~new_new_n21152__ & new_new_n21157__;
  assign new_new_n21159__ = ~pi23 & ~new_new_n21158__;
  assign new_new_n21160__ = pi23 & new_new_n21158__;
  assign new_new_n21161__ = ~new_new_n21159__ & ~new_new_n21160__;
  assign new_new_n21162__ = ~new_new_n21151__ & ~new_new_n21161__;
  assign new_new_n21163__ = ~new_new_n21150__ & ~new_new_n21162__;
  assign new_new_n21164__ = ~new_new_n20685__ & ~new_new_n20686__;
  assign new_new_n21165__ = new_new_n20690__ & new_new_n21164__;
  assign new_new_n21166__ = ~new_new_n20690__ & ~new_new_n21164__;
  assign new_new_n21167__ = ~new_new_n21165__ & ~new_new_n21166__;
  assign new_new_n21168__ = ~new_new_n21163__ & new_new_n21167__;
  assign new_new_n21169__ = new_new_n21163__ & ~new_new_n21167__;
  assign new_new_n21170__ = new_new_n5213__ & ~new_new_n15615__;
  assign new_new_n21171__ = new_new_n5183__ & new_new_n15743__;
  assign new_new_n21172__ = new_new_n5191__ & ~new_new_n15638__;
  assign new_new_n21173__ = new_new_n5215__ & new_new_n19005__;
  assign new_new_n21174__ = ~new_new_n21171__ & ~new_new_n21172__;
  assign new_new_n21175__ = ~new_new_n21170__ & new_new_n21174__;
  assign new_new_n21176__ = ~new_new_n21173__ & new_new_n21175__;
  assign new_new_n21177__ = pi23 & ~new_new_n21176__;
  assign new_new_n21178__ = ~pi23 & new_new_n21176__;
  assign new_new_n21179__ = ~new_new_n21177__ & ~new_new_n21178__;
  assign new_new_n21180__ = ~new_new_n21169__ & new_new_n21179__;
  assign new_new_n21181__ = ~new_new_n21168__ & ~new_new_n21180__;
  assign new_new_n21182__ = ~new_new_n20991__ & new_new_n21181__;
  assign new_new_n21183__ = new_new_n20991__ & ~new_new_n21181__;
  assign new_new_n21184__ = new_new_n5213__ & new_new_n15564__;
  assign new_new_n21185__ = new_new_n5191__ & new_new_n15743__;
  assign new_new_n21186__ = new_new_n5183__ & ~new_new_n15615__;
  assign new_new_n21187__ = new_new_n5215__ & new_new_n18512__;
  assign new_new_n21188__ = ~new_new_n21185__ & ~new_new_n21186__;
  assign new_new_n21189__ = ~new_new_n21184__ & new_new_n21188__;
  assign new_new_n21190__ = ~new_new_n21187__ & new_new_n21189__;
  assign new_new_n21191__ = pi23 & ~new_new_n21190__;
  assign new_new_n21192__ = ~pi23 & new_new_n21190__;
  assign new_new_n21193__ = ~new_new_n21191__ & ~new_new_n21192__;
  assign new_new_n21194__ = ~new_new_n21183__ & ~new_new_n21193__;
  assign new_new_n21195__ = ~new_new_n21182__ & ~new_new_n21194__;
  assign new_new_n21196__ = ~new_new_n20984__ & new_new_n21195__;
  assign new_new_n21197__ = new_new_n5191__ & ~new_new_n15615__;
  assign new_new_n21198__ = new_new_n5183__ & new_new_n15564__;
  assign new_new_n21199__ = ~new_new_n21197__ & ~new_new_n21198__;
  assign new_new_n21200__ = new_new_n5195__ & ~new_new_n20528__;
  assign new_new_n21201__ = pi23 & ~new_new_n21200__;
  assign new_new_n21202__ = pi22 & ~new_new_n15572__;
  assign new_new_n21203__ = ~pi22 & new_new_n15572__;
  assign new_new_n21204__ = ~new_new_n21202__ & ~new_new_n21203__;
  assign new_new_n21205__ = new_new_n5195__ & new_new_n19534__;
  assign new_new_n21206__ = ~new_new_n21204__ & new_new_n21205__;
  assign new_new_n21207__ = ~new_new_n21201__ & ~new_new_n21206__;
  assign new_new_n21208__ = new_new_n21199__ & ~new_new_n21207__;
  assign new_new_n21209__ = new_new_n5195__ & new_new_n20111__;
  assign new_new_n21210__ = new_new_n21199__ & ~new_new_n21209__;
  assign new_new_n21211__ = ~pi23 & ~new_new_n21210__;
  assign new_new_n21212__ = ~new_new_n21208__ & ~new_new_n21211__;
  assign new_new_n21213__ = new_new_n20984__ & ~new_new_n21195__;
  assign new_new_n21214__ = ~new_new_n21212__ & ~new_new_n21213__;
  assign new_new_n21215__ = ~new_new_n21196__ & ~new_new_n21214__;
  assign new_new_n21216__ = ~new_new_n20719__ & ~new_new_n20720__;
  assign new_new_n21217__ = ~new_new_n20276__ & new_new_n20723__;
  assign new_new_n21218__ = new_new_n20276__ & ~new_new_n20723__;
  assign new_new_n21219__ = ~new_new_n21217__ & ~new_new_n21218__;
  assign new_new_n21220__ = new_new_n21216__ & new_new_n21219__;
  assign new_new_n21221__ = ~new_new_n21216__ & ~new_new_n21219__;
  assign new_new_n21222__ = ~new_new_n21220__ & ~new_new_n21221__;
  assign new_new_n21223__ = new_new_n21215__ & ~new_new_n21222__;
  assign new_new_n21224__ = ~new_new_n21215__ & new_new_n21222__;
  assign new_new_n21225__ = new_new_n5213__ & new_new_n15560__;
  assign new_new_n21226__ = new_new_n5183__ & new_new_n15572__;
  assign new_new_n21227__ = new_new_n5191__ & new_new_n15564__;
  assign new_new_n21228__ = new_new_n5215__ & new_new_n18944__;
  assign new_new_n21229__ = ~new_new_n21226__ & ~new_new_n21227__;
  assign new_new_n21230__ = ~new_new_n21225__ & new_new_n21229__;
  assign new_new_n21231__ = ~new_new_n21228__ & new_new_n21230__;
  assign new_new_n21232__ = pi23 & ~new_new_n21231__;
  assign new_new_n21233__ = ~pi23 & new_new_n21231__;
  assign new_new_n21234__ = ~new_new_n21232__ & ~new_new_n21233__;
  assign new_new_n21235__ = ~new_new_n21224__ & ~new_new_n21234__;
  assign new_new_n21236__ = ~new_new_n21223__ & ~new_new_n21235__;
  assign new_new_n21237__ = ~new_new_n20980__ & ~new_new_n21236__;
  assign new_new_n21238__ = new_new_n20980__ & new_new_n21236__;
  assign new_new_n21239__ = ~new_new_n20729__ & ~new_new_n20730__;
  assign new_new_n21240__ = new_new_n20749__ & new_new_n21239__;
  assign new_new_n21241__ = ~new_new_n20749__ & ~new_new_n21239__;
  assign new_new_n21242__ = ~new_new_n21240__ & ~new_new_n21241__;
  assign new_new_n21243__ = ~new_new_n21238__ & ~new_new_n21242__;
  assign new_new_n21244__ = ~new_new_n21237__ & ~new_new_n21243__;
  assign new_new_n21245__ = ~new_new_n20538__ & ~new_new_n20539__;
  assign new_new_n21246__ = new_new_n20751__ & new_new_n21245__;
  assign new_new_n21247__ = ~new_new_n20751__ & ~new_new_n21245__;
  assign new_new_n21248__ = ~new_new_n21246__ & ~new_new_n21247__;
  assign new_new_n21249__ = ~new_new_n21244__ & ~new_new_n21248__;
  assign new_new_n21250__ = new_new_n21244__ & new_new_n21248__;
  assign new_new_n21251__ = new_new_n5191__ & new_new_n15560__;
  assign new_new_n21252__ = new_new_n5183__ & new_new_n15767__;
  assign new_new_n21253__ = new_new_n5213__ & ~new_new_n15533__;
  assign new_new_n21254__ = ~new_new_n21251__ & ~new_new_n21252__;
  assign new_new_n21255__ = ~new_new_n21253__ & new_new_n21254__;
  assign new_new_n21256__ = new_new_n5195__ & new_new_n19893__;
  assign new_new_n21257__ = ~pi23 & ~new_new_n21256__;
  assign new_new_n21258__ = new_new_n5974__ & new_new_n19893__;
  assign new_new_n21259__ = ~new_new_n21257__ & ~new_new_n21258__;
  assign new_new_n21260__ = new_new_n21255__ & ~new_new_n21259__;
  assign new_new_n21261__ = pi23 & ~new_new_n21255__;
  assign new_new_n21262__ = ~new_new_n21260__ & ~new_new_n21261__;
  assign new_new_n21263__ = ~new_new_n21250__ & ~new_new_n21262__;
  assign new_new_n21264__ = ~new_new_n21249__ & ~new_new_n21263__;
  assign new_new_n21265__ = ~new_new_n20968__ & new_new_n21264__;
  assign new_new_n21266__ = ~new_new_n20967__ & ~new_new_n21265__;
  assign new_new_n21267__ = ~new_new_n20776__ & ~new_new_n20777__;
  assign new_new_n21268__ = new_new_n20787__ & new_new_n21267__;
  assign new_new_n21269__ = ~new_new_n20787__ & ~new_new_n21267__;
  assign new_new_n21270__ = ~new_new_n21268__ & ~new_new_n21269__;
  assign new_new_n21271__ = ~new_new_n21266__ & new_new_n21270__;
  assign new_new_n21272__ = new_new_n5183__ & new_new_n15520__;
  assign new_new_n21273__ = new_new_n5191__ & ~new_new_n15533__;
  assign new_new_n21274__ = ~new_new_n21272__ & ~new_new_n21273__;
  assign new_new_n21275__ = new_new_n5195__ & new_new_n18923__;
  assign new_new_n21276__ = new_new_n21274__ & ~new_new_n21275__;
  assign new_new_n21277__ = pi23 & ~new_new_n21276__;
  assign new_new_n21278__ = new_new_n5195__ & ~new_new_n18914__;
  assign new_new_n21279__ = ~pi23 & ~new_new_n21278__;
  assign new_new_n21280__ = ~pi22 & new_new_n15524__;
  assign new_new_n21281__ = pi22 & ~new_new_n15524__;
  assign new_new_n21282__ = new_new_n5195__ & ~new_new_n21280__;
  assign new_new_n21283__ = ~new_new_n21281__ & new_new_n21282__;
  assign new_new_n21284__ = new_new_n18913__ & new_new_n21283__;
  assign new_new_n21285__ = ~new_new_n21279__ & ~new_new_n21284__;
  assign new_new_n21286__ = new_new_n21274__ & ~new_new_n21285__;
  assign new_new_n21287__ = ~new_new_n21277__ & ~new_new_n21286__;
  assign new_new_n21288__ = new_new_n21266__ & ~new_new_n21270__;
  assign new_new_n21289__ = new_new_n21287__ & ~new_new_n21288__;
  assign new_new_n21290__ = ~new_new_n21271__ & ~new_new_n21289__;
  assign new_new_n21291__ = ~new_new_n20790__ & ~new_new_n20791__;
  assign new_new_n21292__ = ~new_new_n20801__ & new_new_n21291__;
  assign new_new_n21293__ = new_new_n20801__ & ~new_new_n21291__;
  assign new_new_n21294__ = ~new_new_n21292__ & ~new_new_n21293__;
  assign new_new_n21295__ = ~new_new_n21290__ & ~new_new_n21294__;
  assign new_new_n21296__ = new_new_n21290__ & new_new_n21294__;
  assign new_new_n21297__ = new_new_n5213__ & ~new_new_n15487__;
  assign new_new_n21298__ = new_new_n5183__ & new_new_n15524__;
  assign new_new_n21299__ = new_new_n5191__ & new_new_n15520__;
  assign new_new_n21300__ = new_new_n5215__ & new_new_n17587__;
  assign new_new_n21301__ = ~new_new_n21298__ & ~new_new_n21299__;
  assign new_new_n21302__ = ~new_new_n21297__ & new_new_n21301__;
  assign new_new_n21303__ = ~new_new_n21300__ & new_new_n21302__;
  assign new_new_n21304__ = ~pi23 & ~new_new_n21303__;
  assign new_new_n21305__ = pi23 & new_new_n21303__;
  assign new_new_n21306__ = ~new_new_n21304__ & ~new_new_n21305__;
  assign new_new_n21307__ = ~new_new_n21296__ & ~new_new_n21306__;
  assign new_new_n21308__ = ~new_new_n21295__ & ~new_new_n21307__;
  assign new_new_n21309__ = new_new_n20950__ & ~new_new_n21308__;
  assign new_new_n21310__ = ~new_new_n20950__ & new_new_n21308__;
  assign new_new_n21311__ = ~new_new_n20804__ & ~new_new_n20805__;
  assign new_new_n21312__ = new_new_n20817__ & new_new_n21311__;
  assign new_new_n21313__ = ~new_new_n20817__ & ~new_new_n21311__;
  assign new_new_n21314__ = ~new_new_n21312__ & ~new_new_n21313__;
  assign new_new_n21315__ = ~new_new_n21310__ & ~new_new_n21314__;
  assign new_new_n21316__ = ~new_new_n21309__ & ~new_new_n21315__;
  assign new_new_n21317__ = ~new_new_n20824__ & ~new_new_n20825__;
  assign new_new_n21318__ = ~new_new_n20837__ & new_new_n21317__;
  assign new_new_n21319__ = new_new_n20837__ & ~new_new_n21317__;
  assign new_new_n21320__ = ~new_new_n21318__ & ~new_new_n21319__;
  assign new_new_n21321__ = ~new_new_n21316__ & new_new_n21320__;
  assign new_new_n21322__ = new_new_n21316__ & ~new_new_n21320__;
  assign new_new_n21323__ = new_new_n6634__ & ~new_new_n15432__;
  assign new_new_n21324__ = new_new_n6629__ & ~new_new_n15439__;
  assign new_new_n21325__ = ~new_new_n6625__ & new_new_n15464__;
  assign new_new_n21326__ = new_new_n6936__ & new_new_n17204__;
  assign new_new_n21327__ = ~new_new_n21324__ & ~new_new_n21325__;
  assign new_new_n21328__ = ~new_new_n21323__ & new_new_n21327__;
  assign new_new_n21329__ = ~new_new_n21326__ & new_new_n21328__;
  assign new_new_n21330__ = ~pi20 & ~new_new_n21329__;
  assign new_new_n21331__ = pi20 & new_new_n21329__;
  assign new_new_n21332__ = ~new_new_n21330__ & ~new_new_n21331__;
  assign new_new_n21333__ = ~new_new_n21322__ & ~new_new_n21332__;
  assign new_new_n21334__ = ~new_new_n21321__ & ~new_new_n21333__;
  assign new_new_n21335__ = new_new_n20933__ & ~new_new_n21334__;
  assign new_new_n21336__ = ~new_new_n20933__ & new_new_n21334__;
  assign new_new_n21337__ = new_new_n7935__ & ~new_new_n15349__;
  assign new_new_n21338__ = new_new_n6964__ & new_new_n15390__;
  assign new_new_n21339__ = new_new_n6968__ & ~new_new_n15398__;
  assign new_new_n21340__ = ~new_new_n21338__ & ~new_new_n21339__;
  assign new_new_n21341__ = ~new_new_n21337__ & new_new_n21340__;
  assign new_new_n21342__ = new_new_n6958__ & ~new_new_n17180__;
  assign new_new_n21343__ = pi17 & ~new_new_n21342__;
  assign new_new_n21344__ = new_new_n7942__ & ~new_new_n17180__;
  assign new_new_n21345__ = ~new_new_n21343__ & ~new_new_n21344__;
  assign new_new_n21346__ = new_new_n21341__ & ~new_new_n21345__;
  assign new_new_n21347__ = ~pi17 & ~new_new_n21341__;
  assign new_new_n21348__ = ~new_new_n21346__ & ~new_new_n21347__;
  assign new_new_n21349__ = ~new_new_n21336__ & ~new_new_n21348__;
  assign new_new_n21350__ = ~new_new_n21335__ & ~new_new_n21349__;
  assign new_new_n21351__ = ~new_new_n20929__ & ~new_new_n21350__;
  assign new_new_n21352__ = ~new_new_n20928__ & ~new_new_n21351__;
  assign new_new_n21353__ = ~new_new_n20905__ & ~new_new_n21352__;
  assign new_new_n21354__ = new_new_n20905__ & new_new_n21352__;
  assign new_new_n21355__ = ~new_new_n20862__ & ~new_new_n20863__;
  assign new_new_n21356__ = new_new_n20867__ & new_new_n21355__;
  assign new_new_n21357__ = ~new_new_n20867__ & ~new_new_n21355__;
  assign new_new_n21358__ = ~new_new_n21356__ & ~new_new_n21357__;
  assign new_new_n21359__ = ~new_new_n21354__ & ~new_new_n21358__;
  assign new_new_n21360__ = ~new_new_n21353__ & ~new_new_n21359__;
  assign new_new_n21361__ = ~new_new_n20466__ & ~new_new_n20467__;
  assign new_new_n21362__ = ~new_new_n20869__ & new_new_n21361__;
  assign new_new_n21363__ = new_new_n20869__ & ~new_new_n21361__;
  assign new_new_n21364__ = ~new_new_n21362__ & ~new_new_n21363__;
  assign new_new_n21365__ = ~new_new_n21360__ & ~new_new_n21364__;
  assign new_new_n21366__ = new_new_n21360__ & new_new_n21364__;
  assign new_new_n21367__ = new_new_n8474__ & new_new_n15905__;
  assign new_new_n21368__ = ~new_new_n8479__ & new_new_n15237__;
  assign new_new_n21369__ = new_new_n8470__ & new_new_n16025__;
  assign new_new_n21370__ = ~new_new_n21367__ & ~new_new_n21368__;
  assign new_new_n21371__ = ~new_new_n21369__ & new_new_n21370__;
  assign new_new_n21372__ = new_new_n8469__ & ~new_new_n15998__;
  assign new_new_n21373__ = pi11 & ~new_new_n21372__;
  assign new_new_n21374__ = new_new_n11368__ & ~new_new_n15998__;
  assign new_new_n21375__ = ~new_new_n21373__ & ~new_new_n21374__;
  assign new_new_n21376__ = new_new_n21371__ & ~new_new_n21375__;
  assign new_new_n21377__ = ~pi11 & ~new_new_n21371__;
  assign new_new_n21378__ = ~new_new_n21376__ & ~new_new_n21377__;
  assign new_new_n21379__ = ~new_new_n21366__ & ~new_new_n21378__;
  assign new_new_n21380__ = ~new_new_n21365__ & ~new_new_n21379__;
  assign new_new_n21381__ = new_new_n20883__ & ~new_new_n21380__;
  assign new_new_n21382__ = ~new_new_n20883__ & new_new_n21380__;
  assign new_new_n21383__ = ~new_new_n21381__ & ~new_new_n21382__;
  assign new_new_n21384__ = ~new_new_n11409__ & new_new_n15905__;
  assign new_new_n21385__ = new_new_n10702__ & ~new_new_n15998__;
  assign new_new_n21386__ = ~new_new_n10697__ & new_new_n16051__;
  assign new_new_n21387__ = new_new_n10694__ & ~new_new_n16056__;
  assign new_new_n21388__ = ~new_new_n21386__ & new_new_n21387__;
  assign new_new_n21389__ = ~new_new_n21384__ & ~new_new_n21385__;
  assign new_new_n21390__ = ~new_new_n21388__ & new_new_n21389__;
  assign new_new_n21391__ = pi08 & ~new_new_n21390__;
  assign new_new_n21392__ = ~pi08 & new_new_n21390__;
  assign new_new_n21393__ = ~new_new_n21391__ & ~new_new_n21392__;
  assign new_new_n21394__ = new_new_n8858__ & new_new_n15244__;
  assign new_new_n21395__ = new_new_n8474__ & ~new_new_n15248__;
  assign new_new_n21396__ = ~new_new_n8479__ & ~new_new_n15314__;
  assign new_new_n21397__ = ~new_new_n21395__ & ~new_new_n21396__;
  assign new_new_n21398__ = ~new_new_n21394__ & new_new_n21397__;
  assign new_new_n21399__ = new_new_n8469__ & new_new_n16378__;
  assign new_new_n21400__ = ~pi11 & ~new_new_n21399__;
  assign new_new_n21401__ = new_new_n11368__ & new_new_n16378__;
  assign new_new_n21402__ = ~new_new_n21400__ & ~new_new_n21401__;
  assign new_new_n21403__ = new_new_n21398__ & ~new_new_n21402__;
  assign new_new_n21404__ = pi11 & ~new_new_n21398__;
  assign new_new_n21405__ = ~new_new_n21403__ & ~new_new_n21404__;
  assign new_new_n21406__ = new_new_n6991__ & ~new_new_n15321__;
  assign new_new_n21407__ = new_new_n6985__ & ~new_new_n15273__;
  assign new_new_n21408__ = ~new_new_n21406__ & ~new_new_n21407__;
  assign new_new_n21409__ = new_new_n6994__ & new_new_n16079__;
  assign new_new_n21410__ = new_new_n21408__ & ~new_new_n21409__;
  assign new_new_n21411__ = pi14 & ~new_new_n21410__;
  assign new_new_n21412__ = new_new_n6994__ & ~new_new_n16088__;
  assign new_new_n21413__ = ~pi14 & new_new_n21408__;
  assign new_new_n21414__ = ~new_new_n21412__ & new_new_n21413__;
  assign new_new_n21415__ = pi13 & new_new_n16078__;
  assign new_new_n21416__ = ~new_new_n20898__ & ~new_new_n21415__;
  assign new_new_n21417__ = new_new_n21412__ & new_new_n21416__;
  assign new_new_n21418__ = ~new_new_n21414__ & ~new_new_n21417__;
  assign new_new_n21419__ = ~new_new_n21411__ & new_new_n21418__;
  assign new_new_n21420__ = new_new_n6968__ & new_new_n15390__;
  assign new_new_n21421__ = new_new_n6964__ & ~new_new_n15362__;
  assign new_new_n21422__ = ~new_new_n21420__ & ~new_new_n21421__;
  assign new_new_n21423__ = new_new_n6958__ & ~new_new_n17364__;
  assign new_new_n21424__ = pi17 & ~new_new_n21423__;
  assign new_new_n21425__ = ~pi16 & new_new_n15398__;
  assign new_new_n21426__ = pi16 & ~new_new_n15398__;
  assign new_new_n21427__ = new_new_n6958__ & ~new_new_n21425__;
  assign new_new_n21428__ = ~new_new_n21426__ & new_new_n21427__;
  assign new_new_n21429__ = new_new_n16956__ & new_new_n21428__;
  assign new_new_n21430__ = ~new_new_n21424__ & ~new_new_n21429__;
  assign new_new_n21431__ = new_new_n21422__ & ~new_new_n21430__;
  assign new_new_n21432__ = new_new_n6958__ & new_new_n17360__;
  assign new_new_n21433__ = new_new_n21422__ & ~new_new_n21432__;
  assign new_new_n21434__ = ~pi17 & ~new_new_n21433__;
  assign new_new_n21435__ = ~new_new_n21431__ & ~new_new_n21434__;
  assign new_new_n21436__ = ~new_new_n21321__ & ~new_new_n21322__;
  assign new_new_n21437__ = new_new_n21332__ & new_new_n21436__;
  assign new_new_n21438__ = ~new_new_n21332__ & ~new_new_n21436__;
  assign new_new_n21439__ = ~new_new_n21437__ & ~new_new_n21438__;
  assign new_new_n21440__ = ~new_new_n21435__ & ~new_new_n21439__;
  assign new_new_n21441__ = new_new_n21435__ & new_new_n21439__;
  assign new_new_n21442__ = new_new_n6629__ & ~new_new_n15471__;
  assign new_new_n21443__ = ~new_new_n6625__ & ~new_new_n15809__;
  assign new_new_n21444__ = new_new_n6634__ & new_new_n15464__;
  assign new_new_n21445__ = ~new_new_n21442__ & ~new_new_n21443__;
  assign new_new_n21446__ = ~new_new_n21444__ & new_new_n21445__;
  assign new_new_n21447__ = new_new_n6631__ & new_new_n15819__;
  assign new_new_n21448__ = pi20 & ~new_new_n21447__;
  assign new_new_n21449__ = new_new_n6640__ & new_new_n15819__;
  assign new_new_n21450__ = ~new_new_n21448__ & ~new_new_n21449__;
  assign new_new_n21451__ = new_new_n21446__ & ~new_new_n21450__;
  assign new_new_n21452__ = ~pi20 & ~new_new_n21446__;
  assign new_new_n21453__ = ~new_new_n21451__ & ~new_new_n21452__;
  assign new_new_n21454__ = new_new_n6629__ & ~new_new_n15809__;
  assign new_new_n21455__ = ~new_new_n6625__ & ~new_new_n15487__;
  assign new_new_n21456__ = new_new_n6634__ & ~new_new_n15471__;
  assign new_new_n21457__ = ~new_new_n21454__ & ~new_new_n21455__;
  assign new_new_n21458__ = ~new_new_n21456__ & new_new_n21457__;
  assign new_new_n21459__ = new_new_n6631__ & ~new_new_n18633__;
  assign new_new_n21460__ = ~pi20 & ~new_new_n21459__;
  assign new_new_n21461__ = new_new_n7015__ & ~new_new_n18633__;
  assign new_new_n21462__ = ~new_new_n21460__ & ~new_new_n21461__;
  assign new_new_n21463__ = new_new_n21458__ & ~new_new_n21462__;
  assign new_new_n21464__ = pi20 & ~new_new_n21458__;
  assign new_new_n21465__ = ~new_new_n21463__ & ~new_new_n21464__;
  assign new_new_n21466__ = new_new_n6634__ & ~new_new_n15487__;
  assign new_new_n21467__ = new_new_n6629__ & new_new_n15524__;
  assign new_new_n21468__ = ~new_new_n6625__ & new_new_n15520__;
  assign new_new_n21469__ = new_new_n6936__ & new_new_n17587__;
  assign new_new_n21470__ = ~new_new_n21467__ & ~new_new_n21468__;
  assign new_new_n21471__ = ~new_new_n21466__ & new_new_n21470__;
  assign new_new_n21472__ = ~new_new_n21469__ & new_new_n21471__;
  assign new_new_n21473__ = ~pi20 & ~new_new_n21472__;
  assign new_new_n21474__ = pi20 & new_new_n21472__;
  assign new_new_n21475__ = ~new_new_n21473__ & ~new_new_n21474__;
  assign new_new_n21476__ = new_new_n6629__ & new_new_n15520__;
  assign new_new_n21477__ = new_new_n15524__ & new_new_n18913__;
  assign new_new_n21478__ = new_new_n6936__ & ~new_new_n18914__;
  assign new_new_n21479__ = ~new_new_n21477__ & new_new_n21478__;
  assign new_new_n21480__ = ~new_new_n6625__ & ~new_new_n15533__;
  assign new_new_n21481__ = new_new_n6634__ & new_new_n15524__;
  assign new_new_n21482__ = ~new_new_n21480__ & ~new_new_n21481__;
  assign new_new_n21483__ = ~new_new_n21476__ & new_new_n21482__;
  assign new_new_n21484__ = ~new_new_n21479__ & new_new_n21483__;
  assign new_new_n21485__ = new_new_n6634__ & new_new_n15520__;
  assign new_new_n21486__ = new_new_n6629__ & ~new_new_n15533__;
  assign new_new_n21487__ = ~new_new_n6625__ & new_new_n15767__;
  assign new_new_n21488__ = new_new_n6936__ & new_new_n19731__;
  assign new_new_n21489__ = ~new_new_n21486__ & ~new_new_n21487__;
  assign new_new_n21490__ = ~new_new_n21485__ & new_new_n21489__;
  assign new_new_n21491__ = ~new_new_n21488__ & new_new_n21490__;
  assign new_new_n21492__ = ~pi20 & ~new_new_n21491__;
  assign new_new_n21493__ = ~new_new_n21237__ & ~new_new_n21238__;
  assign new_new_n21494__ = ~new_new_n21242__ & new_new_n21493__;
  assign new_new_n21495__ = new_new_n21242__ & ~new_new_n21493__;
  assign new_new_n21496__ = ~new_new_n21494__ & ~new_new_n21495__;
  assign new_new_n21497__ = new_new_n21491__ & ~new_new_n21496__;
  assign new_new_n21498__ = ~new_new_n21492__ & ~new_new_n21497__;
  assign new_new_n21499__ = ~new_new_n21484__ & ~new_new_n21498__;
  assign new_new_n21500__ = ~new_new_n21491__ & ~new_new_n21496__;
  assign new_new_n21501__ = new_new_n6629__ & new_new_n15767__;
  assign new_new_n21502__ = new_new_n6936__ & new_new_n19893__;
  assign new_new_n21503__ = ~new_new_n21501__ & ~new_new_n21502__;
  assign new_new_n21504__ = ~new_new_n6625__ & new_new_n15560__;
  assign new_new_n21505__ = new_new_n6634__ & ~new_new_n15533__;
  assign new_new_n21506__ = ~new_new_n21504__ & ~new_new_n21505__;
  assign new_new_n21507__ = new_new_n21503__ & new_new_n21506__;
  assign new_new_n21508__ = pi20 & ~new_new_n21507__;
  assign new_new_n21509__ = new_new_n6625__ & ~new_new_n21505__;
  assign new_new_n21510__ = ~new_new_n6634__ & ~new_new_n15560__;
  assign new_new_n21511__ = ~new_new_n21509__ & ~new_new_n21510__;
  assign new_new_n21512__ = ~pi20 & ~new_new_n21511__;
  assign new_new_n21513__ = new_new_n21503__ & new_new_n21512__;
  assign new_new_n21514__ = ~new_new_n21508__ & ~new_new_n21513__;
  assign new_new_n21515__ = ~new_new_n21168__ & ~new_new_n21169__;
  assign new_new_n21516__ = ~new_new_n21179__ & ~new_new_n21515__;
  assign new_new_n21517__ = new_new_n21179__ & new_new_n21515__;
  assign new_new_n21518__ = ~new_new_n21516__ & ~new_new_n21517__;
  assign new_new_n21519__ = ~new_new_n21150__ & ~new_new_n21151__;
  assign new_new_n21520__ = ~new_new_n21161__ & new_new_n21519__;
  assign new_new_n21521__ = new_new_n21161__ & ~new_new_n21519__;
  assign new_new_n21522__ = ~new_new_n21520__ & ~new_new_n21521__;
  assign new_new_n21523__ = new_new_n6936__ & new_new_n18512__;
  assign new_new_n21524__ = new_new_n6629__ & ~new_new_n15615__;
  assign new_new_n21525__ = ~new_new_n6625__ & new_new_n15743__;
  assign new_new_n21526__ = new_new_n6634__ & new_new_n15564__;
  assign new_new_n21527__ = ~new_new_n21524__ & ~new_new_n21525__;
  assign new_new_n21528__ = ~new_new_n21526__ & new_new_n21527__;
  assign new_new_n21529__ = ~new_new_n21523__ & new_new_n21528__;
  assign new_new_n21530__ = ~pi20 & ~new_new_n21529__;
  assign new_new_n21531__ = pi20 & new_new_n21529__;
  assign new_new_n21532__ = ~new_new_n21530__ & ~new_new_n21531__;
  assign new_new_n21533__ = ~new_new_n21133__ & ~new_new_n21138__;
  assign new_new_n21534__ = new_new_n20611__ & new_new_n20672__;
  assign new_new_n21535__ = ~new_new_n20611__ & ~new_new_n20672__;
  assign new_new_n21536__ = ~new_new_n21534__ & ~new_new_n21535__;
  assign new_new_n21537__ = new_new_n20678__ & ~new_new_n21536__;
  assign new_new_n21538__ = new_new_n20680__ & new_new_n21536__;
  assign new_new_n21539__ = new_new_n20679__ & new_new_n21534__;
  assign new_new_n21540__ = ~new_new_n21537__ & ~new_new_n21539__;
  assign new_new_n21541__ = ~new_new_n21538__ & new_new_n21540__;
  assign new_new_n21542__ = ~new_new_n21533__ & ~new_new_n21541__;
  assign new_new_n21543__ = ~new_new_n20678__ & ~new_new_n21534__;
  assign new_new_n21544__ = ~new_new_n20679__ & ~new_new_n21543__;
  assign new_new_n21545__ = ~new_new_n21537__ & new_new_n21544__;
  assign new_new_n21546__ = new_new_n21533__ & new_new_n21545__;
  assign new_new_n21547__ = ~new_new_n20611__ & new_new_n21132__;
  assign new_new_n21548__ = new_new_n21136__ & new_new_n21547__;
  assign new_new_n21549__ = ~new_new_n21134__ & ~new_new_n21135__;
  assign new_new_n21550__ = ~new_new_n20611__ & new_new_n21549__;
  assign new_new_n21551__ = ~new_new_n21136__ & ~new_new_n21550__;
  assign new_new_n21552__ = new_new_n20210__ & ~new_new_n21551__;
  assign new_new_n21553__ = new_new_n21533__ & new_new_n21552__;
  assign new_new_n21554__ = ~new_new_n21542__ & ~new_new_n21548__;
  assign new_new_n21555__ = ~new_new_n21546__ & ~new_new_n21553__;
  assign new_new_n21556__ = new_new_n21554__ & new_new_n21555__;
  assign new_new_n21557__ = new_new_n21532__ & ~new_new_n21556__;
  assign new_new_n21558__ = ~new_new_n21532__ & new_new_n21556__;
  assign new_new_n21559__ = new_new_n6629__ & ~new_new_n15638__;
  assign new_new_n21560__ = ~new_new_n6625__ & ~new_new_n15582__;
  assign new_new_n21561__ = new_new_n6634__ & new_new_n15743__;
  assign new_new_n21562__ = ~new_new_n21559__ & ~new_new_n21560__;
  assign new_new_n21563__ = ~new_new_n21561__ & new_new_n21562__;
  assign new_new_n21564__ = new_new_n6631__ & new_new_n19494__;
  assign new_new_n21565__ = pi20 & ~new_new_n21564__;
  assign new_new_n21566__ = new_new_n6640__ & new_new_n19494__;
  assign new_new_n21567__ = ~new_new_n21565__ & ~new_new_n21566__;
  assign new_new_n21568__ = new_new_n21563__ & ~new_new_n21567__;
  assign new_new_n21569__ = ~pi20 & ~new_new_n21563__;
  assign new_new_n21570__ = ~new_new_n21568__ & ~new_new_n21569__;
  assign new_new_n21571__ = ~new_new_n21108__ & ~new_new_n21109__;
  assign new_new_n21572__ = ~new_new_n21119__ & new_new_n21571__;
  assign new_new_n21573__ = new_new_n21119__ & ~new_new_n21571__;
  assign new_new_n21574__ = ~new_new_n21572__ & ~new_new_n21573__;
  assign new_new_n21575__ = ~new_new_n21062__ & ~new_new_n21102__;
  assign new_new_n21576__ = new_new_n21062__ & new_new_n21102__;
  assign new_new_n21577__ = ~new_new_n21575__ & ~new_new_n21576__;
  assign new_new_n21578__ = new_new_n21063__ & ~new_new_n21577__;
  assign new_new_n21579__ = new_new_n21078__ & new_new_n21575__;
  assign new_new_n21580__ = ~new_new_n21578__ & ~new_new_n21579__;
  assign new_new_n21581__ = new_new_n21093__ & ~new_new_n21580__;
  assign new_new_n21582__ = ~new_new_n21094__ & new_new_n21577__;
  assign new_new_n21583__ = ~new_new_n21581__ & ~new_new_n21582__;
  assign new_new_n21584__ = new_new_n6936__ & ~new_new_n19118__;
  assign new_new_n21585__ = new_new_n6629__ & ~new_new_n15710__;
  assign new_new_n21586__ = ~new_new_n6625__ & new_new_n15656__;
  assign new_new_n21587__ = new_new_n6634__ & ~new_new_n15647__;
  assign new_new_n21588__ = ~new_new_n21585__ & ~new_new_n21586__;
  assign new_new_n21589__ = ~new_new_n21587__ & new_new_n21588__;
  assign new_new_n21590__ = ~new_new_n21584__ & new_new_n21589__;
  assign new_new_n21591__ = ~pi20 & ~new_new_n21590__;
  assign new_new_n21592__ = pi20 & new_new_n21590__;
  assign new_new_n21593__ = ~new_new_n21591__ & ~new_new_n21592__;
  assign new_new_n21594__ = pi23 & ~new_new_n21067__;
  assign new_new_n21595__ = ~new_new_n21076__ & new_new_n21594__;
  assign new_new_n21596__ = new_new_n21076__ & ~new_new_n21594__;
  assign new_new_n21597__ = ~new_new_n21595__ & ~new_new_n21596__;
  assign new_new_n21598__ = new_new_n6629__ & ~new_new_n15661__;
  assign new_new_n21599__ = ~new_new_n6625__ & new_new_n15668__;
  assign new_new_n21600__ = ~new_new_n21598__ & ~new_new_n21599__;
  assign new_new_n21601__ = new_new_n6631__ & new_new_n20187__;
  assign new_new_n21602__ = new_new_n21600__ & ~new_new_n21601__;
  assign new_new_n21603__ = pi20 & ~new_new_n21602__;
  assign new_new_n21604__ = new_new_n6631__ & ~new_new_n20177__;
  assign new_new_n21605__ = ~pi20 & ~new_new_n21604__;
  assign new_new_n21606__ = ~pi19 & new_new_n15643__;
  assign new_new_n21607__ = pi19 & ~new_new_n15643__;
  assign new_new_n21608__ = new_new_n6631__ & new_new_n20176__;
  assign new_new_n21609__ = ~new_new_n21606__ & new_new_n21608__;
  assign new_new_n21610__ = ~new_new_n21607__ & new_new_n21609__;
  assign new_new_n21611__ = ~new_new_n21605__ & ~new_new_n21610__;
  assign new_new_n21612__ = new_new_n21600__ & ~new_new_n21611__;
  assign new_new_n21613__ = ~new_new_n21603__ & ~new_new_n21612__;
  assign new_new_n21614__ = new_new_n5195__ & ~new_new_n15673__;
  assign new_new_n21615__ = new_new_n6631__ & new_new_n15668__;
  assign new_new_n21616__ = new_new_n15673__ & ~new_new_n21615__;
  assign new_new_n21617__ = new_new_n9921__ & ~new_new_n21616__;
  assign new_new_n21618__ = pi20 & ~new_new_n21617__;
  assign new_new_n21619__ = new_new_n6629__ & new_new_n15668__;
  assign new_new_n21620__ = ~new_new_n6625__ & ~new_new_n15673__;
  assign new_new_n21621__ = ~new_new_n6633__ & new_new_n20195__;
  assign new_new_n21622__ = new_new_n15661__ & ~new_new_n21621__;
  assign new_new_n21623__ = ~new_new_n15661__ & new_new_n21621__;
  assign new_new_n21624__ = new_new_n6631__ & ~new_new_n21622__;
  assign new_new_n21625__ = ~new_new_n21623__ & new_new_n21624__;
  assign new_new_n21626__ = ~new_new_n21620__ & ~new_new_n21625__;
  assign new_new_n21627__ = ~new_new_n21619__ & new_new_n21626__;
  assign new_new_n21628__ = pi20 & ~new_new_n21627__;
  assign new_new_n21629__ = new_new_n6625__ & ~new_new_n15668__;
  assign new_new_n21630__ = new_new_n6629__ & ~new_new_n21629__;
  assign new_new_n21631__ = ~pi20 & ~new_new_n21630__;
  assign new_new_n21632__ = new_new_n21626__ & new_new_n21631__;
  assign new_new_n21633__ = ~new_new_n21628__ & ~new_new_n21632__;
  assign new_new_n21634__ = new_new_n21618__ & new_new_n21633__;
  assign new_new_n21635__ = ~new_new_n21614__ & ~new_new_n21634__;
  assign new_new_n21636__ = new_new_n21613__ & ~new_new_n21635__;
  assign new_new_n21637__ = new_new_n5180__ & new_new_n15674__;
  assign new_new_n21638__ = ~new_new_n5195__ & new_new_n20195__;
  assign new_new_n21639__ = ~new_new_n5179__ & new_new_n15668__;
  assign new_new_n21640__ = new_new_n5182__ & ~new_new_n21639__;
  assign new_new_n21641__ = ~new_new_n5189__ & ~new_new_n20628__;
  assign new_new_n21642__ = ~new_new_n21637__ & new_new_n21641__;
  assign new_new_n21643__ = ~new_new_n21638__ & ~new_new_n21640__;
  assign new_new_n21644__ = new_new_n21642__ & new_new_n21643__;
  assign new_new_n21645__ = ~new_new_n21636__ & ~new_new_n21644__;
  assign new_new_n21646__ = new_new_n21636__ & new_new_n21644__;
  assign new_new_n21647__ = new_new_n6634__ & new_new_n15656__;
  assign new_new_n21648__ = ~new_new_n6625__ & ~new_new_n15661__;
  assign new_new_n21649__ = new_new_n6629__ & new_new_n15643__;
  assign new_new_n21650__ = new_new_n6936__ & new_new_n15687__;
  assign new_new_n21651__ = ~new_new_n21648__ & ~new_new_n21649__;
  assign new_new_n21652__ = ~new_new_n21647__ & new_new_n21651__;
  assign new_new_n21653__ = ~new_new_n21650__ & new_new_n21652__;
  assign new_new_n21654__ = pi20 & ~new_new_n21653__;
  assign new_new_n21655__ = ~pi20 & new_new_n21653__;
  assign new_new_n21656__ = ~new_new_n21654__ & ~new_new_n21655__;
  assign new_new_n21657__ = ~new_new_n21646__ & ~new_new_n21656__;
  assign new_new_n21658__ = ~new_new_n21645__ & ~new_new_n21657__;
  assign new_new_n21659__ = new_new_n21597__ & new_new_n21658__;
  assign new_new_n21660__ = ~new_new_n21597__ & ~new_new_n21658__;
  assign new_new_n21661__ = new_new_n6634__ & ~new_new_n15710__;
  assign new_new_n21662__ = ~new_new_n6625__ & new_new_n15643__;
  assign new_new_n21663__ = new_new_n6629__ & new_new_n15656__;
  assign new_new_n21664__ = new_new_n6936__ & ~new_new_n19466__;
  assign new_new_n21665__ = ~new_new_n21662__ & ~new_new_n21663__;
  assign new_new_n21666__ = ~new_new_n21661__ & new_new_n21665__;
  assign new_new_n21667__ = ~new_new_n21664__ & new_new_n21666__;
  assign new_new_n21668__ = pi20 & ~new_new_n21667__;
  assign new_new_n21669__ = ~pi20 & new_new_n21667__;
  assign new_new_n21670__ = ~new_new_n21668__ & ~new_new_n21669__;
  assign new_new_n21671__ = ~new_new_n21660__ & new_new_n21670__;
  assign new_new_n21672__ = ~new_new_n21659__ & ~new_new_n21671__;
  assign new_new_n21673__ = ~new_new_n21593__ & ~new_new_n21672__;
  assign new_new_n21674__ = new_new_n21593__ & new_new_n21672__;
  assign new_new_n21675__ = ~new_new_n21063__ & ~new_new_n21093__;
  assign new_new_n21676__ = ~new_new_n21094__ & ~new_new_n21675__;
  assign new_new_n21677__ = ~new_new_n21674__ & new_new_n21676__;
  assign new_new_n21678__ = ~new_new_n21063__ & new_new_n21093__;
  assign new_new_n21679__ = new_new_n21078__ & ~new_new_n21678__;
  assign new_new_n21680__ = ~new_new_n21593__ & new_new_n21679__;
  assign new_new_n21681__ = ~new_new_n21673__ & ~new_new_n21680__;
  assign new_new_n21682__ = ~new_new_n21677__ & new_new_n21681__;
  assign new_new_n21683__ = new_new_n21583__ & ~new_new_n21682__;
  assign new_new_n21684__ = ~new_new_n21583__ & new_new_n21682__;
  assign new_new_n21685__ = new_new_n6634__ & ~new_new_n15582__;
  assign new_new_n21686__ = ~new_new_n6625__ & ~new_new_n15710__;
  assign new_new_n21687__ = new_new_n6629__ & ~new_new_n15647__;
  assign new_new_n21688__ = new_new_n6936__ & ~new_new_n15736__;
  assign new_new_n21689__ = ~new_new_n21686__ & ~new_new_n21687__;
  assign new_new_n21690__ = ~new_new_n21685__ & new_new_n21689__;
  assign new_new_n21691__ = ~new_new_n21688__ & new_new_n21690__;
  assign new_new_n21692__ = pi20 & ~new_new_n21691__;
  assign new_new_n21693__ = ~pi20 & new_new_n21691__;
  assign new_new_n21694__ = ~new_new_n21692__ & ~new_new_n21693__;
  assign new_new_n21695__ = ~new_new_n21684__ & new_new_n21694__;
  assign new_new_n21696__ = ~new_new_n21683__ & ~new_new_n21695__;
  assign new_new_n21697__ = new_new_n21574__ & new_new_n21696__;
  assign new_new_n21698__ = ~new_new_n21574__ & ~new_new_n21696__;
  assign new_new_n21699__ = new_new_n6634__ & ~new_new_n15638__;
  assign new_new_n21700__ = ~new_new_n6625__ & ~new_new_n15647__;
  assign new_new_n21701__ = new_new_n6629__ & ~new_new_n15582__;
  assign new_new_n21702__ = new_new_n6936__ & new_new_n19487__;
  assign new_new_n21703__ = ~new_new_n21700__ & ~new_new_n21701__;
  assign new_new_n21704__ = ~new_new_n21699__ & new_new_n21703__;
  assign new_new_n21705__ = ~new_new_n21702__ & new_new_n21704__;
  assign new_new_n21706__ = ~pi20 & ~new_new_n21705__;
  assign new_new_n21707__ = pi20 & new_new_n21705__;
  assign new_new_n21708__ = ~new_new_n21706__ & ~new_new_n21707__;
  assign new_new_n21709__ = ~new_new_n21698__ & new_new_n21708__;
  assign new_new_n21710__ = ~new_new_n21697__ & ~new_new_n21709__;
  assign new_new_n21711__ = ~new_new_n21570__ & new_new_n21710__;
  assign new_new_n21712__ = new_new_n21570__ & ~new_new_n21710__;
  assign new_new_n21713__ = ~new_new_n21122__ & ~new_new_n21123__;
  assign new_new_n21714__ = new_new_n21128__ & new_new_n21713__;
  assign new_new_n21715__ = ~new_new_n21128__ & ~new_new_n21713__;
  assign new_new_n21716__ = ~new_new_n21714__ & ~new_new_n21715__;
  assign new_new_n21717__ = ~new_new_n21712__ & new_new_n21716__;
  assign new_new_n21718__ = ~new_new_n21711__ & ~new_new_n21717__;
  assign new_new_n21719__ = ~new_new_n21033__ & ~new_new_n21034__;
  assign new_new_n21720__ = ~new_new_n21130__ & new_new_n21719__;
  assign new_new_n21721__ = new_new_n21130__ & ~new_new_n21719__;
  assign new_new_n21722__ = ~new_new_n21720__ & ~new_new_n21721__;
  assign new_new_n21723__ = new_new_n21718__ & ~new_new_n21722__;
  assign new_new_n21724__ = ~new_new_n21718__ & new_new_n21722__;
  assign new_new_n21725__ = new_new_n6629__ & new_new_n15743__;
  assign new_new_n21726__ = ~new_new_n6625__ & ~new_new_n15638__;
  assign new_new_n21727__ = new_new_n6634__ & ~new_new_n15615__;
  assign new_new_n21728__ = ~new_new_n21725__ & ~new_new_n21726__;
  assign new_new_n21729__ = ~new_new_n21727__ & new_new_n21728__;
  assign new_new_n21730__ = new_new_n6631__ & new_new_n19005__;
  assign new_new_n21731__ = pi20 & ~new_new_n21730__;
  assign new_new_n21732__ = new_new_n6640__ & new_new_n19005__;
  assign new_new_n21733__ = ~new_new_n21731__ & ~new_new_n21732__;
  assign new_new_n21734__ = new_new_n21729__ & ~new_new_n21733__;
  assign new_new_n21735__ = ~pi20 & ~new_new_n21729__;
  assign new_new_n21736__ = ~new_new_n21734__ & ~new_new_n21735__;
  assign new_new_n21737__ = ~new_new_n21724__ & new_new_n21736__;
  assign new_new_n21738__ = ~new_new_n21723__ & ~new_new_n21737__;
  assign new_new_n21739__ = ~new_new_n21558__ & ~new_new_n21738__;
  assign new_new_n21740__ = ~new_new_n21557__ & ~new_new_n21739__;
  assign new_new_n21741__ = ~new_new_n21522__ & ~new_new_n21740__;
  assign new_new_n21742__ = new_new_n21522__ & new_new_n21740__;
  assign new_new_n21743__ = new_new_n6634__ & new_new_n15572__;
  assign new_new_n21744__ = ~new_new_n6625__ & ~new_new_n15615__;
  assign new_new_n21745__ = new_new_n6629__ & new_new_n15564__;
  assign new_new_n21746__ = new_new_n6936__ & ~new_new_n20114__;
  assign new_new_n21747__ = ~new_new_n21744__ & ~new_new_n21745__;
  assign new_new_n21748__ = ~new_new_n21743__ & new_new_n21747__;
  assign new_new_n21749__ = ~new_new_n21746__ & new_new_n21748__;
  assign new_new_n21750__ = pi20 & ~new_new_n21749__;
  assign new_new_n21751__ = ~pi20 & new_new_n21749__;
  assign new_new_n21752__ = ~new_new_n21750__ & ~new_new_n21751__;
  assign new_new_n21753__ = ~new_new_n21742__ & ~new_new_n21752__;
  assign new_new_n21754__ = ~new_new_n21741__ & ~new_new_n21753__;
  assign new_new_n21755__ = ~new_new_n21518__ & ~new_new_n21754__;
  assign new_new_n21756__ = new_new_n21518__ & new_new_n21754__;
  assign new_new_n21757__ = new_new_n6634__ & new_new_n15560__;
  assign new_new_n21758__ = ~new_new_n6625__ & new_new_n15564__;
  assign new_new_n21759__ = new_new_n6629__ & new_new_n15572__;
  assign new_new_n21760__ = new_new_n6936__ & new_new_n18944__;
  assign new_new_n21761__ = ~new_new_n21758__ & ~new_new_n21759__;
  assign new_new_n21762__ = ~new_new_n21757__ & new_new_n21761__;
  assign new_new_n21763__ = ~new_new_n21760__ & new_new_n21762__;
  assign new_new_n21764__ = ~pi20 & ~new_new_n21763__;
  assign new_new_n21765__ = pi20 & new_new_n21763__;
  assign new_new_n21766__ = ~new_new_n21764__ & ~new_new_n21765__;
  assign new_new_n21767__ = ~new_new_n21756__ & new_new_n21766__;
  assign new_new_n21768__ = ~new_new_n21755__ & ~new_new_n21767__;
  assign new_new_n21769__ = ~new_new_n21182__ & ~new_new_n21183__;
  assign new_new_n21770__ = ~new_new_n21193__ & new_new_n21769__;
  assign new_new_n21771__ = new_new_n21193__ & ~new_new_n21769__;
  assign new_new_n21772__ = ~new_new_n21770__ & ~new_new_n21771__;
  assign new_new_n21773__ = new_new_n21768__ & ~new_new_n21772__;
  assign new_new_n21774__ = ~new_new_n21768__ & new_new_n21772__;
  assign new_new_n21775__ = new_new_n6629__ & new_new_n15560__;
  assign new_new_n21776__ = new_new_n6634__ & new_new_n15767__;
  assign new_new_n21777__ = ~new_new_n6625__ & new_new_n15572__;
  assign new_new_n21778__ = new_new_n6936__ & ~new_new_n18454__;
  assign new_new_n21779__ = ~new_new_n21776__ & ~new_new_n21777__;
  assign new_new_n21780__ = ~new_new_n21775__ & new_new_n21779__;
  assign new_new_n21781__ = ~new_new_n21778__ & new_new_n21780__;
  assign new_new_n21782__ = ~pi20 & ~new_new_n21781__;
  assign new_new_n21783__ = pi20 & new_new_n21781__;
  assign new_new_n21784__ = ~new_new_n21782__ & ~new_new_n21783__;
  assign new_new_n21785__ = ~new_new_n21774__ & ~new_new_n21784__;
  assign new_new_n21786__ = ~new_new_n21773__ & ~new_new_n21785__;
  assign new_new_n21787__ = ~new_new_n21514__ & new_new_n21786__;
  assign new_new_n21788__ = new_new_n21514__ & ~new_new_n21786__;
  assign new_new_n21789__ = ~new_new_n21196__ & ~new_new_n21213__;
  assign new_new_n21790__ = new_new_n21212__ & new_new_n21789__;
  assign new_new_n21791__ = ~new_new_n21212__ & ~new_new_n21789__;
  assign new_new_n21792__ = ~new_new_n21790__ & ~new_new_n21791__;
  assign new_new_n21793__ = ~new_new_n21788__ & new_new_n21792__;
  assign new_new_n21794__ = ~new_new_n21787__ & ~new_new_n21793__;
  assign new_new_n21795__ = ~new_new_n21491__ & ~new_new_n21794__;
  assign new_new_n21796__ = pi20 & ~new_new_n21795__;
  assign new_new_n21797__ = ~new_new_n21500__ & ~new_new_n21796__;
  assign new_new_n21798__ = new_new_n21484__ & ~new_new_n21797__;
  assign new_new_n21799__ = ~pi20 & ~new_new_n21484__;
  assign new_new_n21800__ = new_new_n21496__ & ~new_new_n21799__;
  assign new_new_n21801__ = new_new_n21794__ & ~new_new_n21800__;
  assign new_new_n21802__ = ~new_new_n21499__ & ~new_new_n21801__;
  assign new_new_n21803__ = ~new_new_n21798__ & new_new_n21802__;
  assign new_new_n21804__ = ~new_new_n21223__ & ~new_new_n21224__;
  assign new_new_n21805__ = new_new_n21234__ & new_new_n21804__;
  assign new_new_n21806__ = ~new_new_n21234__ & ~new_new_n21804__;
  assign new_new_n21807__ = ~new_new_n21805__ & ~new_new_n21806__;
  assign new_new_n21808__ = ~new_new_n21803__ & new_new_n21807__;
  assign new_new_n21809__ = pi20 & ~new_new_n21496__;
  assign new_new_n21810__ = pi20 & new_new_n21491__;
  assign new_new_n21811__ = ~new_new_n21500__ & ~new_new_n21810__;
  assign new_new_n21812__ = new_new_n21794__ & ~new_new_n21811__;
  assign new_new_n21813__ = ~new_new_n21809__ & ~new_new_n21812__;
  assign new_new_n21814__ = new_new_n21484__ & ~new_new_n21813__;
  assign new_new_n21815__ = ~pi20 & ~new_new_n21496__;
  assign new_new_n21816__ = ~new_new_n21498__ & new_new_n21794__;
  assign new_new_n21817__ = ~new_new_n21815__ & ~new_new_n21816__;
  assign new_new_n21818__ = ~new_new_n21484__ & ~new_new_n21817__;
  assign new_new_n21819__ = ~new_new_n21814__ & ~new_new_n21818__;
  assign new_new_n21820__ = ~new_new_n21808__ & new_new_n21819__;
  assign new_new_n21821__ = new_new_n21475__ & new_new_n21820__;
  assign new_new_n21822__ = ~new_new_n21475__ & ~new_new_n21820__;
  assign new_new_n21823__ = ~new_new_n21249__ & ~new_new_n21250__;
  assign new_new_n21824__ = new_new_n21262__ & ~new_new_n21823__;
  assign new_new_n21825__ = ~new_new_n21262__ & new_new_n21823__;
  assign new_new_n21826__ = ~new_new_n21824__ & ~new_new_n21825__;
  assign new_new_n21827__ = ~new_new_n21822__ & new_new_n21826__;
  assign new_new_n21828__ = ~new_new_n21821__ & ~new_new_n21827__;
  assign new_new_n21829__ = ~new_new_n20967__ & ~new_new_n20968__;
  assign new_new_n21830__ = new_new_n21264__ & new_new_n21829__;
  assign new_new_n21831__ = ~new_new_n21264__ & ~new_new_n21829__;
  assign new_new_n21832__ = ~new_new_n21830__ & ~new_new_n21831__;
  assign new_new_n21833__ = ~new_new_n21828__ & ~new_new_n21832__;
  assign new_new_n21834__ = new_new_n21828__ & new_new_n21832__;
  assign new_new_n21835__ = new_new_n6634__ & ~new_new_n15809__;
  assign new_new_n21836__ = ~new_new_n6625__ & new_new_n15524__;
  assign new_new_n21837__ = new_new_n6629__ & ~new_new_n15487__;
  assign new_new_n21838__ = new_new_n6936__ & new_new_n18020__;
  assign new_new_n21839__ = ~new_new_n21836__ & ~new_new_n21837__;
  assign new_new_n21840__ = ~new_new_n21835__ & new_new_n21839__;
  assign new_new_n21841__ = ~new_new_n21838__ & new_new_n21840__;
  assign new_new_n21842__ = pi20 & ~new_new_n21841__;
  assign new_new_n21843__ = ~pi20 & new_new_n21841__;
  assign new_new_n21844__ = ~new_new_n21842__ & ~new_new_n21843__;
  assign new_new_n21845__ = ~new_new_n21834__ & ~new_new_n21844__;
  assign new_new_n21846__ = ~new_new_n21833__ & ~new_new_n21845__;
  assign new_new_n21847__ = ~new_new_n21465__ & ~new_new_n21846__;
  assign new_new_n21848__ = new_new_n21465__ & new_new_n21846__;
  assign new_new_n21849__ = ~new_new_n21271__ & ~new_new_n21288__;
  assign new_new_n21850__ = new_new_n21287__ & new_new_n21849__;
  assign new_new_n21851__ = ~new_new_n21287__ & ~new_new_n21849__;
  assign new_new_n21852__ = ~new_new_n21850__ & ~new_new_n21851__;
  assign new_new_n21853__ = ~new_new_n21848__ & ~new_new_n21852__;
  assign new_new_n21854__ = ~new_new_n21847__ & ~new_new_n21853__;
  assign new_new_n21855__ = new_new_n21453__ & ~new_new_n21854__;
  assign new_new_n21856__ = ~new_new_n21453__ & new_new_n21854__;
  assign new_new_n21857__ = ~new_new_n21295__ & ~new_new_n21296__;
  assign new_new_n21858__ = ~new_new_n21306__ & new_new_n21857__;
  assign new_new_n21859__ = new_new_n21306__ & ~new_new_n21857__;
  assign new_new_n21860__ = ~new_new_n21858__ & ~new_new_n21859__;
  assign new_new_n21861__ = ~new_new_n21856__ & ~new_new_n21860__;
  assign new_new_n21862__ = ~new_new_n21855__ & ~new_new_n21861__;
  assign new_new_n21863__ = ~new_new_n21309__ & ~new_new_n21310__;
  assign new_new_n21864__ = ~new_new_n21314__ & new_new_n21863__;
  assign new_new_n21865__ = new_new_n21314__ & ~new_new_n21863__;
  assign new_new_n21866__ = ~new_new_n21864__ & ~new_new_n21865__;
  assign new_new_n21867__ = ~new_new_n21862__ & ~new_new_n21866__;
  assign new_new_n21868__ = new_new_n21862__ & new_new_n21866__;
  assign new_new_n21869__ = new_new_n6629__ & new_new_n15464__;
  assign new_new_n21870__ = ~new_new_n6625__ & ~new_new_n15471__;
  assign new_new_n21871__ = new_new_n6634__ & ~new_new_n15439__;
  assign new_new_n21872__ = ~new_new_n21869__ & ~new_new_n21870__;
  assign new_new_n21873__ = ~new_new_n21871__ & new_new_n21872__;
  assign new_new_n21874__ = new_new_n6631__ & ~new_new_n17240__;
  assign new_new_n21875__ = ~pi20 & ~new_new_n21874__;
  assign new_new_n21876__ = new_new_n7015__ & ~new_new_n17240__;
  assign new_new_n21877__ = ~new_new_n21875__ & ~new_new_n21876__;
  assign new_new_n21878__ = new_new_n21873__ & ~new_new_n21877__;
  assign new_new_n21879__ = pi20 & ~new_new_n21873__;
  assign new_new_n21880__ = ~new_new_n21878__ & ~new_new_n21879__;
  assign new_new_n21881__ = ~new_new_n21868__ & ~new_new_n21880__;
  assign new_new_n21882__ = ~new_new_n21867__ & ~new_new_n21881__;
  assign new_new_n21883__ = ~new_new_n21441__ & new_new_n21882__;
  assign new_new_n21884__ = ~new_new_n21440__ & ~new_new_n21883__;
  assign new_new_n21885__ = ~new_new_n21419__ & new_new_n21884__;
  assign new_new_n21886__ = new_new_n21419__ & ~new_new_n21884__;
  assign new_new_n21887__ = ~new_new_n21885__ & ~new_new_n21886__;
  assign new_new_n21888__ = ~new_new_n21335__ & ~new_new_n21336__;
  assign new_new_n21889__ = ~new_new_n21348__ & new_new_n21888__;
  assign new_new_n21890__ = new_new_n21348__ & ~new_new_n21888__;
  assign new_new_n21891__ = ~new_new_n21889__ & ~new_new_n21890__;
  assign new_new_n21892__ = new_new_n21887__ & ~new_new_n21891__;
  assign new_new_n21893__ = ~new_new_n21887__ & new_new_n21891__;
  assign new_new_n21894__ = ~new_new_n21892__ & ~new_new_n21893__;
  assign new_new_n21895__ = new_new_n21405__ & ~new_new_n21894__;
  assign new_new_n21896__ = ~new_new_n21405__ & new_new_n21894__;
  assign new_new_n21897__ = ~new_new_n21855__ & ~new_new_n21856__;
  assign new_new_n21898__ = ~new_new_n21860__ & new_new_n21897__;
  assign new_new_n21899__ = new_new_n21860__ & ~new_new_n21897__;
  assign new_new_n21900__ = ~new_new_n21898__ & ~new_new_n21899__;
  assign new_new_n21901__ = new_new_n7935__ & ~new_new_n15432__;
  assign new_new_n21902__ = new_new_n6964__ & new_new_n15464__;
  assign new_new_n21903__ = new_new_n6968__ & ~new_new_n15439__;
  assign new_new_n21904__ = ~new_new_n21902__ & ~new_new_n21903__;
  assign new_new_n21905__ = ~new_new_n21901__ & new_new_n21904__;
  assign new_new_n21906__ = new_new_n6958__ & new_new_n17204__;
  assign new_new_n21907__ = ~pi17 & ~new_new_n21906__;
  assign new_new_n21908__ = new_new_n8160__ & new_new_n17204__;
  assign new_new_n21909__ = ~new_new_n21907__ & ~new_new_n21908__;
  assign new_new_n21910__ = new_new_n21905__ & ~new_new_n21909__;
  assign new_new_n21911__ = pi17 & ~new_new_n21905__;
  assign new_new_n21912__ = ~new_new_n21910__ & ~new_new_n21911__;
  assign new_new_n21913__ = new_new_n6959__ & ~new_new_n17240__;
  assign new_new_n21914__ = new_new_n6964__ & ~new_new_n15471__;
  assign new_new_n21915__ = new_new_n6968__ & new_new_n15464__;
  assign new_new_n21916__ = ~new_new_n21914__ & ~new_new_n21915__;
  assign new_new_n21917__ = ~new_new_n21913__ & new_new_n21916__;
  assign new_new_n21918__ = new_new_n6958__ & ~new_new_n15439__;
  assign new_new_n21919__ = pi17 & ~new_new_n21918__;
  assign new_new_n21920__ = new_new_n8160__ & ~new_new_n15439__;
  assign new_new_n21921__ = ~new_new_n21919__ & ~new_new_n21920__;
  assign new_new_n21922__ = new_new_n21917__ & ~new_new_n21921__;
  assign new_new_n21923__ = ~pi17 & ~new_new_n21917__;
  assign new_new_n21924__ = ~new_new_n21922__ & ~new_new_n21923__;
  assign new_new_n21925__ = ~new_new_n21833__ & ~new_new_n21834__;
  assign new_new_n21926__ = ~new_new_n21844__ & new_new_n21925__;
  assign new_new_n21927__ = new_new_n21844__ & ~new_new_n21925__;
  assign new_new_n21928__ = ~new_new_n21926__ & ~new_new_n21927__;
  assign new_new_n21929__ = ~new_new_n21924__ & ~new_new_n21928__;
  assign new_new_n21930__ = new_new_n21924__ & new_new_n21928__;
  assign new_new_n21931__ = new_new_n7935__ & new_new_n15464__;
  assign new_new_n21932__ = new_new_n6968__ & ~new_new_n15471__;
  assign new_new_n21933__ = new_new_n6959__ & new_new_n15819__;
  assign new_new_n21934__ = ~new_new_n21931__ & ~new_new_n21932__;
  assign new_new_n21935__ = ~new_new_n21933__ & new_new_n21934__;
  assign new_new_n21936__ = new_new_n10337__ & ~new_new_n15809__;
  assign new_new_n21937__ = pi17 & ~new_new_n21936__;
  assign new_new_n21938__ = new_new_n10340__ & ~new_new_n15809__;
  assign new_new_n21939__ = ~pi17 & ~new_new_n21938__;
  assign new_new_n21940__ = pi14 & ~new_new_n21939__;
  assign new_new_n21941__ = ~new_new_n21937__ & ~new_new_n21940__;
  assign new_new_n21942__ = new_new_n21935__ & ~new_new_n21941__;
  assign new_new_n21943__ = ~pi17 & ~new_new_n21935__;
  assign new_new_n21944__ = ~new_new_n21942__ & ~new_new_n21943__;
  assign new_new_n21945__ = ~new_new_n21821__ & ~new_new_n21822__;
  assign new_new_n21946__ = new_new_n21826__ & new_new_n21945__;
  assign new_new_n21947__ = ~new_new_n21826__ & ~new_new_n21945__;
  assign new_new_n21948__ = ~new_new_n21946__ & ~new_new_n21947__;
  assign new_new_n21949__ = ~new_new_n21944__ & ~new_new_n21948__;
  assign new_new_n21950__ = new_new_n21944__ & new_new_n21948__;
  assign new_new_n21951__ = ~new_new_n21794__ & ~new_new_n21807__;
  assign new_new_n21952__ = ~pi20 & new_new_n21496__;
  assign new_new_n21953__ = ~new_new_n21809__ & ~new_new_n21952__;
  assign new_new_n21954__ = ~new_new_n21484__ & new_new_n21953__;
  assign new_new_n21955__ = new_new_n21484__ & ~new_new_n21953__;
  assign new_new_n21956__ = ~new_new_n21954__ & ~new_new_n21955__;
  assign new_new_n21957__ = new_new_n21951__ & ~new_new_n21956__;
  assign new_new_n21958__ = new_new_n21794__ & new_new_n21807__;
  assign new_new_n21959__ = ~new_new_n21951__ & ~new_new_n21958__;
  assign new_new_n21960__ = new_new_n21491__ & new_new_n21496__;
  assign new_new_n21961__ = ~new_new_n21500__ & ~new_new_n21960__;
  assign new_new_n21962__ = new_new_n21484__ & new_new_n21961__;
  assign new_new_n21963__ = ~new_new_n21484__ & ~new_new_n21961__;
  assign new_new_n21964__ = ~new_new_n21962__ & ~new_new_n21963__;
  assign new_new_n21965__ = new_new_n21959__ & new_new_n21964__;
  assign new_new_n21966__ = new_new_n21956__ & new_new_n21958__;
  assign new_new_n21967__ = ~new_new_n21957__ & ~new_new_n21965__;
  assign new_new_n21968__ = ~new_new_n21966__ & new_new_n21967__;
  assign new_new_n21969__ = ~new_new_n21787__ & ~new_new_n21788__;
  assign new_new_n21970__ = ~new_new_n21792__ & new_new_n21969__;
  assign new_new_n21971__ = new_new_n21792__ & ~new_new_n21969__;
  assign new_new_n21972__ = ~new_new_n21970__ & ~new_new_n21971__;
  assign new_new_n21973__ = new_new_n7935__ & ~new_new_n15487__;
  assign new_new_n21974__ = new_new_n6968__ & new_new_n15524__;
  assign new_new_n21975__ = new_new_n6964__ & new_new_n15520__;
  assign new_new_n21976__ = new_new_n6959__ & new_new_n17587__;
  assign new_new_n21977__ = ~new_new_n21974__ & ~new_new_n21975__;
  assign new_new_n21978__ = ~new_new_n21973__ & new_new_n21977__;
  assign new_new_n21979__ = ~new_new_n21976__ & new_new_n21978__;
  assign new_new_n21980__ = pi17 & ~new_new_n21972__;
  assign new_new_n21981__ = ~pi17 & new_new_n21972__;
  assign new_new_n21982__ = ~new_new_n21980__ & ~new_new_n21981__;
  assign new_new_n21983__ = new_new_n21979__ & new_new_n21982__;
  assign new_new_n21984__ = ~new_new_n21979__ & ~new_new_n21982__;
  assign new_new_n21985__ = ~new_new_n21983__ & ~new_new_n21984__;
  assign new_new_n21986__ = ~new_new_n21972__ & ~new_new_n21985__;
  assign new_new_n21987__ = new_new_n6968__ & new_new_n15520__;
  assign new_new_n21988__ = new_new_n6964__ & ~new_new_n15533__;
  assign new_new_n21989__ = ~new_new_n21987__ & ~new_new_n21988__;
  assign new_new_n21990__ = new_new_n6958__ & new_new_n18923__;
  assign new_new_n21991__ = new_new_n21989__ & ~new_new_n21990__;
  assign new_new_n21992__ = pi17 & ~new_new_n21991__;
  assign new_new_n21993__ = new_new_n6958__ & ~new_new_n18914__;
  assign new_new_n21994__ = ~pi17 & ~new_new_n21993__;
  assign new_new_n21995__ = ~pi16 & new_new_n15524__;
  assign new_new_n21996__ = pi16 & ~new_new_n15524__;
  assign new_new_n21997__ = new_new_n6958__ & ~new_new_n21995__;
  assign new_new_n21998__ = ~new_new_n21996__ & new_new_n21997__;
  assign new_new_n21999__ = new_new_n18913__ & new_new_n21998__;
  assign new_new_n22000__ = ~new_new_n21994__ & ~new_new_n21999__;
  assign new_new_n22001__ = new_new_n21989__ & ~new_new_n22000__;
  assign new_new_n22002__ = ~new_new_n21992__ & ~new_new_n22001__;
  assign new_new_n22003__ = ~new_new_n21773__ & ~new_new_n21774__;
  assign new_new_n22004__ = new_new_n21784__ & new_new_n22003__;
  assign new_new_n22005__ = ~new_new_n21784__ & ~new_new_n22003__;
  assign new_new_n22006__ = ~new_new_n22004__ & ~new_new_n22005__;
  assign new_new_n22007__ = new_new_n22002__ & ~new_new_n22006__;
  assign new_new_n22008__ = ~new_new_n22002__ & new_new_n22006__;
  assign new_new_n22009__ = ~new_new_n21741__ & ~new_new_n21742__;
  assign new_new_n22010__ = ~new_new_n21752__ & new_new_n22009__;
  assign new_new_n22011__ = new_new_n21752__ & ~new_new_n22009__;
  assign new_new_n22012__ = ~new_new_n22010__ & ~new_new_n22011__;
  assign new_new_n22013__ = ~new_new_n21557__ & ~new_new_n21558__;
  assign new_new_n22014__ = ~new_new_n21738__ & new_new_n22013__;
  assign new_new_n22015__ = new_new_n21738__ & ~new_new_n22013__;
  assign new_new_n22016__ = ~new_new_n22014__ & ~new_new_n22015__;
  assign new_new_n22017__ = new_new_n6959__ & new_new_n18944__;
  assign new_new_n22018__ = new_new_n6964__ & new_new_n15564__;
  assign new_new_n22019__ = new_new_n6968__ & new_new_n15572__;
  assign new_new_n22020__ = ~new_new_n22018__ & ~new_new_n22019__;
  assign new_new_n22021__ = ~new_new_n22017__ & new_new_n22020__;
  assign new_new_n22022__ = new_new_n6958__ & new_new_n15560__;
  assign new_new_n22023__ = pi17 & ~new_new_n22022__;
  assign new_new_n22024__ = new_new_n8160__ & new_new_n15560__;
  assign new_new_n22025__ = ~new_new_n22023__ & ~new_new_n22024__;
  assign new_new_n22026__ = new_new_n22021__ & ~new_new_n22025__;
  assign new_new_n22027__ = ~pi17 & ~new_new_n22021__;
  assign new_new_n22028__ = ~new_new_n22026__ & ~new_new_n22027__;
  assign new_new_n22029__ = ~new_new_n21711__ & ~new_new_n21712__;
  assign new_new_n22030__ = new_new_n21716__ & new_new_n22029__;
  assign new_new_n22031__ = ~new_new_n21716__ & ~new_new_n22029__;
  assign new_new_n22032__ = ~new_new_n22030__ & ~new_new_n22031__;
  assign new_new_n22033__ = new_new_n6968__ & ~new_new_n15615__;
  assign new_new_n22034__ = new_new_n6964__ & new_new_n15743__;
  assign new_new_n22035__ = new_new_n7935__ & new_new_n15564__;
  assign new_new_n22036__ = ~new_new_n22033__ & ~new_new_n22034__;
  assign new_new_n22037__ = ~new_new_n22035__ & new_new_n22036__;
  assign new_new_n22038__ = new_new_n6958__ & new_new_n18512__;
  assign new_new_n22039__ = pi17 & ~new_new_n22038__;
  assign new_new_n22040__ = new_new_n7942__ & new_new_n18512__;
  assign new_new_n22041__ = ~new_new_n22039__ & ~new_new_n22040__;
  assign new_new_n22042__ = new_new_n22037__ & ~new_new_n22041__;
  assign new_new_n22043__ = ~pi17 & ~new_new_n22037__;
  assign new_new_n22044__ = ~new_new_n22042__ & ~new_new_n22043__;
  assign new_new_n22045__ = ~new_new_n21683__ & ~new_new_n21684__;
  assign new_new_n22046__ = new_new_n21694__ & new_new_n22045__;
  assign new_new_n22047__ = ~new_new_n21694__ & ~new_new_n22045__;
  assign new_new_n22048__ = ~new_new_n22046__ & ~new_new_n22047__;
  assign new_new_n22049__ = ~new_new_n21673__ & ~new_new_n21674__;
  assign new_new_n22050__ = ~new_new_n21676__ & ~new_new_n21680__;
  assign new_new_n22051__ = new_new_n22049__ & ~new_new_n22050__;
  assign new_new_n22052__ = ~new_new_n21676__ & ~new_new_n21679__;
  assign new_new_n22053__ = ~new_new_n22049__ & new_new_n22052__;
  assign new_new_n22054__ = ~new_new_n22051__ & ~new_new_n22053__;
  assign new_new_n22055__ = ~new_new_n21659__ & ~new_new_n21660__;
  assign new_new_n22056__ = new_new_n21670__ & new_new_n22055__;
  assign new_new_n22057__ = ~new_new_n21670__ & ~new_new_n22055__;
  assign new_new_n22058__ = ~new_new_n22056__ & ~new_new_n22057__;
  assign new_new_n22059__ = new_new_n7935__ & ~new_new_n15582__;
  assign new_new_n22060__ = new_new_n6964__ & ~new_new_n15710__;
  assign new_new_n22061__ = new_new_n6968__ & ~new_new_n15647__;
  assign new_new_n22062__ = ~new_new_n22060__ & ~new_new_n22061__;
  assign new_new_n22063__ = ~new_new_n22059__ & new_new_n22062__;
  assign new_new_n22064__ = new_new_n6958__ & ~new_new_n15736__;
  assign new_new_n22065__ = pi17 & ~new_new_n22064__;
  assign new_new_n22066__ = new_new_n7942__ & ~new_new_n15736__;
  assign new_new_n22067__ = ~new_new_n22065__ & ~new_new_n22066__;
  assign new_new_n22068__ = new_new_n22063__ & ~new_new_n22067__;
  assign new_new_n22069__ = ~pi17 & ~new_new_n22063__;
  assign new_new_n22070__ = ~new_new_n22068__ & ~new_new_n22069__;
  assign new_new_n22071__ = new_new_n6631__ & ~new_new_n15673__;
  assign new_new_n22072__ = new_new_n6963__ & ~new_new_n20628__;
  assign new_new_n22073__ = new_new_n6958__ & ~new_new_n15661__;
  assign new_new_n22074__ = ~new_new_n6964__ & ~new_new_n22073__;
  assign new_new_n22075__ = ~new_new_n15673__ & ~new_new_n22074__;
  assign new_new_n22076__ = new_new_n6955__ & new_new_n15668__;
  assign new_new_n22077__ = new_new_n15661__ & ~new_new_n22076__;
  assign new_new_n22078__ = ~new_new_n15679__ & new_new_n22076__;
  assign new_new_n22079__ = new_new_n6958__ & ~new_new_n22077__;
  assign new_new_n22080__ = ~new_new_n22078__ & new_new_n22079__;
  assign new_new_n22081__ = ~new_new_n22075__ & ~new_new_n22080__;
  assign new_new_n22082__ = pi17 & ~new_new_n22072__;
  assign new_new_n22083__ = new_new_n22081__ & new_new_n22082__;
  assign new_new_n22084__ = ~new_new_n22071__ & ~new_new_n22083__;
  assign new_new_n22085__ = new_new_n7935__ & new_new_n15643__;
  assign new_new_n22086__ = new_new_n6959__ & new_new_n20646__;
  assign new_new_n22087__ = new_new_n6968__ & ~new_new_n15661__;
  assign new_new_n22088__ = ~new_new_n22085__ & ~new_new_n22087__;
  assign new_new_n22089__ = ~new_new_n22086__ & new_new_n22088__;
  assign new_new_n22090__ = new_new_n10337__ & new_new_n15668__;
  assign new_new_n22091__ = pi17 & ~new_new_n22090__;
  assign new_new_n22092__ = new_new_n10340__ & new_new_n15668__;
  assign new_new_n22093__ = ~pi17 & ~new_new_n22092__;
  assign new_new_n22094__ = pi14 & ~new_new_n22093__;
  assign new_new_n22095__ = ~new_new_n22091__ & ~new_new_n22094__;
  assign new_new_n22096__ = new_new_n22089__ & ~new_new_n22095__;
  assign new_new_n22097__ = ~pi17 & ~new_new_n22089__;
  assign new_new_n22098__ = ~new_new_n22096__ & ~new_new_n22097__;
  assign new_new_n22099__ = ~new_new_n22084__ & ~new_new_n22098__;
  assign new_new_n22100__ = new_new_n6627__ & new_new_n15674__;
  assign new_new_n22101__ = ~new_new_n6631__ & new_new_n20195__;
  assign new_new_n22102__ = ~new_new_n6622__ & new_new_n15668__;
  assign new_new_n22103__ = new_new_n6628__ & ~new_new_n22102__;
  assign new_new_n22104__ = ~new_new_n9920__ & ~new_new_n20628__;
  assign new_new_n22105__ = ~new_new_n22100__ & new_new_n22104__;
  assign new_new_n22106__ = ~new_new_n22101__ & ~new_new_n22103__;
  assign new_new_n22107__ = new_new_n22105__ & new_new_n22106__;
  assign new_new_n22108__ = new_new_n22099__ & new_new_n22107__;
  assign new_new_n22109__ = ~new_new_n22099__ & ~new_new_n22107__;
  assign new_new_n22110__ = new_new_n7935__ & new_new_n15656__;
  assign new_new_n22111__ = new_new_n6968__ & new_new_n15643__;
  assign new_new_n22112__ = new_new_n6964__ & ~new_new_n15661__;
  assign new_new_n22113__ = new_new_n6959__ & new_new_n15687__;
  assign new_new_n22114__ = ~new_new_n22111__ & ~new_new_n22112__;
  assign new_new_n22115__ = ~new_new_n22110__ & new_new_n22114__;
  assign new_new_n22116__ = ~new_new_n22113__ & new_new_n22115__;
  assign new_new_n22117__ = ~pi17 & ~new_new_n22116__;
  assign new_new_n22118__ = pi17 & new_new_n22116__;
  assign new_new_n22119__ = ~new_new_n22117__ & ~new_new_n22118__;
  assign new_new_n22120__ = ~new_new_n22109__ & ~new_new_n22119__;
  assign new_new_n22121__ = ~new_new_n22108__ & ~new_new_n22120__;
  assign new_new_n22122__ = new_new_n21618__ & ~new_new_n21633__;
  assign new_new_n22123__ = ~new_new_n21618__ & new_new_n21633__;
  assign new_new_n22124__ = ~new_new_n22122__ & ~new_new_n22123__;
  assign new_new_n22125__ = new_new_n22121__ & new_new_n22124__;
  assign new_new_n22126__ = new_new_n7935__ & ~new_new_n15710__;
  assign new_new_n22127__ = new_new_n6964__ & new_new_n15643__;
  assign new_new_n22128__ = new_new_n6968__ & new_new_n15656__;
  assign new_new_n22129__ = ~new_new_n22127__ & ~new_new_n22128__;
  assign new_new_n22130__ = ~new_new_n22126__ & new_new_n22129__;
  assign new_new_n22131__ = new_new_n6958__ & ~new_new_n19466__;
  assign new_new_n22132__ = ~pi17 & ~new_new_n22131__;
  assign new_new_n22133__ = new_new_n8160__ & ~new_new_n19466__;
  assign new_new_n22134__ = ~new_new_n22132__ & ~new_new_n22133__;
  assign new_new_n22135__ = new_new_n22130__ & ~new_new_n22134__;
  assign new_new_n22136__ = pi17 & ~new_new_n22130__;
  assign new_new_n22137__ = ~new_new_n22135__ & ~new_new_n22136__;
  assign new_new_n22138__ = ~new_new_n22125__ & new_new_n22137__;
  assign new_new_n22139__ = new_new_n21617__ & new_new_n21633__;
  assign new_new_n22140__ = ~new_new_n22121__ & new_new_n22139__;
  assign new_new_n22141__ = ~new_new_n22138__ & ~new_new_n22140__;
  assign new_new_n22142__ = ~pi21 & ~new_new_n15673__;
  assign new_new_n22143__ = ~new_new_n21617__ & new_new_n22142__;
  assign new_new_n22144__ = new_new_n21633__ & new_new_n22143__;
  assign new_new_n22145__ = ~new_new_n21635__ & new_new_n22144__;
  assign new_new_n22146__ = ~new_new_n21613__ & new_new_n21635__;
  assign new_new_n22147__ = ~new_new_n21636__ & ~new_new_n22146__;
  assign new_new_n22148__ = ~new_new_n22145__ & ~new_new_n22147__;
  assign new_new_n22149__ = ~new_new_n22141__ & ~new_new_n22148__;
  assign new_new_n22150__ = new_new_n22141__ & new_new_n22148__;
  assign new_new_n22151__ = new_new_n6959__ & ~new_new_n19118__;
  assign new_new_n22152__ = new_new_n6964__ & new_new_n15656__;
  assign new_new_n22153__ = new_new_n6968__ & ~new_new_n15710__;
  assign new_new_n22154__ = new_new_n7935__ & ~new_new_n15647__;
  assign new_new_n22155__ = ~new_new_n22152__ & ~new_new_n22153__;
  assign new_new_n22156__ = ~new_new_n22154__ & new_new_n22155__;
  assign new_new_n22157__ = ~new_new_n22151__ & new_new_n22156__;
  assign new_new_n22158__ = pi17 & ~new_new_n22157__;
  assign new_new_n22159__ = ~pi17 & new_new_n22157__;
  assign new_new_n22160__ = ~new_new_n22158__ & ~new_new_n22159__;
  assign new_new_n22161__ = ~new_new_n22150__ & new_new_n22160__;
  assign new_new_n22162__ = ~new_new_n22149__ & ~new_new_n22161__;
  assign new_new_n22163__ = ~new_new_n22070__ & ~new_new_n22162__;
  assign new_new_n22164__ = new_new_n22070__ & new_new_n22162__;
  assign new_new_n22165__ = ~new_new_n21645__ & ~new_new_n21646__;
  assign new_new_n22166__ = new_new_n21656__ & ~new_new_n22165__;
  assign new_new_n22167__ = ~new_new_n21656__ & new_new_n22165__;
  assign new_new_n22168__ = ~new_new_n22166__ & ~new_new_n22167__;
  assign new_new_n22169__ = ~new_new_n22164__ & ~new_new_n22168__;
  assign new_new_n22170__ = ~new_new_n22163__ & ~new_new_n22169__;
  assign new_new_n22171__ = new_new_n22058__ & ~new_new_n22170__;
  assign new_new_n22172__ = ~new_new_n22058__ & new_new_n22170__;
  assign new_new_n22173__ = new_new_n6959__ & new_new_n19487__;
  assign new_new_n22174__ = new_new_n6964__ & ~new_new_n15647__;
  assign new_new_n22175__ = new_new_n6968__ & ~new_new_n15582__;
  assign new_new_n22176__ = ~new_new_n22174__ & ~new_new_n22175__;
  assign new_new_n22177__ = ~new_new_n22173__ & new_new_n22176__;
  assign new_new_n22178__ = new_new_n6958__ & ~new_new_n15638__;
  assign new_new_n22179__ = ~pi17 & ~new_new_n22178__;
  assign new_new_n22180__ = new_new_n7942__ & ~new_new_n15638__;
  assign new_new_n22181__ = ~new_new_n22179__ & ~new_new_n22180__;
  assign new_new_n22182__ = new_new_n22177__ & ~new_new_n22181__;
  assign new_new_n22183__ = pi17 & ~new_new_n22177__;
  assign new_new_n22184__ = ~new_new_n22182__ & ~new_new_n22183__;
  assign new_new_n22185__ = ~new_new_n22172__ & new_new_n22184__;
  assign new_new_n22186__ = ~new_new_n22171__ & ~new_new_n22185__;
  assign new_new_n22187__ = ~new_new_n22054__ & new_new_n22186__;
  assign new_new_n22188__ = new_new_n22054__ & ~new_new_n22186__;
  assign new_new_n22189__ = new_new_n6959__ & new_new_n19494__;
  assign new_new_n22190__ = new_new_n6964__ & ~new_new_n15582__;
  assign new_new_n22191__ = new_new_n6968__ & ~new_new_n15638__;
  assign new_new_n22192__ = new_new_n7935__ & new_new_n15743__;
  assign new_new_n22193__ = ~new_new_n22190__ & ~new_new_n22191__;
  assign new_new_n22194__ = ~new_new_n22192__ & new_new_n22193__;
  assign new_new_n22195__ = ~new_new_n22189__ & new_new_n22194__;
  assign new_new_n22196__ = pi17 & ~new_new_n22195__;
  assign new_new_n22197__ = ~pi17 & new_new_n22195__;
  assign new_new_n22198__ = ~new_new_n22196__ & ~new_new_n22197__;
  assign new_new_n22199__ = ~new_new_n22188__ & ~new_new_n22198__;
  assign new_new_n22200__ = ~new_new_n22187__ & ~new_new_n22199__;
  assign new_new_n22201__ = ~new_new_n22048__ & ~new_new_n22200__;
  assign new_new_n22202__ = new_new_n22048__ & new_new_n22200__;
  assign new_new_n22203__ = new_new_n7935__ & ~new_new_n15615__;
  assign new_new_n22204__ = new_new_n6968__ & new_new_n15743__;
  assign new_new_n22205__ = new_new_n6964__ & ~new_new_n15638__;
  assign new_new_n22206__ = new_new_n6959__ & new_new_n19005__;
  assign new_new_n22207__ = ~new_new_n22204__ & ~new_new_n22205__;
  assign new_new_n22208__ = ~new_new_n22203__ & new_new_n22207__;
  assign new_new_n22209__ = ~new_new_n22206__ & new_new_n22208__;
  assign new_new_n22210__ = pi17 & ~new_new_n22209__;
  assign new_new_n22211__ = ~pi17 & new_new_n22209__;
  assign new_new_n22212__ = ~new_new_n22210__ & ~new_new_n22211__;
  assign new_new_n22213__ = ~new_new_n22202__ & ~new_new_n22212__;
  assign new_new_n22214__ = ~new_new_n22201__ & ~new_new_n22213__;
  assign new_new_n22215__ = new_new_n22044__ & ~new_new_n22214__;
  assign new_new_n22216__ = ~new_new_n22044__ & new_new_n22214__;
  assign new_new_n22217__ = pi20 & new_new_n21574__;
  assign new_new_n22218__ = ~pi20 & ~new_new_n21574__;
  assign new_new_n22219__ = ~new_new_n22217__ & ~new_new_n22218__;
  assign new_new_n22220__ = ~new_new_n21696__ & new_new_n21705__;
  assign new_new_n22221__ = new_new_n21696__ & ~new_new_n21705__;
  assign new_new_n22222__ = ~new_new_n22220__ & ~new_new_n22221__;
  assign new_new_n22223__ = new_new_n22219__ & new_new_n22222__;
  assign new_new_n22224__ = ~new_new_n22219__ & ~new_new_n22222__;
  assign new_new_n22225__ = ~new_new_n22223__ & ~new_new_n22224__;
  assign new_new_n22226__ = ~new_new_n22216__ & ~new_new_n22225__;
  assign new_new_n22227__ = ~new_new_n22215__ & ~new_new_n22226__;
  assign new_new_n22228__ = ~new_new_n22032__ & ~new_new_n22227__;
  assign new_new_n22229__ = new_new_n22032__ & new_new_n22227__;
  assign new_new_n22230__ = new_new_n7935__ & new_new_n15572__;
  assign new_new_n22231__ = new_new_n6964__ & ~new_new_n15615__;
  assign new_new_n22232__ = new_new_n6968__ & new_new_n15564__;
  assign new_new_n22233__ = ~new_new_n22231__ & ~new_new_n22232__;
  assign new_new_n22234__ = ~new_new_n22230__ & new_new_n22233__;
  assign new_new_n22235__ = new_new_n6958__ & ~new_new_n20114__;
  assign new_new_n22236__ = pi17 & ~new_new_n22235__;
  assign new_new_n22237__ = new_new_n7942__ & ~new_new_n20114__;
  assign new_new_n22238__ = ~new_new_n22236__ & ~new_new_n22237__;
  assign new_new_n22239__ = new_new_n22234__ & ~new_new_n22238__;
  assign new_new_n22240__ = ~pi17 & ~new_new_n22234__;
  assign new_new_n22241__ = ~new_new_n22239__ & ~new_new_n22240__;
  assign new_new_n22242__ = ~new_new_n22229__ & new_new_n22241__;
  assign new_new_n22243__ = ~new_new_n22228__ & ~new_new_n22242__;
  assign new_new_n22244__ = new_new_n22028__ & ~new_new_n22243__;
  assign new_new_n22245__ = ~new_new_n22028__ & new_new_n22243__;
  assign new_new_n22246__ = ~new_new_n21723__ & ~new_new_n21724__;
  assign new_new_n22247__ = ~new_new_n21736__ & new_new_n22246__;
  assign new_new_n22248__ = new_new_n21736__ & ~new_new_n22246__;
  assign new_new_n22249__ = ~new_new_n22247__ & ~new_new_n22248__;
  assign new_new_n22250__ = ~new_new_n22245__ & ~new_new_n22249__;
  assign new_new_n22251__ = ~new_new_n22244__ & ~new_new_n22250__;
  assign new_new_n22252__ = ~new_new_n22016__ & new_new_n22251__;
  assign new_new_n22253__ = new_new_n22016__ & ~new_new_n22251__;
  assign new_new_n22254__ = new_new_n6968__ & new_new_n15560__;
  assign new_new_n22255__ = new_new_n6964__ & new_new_n15572__;
  assign new_new_n22256__ = new_new_n7935__ & new_new_n15767__;
  assign new_new_n22257__ = ~new_new_n22255__ & ~new_new_n22256__;
  assign new_new_n22258__ = ~new_new_n22254__ & new_new_n22257__;
  assign new_new_n22259__ = new_new_n6958__ & ~new_new_n18454__;
  assign new_new_n22260__ = pi17 & ~new_new_n22259__;
  assign new_new_n22261__ = new_new_n7942__ & ~new_new_n18454__;
  assign new_new_n22262__ = ~new_new_n22260__ & ~new_new_n22261__;
  assign new_new_n22263__ = new_new_n22258__ & ~new_new_n22262__;
  assign new_new_n22264__ = ~pi17 & ~new_new_n22258__;
  assign new_new_n22265__ = ~new_new_n22263__ & ~new_new_n22264__;
  assign new_new_n22266__ = ~new_new_n22253__ & ~new_new_n22265__;
  assign new_new_n22267__ = ~new_new_n22252__ & ~new_new_n22266__;
  assign new_new_n22268__ = ~new_new_n22012__ & ~new_new_n22267__;
  assign new_new_n22269__ = new_new_n22012__ & new_new_n22267__;
  assign new_new_n22270__ = ~new_new_n22268__ & ~new_new_n22269__;
  assign new_new_n22271__ = new_new_n7935__ & ~new_new_n15533__;
  assign new_new_n22272__ = new_new_n6968__ & new_new_n15767__;
  assign new_new_n22273__ = new_new_n6964__ & new_new_n15560__;
  assign new_new_n22274__ = new_new_n6959__ & new_new_n19893__;
  assign new_new_n22275__ = ~new_new_n22272__ & ~new_new_n22273__;
  assign new_new_n22276__ = ~new_new_n22271__ & new_new_n22275__;
  assign new_new_n22277__ = ~new_new_n22274__ & new_new_n22276__;
  assign new_new_n22278__ = pi17 & ~new_new_n22277__;
  assign new_new_n22279__ = ~pi17 & new_new_n22277__;
  assign new_new_n22280__ = ~new_new_n22278__ & ~new_new_n22279__;
  assign new_new_n22281__ = new_new_n22270__ & new_new_n22280__;
  assign new_new_n22282__ = ~new_new_n22268__ & ~new_new_n22281__;
  assign new_new_n22283__ = ~new_new_n21755__ & ~new_new_n21756__;
  assign new_new_n22284__ = ~new_new_n21766__ & new_new_n22283__;
  assign new_new_n22285__ = new_new_n21766__ & ~new_new_n22283__;
  assign new_new_n22286__ = ~new_new_n22284__ & ~new_new_n22285__;
  assign new_new_n22287__ = new_new_n22282__ & ~new_new_n22286__;
  assign new_new_n22288__ = ~new_new_n22282__ & new_new_n22286__;
  assign new_new_n22289__ = new_new_n7935__ & new_new_n15520__;
  assign new_new_n22290__ = new_new_n6964__ & new_new_n15767__;
  assign new_new_n22291__ = new_new_n6968__ & ~new_new_n15533__;
  assign new_new_n22292__ = ~new_new_n22290__ & ~new_new_n22291__;
  assign new_new_n22293__ = ~new_new_n22289__ & new_new_n22292__;
  assign new_new_n22294__ = new_new_n6958__ & new_new_n19731__;
  assign new_new_n22295__ = pi17 & ~new_new_n22294__;
  assign new_new_n22296__ = new_new_n7942__ & new_new_n19731__;
  assign new_new_n22297__ = ~new_new_n22295__ & ~new_new_n22296__;
  assign new_new_n22298__ = new_new_n22293__ & ~new_new_n22297__;
  assign new_new_n22299__ = ~pi17 & ~new_new_n22293__;
  assign new_new_n22300__ = ~new_new_n22298__ & ~new_new_n22299__;
  assign new_new_n22301__ = ~new_new_n22288__ & new_new_n22300__;
  assign new_new_n22302__ = ~new_new_n22287__ & ~new_new_n22301__;
  assign new_new_n22303__ = ~new_new_n22008__ & new_new_n22302__;
  assign new_new_n22304__ = ~new_new_n22007__ & ~new_new_n22303__;
  assign new_new_n22305__ = new_new_n21985__ & new_new_n22304__;
  assign new_new_n22306__ = ~new_new_n21986__ & ~new_new_n22305__;
  assign new_new_n22307__ = new_new_n7935__ & ~new_new_n15809__;
  assign new_new_n22308__ = new_new_n6964__ & new_new_n15524__;
  assign new_new_n22309__ = new_new_n6968__ & ~new_new_n15487__;
  assign new_new_n22310__ = ~new_new_n22308__ & ~new_new_n22309__;
  assign new_new_n22311__ = ~new_new_n22307__ & new_new_n22310__;
  assign new_new_n22312__ = new_new_n6958__ & new_new_n18020__;
  assign new_new_n22313__ = ~pi17 & ~new_new_n22312__;
  assign new_new_n22314__ = new_new_n8160__ & new_new_n18020__;
  assign new_new_n22315__ = ~new_new_n22313__ & ~new_new_n22314__;
  assign new_new_n22316__ = new_new_n22311__ & ~new_new_n22315__;
  assign new_new_n22317__ = pi17 & ~new_new_n22311__;
  assign new_new_n22318__ = ~new_new_n22316__ & ~new_new_n22317__;
  assign new_new_n22319__ = new_new_n22306__ & new_new_n22318__;
  assign new_new_n22320__ = ~new_new_n22306__ & ~new_new_n22318__;
  assign new_new_n22321__ = ~new_new_n21492__ & ~new_new_n21810__;
  assign new_new_n22322__ = ~new_new_n21959__ & ~new_new_n22321__;
  assign new_new_n22323__ = new_new_n21959__ & new_new_n22321__;
  assign new_new_n22324__ = ~new_new_n22322__ & ~new_new_n22323__;
  assign new_new_n22325__ = ~new_new_n22320__ & ~new_new_n22324__;
  assign new_new_n22326__ = ~new_new_n22319__ & ~new_new_n22325__;
  assign new_new_n22327__ = new_new_n21968__ & ~new_new_n22326__;
  assign new_new_n22328__ = ~new_new_n21968__ & new_new_n22326__;
  assign new_new_n22329__ = new_new_n6964__ & ~new_new_n15487__;
  assign new_new_n22330__ = new_new_n6959__ & ~new_new_n18633__;
  assign new_new_n22331__ = ~new_new_n22329__ & ~new_new_n22330__;
  assign new_new_n22332__ = new_new_n6968__ & ~new_new_n15809__;
  assign new_new_n22333__ = new_new_n7935__ & ~new_new_n15471__;
  assign new_new_n22334__ = ~new_new_n22332__ & ~new_new_n22333__;
  assign new_new_n22335__ = new_new_n22331__ & new_new_n22334__;
  assign new_new_n22336__ = ~pi17 & ~new_new_n22335__;
  assign new_new_n22337__ = ~new_new_n6968__ & new_new_n15471__;
  assign new_new_n22338__ = new_new_n7935__ & ~new_new_n22337__;
  assign new_new_n22339__ = pi17 & ~new_new_n22332__;
  assign new_new_n22340__ = ~new_new_n22338__ & new_new_n22339__;
  assign new_new_n22341__ = new_new_n22331__ & new_new_n22340__;
  assign new_new_n22342__ = ~new_new_n22336__ & ~new_new_n22341__;
  assign new_new_n22343__ = ~new_new_n22328__ & ~new_new_n22342__;
  assign new_new_n22344__ = ~new_new_n22327__ & ~new_new_n22343__;
  assign new_new_n22345__ = ~new_new_n21950__ & ~new_new_n22344__;
  assign new_new_n22346__ = ~new_new_n21949__ & ~new_new_n22345__;
  assign new_new_n22347__ = ~new_new_n21930__ & ~new_new_n22346__;
  assign new_new_n22348__ = ~new_new_n21929__ & ~new_new_n22347__;
  assign new_new_n22349__ = new_new_n21912__ & ~new_new_n22348__;
  assign new_new_n22350__ = ~new_new_n21912__ & new_new_n22348__;
  assign new_new_n22351__ = ~new_new_n21847__ & ~new_new_n21848__;
  assign new_new_n22352__ = ~new_new_n21852__ & new_new_n22351__;
  assign new_new_n22353__ = new_new_n21852__ & ~new_new_n22351__;
  assign new_new_n22354__ = ~new_new_n22352__ & ~new_new_n22353__;
  assign new_new_n22355__ = ~new_new_n22350__ & ~new_new_n22354__;
  assign new_new_n22356__ = ~new_new_n22349__ & ~new_new_n22355__;
  assign new_new_n22357__ = new_new_n21900__ & new_new_n22356__;
  assign new_new_n22358__ = ~new_new_n21900__ & ~new_new_n22356__;
  assign new_new_n22359__ = new_new_n7935__ & ~new_new_n15362__;
  assign new_new_n22360__ = new_new_n6968__ & ~new_new_n15432__;
  assign new_new_n22361__ = new_new_n6959__ & new_new_n16771__;
  assign new_new_n22362__ = ~new_new_n22359__ & ~new_new_n22360__;
  assign new_new_n22363__ = ~new_new_n22361__ & new_new_n22362__;
  assign new_new_n22364__ = new_new_n10337__ & ~new_new_n15439__;
  assign new_new_n22365__ = pi17 & ~new_new_n22364__;
  assign new_new_n22366__ = new_new_n10340__ & ~new_new_n15439__;
  assign new_new_n22367__ = ~pi17 & ~new_new_n22366__;
  assign new_new_n22368__ = pi14 & ~new_new_n22367__;
  assign new_new_n22369__ = ~new_new_n22365__ & ~new_new_n22368__;
  assign new_new_n22370__ = new_new_n22363__ & ~new_new_n22369__;
  assign new_new_n22371__ = ~pi17 & ~new_new_n22363__;
  assign new_new_n22372__ = ~new_new_n22370__ & ~new_new_n22371__;
  assign new_new_n22373__ = ~new_new_n22358__ & new_new_n22372__;
  assign new_new_n22374__ = ~new_new_n22357__ & ~new_new_n22373__;
  assign new_new_n22375__ = ~new_new_n21867__ & ~new_new_n21868__;
  assign new_new_n22376__ = new_new_n6964__ & ~new_new_n15432__;
  assign new_new_n22377__ = new_new_n6968__ & ~new_new_n15362__;
  assign new_new_n22378__ = ~new_new_n22376__ & ~new_new_n22377__;
  assign new_new_n22379__ = new_new_n6958__ & ~new_new_n17918__;
  assign new_new_n22380__ = pi17 & ~new_new_n22379__;
  assign new_new_n22381__ = pi16 & new_new_n15390__;
  assign new_new_n22382__ = ~pi16 & ~new_new_n15390__;
  assign new_new_n22383__ = new_new_n6958__ & new_new_n15829__;
  assign new_new_n22384__ = ~new_new_n22381__ & ~new_new_n22382__;
  assign new_new_n22385__ = new_new_n22383__ & new_new_n22384__;
  assign new_new_n22386__ = ~new_new_n22380__ & ~new_new_n22385__;
  assign new_new_n22387__ = new_new_n22378__ & ~new_new_n22386__;
  assign new_new_n22388__ = new_new_n6958__ & new_new_n17914__;
  assign new_new_n22389__ = new_new_n22378__ & ~new_new_n22388__;
  assign new_new_n22390__ = ~pi17 & ~new_new_n22389__;
  assign new_new_n22391__ = ~new_new_n22387__ & ~new_new_n22390__;
  assign new_new_n22392__ = new_new_n22375__ & ~new_new_n22391__;
  assign new_new_n22393__ = ~new_new_n22375__ & new_new_n22391__;
  assign new_new_n22394__ = ~new_new_n22392__ & ~new_new_n22393__;
  assign new_new_n22395__ = new_new_n21880__ & new_new_n22394__;
  assign new_new_n22396__ = ~new_new_n21880__ & ~new_new_n22394__;
  assign new_new_n22397__ = ~new_new_n22395__ & ~new_new_n22396__;
  assign new_new_n22398__ = ~new_new_n22374__ & new_new_n22397__;
  assign new_new_n22399__ = new_new_n22391__ & ~new_new_n22397__;
  assign new_new_n22400__ = ~new_new_n22398__ & ~new_new_n22399__;
  assign new_new_n22401__ = ~new_new_n21440__ & ~new_new_n21441__;
  assign new_new_n22402__ = new_new_n21882__ & ~new_new_n22401__;
  assign new_new_n22403__ = ~new_new_n21882__ & new_new_n22401__;
  assign new_new_n22404__ = ~new_new_n22402__ & ~new_new_n22403__;
  assign new_new_n22405__ = new_new_n22400__ & ~new_new_n22404__;
  assign new_new_n22406__ = ~new_new_n22400__ & new_new_n22404__;
  assign new_new_n22407__ = new_new_n6991__ & ~new_new_n15349__;
  assign new_new_n22408__ = new_new_n6985__ & ~new_new_n15321__;
  assign new_new_n22409__ = ~new_new_n22407__ & ~new_new_n22408__;
  assign new_new_n22410__ = new_new_n6994__ & ~new_new_n15273__;
  assign new_new_n22411__ = ~new_new_n17103__ & new_new_n22410__;
  assign new_new_n22412__ = new_new_n22409__ & ~new_new_n22411__;
  assign new_new_n22413__ = pi14 & ~new_new_n22412__;
  assign new_new_n22414__ = ~pi13 & ~new_new_n15273__;
  assign new_new_n22415__ = new_new_n15273__ & new_new_n17103__;
  assign new_new_n22416__ = new_new_n6994__ & ~new_new_n22415__;
  assign new_new_n22417__ = pi13 & ~new_new_n17103__;
  assign new_new_n22418__ = ~new_new_n22414__ & ~new_new_n22417__;
  assign new_new_n22419__ = new_new_n22416__ & new_new_n22418__;
  assign new_new_n22420__ = ~pi14 & new_new_n22409__;
  assign new_new_n22421__ = ~new_new_n22416__ & new_new_n22420__;
  assign new_new_n22422__ = ~new_new_n22413__ & ~new_new_n22419__;
  assign new_new_n22423__ = ~new_new_n22421__ & new_new_n22422__;
  assign new_new_n22424__ = ~new_new_n22406__ & new_new_n22423__;
  assign new_new_n22425__ = ~new_new_n22405__ & ~new_new_n22424__;
  assign new_new_n22426__ = ~new_new_n21896__ & ~new_new_n22425__;
  assign new_new_n22427__ = ~new_new_n21895__ & ~new_new_n22426__;
  assign new_new_n22428__ = new_new_n21393__ & ~new_new_n22427__;
  assign new_new_n22429__ = ~new_new_n21393__ & new_new_n22427__;
  assign new_new_n22430__ = ~new_new_n22428__ & ~new_new_n22429__;
  assign new_new_n22431__ = ~new_new_n21886__ & ~new_new_n21891__;
  assign new_new_n22432__ = ~new_new_n21885__ & ~new_new_n22431__;
  assign new_new_n22433__ = ~new_new_n20928__ & ~new_new_n20929__;
  assign new_new_n22434__ = ~new_new_n21350__ & new_new_n22433__;
  assign new_new_n22435__ = new_new_n21350__ & ~new_new_n22433__;
  assign new_new_n22436__ = ~new_new_n22434__ & ~new_new_n22435__;
  assign new_new_n22437__ = new_new_n22432__ & new_new_n22436__;
  assign new_new_n22438__ = ~new_new_n22432__ & ~new_new_n22436__;
  assign new_new_n22439__ = ~new_new_n22437__ & ~new_new_n22438__;
  assign new_new_n22440__ = new_new_n8474__ & new_new_n15244__;
  assign new_new_n22441__ = ~new_new_n8479__ & ~new_new_n15248__;
  assign new_new_n22442__ = new_new_n8858__ & new_new_n15237__;
  assign new_new_n22443__ = ~new_new_n22440__ & ~new_new_n22441__;
  assign new_new_n22444__ = ~new_new_n22442__ & new_new_n22443__;
  assign new_new_n22445__ = new_new_n8469__ & ~new_new_n16603__;
  assign new_new_n22446__ = pi11 & ~new_new_n22445__;
  assign new_new_n22447__ = new_new_n11530__ & ~new_new_n16603__;
  assign new_new_n22448__ = ~new_new_n22446__ & ~new_new_n22447__;
  assign new_new_n22449__ = new_new_n22444__ & ~new_new_n22448__;
  assign new_new_n22450__ = ~pi11 & ~new_new_n22444__;
  assign new_new_n22451__ = ~new_new_n22449__ & ~new_new_n22450__;
  assign new_new_n22452__ = new_new_n22439__ & ~new_new_n22451__;
  assign new_new_n22453__ = ~new_new_n22439__ & new_new_n22451__;
  assign new_new_n22454__ = ~new_new_n22452__ & ~new_new_n22453__;
  assign new_new_n22455__ = new_new_n22430__ & ~new_new_n22454__;
  assign new_new_n22456__ = ~new_new_n22430__ & new_new_n22454__;
  assign new_new_n22457__ = ~new_new_n22455__ & ~new_new_n22456__;
  assign new_new_n22458__ = new_new_n6985__ & ~new_new_n15349__;
  assign new_new_n22459__ = new_new_n6991__ & ~new_new_n15398__;
  assign new_new_n22460__ = ~new_new_n22458__ & ~new_new_n22459__;
  assign new_new_n22461__ = new_new_n6994__ & ~new_new_n15321__;
  assign new_new_n22462__ = new_new_n16458__ & new_new_n22461__;
  assign new_new_n22463__ = new_new_n22460__ & ~new_new_n22462__;
  assign new_new_n22464__ = pi14 & ~new_new_n22463__;
  assign new_new_n22465__ = pi13 & new_new_n16458__;
  assign new_new_n22466__ = new_new_n15321__ & ~new_new_n16458__;
  assign new_new_n22467__ = new_new_n6994__ & ~new_new_n22466__;
  assign new_new_n22468__ = ~pi13 & ~new_new_n15321__;
  assign new_new_n22469__ = ~new_new_n22465__ & ~new_new_n22468__;
  assign new_new_n22470__ = new_new_n22467__ & new_new_n22469__;
  assign new_new_n22471__ = ~pi14 & new_new_n22460__;
  assign new_new_n22472__ = ~new_new_n22467__ & new_new_n22471__;
  assign new_new_n22473__ = ~new_new_n22464__ & ~new_new_n22470__;
  assign new_new_n22474__ = ~new_new_n22472__ & new_new_n22473__;
  assign new_new_n22475__ = new_new_n6991__ & new_new_n15390__;
  assign new_new_n22476__ = new_new_n6985__ & ~new_new_n15398__;
  assign new_new_n22477__ = ~new_new_n22475__ & ~new_new_n22476__;
  assign new_new_n22478__ = new_new_n6994__ & ~new_new_n15349__;
  assign new_new_n22479__ = ~new_new_n17180__ & new_new_n22478__;
  assign new_new_n22480__ = new_new_n22477__ & ~new_new_n22479__;
  assign new_new_n22481__ = ~pi14 & ~new_new_n22480__;
  assign new_new_n22482__ = pi13 & ~new_new_n15349__;
  assign new_new_n22483__ = ~pi13 & ~new_new_n17180__;
  assign new_new_n22484__ = new_new_n15349__ & new_new_n17179__;
  assign new_new_n22485__ = new_new_n6994__ & ~new_new_n22484__;
  assign new_new_n22486__ = ~new_new_n22482__ & ~new_new_n22483__;
  assign new_new_n22487__ = new_new_n22485__ & new_new_n22486__;
  assign new_new_n22488__ = pi14 & new_new_n22477__;
  assign new_new_n22489__ = ~new_new_n22485__ & new_new_n22488__;
  assign new_new_n22490__ = ~new_new_n22481__ & ~new_new_n22489__;
  assign new_new_n22491__ = ~new_new_n22487__ & new_new_n22490__;
  assign new_new_n22492__ = new_new_n6991__ & ~new_new_n15432__;
  assign new_new_n22493__ = new_new_n6985__ & ~new_new_n15362__;
  assign new_new_n22494__ = ~new_new_n22492__ & ~new_new_n22493__;
  assign new_new_n22495__ = new_new_n6994__ & ~new_new_n17918__;
  assign new_new_n22496__ = pi14 & ~new_new_n22495__;
  assign new_new_n22497__ = ~new_new_n15828__ & new_new_n16954__;
  assign new_new_n22498__ = new_new_n8388__ & new_new_n22497__;
  assign new_new_n22499__ = ~new_new_n22496__ & ~new_new_n22498__;
  assign new_new_n22500__ = new_new_n22494__ & ~new_new_n22499__;
  assign new_new_n22501__ = new_new_n6994__ & new_new_n17914__;
  assign new_new_n22502__ = new_new_n22494__ & ~new_new_n22501__;
  assign new_new_n22503__ = ~pi14 & ~new_new_n22502__;
  assign new_new_n22504__ = new_new_n8820__ & ~new_new_n15826__;
  assign new_new_n22505__ = new_new_n16955__ & new_new_n22504__;
  assign new_new_n22506__ = ~new_new_n22503__ & ~new_new_n22505__;
  assign new_new_n22507__ = ~new_new_n22500__ & new_new_n22506__;
  assign new_new_n22508__ = ~new_new_n21929__ & ~new_new_n21930__;
  assign new_new_n22509__ = new_new_n6991__ & ~new_new_n15439__;
  assign new_new_n22510__ = new_new_n6985__ & ~new_new_n15432__;
  assign new_new_n22511__ = ~new_new_n22509__ & ~new_new_n22510__;
  assign new_new_n22512__ = new_new_n6994__ & ~new_new_n15362__;
  assign new_new_n22513__ = ~new_new_n16768__ & new_new_n22512__;
  assign new_new_n22514__ = new_new_n22511__ & ~new_new_n22513__;
  assign new_new_n22515__ = pi14 & ~new_new_n22514__;
  assign new_new_n22516__ = ~pi13 & ~new_new_n15362__;
  assign new_new_n22517__ = pi13 & new_new_n15362__;
  assign new_new_n22518__ = new_new_n6994__ & ~new_new_n22516__;
  assign new_new_n22519__ = ~new_new_n22517__ & new_new_n22518__;
  assign new_new_n22520__ = new_new_n16768__ & new_new_n22519__;
  assign new_new_n22521__ = new_new_n6994__ & ~new_new_n16769__;
  assign new_new_n22522__ = ~pi14 & new_new_n22511__;
  assign new_new_n22523__ = ~new_new_n22521__ & new_new_n22522__;
  assign new_new_n22524__ = ~new_new_n22515__ & ~new_new_n22520__;
  assign new_new_n22525__ = ~new_new_n22523__ & new_new_n22524__;
  assign new_new_n22526__ = ~new_new_n21949__ & ~new_new_n21950__;
  assign new_new_n22527__ = new_new_n22344__ & ~new_new_n22526__;
  assign new_new_n22528__ = ~new_new_n22344__ & new_new_n22526__;
  assign new_new_n22529__ = ~new_new_n22527__ & ~new_new_n22528__;
  assign new_new_n22530__ = ~new_new_n22525__ & ~new_new_n22529__;
  assign new_new_n22531__ = new_new_n22525__ & new_new_n22529__;
  assign new_new_n22532__ = ~new_new_n22327__ & ~new_new_n22328__;
  assign new_new_n22533__ = ~new_new_n22342__ & new_new_n22532__;
  assign new_new_n22534__ = new_new_n22342__ & ~new_new_n22532__;
  assign new_new_n22535__ = ~new_new_n22533__ & ~new_new_n22534__;
  assign new_new_n22536__ = new_new_n6991__ & ~new_new_n15471__;
  assign new_new_n22537__ = new_new_n6985__ & new_new_n15464__;
  assign new_new_n22538__ = ~new_new_n22536__ & ~new_new_n22537__;
  assign new_new_n22539__ = new_new_n6994__ & ~new_new_n15439__;
  assign new_new_n22540__ = ~new_new_n17240__ & new_new_n22539__;
  assign new_new_n22541__ = new_new_n22538__ & ~new_new_n22540__;
  assign new_new_n22542__ = pi14 & ~new_new_n22541__;
  assign new_new_n22543__ = ~pi13 & ~new_new_n15439__;
  assign new_new_n22544__ = pi13 & ~new_new_n17240__;
  assign new_new_n22545__ = new_new_n15439__ & new_new_n17239__;
  assign new_new_n22546__ = new_new_n6994__ & ~new_new_n22545__;
  assign new_new_n22547__ = ~new_new_n22543__ & ~new_new_n22544__;
  assign new_new_n22548__ = new_new_n22546__ & new_new_n22547__;
  assign new_new_n22549__ = ~pi14 & new_new_n22538__;
  assign new_new_n22550__ = ~new_new_n22546__ & new_new_n22549__;
  assign new_new_n22551__ = ~new_new_n22542__ & ~new_new_n22550__;
  assign new_new_n22552__ = ~new_new_n22548__ & new_new_n22551__;
  assign new_new_n22553__ = new_new_n21794__ & ~new_new_n22306__;
  assign new_new_n22554__ = ~new_new_n21794__ & new_new_n22306__;
  assign new_new_n22555__ = ~new_new_n22553__ & ~new_new_n22554__;
  assign new_new_n22556__ = new_new_n21807__ & new_new_n22555__;
  assign new_new_n22557__ = ~new_new_n21807__ & ~new_new_n22555__;
  assign new_new_n22558__ = ~new_new_n22556__ & ~new_new_n22557__;
  assign new_new_n22559__ = new_new_n22321__ & ~new_new_n22558__;
  assign new_new_n22560__ = ~new_new_n22321__ & new_new_n22558__;
  assign new_new_n22561__ = ~new_new_n22559__ & ~new_new_n22560__;
  assign new_new_n22562__ = new_new_n22318__ & new_new_n22561__;
  assign new_new_n22563__ = ~new_new_n22318__ & ~new_new_n22561__;
  assign new_new_n22564__ = ~new_new_n22562__ & ~new_new_n22563__;
  assign new_new_n22565__ = ~new_new_n22552__ & new_new_n22564__;
  assign new_new_n22566__ = new_new_n22552__ & ~new_new_n22564__;
  assign new_new_n22567__ = new_new_n6991__ & ~new_new_n15809__;
  assign new_new_n22568__ = new_new_n6985__ & ~new_new_n15471__;
  assign new_new_n22569__ = ~new_new_n22567__ & ~new_new_n22568__;
  assign new_new_n22570__ = new_new_n6994__ & new_new_n15464__;
  assign new_new_n22571__ = new_new_n15819__ & new_new_n22570__;
  assign new_new_n22572__ = new_new_n22569__ & ~new_new_n22571__;
  assign new_new_n22573__ = ~pi14 & ~new_new_n22572__;
  assign new_new_n22574__ = pi13 & new_new_n15464__;
  assign new_new_n22575__ = ~new_new_n15464__ & ~new_new_n15819__;
  assign new_new_n22576__ = new_new_n6994__ & ~new_new_n22575__;
  assign new_new_n22577__ = ~pi13 & new_new_n15819__;
  assign new_new_n22578__ = ~new_new_n22574__ & ~new_new_n22577__;
  assign new_new_n22579__ = new_new_n22576__ & new_new_n22578__;
  assign new_new_n22580__ = pi14 & new_new_n22569__;
  assign new_new_n22581__ = ~new_new_n22576__ & new_new_n22580__;
  assign new_new_n22582__ = ~new_new_n22573__ & ~new_new_n22579__;
  assign new_new_n22583__ = ~new_new_n22581__ & new_new_n22582__;
  assign new_new_n22584__ = ~new_new_n22007__ & ~new_new_n22008__;
  assign new_new_n22585__ = ~new_new_n22302__ & new_new_n22584__;
  assign new_new_n22586__ = new_new_n22302__ & ~new_new_n22584__;
  assign new_new_n22587__ = ~new_new_n22585__ & ~new_new_n22586__;
  assign new_new_n22588__ = new_new_n6985__ & ~new_new_n15487__;
  assign new_new_n22589__ = new_new_n6991__ & new_new_n15524__;
  assign new_new_n22590__ = ~new_new_n22588__ & ~new_new_n22589__;
  assign new_new_n22591__ = new_new_n6994__ & ~new_new_n15809__;
  assign new_new_n22592__ = new_new_n18020__ & new_new_n22591__;
  assign new_new_n22593__ = new_new_n22590__ & ~new_new_n22592__;
  assign new_new_n22594__ = pi14 & ~new_new_n22593__;
  assign new_new_n22595__ = ~pi13 & ~new_new_n20943__;
  assign new_new_n22596__ = pi13 & ~new_new_n18018__;
  assign new_new_n22597__ = new_new_n6994__ & ~new_new_n22595__;
  assign new_new_n22598__ = ~new_new_n22596__ & new_new_n22597__;
  assign new_new_n22599__ = new_new_n6994__ & ~new_new_n18019__;
  assign new_new_n22600__ = ~pi14 & new_new_n22590__;
  assign new_new_n22601__ = ~new_new_n22599__ & new_new_n22600__;
  assign new_new_n22602__ = ~new_new_n22598__ & ~new_new_n22601__;
  assign new_new_n22603__ = ~new_new_n22594__ & new_new_n22602__;
  assign new_new_n22604__ = new_new_n6985__ & new_new_n15520__;
  assign new_new_n22605__ = new_new_n6991__ & ~new_new_n15533__;
  assign new_new_n22606__ = ~new_new_n22604__ & ~new_new_n22605__;
  assign new_new_n22607__ = new_new_n6994__ & ~new_new_n18914__;
  assign new_new_n22608__ = pi14 & ~new_new_n22607__;
  assign new_new_n22609__ = new_new_n8388__ & new_new_n21477__;
  assign new_new_n22610__ = ~new_new_n22608__ & ~new_new_n22609__;
  assign new_new_n22611__ = new_new_n22606__ & ~new_new_n22610__;
  assign new_new_n22612__ = new_new_n6994__ & new_new_n18923__;
  assign new_new_n22613__ = new_new_n22606__ & ~new_new_n22612__;
  assign new_new_n22614__ = ~pi14 & ~new_new_n22613__;
  assign new_new_n22615__ = new_new_n8820__ & ~new_new_n15524__;
  assign new_new_n22616__ = new_new_n18913__ & new_new_n22615__;
  assign new_new_n22617__ = ~new_new_n22614__ & ~new_new_n22616__;
  assign new_new_n22618__ = ~new_new_n22611__ & new_new_n22617__;
  assign new_new_n22619__ = ~pi13 & new_new_n19730__;
  assign new_new_n22620__ = pi13 & ~new_new_n15520__;
  assign new_new_n22621__ = new_new_n19731__ & new_new_n22620__;
  assign new_new_n22622__ = ~new_new_n22619__ & ~new_new_n22621__;
  assign new_new_n22623__ = new_new_n6994__ & ~new_new_n22622__;
  assign new_new_n22624__ = new_new_n6991__ & new_new_n15767__;
  assign new_new_n22625__ = new_new_n6985__ & ~new_new_n15533__;
  assign new_new_n22626__ = ~new_new_n22624__ & ~new_new_n22625__;
  assign new_new_n22627__ = new_new_n6994__ & new_new_n15520__;
  assign new_new_n22628__ = new_new_n19731__ & new_new_n22627__;
  assign new_new_n22629__ = new_new_n22626__ & ~new_new_n22628__;
  assign new_new_n22630__ = ~pi14 & ~new_new_n22629__;
  assign new_new_n22631__ = new_new_n6994__ & ~new_new_n18432__;
  assign new_new_n22632__ = pi14 & new_new_n22626__;
  assign new_new_n22633__ = ~new_new_n22631__ & new_new_n22632__;
  assign new_new_n22634__ = ~new_new_n22623__ & ~new_new_n22633__;
  assign new_new_n22635__ = ~new_new_n22630__ & new_new_n22634__;
  assign new_new_n22636__ = new_new_n6991__ & new_new_n15560__;
  assign new_new_n22637__ = new_new_n6985__ & new_new_n15767__;
  assign new_new_n22638__ = ~new_new_n22636__ & ~new_new_n22637__;
  assign new_new_n22639__ = new_new_n6994__ & ~new_new_n15533__;
  assign new_new_n22640__ = new_new_n19893__ & new_new_n22639__;
  assign new_new_n22641__ = new_new_n22638__ & ~new_new_n22640__;
  assign new_new_n22642__ = pi14 & ~new_new_n22641__;
  assign new_new_n22643__ = ~pi13 & ~new_new_n15533__;
  assign new_new_n22644__ = pi13 & new_new_n15533__;
  assign new_new_n22645__ = new_new_n6994__ & ~new_new_n22643__;
  assign new_new_n22646__ = ~new_new_n22644__ & new_new_n22645__;
  assign new_new_n22647__ = new_new_n19890__ & new_new_n22646__;
  assign new_new_n22648__ = new_new_n6994__ & ~new_new_n19892__;
  assign new_new_n22649__ = ~pi14 & new_new_n22638__;
  assign new_new_n22650__ = ~new_new_n22648__ & new_new_n22649__;
  assign new_new_n22651__ = ~new_new_n22647__ & ~new_new_n22650__;
  assign new_new_n22652__ = ~new_new_n22642__ & new_new_n22651__;
  assign new_new_n22653__ = new_new_n6991__ & new_new_n15572__;
  assign new_new_n22654__ = new_new_n6985__ & new_new_n15560__;
  assign new_new_n22655__ = ~new_new_n22653__ & ~new_new_n22654__;
  assign new_new_n22656__ = new_new_n6994__ & new_new_n15767__;
  assign new_new_n22657__ = ~new_new_n18454__ & new_new_n22656__;
  assign new_new_n22658__ = new_new_n22655__ & ~new_new_n22657__;
  assign new_new_n22659__ = ~pi14 & ~new_new_n22658__;
  assign new_new_n22660__ = pi13 & new_new_n15767__;
  assign new_new_n22661__ = ~new_new_n15767__ & new_new_n18454__;
  assign new_new_n22662__ = new_new_n6994__ & ~new_new_n22661__;
  assign new_new_n22663__ = ~pi13 & ~new_new_n18454__;
  assign new_new_n22664__ = ~new_new_n22660__ & ~new_new_n22663__;
  assign new_new_n22665__ = new_new_n22662__ & new_new_n22664__;
  assign new_new_n22666__ = pi14 & new_new_n22655__;
  assign new_new_n22667__ = ~new_new_n22662__ & new_new_n22666__;
  assign new_new_n22668__ = ~new_new_n22659__ & ~new_new_n22665__;
  assign new_new_n22669__ = ~new_new_n22667__ & new_new_n22668__;
  assign new_new_n22670__ = ~new_new_n22215__ & ~new_new_n22216__;
  assign new_new_n22671__ = new_new_n22225__ & new_new_n22670__;
  assign new_new_n22672__ = ~new_new_n22225__ & ~new_new_n22670__;
  assign new_new_n22673__ = ~new_new_n22671__ & ~new_new_n22672__;
  assign new_new_n22674__ = new_new_n22669__ & ~new_new_n22673__;
  assign new_new_n22675__ = ~new_new_n22669__ & new_new_n22673__;
  assign new_new_n22676__ = new_new_n6991__ & ~new_new_n15638__;
  assign new_new_n22677__ = new_new_n6985__ & new_new_n15743__;
  assign new_new_n22678__ = ~new_new_n22676__ & ~new_new_n22677__;
  assign new_new_n22679__ = new_new_n6994__ & ~new_new_n15615__;
  assign new_new_n22680__ = new_new_n19005__ & new_new_n22679__;
  assign new_new_n22681__ = new_new_n22678__ & ~new_new_n22680__;
  assign new_new_n22682__ = ~pi14 & ~new_new_n22681__;
  assign new_new_n22683__ = ~pi13 & new_new_n19005__;
  assign new_new_n22684__ = new_new_n15615__ & ~new_new_n19005__;
  assign new_new_n22685__ = new_new_n6994__ & ~new_new_n22684__;
  assign new_new_n22686__ = pi13 & ~new_new_n15615__;
  assign new_new_n22687__ = ~new_new_n22683__ & ~new_new_n22686__;
  assign new_new_n22688__ = new_new_n22685__ & new_new_n22687__;
  assign new_new_n22689__ = pi14 & new_new_n22678__;
  assign new_new_n22690__ = ~new_new_n22685__ & new_new_n22689__;
  assign new_new_n22691__ = ~new_new_n22682__ & ~new_new_n22688__;
  assign new_new_n22692__ = ~new_new_n22690__ & new_new_n22691__;
  assign new_new_n22693__ = new_new_n6991__ & ~new_new_n15582__;
  assign new_new_n22694__ = new_new_n6985__ & ~new_new_n15638__;
  assign new_new_n22695__ = ~new_new_n22693__ & ~new_new_n22694__;
  assign new_new_n22696__ = new_new_n6994__ & new_new_n15743__;
  assign new_new_n22697__ = ~new_new_n19491__ & new_new_n22696__;
  assign new_new_n22698__ = new_new_n22695__ & ~new_new_n22697__;
  assign new_new_n22699__ = pi14 & ~new_new_n22698__;
  assign new_new_n22700__ = new_new_n6994__ & ~new_new_n19492__;
  assign new_new_n22701__ = pi13 & new_new_n19494__;
  assign new_new_n22702__ = ~pi13 & new_new_n15743__;
  assign new_new_n22703__ = new_new_n22700__ & ~new_new_n22702__;
  assign new_new_n22704__ = ~new_new_n22701__ & new_new_n22703__;
  assign new_new_n22705__ = ~pi14 & new_new_n22695__;
  assign new_new_n22706__ = ~new_new_n22700__ & new_new_n22705__;
  assign new_new_n22707__ = ~new_new_n22699__ & ~new_new_n22706__;
  assign new_new_n22708__ = ~new_new_n22704__ & new_new_n22707__;
  assign new_new_n22709__ = ~new_new_n22149__ & ~new_new_n22150__;
  assign new_new_n22710__ = new_new_n22160__ & new_new_n22709__;
  assign new_new_n22711__ = ~new_new_n22160__ & ~new_new_n22709__;
  assign new_new_n22712__ = ~new_new_n22710__ & ~new_new_n22711__;
  assign new_new_n22713__ = ~new_new_n22708__ & ~new_new_n22712__;
  assign new_new_n22714__ = new_new_n22708__ & new_new_n22712__;
  assign new_new_n22715__ = new_new_n22121__ & ~new_new_n22137__;
  assign new_new_n22716__ = new_new_n22141__ & ~new_new_n22715__;
  assign new_new_n22717__ = ~new_new_n22121__ & new_new_n22137__;
  assign new_new_n22718__ = ~new_new_n22715__ & ~new_new_n22717__;
  assign new_new_n22719__ = ~new_new_n22124__ & ~new_new_n22718__;
  assign new_new_n22720__ = new_new_n22122__ & ~new_new_n22137__;
  assign new_new_n22721__ = ~new_new_n22716__ & ~new_new_n22720__;
  assign new_new_n22722__ = ~new_new_n22719__ & new_new_n22721__;
  assign new_new_n22723__ = new_new_n6991__ & ~new_new_n15710__;
  assign new_new_n22724__ = new_new_n6985__ & ~new_new_n15647__;
  assign new_new_n22725__ = ~new_new_n22723__ & ~new_new_n22724__;
  assign new_new_n22726__ = new_new_n6994__ & new_new_n19058__;
  assign new_new_n22727__ = new_new_n22725__ & ~new_new_n22726__;
  assign new_new_n22728__ = pi14 & ~new_new_n22727__;
  assign new_new_n22729__ = ~pi13 & ~new_new_n15582__;
  assign new_new_n22730__ = new_new_n6994__ & ~new_new_n19052__;
  assign new_new_n22731__ = pi13 & ~new_new_n15736__;
  assign new_new_n22732__ = ~new_new_n22729__ & ~new_new_n22731__;
  assign new_new_n22733__ = new_new_n22730__ & new_new_n22732__;
  assign new_new_n22734__ = ~pi14 & new_new_n22725__;
  assign new_new_n22735__ = ~new_new_n22730__ & new_new_n22734__;
  assign new_new_n22736__ = ~new_new_n22733__ & ~new_new_n22735__;
  assign new_new_n22737__ = ~new_new_n22728__ & new_new_n22736__;
  assign new_new_n22738__ = ~new_new_n22108__ & ~new_new_n22109__;
  assign new_new_n22739__ = new_new_n22119__ & ~new_new_n22738__;
  assign new_new_n22740__ = ~new_new_n22119__ & new_new_n22738__;
  assign new_new_n22741__ = ~new_new_n22739__ & ~new_new_n22740__;
  assign new_new_n22742__ = new_new_n22737__ & new_new_n22741__;
  assign new_new_n22743__ = ~new_new_n22737__ & ~new_new_n22741__;
  assign new_new_n22744__ = new_new_n6985__ & ~new_new_n15710__;
  assign new_new_n22745__ = new_new_n6991__ & new_new_n15656__;
  assign new_new_n22746__ = ~new_new_n22744__ & ~new_new_n22745__;
  assign new_new_n22747__ = new_new_n6994__ & ~new_new_n15647__;
  assign new_new_n22748__ = ~new_new_n19118__ & new_new_n22747__;
  assign new_new_n22749__ = new_new_n22746__ & ~new_new_n22748__;
  assign new_new_n22750__ = ~pi14 & ~new_new_n22749__;
  assign new_new_n22751__ = pi13 & ~new_new_n15647__;
  assign new_new_n22752__ = ~pi13 & ~new_new_n19118__;
  assign new_new_n22753__ = new_new_n15647__ & new_new_n19117__;
  assign new_new_n22754__ = new_new_n6994__ & ~new_new_n22753__;
  assign new_new_n22755__ = ~new_new_n22751__ & ~new_new_n22752__;
  assign new_new_n22756__ = new_new_n22754__ & new_new_n22755__;
  assign new_new_n22757__ = pi14 & new_new_n22746__;
  assign new_new_n22758__ = ~new_new_n22754__ & new_new_n22757__;
  assign new_new_n22759__ = ~new_new_n22750__ & ~new_new_n22758__;
  assign new_new_n22760__ = ~new_new_n22756__ & new_new_n22759__;
  assign new_new_n22761__ = new_new_n6991__ & new_new_n15643__;
  assign new_new_n22762__ = new_new_n6985__ & new_new_n15656__;
  assign new_new_n22763__ = ~new_new_n22761__ & ~new_new_n22762__;
  assign new_new_n22764__ = ~new_new_n15710__ & ~new_new_n19466__;
  assign new_new_n22765__ = new_new_n6994__ & new_new_n22764__;
  assign new_new_n22766__ = new_new_n22763__ & ~new_new_n22765__;
  assign new_new_n22767__ = pi14 & ~new_new_n22766__;
  assign new_new_n22768__ = new_new_n15710__ & ~new_new_n19466__;
  assign new_new_n22769__ = ~pi13 & ~new_new_n22768__;
  assign new_new_n22770__ = ~new_new_n15710__ & new_new_n19466__;
  assign new_new_n22771__ = pi13 & ~new_new_n22770__;
  assign new_new_n22772__ = new_new_n6994__ & ~new_new_n22769__;
  assign new_new_n22773__ = ~new_new_n22771__ & new_new_n22772__;
  assign new_new_n22774__ = new_new_n15710__ & new_new_n19466__;
  assign new_new_n22775__ = new_new_n6994__ & ~new_new_n22774__;
  assign new_new_n22776__ = ~pi14 & new_new_n22763__;
  assign new_new_n22777__ = ~new_new_n22775__ & new_new_n22776__;
  assign new_new_n22778__ = ~new_new_n22767__ & ~new_new_n22777__;
  assign new_new_n22779__ = ~new_new_n22773__ & new_new_n22778__;
  assign new_new_n22780__ = pi17 & new_new_n6958__;
  assign new_new_n22781__ = ~new_new_n6968__ & ~new_new_n22780__;
  assign new_new_n22782__ = pi17 & ~new_new_n15673__;
  assign new_new_n22783__ = ~new_new_n15668__ & ~new_new_n22782__;
  assign new_new_n22784__ = ~new_new_n6958__ & new_new_n22782__;
  assign new_new_n22785__ = new_new_n15668__ & new_new_n22784__;
  assign new_new_n22786__ = ~new_new_n22781__ & ~new_new_n22783__;
  assign new_new_n22787__ = ~new_new_n22785__ & new_new_n22786__;
  assign new_new_n22788__ = new_new_n22081__ & ~new_new_n22787__;
  assign new_new_n22789__ = new_new_n6968__ & ~new_new_n15674__;
  assign new_new_n22790__ = ~new_new_n20628__ & new_new_n22780__;
  assign new_new_n22791__ = ~new_new_n22789__ & new_new_n22790__;
  assign new_new_n22792__ = ~new_new_n22081__ & new_new_n22791__;
  assign new_new_n22793__ = ~new_new_n22788__ & ~new_new_n22792__;
  assign new_new_n22794__ = new_new_n22779__ & new_new_n22793__;
  assign new_new_n22795__ = new_new_n6991__ & new_new_n15668__;
  assign new_new_n22796__ = new_new_n6985__ & ~new_new_n15661__;
  assign new_new_n22797__ = ~new_new_n22795__ & ~new_new_n22796__;
  assign new_new_n22798__ = new_new_n6994__ & ~new_new_n20177__;
  assign new_new_n22799__ = ~pi14 & ~new_new_n22798__;
  assign new_new_n22800__ = new_new_n8820__ & new_new_n21085__;
  assign new_new_n22801__ = ~new_new_n22799__ & ~new_new_n22800__;
  assign new_new_n22802__ = new_new_n22797__ & ~new_new_n22801__;
  assign new_new_n22803__ = new_new_n6994__ & new_new_n20187__;
  assign new_new_n22804__ = new_new_n22797__ & ~new_new_n22803__;
  assign new_new_n22805__ = pi14 & ~new_new_n22804__;
  assign new_new_n22806__ = new_new_n8388__ & ~new_new_n15643__;
  assign new_new_n22807__ = new_new_n20176__ & new_new_n22806__;
  assign new_new_n22808__ = ~new_new_n22805__ & ~new_new_n22807__;
  assign new_new_n22809__ = ~new_new_n22802__ & new_new_n22808__;
  assign new_new_n22810__ = new_new_n6991__ & ~new_new_n15673__;
  assign new_new_n22811__ = new_new_n6985__ & new_new_n15668__;
  assign new_new_n22812__ = ~new_new_n22810__ & ~new_new_n22811__;
  assign new_new_n22813__ = new_new_n6994__ & ~new_new_n20196__;
  assign new_new_n22814__ = pi14 & ~new_new_n22813__;
  assign new_new_n22815__ = new_new_n8388__ & new_new_n20195__;
  assign new_new_n22816__ = ~new_new_n15661__ & new_new_n22815__;
  assign new_new_n22817__ = ~new_new_n22814__ & ~new_new_n22816__;
  assign new_new_n22818__ = new_new_n22812__ & ~new_new_n22817__;
  assign new_new_n22819__ = new_new_n6994__ & new_new_n20206__;
  assign new_new_n22820__ = new_new_n22812__ & ~new_new_n22819__;
  assign new_new_n22821__ = ~pi14 & ~new_new_n22820__;
  assign new_new_n22822__ = new_new_n8820__ & new_new_n15668__;
  assign new_new_n22823__ = new_new_n15679__ & new_new_n22822__;
  assign new_new_n22824__ = ~new_new_n22821__ & ~new_new_n22823__;
  assign new_new_n22825__ = ~new_new_n22818__ & new_new_n22824__;
  assign new_new_n22826__ = new_new_n6994__ & ~new_new_n20628__;
  assign new_new_n22827__ = ~new_new_n15673__ & new_new_n19825__;
  assign new_new_n22828__ = pi14 & ~new_new_n22827__;
  assign new_new_n22829__ = ~new_new_n22826__ & new_new_n22828__;
  assign new_new_n22830__ = ~new_new_n22825__ & new_new_n22829__;
  assign new_new_n22831__ = new_new_n6958__ & ~new_new_n15673__;
  assign new_new_n22832__ = ~new_new_n22830__ & ~new_new_n22831__;
  assign new_new_n22833__ = new_new_n22809__ & ~new_new_n22832__;
  assign new_new_n22834__ = new_new_n6991__ & ~new_new_n15661__;
  assign new_new_n22835__ = new_new_n6985__ & new_new_n15643__;
  assign new_new_n22836__ = ~new_new_n22834__ & ~new_new_n22835__;
  assign new_new_n22837__ = new_new_n6994__ & new_new_n15656__;
  assign new_new_n22838__ = new_new_n15687__ & new_new_n22837__;
  assign new_new_n22839__ = new_new_n22836__ & ~new_new_n22838__;
  assign new_new_n22840__ = pi14 & ~new_new_n22839__;
  assign new_new_n22841__ = pi13 & new_new_n15686__;
  assign new_new_n22842__ = ~pi13 & ~new_new_n15656__;
  assign new_new_n22843__ = new_new_n15677__ & new_new_n22842__;
  assign new_new_n22844__ = ~new_new_n22841__ & ~new_new_n22843__;
  assign new_new_n22845__ = new_new_n6994__ & ~new_new_n22844__;
  assign new_new_n22846__ = new_new_n6994__ & ~new_new_n15678__;
  assign new_new_n22847__ = ~pi14 & new_new_n22836__;
  assign new_new_n22848__ = ~new_new_n22846__ & new_new_n22847__;
  assign new_new_n22849__ = ~new_new_n22845__ & ~new_new_n22848__;
  assign new_new_n22850__ = ~new_new_n22840__ & new_new_n22849__;
  assign new_new_n22851__ = new_new_n22833__ & new_new_n22850__;
  assign new_new_n22852__ = new_new_n6958__ & new_new_n15668__;
  assign new_new_n22853__ = new_new_n15673__ & ~new_new_n22852__;
  assign new_new_n22854__ = new_new_n6966__ & new_new_n15674__;
  assign new_new_n22855__ = ~new_new_n6956__ & new_new_n15668__;
  assign new_new_n22856__ = new_new_n6967__ & ~new_new_n22855__;
  assign new_new_n22857__ = ~new_new_n6962__ & ~new_new_n22853__;
  assign new_new_n22858__ = ~new_new_n22854__ & ~new_new_n22856__;
  assign new_new_n22859__ = new_new_n22857__ & new_new_n22858__;
  assign new_new_n22860__ = ~new_new_n22851__ & ~new_new_n22859__;
  assign new_new_n22861__ = ~new_new_n22779__ & ~new_new_n22793__;
  assign new_new_n22862__ = ~new_new_n22833__ & ~new_new_n22850__;
  assign new_new_n22863__ = ~new_new_n22860__ & ~new_new_n22862__;
  assign new_new_n22864__ = ~new_new_n22861__ & new_new_n22863__;
  assign new_new_n22865__ = ~new_new_n22794__ & ~new_new_n22864__;
  assign new_new_n22866__ = ~new_new_n22760__ & ~new_new_n22865__;
  assign new_new_n22867__ = new_new_n22760__ & new_new_n22865__;
  assign new_new_n22868__ = new_new_n22084__ & new_new_n22098__;
  assign new_new_n22869__ = ~new_new_n22099__ & ~new_new_n22868__;
  assign new_new_n22870__ = new_new_n22071__ & new_new_n22083__;
  assign new_new_n22871__ = ~new_new_n22869__ & ~new_new_n22870__;
  assign new_new_n22872__ = ~new_new_n22867__ & ~new_new_n22871__;
  assign new_new_n22873__ = ~new_new_n22866__ & ~new_new_n22872__;
  assign new_new_n22874__ = ~new_new_n22743__ & ~new_new_n22873__;
  assign new_new_n22875__ = ~new_new_n22742__ & ~new_new_n22874__;
  assign new_new_n22876__ = new_new_n22722__ & new_new_n22875__;
  assign new_new_n22877__ = ~new_new_n22722__ & ~new_new_n22875__;
  assign new_new_n22878__ = new_new_n6991__ & ~new_new_n15647__;
  assign new_new_n22879__ = new_new_n6985__ & ~new_new_n15582__;
  assign new_new_n22880__ = ~new_new_n22878__ & ~new_new_n22879__;
  assign new_new_n22881__ = new_new_n6994__ & ~new_new_n15638__;
  assign new_new_n22882__ = new_new_n19487__ & new_new_n22881__;
  assign new_new_n22883__ = new_new_n22880__ & ~new_new_n22882__;
  assign new_new_n22884__ = pi14 & ~new_new_n22883__;
  assign new_new_n22885__ = pi13 & new_new_n19487__;
  assign new_new_n22886__ = new_new_n6994__ & ~new_new_n19488__;
  assign new_new_n22887__ = ~pi13 & ~new_new_n15638__;
  assign new_new_n22888__ = ~new_new_n22885__ & ~new_new_n22887__;
  assign new_new_n22889__ = new_new_n22886__ & new_new_n22888__;
  assign new_new_n22890__ = ~pi14 & new_new_n22880__;
  assign new_new_n22891__ = ~new_new_n22886__ & new_new_n22890__;
  assign new_new_n22892__ = ~new_new_n22884__ & ~new_new_n22889__;
  assign new_new_n22893__ = ~new_new_n22891__ & new_new_n22892__;
  assign new_new_n22894__ = ~new_new_n22877__ & ~new_new_n22893__;
  assign new_new_n22895__ = ~new_new_n22876__ & ~new_new_n22894__;
  assign new_new_n22896__ = ~new_new_n22714__ & ~new_new_n22895__;
  assign new_new_n22897__ = ~new_new_n22713__ & ~new_new_n22896__;
  assign new_new_n22898__ = ~new_new_n22692__ & new_new_n22897__;
  assign new_new_n22899__ = new_new_n22692__ & ~new_new_n22897__;
  assign new_new_n22900__ = ~new_new_n22163__ & ~new_new_n22164__;
  assign new_new_n22901__ = new_new_n22168__ & ~new_new_n22900__;
  assign new_new_n22902__ = ~new_new_n22168__ & new_new_n22900__;
  assign new_new_n22903__ = ~new_new_n22901__ & ~new_new_n22902__;
  assign new_new_n22904__ = ~new_new_n22899__ & new_new_n22903__;
  assign new_new_n22905__ = ~new_new_n22898__ & ~new_new_n22904__;
  assign new_new_n22906__ = ~new_new_n22171__ & ~new_new_n22172__;
  assign new_new_n22907__ = new_new_n6985__ & ~new_new_n15615__;
  assign new_new_n22908__ = new_new_n6991__ & new_new_n15743__;
  assign new_new_n22909__ = ~new_new_n22907__ & ~new_new_n22908__;
  assign new_new_n22910__ = new_new_n6994__ & new_new_n15564__;
  assign new_new_n22911__ = new_new_n18512__ & new_new_n22910__;
  assign new_new_n22912__ = new_new_n22909__ & ~new_new_n22911__;
  assign new_new_n22913__ = ~pi14 & ~new_new_n22912__;
  assign new_new_n22914__ = new_new_n6994__ & ~new_new_n20738__;
  assign new_new_n22915__ = pi14 & new_new_n22909__;
  assign new_new_n22916__ = ~new_new_n22914__ & new_new_n22915__;
  assign new_new_n22917__ = ~pi13 & ~new_new_n20743__;
  assign new_new_n22918__ = pi13 & ~new_new_n20741__;
  assign new_new_n22919__ = new_new_n6994__ & ~new_new_n22917__;
  assign new_new_n22920__ = ~new_new_n22918__ & new_new_n22919__;
  assign new_new_n22921__ = ~new_new_n22913__ & ~new_new_n22916__;
  assign new_new_n22922__ = ~new_new_n22920__ & new_new_n22921__;
  assign new_new_n22923__ = new_new_n22906__ & ~new_new_n22922__;
  assign new_new_n22924__ = ~new_new_n22906__ & new_new_n22922__;
  assign new_new_n22925__ = ~new_new_n22923__ & ~new_new_n22924__;
  assign new_new_n22926__ = new_new_n22184__ & new_new_n22925__;
  assign new_new_n22927__ = ~new_new_n22184__ & ~new_new_n22925__;
  assign new_new_n22928__ = ~new_new_n22926__ & ~new_new_n22927__;
  assign new_new_n22929__ = new_new_n22905__ & new_new_n22928__;
  assign new_new_n22930__ = new_new_n22922__ & ~new_new_n22928__;
  assign new_new_n22931__ = ~new_new_n22929__ & ~new_new_n22930__;
  assign new_new_n22932__ = ~new_new_n22187__ & ~new_new_n22188__;
  assign new_new_n22933__ = new_new_n22198__ & new_new_n22932__;
  assign new_new_n22934__ = ~new_new_n22198__ & ~new_new_n22932__;
  assign new_new_n22935__ = ~new_new_n22933__ & ~new_new_n22934__;
  assign new_new_n22936__ = ~new_new_n22931__ & ~new_new_n22935__;
  assign new_new_n22937__ = new_new_n22931__ & new_new_n22935__;
  assign new_new_n22938__ = new_new_n8820__ & new_new_n20113__;
  assign new_new_n22939__ = new_new_n6991__ & ~new_new_n15615__;
  assign new_new_n22940__ = new_new_n6985__ & new_new_n15564__;
  assign new_new_n22941__ = ~new_new_n22939__ & ~new_new_n22940__;
  assign new_new_n22942__ = new_new_n6994__ & ~new_new_n20528__;
  assign new_new_n22943__ = pi14 & ~new_new_n22942__;
  assign new_new_n22944__ = new_new_n8388__ & new_new_n15572__;
  assign new_new_n22945__ = new_new_n19534__ & new_new_n22944__;
  assign new_new_n22946__ = ~new_new_n22943__ & ~new_new_n22945__;
  assign new_new_n22947__ = new_new_n22941__ & ~new_new_n22946__;
  assign new_new_n22948__ = new_new_n6994__ & new_new_n20111__;
  assign new_new_n22949__ = new_new_n22941__ & ~new_new_n22948__;
  assign new_new_n22950__ = ~pi14 & ~new_new_n22949__;
  assign new_new_n22951__ = ~new_new_n22938__ & ~new_new_n22950__;
  assign new_new_n22952__ = ~new_new_n22947__ & new_new_n22951__;
  assign new_new_n22953__ = ~new_new_n22937__ & new_new_n22952__;
  assign new_new_n22954__ = ~new_new_n22936__ & ~new_new_n22953__;
  assign new_new_n22955__ = ~new_new_n22201__ & ~new_new_n22202__;
  assign new_new_n22956__ = new_new_n22212__ & ~new_new_n22955__;
  assign new_new_n22957__ = ~new_new_n22212__ & new_new_n22955__;
  assign new_new_n22958__ = ~new_new_n22956__ & ~new_new_n22957__;
  assign new_new_n22959__ = ~new_new_n22954__ & new_new_n22958__;
  assign new_new_n22960__ = new_new_n22954__ & ~new_new_n22958__;
  assign new_new_n22961__ = ~pi13 & new_new_n18943__;
  assign new_new_n22962__ = pi13 & ~new_new_n15560__;
  assign new_new_n22963__ = new_new_n18944__ & new_new_n22962__;
  assign new_new_n22964__ = ~new_new_n22961__ & ~new_new_n22963__;
  assign new_new_n22965__ = new_new_n6994__ & ~new_new_n22964__;
  assign new_new_n22966__ = new_new_n6991__ & new_new_n15564__;
  assign new_new_n22967__ = new_new_n6985__ & new_new_n15572__;
  assign new_new_n22968__ = ~new_new_n22966__ & ~new_new_n22967__;
  assign new_new_n22969__ = new_new_n6994__ & new_new_n15560__;
  assign new_new_n22970__ = new_new_n18944__ & new_new_n22969__;
  assign new_new_n22971__ = new_new_n22968__ & ~new_new_n22970__;
  assign new_new_n22972__ = ~pi14 & ~new_new_n22971__;
  assign new_new_n22973__ = new_new_n6994__ & new_new_n18939__;
  assign new_new_n22974__ = pi14 & new_new_n22968__;
  assign new_new_n22975__ = ~new_new_n22973__ & new_new_n22974__;
  assign new_new_n22976__ = ~new_new_n22965__ & ~new_new_n22975__;
  assign new_new_n22977__ = ~new_new_n22972__ & new_new_n22976__;
  assign new_new_n22978__ = ~new_new_n22960__ & new_new_n22977__;
  assign new_new_n22979__ = ~new_new_n22959__ & ~new_new_n22978__;
  assign new_new_n22980__ = ~new_new_n22675__ & ~new_new_n22979__;
  assign new_new_n22981__ = ~new_new_n22674__ & ~new_new_n22980__;
  assign new_new_n22982__ = ~new_new_n22652__ & ~new_new_n22981__;
  assign new_new_n22983__ = new_new_n22652__ & new_new_n22981__;
  assign new_new_n22984__ = ~new_new_n22228__ & ~new_new_n22229__;
  assign new_new_n22985__ = ~new_new_n22241__ & new_new_n22984__;
  assign new_new_n22986__ = new_new_n22241__ & ~new_new_n22984__;
  assign new_new_n22987__ = ~new_new_n22985__ & ~new_new_n22986__;
  assign new_new_n22988__ = ~new_new_n22983__ & ~new_new_n22987__;
  assign new_new_n22989__ = ~new_new_n22982__ & ~new_new_n22988__;
  assign new_new_n22990__ = ~new_new_n22635__ & new_new_n22989__;
  assign new_new_n22991__ = new_new_n22635__ & ~new_new_n22989__;
  assign new_new_n22992__ = ~new_new_n22244__ & ~new_new_n22245__;
  assign new_new_n22993__ = ~new_new_n22249__ & new_new_n22992__;
  assign new_new_n22994__ = new_new_n22249__ & ~new_new_n22992__;
  assign new_new_n22995__ = ~new_new_n22993__ & ~new_new_n22994__;
  assign new_new_n22996__ = ~new_new_n22991__ & ~new_new_n22995__;
  assign new_new_n22997__ = ~new_new_n22990__ & ~new_new_n22996__;
  assign new_new_n22998__ = new_new_n22618__ & new_new_n22997__;
  assign new_new_n22999__ = ~new_new_n22618__ & ~new_new_n22997__;
  assign new_new_n23000__ = ~new_new_n22252__ & ~new_new_n22253__;
  assign new_new_n23001__ = ~new_new_n22265__ & new_new_n23000__;
  assign new_new_n23002__ = new_new_n22265__ & ~new_new_n23000__;
  assign new_new_n23003__ = ~new_new_n23001__ & ~new_new_n23002__;
  assign new_new_n23004__ = ~new_new_n22999__ & ~new_new_n23003__;
  assign new_new_n23005__ = ~new_new_n22998__ & ~new_new_n23004__;
  assign new_new_n23006__ = new_new_n6991__ & new_new_n15520__;
  assign new_new_n23007__ = new_new_n6985__ & new_new_n15524__;
  assign new_new_n23008__ = ~new_new_n23006__ & ~new_new_n23007__;
  assign new_new_n23009__ = new_new_n6994__ & ~new_new_n15487__;
  assign new_new_n23010__ = new_new_n17587__ & new_new_n23009__;
  assign new_new_n23011__ = new_new_n23008__ & ~new_new_n23010__;
  assign new_new_n23012__ = pi14 & ~new_new_n23011__;
  assign new_new_n23013__ = pi13 & new_new_n17587__;
  assign new_new_n23014__ = new_new_n15487__ & ~new_new_n17587__;
  assign new_new_n23015__ = new_new_n6994__ & ~new_new_n23014__;
  assign new_new_n23016__ = ~pi13 & ~new_new_n15487__;
  assign new_new_n23017__ = ~new_new_n23013__ & ~new_new_n23016__;
  assign new_new_n23018__ = new_new_n23015__ & new_new_n23017__;
  assign new_new_n23019__ = ~pi14 & new_new_n23008__;
  assign new_new_n23020__ = ~new_new_n23015__ & new_new_n23019__;
  assign new_new_n23021__ = ~new_new_n23012__ & ~new_new_n23018__;
  assign new_new_n23022__ = ~new_new_n23020__ & new_new_n23021__;
  assign new_new_n23023__ = ~new_new_n23005__ & ~new_new_n23022__;
  assign new_new_n23024__ = new_new_n23005__ & new_new_n23022__;
  assign new_new_n23025__ = ~new_new_n22270__ & ~new_new_n22280__;
  assign new_new_n23026__ = ~new_new_n22281__ & ~new_new_n23025__;
  assign new_new_n23027__ = ~new_new_n23024__ & ~new_new_n23026__;
  assign new_new_n23028__ = ~new_new_n23023__ & ~new_new_n23027__;
  assign new_new_n23029__ = new_new_n22603__ & new_new_n23028__;
  assign new_new_n23030__ = ~new_new_n22603__ & ~new_new_n23028__;
  assign new_new_n23031__ = ~new_new_n22287__ & ~new_new_n22288__;
  assign new_new_n23032__ = ~new_new_n22300__ & new_new_n23031__;
  assign new_new_n23033__ = new_new_n22300__ & ~new_new_n23031__;
  assign new_new_n23034__ = ~new_new_n23032__ & ~new_new_n23033__;
  assign new_new_n23035__ = ~new_new_n23030__ & new_new_n23034__;
  assign new_new_n23036__ = ~new_new_n23029__ & ~new_new_n23035__;
  assign new_new_n23037__ = ~new_new_n22587__ & ~new_new_n23036__;
  assign new_new_n23038__ = new_new_n22587__ & new_new_n23036__;
  assign new_new_n23039__ = new_new_n6985__ & ~new_new_n15809__;
  assign new_new_n23040__ = new_new_n6991__ & ~new_new_n15487__;
  assign new_new_n23041__ = ~new_new_n23039__ & ~new_new_n23040__;
  assign new_new_n23042__ = new_new_n6994__ & new_new_n18631__;
  assign new_new_n23043__ = new_new_n23041__ & ~new_new_n23042__;
  assign new_new_n23044__ = ~pi14 & ~new_new_n23043__;
  assign new_new_n23045__ = ~pi13 & new_new_n15471__;
  assign new_new_n23046__ = pi13 & ~new_new_n15471__;
  assign new_new_n23047__ = new_new_n6994__ & ~new_new_n23045__;
  assign new_new_n23048__ = ~new_new_n23046__ & new_new_n23047__;
  assign new_new_n23049__ = new_new_n18630__ & new_new_n23048__;
  assign new_new_n23050__ = new_new_n15471__ & ~new_new_n18630__;
  assign new_new_n23051__ = new_new_n6994__ & ~new_new_n23050__;
  assign new_new_n23052__ = pi14 & new_new_n23041__;
  assign new_new_n23053__ = ~new_new_n23051__ & new_new_n23052__;
  assign new_new_n23054__ = ~new_new_n23049__ & ~new_new_n23053__;
  assign new_new_n23055__ = ~new_new_n23044__ & new_new_n23054__;
  assign new_new_n23056__ = ~new_new_n23038__ & ~new_new_n23055__;
  assign new_new_n23057__ = ~new_new_n23037__ & ~new_new_n23056__;
  assign new_new_n23058__ = ~new_new_n21985__ & ~new_new_n22304__;
  assign new_new_n23059__ = ~new_new_n22305__ & ~new_new_n23058__;
  assign new_new_n23060__ = new_new_n23057__ & new_new_n23059__;
  assign new_new_n23061__ = ~new_new_n22583__ & ~new_new_n23060__;
  assign new_new_n23062__ = ~new_new_n23057__ & ~new_new_n23059__;
  assign new_new_n23063__ = ~new_new_n23061__ & ~new_new_n23062__;
  assign new_new_n23064__ = ~new_new_n22566__ & new_new_n23063__;
  assign new_new_n23065__ = ~new_new_n22565__ & ~new_new_n23064__;
  assign new_new_n23066__ = ~new_new_n22535__ & ~new_new_n23065__;
  assign new_new_n23067__ = new_new_n22535__ & new_new_n23065__;
  assign new_new_n23068__ = new_new_n6991__ & new_new_n15464__;
  assign new_new_n23069__ = new_new_n6985__ & ~new_new_n15439__;
  assign new_new_n23070__ = ~new_new_n23068__ & ~new_new_n23069__;
  assign new_new_n23071__ = new_new_n6994__ & ~new_new_n15432__;
  assign new_new_n23072__ = new_new_n17204__ & new_new_n23071__;
  assign new_new_n23073__ = new_new_n23070__ & ~new_new_n23072__;
  assign new_new_n23074__ = pi14 & ~new_new_n23073__;
  assign new_new_n23075__ = new_new_n15432__ & ~new_new_n17204__;
  assign new_new_n23076__ = new_new_n6994__ & ~new_new_n23075__;
  assign new_new_n23077__ = ~pi13 & ~new_new_n15432__;
  assign new_new_n23078__ = pi13 & new_new_n17204__;
  assign new_new_n23079__ = ~new_new_n23077__ & ~new_new_n23078__;
  assign new_new_n23080__ = new_new_n23076__ & new_new_n23079__;
  assign new_new_n23081__ = ~pi14 & new_new_n23070__;
  assign new_new_n23082__ = ~new_new_n23076__ & new_new_n23081__;
  assign new_new_n23083__ = ~new_new_n23074__ & ~new_new_n23080__;
  assign new_new_n23084__ = ~new_new_n23082__ & new_new_n23083__;
  assign new_new_n23085__ = ~new_new_n23067__ & ~new_new_n23084__;
  assign new_new_n23086__ = ~new_new_n23066__ & ~new_new_n23085__;
  assign new_new_n23087__ = ~new_new_n22531__ & ~new_new_n23086__;
  assign new_new_n23088__ = ~new_new_n22530__ & ~new_new_n23087__;
  assign new_new_n23089__ = new_new_n22508__ & ~new_new_n23088__;
  assign new_new_n23090__ = ~new_new_n22508__ & new_new_n23088__;
  assign new_new_n23091__ = ~new_new_n23089__ & ~new_new_n23090__;
  assign new_new_n23092__ = new_new_n22346__ & new_new_n23091__;
  assign new_new_n23093__ = ~new_new_n22346__ & ~new_new_n23091__;
  assign new_new_n23094__ = ~new_new_n23092__ & ~new_new_n23093__;
  assign new_new_n23095__ = new_new_n22507__ & new_new_n23094__;
  assign new_new_n23096__ = ~new_new_n23088__ & ~new_new_n23094__;
  assign new_new_n23097__ = ~new_new_n23095__ & ~new_new_n23096__;
  assign new_new_n23098__ = ~new_new_n22349__ & ~new_new_n22350__;
  assign new_new_n23099__ = new_new_n22354__ & ~new_new_n23098__;
  assign new_new_n23100__ = ~new_new_n22354__ & new_new_n23098__;
  assign new_new_n23101__ = ~new_new_n23099__ & ~new_new_n23100__;
  assign new_new_n23102__ = new_new_n23097__ & new_new_n23101__;
  assign new_new_n23103__ = ~new_new_n23097__ & ~new_new_n23101__;
  assign new_new_n23104__ = new_new_n6985__ & new_new_n15390__;
  assign new_new_n23105__ = new_new_n6991__ & ~new_new_n15362__;
  assign new_new_n23106__ = ~new_new_n23104__ & ~new_new_n23105__;
  assign new_new_n23107__ = new_new_n6994__ & ~new_new_n17364__;
  assign new_new_n23108__ = pi14 & ~new_new_n23107__;
  assign new_new_n23109__ = new_new_n6994__ & new_new_n16956__;
  assign new_new_n23110__ = ~pi13 & ~new_new_n15398__;
  assign new_new_n23111__ = new_new_n23109__ & new_new_n23110__;
  assign new_new_n23112__ = ~new_new_n23108__ & ~new_new_n23111__;
  assign new_new_n23113__ = new_new_n23106__ & ~new_new_n23112__;
  assign new_new_n23114__ = new_new_n6994__ & new_new_n17360__;
  assign new_new_n23115__ = new_new_n23106__ & ~new_new_n23114__;
  assign new_new_n23116__ = ~pi14 & ~new_new_n23115__;
  assign new_new_n23117__ = pi13 & new_new_n15398__;
  assign new_new_n23118__ = new_new_n23109__ & new_new_n23117__;
  assign new_new_n23119__ = ~new_new_n23116__ & ~new_new_n23118__;
  assign new_new_n23120__ = ~new_new_n23113__ & new_new_n23119__;
  assign new_new_n23121__ = ~new_new_n23103__ & ~new_new_n23120__;
  assign new_new_n23122__ = ~new_new_n23102__ & ~new_new_n23121__;
  assign new_new_n23123__ = ~new_new_n22491__ & ~new_new_n23122__;
  assign new_new_n23124__ = new_new_n22491__ & new_new_n23122__;
  assign new_new_n23125__ = ~new_new_n22357__ & ~new_new_n22358__;
  assign new_new_n23126__ = new_new_n22372__ & new_new_n23125__;
  assign new_new_n23127__ = ~new_new_n22372__ & ~new_new_n23125__;
  assign new_new_n23128__ = ~new_new_n23126__ & ~new_new_n23127__;
  assign new_new_n23129__ = ~new_new_n23124__ & ~new_new_n23128__;
  assign new_new_n23130__ = ~new_new_n23123__ & ~new_new_n23129__;
  assign new_new_n23131__ = new_new_n22474__ & ~new_new_n23130__;
  assign new_new_n23132__ = ~new_new_n22474__ & new_new_n23130__;
  assign new_new_n23133__ = new_new_n22374__ & ~new_new_n22397__;
  assign new_new_n23134__ = ~new_new_n22398__ & ~new_new_n23133__;
  assign new_new_n23135__ = ~new_new_n23132__ & ~new_new_n23134__;
  assign new_new_n23136__ = ~new_new_n23131__ & ~new_new_n23135__;
  assign new_new_n23137__ = ~new_new_n22405__ & ~new_new_n22406__;
  assign new_new_n23138__ = ~new_new_n22423__ & new_new_n23137__;
  assign new_new_n23139__ = new_new_n22423__ & ~new_new_n23137__;
  assign new_new_n23140__ = ~new_new_n23138__ & ~new_new_n23139__;
  assign new_new_n23141__ = new_new_n23136__ & new_new_n23140__;
  assign new_new_n23142__ = new_new_n8474__ & ~new_new_n15314__;
  assign new_new_n23143__ = ~new_new_n8479__ & new_new_n15285__;
  assign new_new_n23144__ = new_new_n8470__ & new_new_n16725__;
  assign new_new_n23145__ = ~new_new_n23142__ & ~new_new_n23143__;
  assign new_new_n23146__ = ~new_new_n23144__ & new_new_n23145__;
  assign new_new_n23147__ = new_new_n8469__ & ~new_new_n15248__;
  assign new_new_n23148__ = pi11 & ~new_new_n23147__;
  assign new_new_n23149__ = new_new_n11368__ & ~new_new_n15248__;
  assign new_new_n23150__ = ~new_new_n23148__ & ~new_new_n23149__;
  assign new_new_n23151__ = new_new_n23146__ & ~new_new_n23150__;
  assign new_new_n23152__ = ~pi11 & ~new_new_n23146__;
  assign new_new_n23153__ = ~new_new_n23151__ & ~new_new_n23152__;
  assign new_new_n23154__ = ~new_new_n23136__ & ~new_new_n23140__;
  assign new_new_n23155__ = ~new_new_n23141__ & ~new_new_n23154__;
  assign new_new_n23156__ = new_new_n23153__ & new_new_n23155__;
  assign new_new_n23157__ = ~new_new_n23141__ & ~new_new_n23156__;
  assign new_new_n23158__ = ~new_new_n21895__ & ~new_new_n21896__;
  assign new_new_n23159__ = ~new_new_n22425__ & new_new_n23158__;
  assign new_new_n23160__ = new_new_n22425__ & ~new_new_n23158__;
  assign new_new_n23161__ = ~new_new_n23159__ & ~new_new_n23160__;
  assign new_new_n23162__ = ~new_new_n23157__ & ~new_new_n23161__;
  assign new_new_n23163__ = new_new_n23157__ & new_new_n23161__;
  assign new_new_n23164__ = new_new_n10698__ & ~new_new_n15998__;
  assign new_new_n23165__ = new_new_n10702__ & new_new_n15905__;
  assign new_new_n23166__ = ~new_new_n11409__ & new_new_n15237__;
  assign new_new_n23167__ = new_new_n11378__ & new_new_n16025__;
  assign new_new_n23168__ = ~new_new_n23165__ & ~new_new_n23166__;
  assign new_new_n23169__ = ~new_new_n23164__ & new_new_n23168__;
  assign new_new_n23170__ = ~new_new_n23167__ & new_new_n23169__;
  assign new_new_n23171__ = pi08 & ~new_new_n23170__;
  assign new_new_n23172__ = ~pi08 & new_new_n23170__;
  assign new_new_n23173__ = ~new_new_n23171__ & ~new_new_n23172__;
  assign new_new_n23174__ = ~new_new_n23163__ & ~new_new_n23173__;
  assign new_new_n23175__ = ~new_new_n23162__ & ~new_new_n23174__;
  assign new_new_n23176__ = new_new_n22457__ & ~new_new_n23175__;
  assign new_new_n23177__ = ~new_new_n22457__ & new_new_n23175__;
  assign new_new_n23178__ = ~pi05 & ~new_new_n12830__;
  assign new_new_n23179__ = ~new_new_n12828__ & ~new_new_n23178__;
  assign new_new_n23180__ = ~new_new_n23177__ & new_new_n23179__;
  assign new_new_n23181__ = ~new_new_n23176__ & ~new_new_n23180__;
  assign new_new_n23182__ = new_new_n11378__ & ~new_new_n15917__;
  assign new_new_n23183__ = ~new_new_n11409__ & new_new_n15244__;
  assign new_new_n23184__ = new_new_n10702__ & new_new_n15237__;
  assign new_new_n23185__ = ~new_new_n23183__ & ~new_new_n23184__;
  assign new_new_n23186__ = ~new_new_n23182__ & new_new_n23185__;
  assign new_new_n23187__ = new_new_n10694__ & new_new_n15905__;
  assign new_new_n23188__ = pi08 & ~new_new_n23187__;
  assign new_new_n23189__ = new_new_n12121__ & new_new_n15905__;
  assign new_new_n23190__ = ~new_new_n23188__ & ~new_new_n23189__;
  assign new_new_n23191__ = new_new_n23186__ & ~new_new_n23190__;
  assign new_new_n23192__ = ~pi08 & ~new_new_n23186__;
  assign new_new_n23193__ = ~new_new_n23191__ & ~new_new_n23192__;
  assign new_new_n23194__ = new_new_n8474__ & new_new_n15285__;
  assign new_new_n23195__ = ~new_new_n8479__ & ~new_new_n15273__;
  assign new_new_n23196__ = new_new_n8858__ & ~new_new_n15314__;
  assign new_new_n23197__ = ~new_new_n23194__ & ~new_new_n23195__;
  assign new_new_n23198__ = ~new_new_n23196__ & new_new_n23197__;
  assign new_new_n23199__ = new_new_n8469__ & new_new_n17140__;
  assign new_new_n23200__ = pi11 & ~new_new_n23199__;
  assign new_new_n23201__ = new_new_n11530__ & new_new_n17140__;
  assign new_new_n23202__ = ~new_new_n23200__ & ~new_new_n23201__;
  assign new_new_n23203__ = new_new_n23198__ & ~new_new_n23202__;
  assign new_new_n23204__ = ~pi11 & ~new_new_n23198__;
  assign new_new_n23205__ = ~new_new_n23203__ & ~new_new_n23204__;
  assign new_new_n23206__ = ~new_new_n23123__ & ~new_new_n23124__;
  assign new_new_n23207__ = ~new_new_n23128__ & new_new_n23206__;
  assign new_new_n23208__ = new_new_n23128__ & ~new_new_n23206__;
  assign new_new_n23209__ = ~new_new_n23207__ & ~new_new_n23208__;
  assign new_new_n23210__ = ~new_new_n23102__ & ~new_new_n23103__;
  assign new_new_n23211__ = new_new_n23120__ & new_new_n23210__;
  assign new_new_n23212__ = ~new_new_n23120__ & ~new_new_n23210__;
  assign new_new_n23213__ = ~new_new_n23211__ & ~new_new_n23212__;
  assign new_new_n23214__ = ~new_new_n22507__ & ~new_new_n23094__;
  assign new_new_n23215__ = ~new_new_n23095__ & ~new_new_n23214__;
  assign new_new_n23216__ = new_new_n8858__ & ~new_new_n15321__;
  assign new_new_n23217__ = ~new_new_n8479__ & ~new_new_n15398__;
  assign new_new_n23218__ = new_new_n8474__ & ~new_new_n15349__;
  assign new_new_n23219__ = ~new_new_n23217__ & ~new_new_n23218__;
  assign new_new_n23220__ = ~new_new_n23216__ & new_new_n23219__;
  assign new_new_n23221__ = new_new_n8469__ & new_new_n16458__;
  assign new_new_n23222__ = ~pi11 & ~new_new_n23221__;
  assign new_new_n23223__ = new_new_n11368__ & new_new_n16458__;
  assign new_new_n23224__ = ~new_new_n23222__ & ~new_new_n23223__;
  assign new_new_n23225__ = new_new_n23220__ & ~new_new_n23224__;
  assign new_new_n23226__ = pi11 & ~new_new_n23220__;
  assign new_new_n23227__ = ~new_new_n23225__ & ~new_new_n23226__;
  assign new_new_n23228__ = new_new_n23215__ & ~new_new_n23227__;
  assign new_new_n23229__ = ~new_new_n23215__ & new_new_n23227__;
  assign new_new_n23230__ = ~new_new_n22530__ & ~new_new_n22531__;
  assign new_new_n23231__ = new_new_n23086__ & new_new_n23230__;
  assign new_new_n23232__ = ~new_new_n23086__ & ~new_new_n23230__;
  assign new_new_n23233__ = ~new_new_n23231__ & ~new_new_n23232__;
  assign new_new_n23234__ = new_new_n8474__ & new_new_n15390__;
  assign new_new_n23235__ = ~new_new_n8479__ & ~new_new_n15362__;
  assign new_new_n23236__ = ~new_new_n23234__ & ~new_new_n23235__;
  assign new_new_n23237__ = new_new_n8469__ & ~new_new_n17364__;
  assign new_new_n23238__ = pi11 & ~new_new_n23237__;
  assign new_new_n23239__ = ~pi10 & new_new_n15398__;
  assign new_new_n23240__ = pi10 & ~new_new_n15398__;
  assign new_new_n23241__ = new_new_n8469__ & ~new_new_n23239__;
  assign new_new_n23242__ = ~new_new_n23240__ & new_new_n23241__;
  assign new_new_n23243__ = new_new_n16956__ & new_new_n23242__;
  assign new_new_n23244__ = ~new_new_n23238__ & ~new_new_n23243__;
  assign new_new_n23245__ = new_new_n23236__ & ~new_new_n23244__;
  assign new_new_n23246__ = new_new_n8469__ & new_new_n17360__;
  assign new_new_n23247__ = new_new_n23236__ & ~new_new_n23246__;
  assign new_new_n23248__ = ~pi11 & ~new_new_n23247__;
  assign new_new_n23249__ = ~new_new_n23245__ & ~new_new_n23248__;
  assign new_new_n23250__ = ~new_new_n8479__ & ~new_new_n15432__;
  assign new_new_n23251__ = new_new_n8474__ & ~new_new_n15362__;
  assign new_new_n23252__ = ~new_new_n23250__ & ~new_new_n23251__;
  assign new_new_n23253__ = new_new_n8469__ & new_new_n17914__;
  assign new_new_n23254__ = new_new_n23252__ & ~new_new_n23253__;
  assign new_new_n23255__ = pi11 & ~new_new_n23254__;
  assign new_new_n23256__ = new_new_n8469__ & ~new_new_n17918__;
  assign new_new_n23257__ = ~pi11 & ~new_new_n23256__;
  assign new_new_n23258__ = ~pi10 & new_new_n15390__;
  assign new_new_n23259__ = pi10 & ~new_new_n15390__;
  assign new_new_n23260__ = new_new_n8469__ & new_new_n15829__;
  assign new_new_n23261__ = ~new_new_n23258__ & ~new_new_n23259__;
  assign new_new_n23262__ = new_new_n23260__ & new_new_n23261__;
  assign new_new_n23263__ = ~new_new_n23257__ & ~new_new_n23262__;
  assign new_new_n23264__ = new_new_n23252__ & ~new_new_n23263__;
  assign new_new_n23265__ = ~new_new_n23255__ & ~new_new_n23264__;
  assign new_new_n23266__ = ~new_new_n22565__ & ~new_new_n22566__;
  assign new_new_n23267__ = new_new_n23063__ & new_new_n23266__;
  assign new_new_n23268__ = ~new_new_n23063__ & ~new_new_n23266__;
  assign new_new_n23269__ = ~new_new_n23267__ & ~new_new_n23268__;
  assign new_new_n23270__ = new_new_n23265__ & ~new_new_n23269__;
  assign new_new_n23271__ = ~new_new_n23265__ & new_new_n23269__;
  assign new_new_n23272__ = new_new_n8474__ & ~new_new_n15432__;
  assign new_new_n23273__ = ~new_new_n8479__ & ~new_new_n15439__;
  assign new_new_n23274__ = new_new_n8470__ & new_new_n16771__;
  assign new_new_n23275__ = ~new_new_n23272__ & ~new_new_n23273__;
  assign new_new_n23276__ = ~new_new_n23274__ & new_new_n23275__;
  assign new_new_n23277__ = new_new_n8469__ & ~new_new_n15362__;
  assign new_new_n23278__ = pi11 & ~new_new_n23277__;
  assign new_new_n23279__ = new_new_n11368__ & ~new_new_n15362__;
  assign new_new_n23280__ = ~new_new_n23278__ & ~new_new_n23279__;
  assign new_new_n23281__ = new_new_n23276__ & ~new_new_n23280__;
  assign new_new_n23282__ = ~pi11 & ~new_new_n23276__;
  assign new_new_n23283__ = ~new_new_n23281__ & ~new_new_n23282__;
  assign new_new_n23284__ = new_new_n8474__ & ~new_new_n15439__;
  assign new_new_n23285__ = ~new_new_n8479__ & new_new_n15464__;
  assign new_new_n23286__ = new_new_n8858__ & ~new_new_n15432__;
  assign new_new_n23287__ = ~new_new_n23284__ & ~new_new_n23285__;
  assign new_new_n23288__ = ~new_new_n23286__ & new_new_n23287__;
  assign new_new_n23289__ = new_new_n8469__ & new_new_n17204__;
  assign new_new_n23290__ = ~pi11 & ~new_new_n23289__;
  assign new_new_n23291__ = new_new_n11368__ & new_new_n17204__;
  assign new_new_n23292__ = ~new_new_n23290__ & ~new_new_n23291__;
  assign new_new_n23293__ = new_new_n23288__ & ~new_new_n23292__;
  assign new_new_n23294__ = pi11 & ~new_new_n23288__;
  assign new_new_n23295__ = ~new_new_n23293__ & ~new_new_n23294__;
  assign new_new_n23296__ = ~new_new_n23029__ & ~new_new_n23030__;
  assign new_new_n23297__ = ~new_new_n23034__ & new_new_n23296__;
  assign new_new_n23298__ = new_new_n23034__ & ~new_new_n23296__;
  assign new_new_n23299__ = ~new_new_n23297__ & ~new_new_n23298__;
  assign new_new_n23300__ = new_new_n8474__ & ~new_new_n15471__;
  assign new_new_n23301__ = ~new_new_n8479__ & ~new_new_n15809__;
  assign new_new_n23302__ = new_new_n8858__ & new_new_n15464__;
  assign new_new_n23303__ = ~new_new_n23300__ & ~new_new_n23301__;
  assign new_new_n23304__ = ~new_new_n23302__ & new_new_n23303__;
  assign new_new_n23305__ = new_new_n8469__ & new_new_n15819__;
  assign new_new_n23306__ = ~pi11 & ~new_new_n23305__;
  assign new_new_n23307__ = new_new_n11368__ & new_new_n15819__;
  assign new_new_n23308__ = ~new_new_n23306__ & ~new_new_n23307__;
  assign new_new_n23309__ = new_new_n23304__ & ~new_new_n23308__;
  assign new_new_n23310__ = pi11 & ~new_new_n23304__;
  assign new_new_n23311__ = ~new_new_n23309__ & ~new_new_n23310__;
  assign new_new_n23312__ = ~new_new_n23023__ & ~new_new_n23024__;
  assign new_new_n23313__ = ~new_new_n23026__ & new_new_n23312__;
  assign new_new_n23314__ = new_new_n23026__ & ~new_new_n23312__;
  assign new_new_n23315__ = ~new_new_n23313__ & ~new_new_n23314__;
  assign new_new_n23316__ = new_new_n23311__ & ~new_new_n23315__;
  assign new_new_n23317__ = ~new_new_n23311__ & new_new_n23315__;
  assign new_new_n23318__ = ~new_new_n22998__ & ~new_new_n22999__;
  assign new_new_n23319__ = ~new_new_n23003__ & new_new_n23318__;
  assign new_new_n23320__ = new_new_n23003__ & ~new_new_n23318__;
  assign new_new_n23321__ = ~new_new_n23319__ & ~new_new_n23320__;
  assign new_new_n23322__ = new_new_n8858__ & ~new_new_n15487__;
  assign new_new_n23323__ = new_new_n8474__ & new_new_n15524__;
  assign new_new_n23324__ = ~new_new_n8479__ & new_new_n15520__;
  assign new_new_n23325__ = ~new_new_n23323__ & ~new_new_n23324__;
  assign new_new_n23326__ = ~new_new_n23322__ & new_new_n23325__;
  assign new_new_n23327__ = new_new_n8469__ & new_new_n17587__;
  assign new_new_n23328__ = pi11 & ~new_new_n23327__;
  assign new_new_n23329__ = new_new_n11530__ & new_new_n17587__;
  assign new_new_n23330__ = ~new_new_n23328__ & ~new_new_n23329__;
  assign new_new_n23331__ = new_new_n23326__ & ~new_new_n23330__;
  assign new_new_n23332__ = ~pi11 & ~new_new_n23326__;
  assign new_new_n23333__ = ~new_new_n23331__ & ~new_new_n23332__;
  assign new_new_n23334__ = ~new_new_n22982__ & ~new_new_n22983__;
  assign new_new_n23335__ = ~new_new_n22987__ & new_new_n23334__;
  assign new_new_n23336__ = new_new_n22987__ & ~new_new_n23334__;
  assign new_new_n23337__ = ~new_new_n23335__ & ~new_new_n23336__;
  assign new_new_n23338__ = ~new_new_n23333__ & ~new_new_n23337__;
  assign new_new_n23339__ = new_new_n23333__ & new_new_n23337__;
  assign new_new_n23340__ = ~new_new_n22674__ & ~new_new_n22675__;
  assign new_new_n23341__ = ~new_new_n22979__ & new_new_n23340__;
  assign new_new_n23342__ = new_new_n22979__ & ~new_new_n23340__;
  assign new_new_n23343__ = ~new_new_n23341__ & ~new_new_n23342__;
  assign new_new_n23344__ = new_new_n8474__ & ~new_new_n15533__;
  assign new_new_n23345__ = ~new_new_n8479__ & new_new_n15767__;
  assign new_new_n23346__ = new_new_n8858__ & new_new_n15520__;
  assign new_new_n23347__ = ~new_new_n23344__ & ~new_new_n23345__;
  assign new_new_n23348__ = ~new_new_n23346__ & new_new_n23347__;
  assign new_new_n23349__ = new_new_n8469__ & new_new_n19731__;
  assign new_new_n23350__ = ~pi11 & ~new_new_n23349__;
  assign new_new_n23351__ = new_new_n11368__ & new_new_n19731__;
  assign new_new_n23352__ = ~new_new_n23350__ & ~new_new_n23351__;
  assign new_new_n23353__ = new_new_n23348__ & ~new_new_n23352__;
  assign new_new_n23354__ = pi11 & ~new_new_n23348__;
  assign new_new_n23355__ = ~new_new_n23353__ & ~new_new_n23354__;
  assign new_new_n23356__ = new_new_n8858__ & ~new_new_n15533__;
  assign new_new_n23357__ = ~new_new_n8479__ & new_new_n15560__;
  assign new_new_n23358__ = new_new_n8474__ & new_new_n15767__;
  assign new_new_n23359__ = new_new_n8470__ & new_new_n19893__;
  assign new_new_n23360__ = ~new_new_n23357__ & ~new_new_n23358__;
  assign new_new_n23361__ = ~new_new_n23356__ & new_new_n23360__;
  assign new_new_n23362__ = ~new_new_n23359__ & new_new_n23361__;
  assign new_new_n23363__ = pi11 & ~new_new_n23362__;
  assign new_new_n23364__ = ~pi11 & new_new_n23362__;
  assign new_new_n23365__ = ~new_new_n23363__ & ~new_new_n23364__;
  assign new_new_n23366__ = new_new_n8474__ & new_new_n15564__;
  assign new_new_n23367__ = ~new_new_n8479__ & ~new_new_n15615__;
  assign new_new_n23368__ = new_new_n8858__ & new_new_n15572__;
  assign new_new_n23369__ = ~new_new_n23366__ & ~new_new_n23367__;
  assign new_new_n23370__ = ~new_new_n23368__ & new_new_n23369__;
  assign new_new_n23371__ = new_new_n8469__ & ~new_new_n20114__;
  assign new_new_n23372__ = ~pi11 & ~new_new_n23371__;
  assign new_new_n23373__ = new_new_n11368__ & ~new_new_n20114__;
  assign new_new_n23374__ = ~new_new_n23372__ & ~new_new_n23373__;
  assign new_new_n23375__ = new_new_n23370__ & ~new_new_n23374__;
  assign new_new_n23376__ = pi11 & ~new_new_n23370__;
  assign new_new_n23377__ = ~new_new_n23375__ & ~new_new_n23376__;
  assign new_new_n23378__ = ~new_new_n22713__ & ~new_new_n22714__;
  assign new_new_n23379__ = new_new_n22895__ & ~new_new_n23378__;
  assign new_new_n23380__ = ~new_new_n22895__ & new_new_n23378__;
  assign new_new_n23381__ = ~new_new_n23379__ & ~new_new_n23380__;
  assign new_new_n23382__ = ~new_new_n23377__ & new_new_n23381__;
  assign new_new_n23383__ = new_new_n23377__ & ~new_new_n23381__;
  assign new_new_n23384__ = new_new_n8474__ & ~new_new_n15615__;
  assign new_new_n23385__ = ~new_new_n8479__ & new_new_n15743__;
  assign new_new_n23386__ = new_new_n8470__ & new_new_n18512__;
  assign new_new_n23387__ = ~new_new_n23384__ & ~new_new_n23385__;
  assign new_new_n23388__ = ~new_new_n23386__ & new_new_n23387__;
  assign new_new_n23389__ = new_new_n8469__ & new_new_n15564__;
  assign new_new_n23390__ = pi11 & ~new_new_n23389__;
  assign new_new_n23391__ = new_new_n11368__ & new_new_n15564__;
  assign new_new_n23392__ = ~new_new_n23390__ & ~new_new_n23391__;
  assign new_new_n23393__ = new_new_n23388__ & ~new_new_n23392__;
  assign new_new_n23394__ = ~pi11 & ~new_new_n23388__;
  assign new_new_n23395__ = ~new_new_n23393__ & ~new_new_n23394__;
  assign new_new_n23396__ = ~new_new_n22742__ & ~new_new_n22743__;
  assign new_new_n23397__ = ~new_new_n22873__ & new_new_n23396__;
  assign new_new_n23398__ = new_new_n22873__ & ~new_new_n23396__;
  assign new_new_n23399__ = ~new_new_n23397__ & ~new_new_n23398__;
  assign new_new_n23400__ = new_new_n8474__ & ~new_new_n15638__;
  assign new_new_n23401__ = ~new_new_n8479__ & ~new_new_n15582__;
  assign new_new_n23402__ = new_new_n8470__ & new_new_n19494__;
  assign new_new_n23403__ = ~new_new_n23400__ & ~new_new_n23401__;
  assign new_new_n23404__ = ~new_new_n23402__ & new_new_n23403__;
  assign new_new_n23405__ = new_new_n8469__ & new_new_n15743__;
  assign new_new_n23406__ = pi11 & ~new_new_n23405__;
  assign new_new_n23407__ = new_new_n11368__ & new_new_n15743__;
  assign new_new_n23408__ = ~new_new_n23406__ & ~new_new_n23407__;
  assign new_new_n23409__ = new_new_n23404__ & ~new_new_n23408__;
  assign new_new_n23410__ = ~pi11 & ~new_new_n23404__;
  assign new_new_n23411__ = ~new_new_n23409__ & ~new_new_n23410__;
  assign new_new_n23412__ = ~new_new_n22866__ & ~new_new_n22867__;
  assign new_new_n23413__ = new_new_n22871__ & ~new_new_n23412__;
  assign new_new_n23414__ = ~new_new_n22871__ & new_new_n23412__;
  assign new_new_n23415__ = ~new_new_n23413__ & ~new_new_n23414__;
  assign new_new_n23416__ = ~new_new_n23411__ & new_new_n23415__;
  assign new_new_n23417__ = new_new_n23411__ & ~new_new_n23415__;
  assign new_new_n23418__ = new_new_n8474__ & ~new_new_n15582__;
  assign new_new_n23419__ = ~new_new_n8479__ & ~new_new_n15647__;
  assign new_new_n23420__ = new_new_n8470__ & new_new_n19487__;
  assign new_new_n23421__ = ~new_new_n23418__ & ~new_new_n23419__;
  assign new_new_n23422__ = ~new_new_n23420__ & new_new_n23421__;
  assign new_new_n23423__ = new_new_n8469__ & ~new_new_n15638__;
  assign new_new_n23424__ = pi11 & ~new_new_n23423__;
  assign new_new_n23425__ = new_new_n11368__ & ~new_new_n15638__;
  assign new_new_n23426__ = ~new_new_n23424__ & ~new_new_n23425__;
  assign new_new_n23427__ = new_new_n23422__ & ~new_new_n23426__;
  assign new_new_n23428__ = ~pi11 & ~new_new_n23422__;
  assign new_new_n23429__ = ~new_new_n23427__ & ~new_new_n23428__;
  assign new_new_n23430__ = ~new_new_n22851__ & ~new_new_n22862__;
  assign new_new_n23431__ = new_new_n22859__ & ~new_new_n23430__;
  assign new_new_n23432__ = ~new_new_n22859__ & new_new_n23430__;
  assign new_new_n23433__ = ~new_new_n23431__ & ~new_new_n23432__;
  assign new_new_n23434__ = ~new_new_n22809__ & new_new_n22832__;
  assign new_new_n23435__ = ~new_new_n22833__ & ~new_new_n23434__;
  assign new_new_n23436__ = new_new_n22830__ & new_new_n22831__;
  assign new_new_n23437__ = ~new_new_n23435__ & ~new_new_n23436__;
  assign new_new_n23438__ = ~new_new_n8479__ & new_new_n15643__;
  assign new_new_n23439__ = new_new_n8474__ & new_new_n15656__;
  assign new_new_n23440__ = ~new_new_n23438__ & ~new_new_n23439__;
  assign new_new_n23441__ = new_new_n8469__ & new_new_n22764__;
  assign new_new_n23442__ = new_new_n23440__ & ~new_new_n23441__;
  assign new_new_n23443__ = pi11 & ~new_new_n23442__;
  assign new_new_n23444__ = new_new_n8469__ & ~new_new_n22774__;
  assign new_new_n23445__ = ~pi11 & ~new_new_n23444__;
  assign new_new_n23446__ = ~pi10 & ~new_new_n22768__;
  assign new_new_n23447__ = pi10 & ~new_new_n22770__;
  assign new_new_n23448__ = new_new_n8469__ & ~new_new_n23446__;
  assign new_new_n23449__ = ~new_new_n23447__ & new_new_n23448__;
  assign new_new_n23450__ = ~new_new_n23445__ & ~new_new_n23449__;
  assign new_new_n23451__ = new_new_n23440__ & ~new_new_n23450__;
  assign new_new_n23452__ = ~new_new_n23443__ & ~new_new_n23451__;
  assign new_new_n23453__ = new_new_n8474__ & ~new_new_n15661__;
  assign new_new_n23454__ = ~new_new_n8479__ & new_new_n15668__;
  assign new_new_n23455__ = ~new_new_n23453__ & ~new_new_n23454__;
  assign new_new_n23456__ = new_new_n8469__ & ~new_new_n20177__;
  assign new_new_n23457__ = pi11 & ~new_new_n23456__;
  assign new_new_n23458__ = pi10 & ~new_new_n15643__;
  assign new_new_n23459__ = ~pi10 & new_new_n15643__;
  assign new_new_n23460__ = ~new_new_n23458__ & ~new_new_n23459__;
  assign new_new_n23461__ = new_new_n8469__ & new_new_n20176__;
  assign new_new_n23462__ = ~new_new_n23460__ & new_new_n23461__;
  assign new_new_n23463__ = ~new_new_n23457__ & ~new_new_n23462__;
  assign new_new_n23464__ = new_new_n23455__ & ~new_new_n23463__;
  assign new_new_n23465__ = new_new_n8469__ & new_new_n20187__;
  assign new_new_n23466__ = new_new_n23455__ & ~new_new_n23465__;
  assign new_new_n23467__ = ~pi11 & ~new_new_n23466__;
  assign new_new_n23468__ = ~new_new_n23464__ & ~new_new_n23467__;
  assign new_new_n23469__ = new_new_n6994__ & ~new_new_n15673__;
  assign new_new_n23470__ = ~new_new_n8469__ & ~new_new_n8474__;
  assign new_new_n23471__ = ~new_new_n20628__ & ~new_new_n23470__;
  assign new_new_n23472__ = new_new_n8469__ & ~new_new_n15661__;
  assign new_new_n23473__ = new_new_n8479__ & ~new_new_n23472__;
  assign new_new_n23474__ = ~new_new_n15673__ & ~new_new_n23473__;
  assign new_new_n23475__ = ~new_new_n8468__ & new_new_n15668__;
  assign new_new_n23476__ = ~new_new_n15679__ & new_new_n23475__;
  assign new_new_n23477__ = new_new_n15661__ & ~new_new_n23475__;
  assign new_new_n23478__ = new_new_n8469__ & ~new_new_n23477__;
  assign new_new_n23479__ = ~new_new_n23476__ & new_new_n23478__;
  assign new_new_n23480__ = ~new_new_n23474__ & ~new_new_n23479__;
  assign new_new_n23481__ = pi11 & ~new_new_n23471__;
  assign new_new_n23482__ = new_new_n23480__ & new_new_n23481__;
  assign new_new_n23483__ = ~new_new_n23469__ & ~new_new_n23482__;
  assign new_new_n23484__ = ~new_new_n23468__ & ~new_new_n23483__;
  assign new_new_n23485__ = pi11 & new_new_n19823__;
  assign new_new_n23486__ = new_new_n6982__ & new_new_n15674__;
  assign new_new_n23487__ = ~new_new_n6994__ & new_new_n20195__;
  assign new_new_n23488__ = ~new_new_n6981__ & new_new_n15668__;
  assign new_new_n23489__ = new_new_n6984__ & ~new_new_n23488__;
  assign new_new_n23490__ = ~new_new_n20628__ & ~new_new_n23485__;
  assign new_new_n23491__ = ~new_new_n23486__ & new_new_n23490__;
  assign new_new_n23492__ = ~new_new_n23487__ & ~new_new_n23489__;
  assign new_new_n23493__ = new_new_n23491__ & new_new_n23492__;
  assign new_new_n23494__ = ~new_new_n23484__ & ~new_new_n23493__;
  assign new_new_n23495__ = new_new_n23484__ & new_new_n23493__;
  assign new_new_n23496__ = new_new_n8858__ & new_new_n15656__;
  assign new_new_n23497__ = ~new_new_n8479__ & ~new_new_n15661__;
  assign new_new_n23498__ = new_new_n8474__ & new_new_n15643__;
  assign new_new_n23499__ = new_new_n8470__ & new_new_n15687__;
  assign new_new_n23500__ = ~new_new_n23497__ & ~new_new_n23498__;
  assign new_new_n23501__ = ~new_new_n23496__ & new_new_n23500__;
  assign new_new_n23502__ = ~new_new_n23499__ & new_new_n23501__;
  assign new_new_n23503__ = pi11 & ~new_new_n23502__;
  assign new_new_n23504__ = ~pi11 & new_new_n23502__;
  assign new_new_n23505__ = ~new_new_n23503__ & ~new_new_n23504__;
  assign new_new_n23506__ = ~new_new_n23495__ & ~new_new_n23505__;
  assign new_new_n23507__ = ~new_new_n23494__ & ~new_new_n23506__;
  assign new_new_n23508__ = ~new_new_n23452__ & ~new_new_n23507__;
  assign new_new_n23509__ = new_new_n23452__ & new_new_n23507__;
  assign new_new_n23510__ = new_new_n22825__ & ~new_new_n22829__;
  assign new_new_n23511__ = new_new_n10998__ & ~new_new_n20628__;
  assign new_new_n23512__ = pi14 & ~new_new_n23511__;
  assign new_new_n23513__ = ~new_new_n22825__ & new_new_n23512__;
  assign new_new_n23514__ = ~new_new_n23510__ & ~new_new_n23513__;
  assign new_new_n23515__ = ~new_new_n23509__ & ~new_new_n23514__;
  assign new_new_n23516__ = ~new_new_n23508__ & ~new_new_n23515__;
  assign new_new_n23517__ = new_new_n23437__ & ~new_new_n23516__;
  assign new_new_n23518__ = ~new_new_n23437__ & new_new_n23516__;
  assign new_new_n23519__ = new_new_n8474__ & ~new_new_n15710__;
  assign new_new_n23520__ = ~new_new_n8479__ & new_new_n15656__;
  assign new_new_n23521__ = new_new_n8858__ & ~new_new_n15647__;
  assign new_new_n23522__ = new_new_n8470__ & ~new_new_n19118__;
  assign new_new_n23523__ = ~new_new_n23519__ & ~new_new_n23520__;
  assign new_new_n23524__ = ~new_new_n23521__ & new_new_n23523__;
  assign new_new_n23525__ = ~new_new_n23522__ & new_new_n23524__;
  assign new_new_n23526__ = pi11 & ~new_new_n23525__;
  assign new_new_n23527__ = ~pi11 & new_new_n23525__;
  assign new_new_n23528__ = ~new_new_n23526__ & ~new_new_n23527__;
  assign new_new_n23529__ = ~new_new_n23518__ & ~new_new_n23528__;
  assign new_new_n23530__ = ~new_new_n23517__ & ~new_new_n23529__;
  assign new_new_n23531__ = ~new_new_n23433__ & new_new_n23530__;
  assign new_new_n23532__ = new_new_n23433__ & ~new_new_n23530__;
  assign new_new_n23533__ = new_new_n8858__ & ~new_new_n15582__;
  assign new_new_n23534__ = ~new_new_n8479__ & ~new_new_n15710__;
  assign new_new_n23535__ = new_new_n8474__ & ~new_new_n15647__;
  assign new_new_n23536__ = new_new_n8470__ & ~new_new_n15736__;
  assign new_new_n23537__ = ~new_new_n23534__ & ~new_new_n23535__;
  assign new_new_n23538__ = ~new_new_n23533__ & new_new_n23537__;
  assign new_new_n23539__ = ~new_new_n23536__ & new_new_n23538__;
  assign new_new_n23540__ = ~pi11 & ~new_new_n23539__;
  assign new_new_n23541__ = pi11 & new_new_n23539__;
  assign new_new_n23542__ = ~new_new_n23540__ & ~new_new_n23541__;
  assign new_new_n23543__ = ~new_new_n23532__ & ~new_new_n23542__;
  assign new_new_n23544__ = ~new_new_n23531__ & ~new_new_n23543__;
  assign new_new_n23545__ = ~new_new_n23429__ & ~new_new_n23544__;
  assign new_new_n23546__ = new_new_n23429__ & new_new_n23544__;
  assign new_new_n23547__ = ~new_new_n22794__ & new_new_n22864__;
  assign new_new_n23548__ = ~new_new_n22833__ & new_new_n22861__;
  assign new_new_n23549__ = new_new_n22794__ & ~new_new_n22859__;
  assign new_new_n23550__ = ~new_new_n23548__ & ~new_new_n23549__;
  assign new_new_n23551__ = ~new_new_n22850__ & ~new_new_n23550__;
  assign new_new_n23552__ = new_new_n22794__ & ~new_new_n22833__;
  assign new_new_n23553__ = ~new_new_n22859__ & new_new_n22861__;
  assign new_new_n23554__ = ~new_new_n23552__ & ~new_new_n23553__;
  assign new_new_n23555__ = ~new_new_n23433__ & ~new_new_n23554__;
  assign new_new_n23556__ = ~new_new_n23547__ & ~new_new_n23551__;
  assign new_new_n23557__ = ~new_new_n23555__ & new_new_n23556__;
  assign new_new_n23558__ = ~new_new_n23546__ & new_new_n23557__;
  assign new_new_n23559__ = ~new_new_n23545__ & ~new_new_n23558__;
  assign new_new_n23560__ = ~new_new_n23417__ & ~new_new_n23559__;
  assign new_new_n23561__ = ~new_new_n23416__ & ~new_new_n23560__;
  assign new_new_n23562__ = ~new_new_n23399__ & new_new_n23561__;
  assign new_new_n23563__ = new_new_n23399__ & ~new_new_n23561__;
  assign new_new_n23564__ = new_new_n8858__ & ~new_new_n15615__;
  assign new_new_n23565__ = ~new_new_n8479__ & ~new_new_n15638__;
  assign new_new_n23566__ = new_new_n8474__ & new_new_n15743__;
  assign new_new_n23567__ = new_new_n8470__ & new_new_n19005__;
  assign new_new_n23568__ = ~new_new_n23565__ & ~new_new_n23566__;
  assign new_new_n23569__ = ~new_new_n23564__ & new_new_n23568__;
  assign new_new_n23570__ = ~new_new_n23567__ & new_new_n23569__;
  assign new_new_n23571__ = pi11 & ~new_new_n23570__;
  assign new_new_n23572__ = ~pi11 & new_new_n23570__;
  assign new_new_n23573__ = ~new_new_n23571__ & ~new_new_n23572__;
  assign new_new_n23574__ = ~new_new_n23563__ & ~new_new_n23573__;
  assign new_new_n23575__ = ~new_new_n23562__ & ~new_new_n23574__;
  assign new_new_n23576__ = new_new_n23395__ & ~new_new_n23575__;
  assign new_new_n23577__ = ~new_new_n23395__ & new_new_n23575__;
  assign new_new_n23578__ = ~new_new_n22876__ & ~new_new_n22877__;
  assign new_new_n23579__ = ~new_new_n22893__ & new_new_n23578__;
  assign new_new_n23580__ = new_new_n22893__ & ~new_new_n23578__;
  assign new_new_n23581__ = ~new_new_n23579__ & ~new_new_n23580__;
  assign new_new_n23582__ = ~new_new_n23577__ & new_new_n23581__;
  assign new_new_n23583__ = ~new_new_n23576__ & ~new_new_n23582__;
  assign new_new_n23584__ = ~new_new_n23383__ & ~new_new_n23583__;
  assign new_new_n23585__ = ~new_new_n23382__ & ~new_new_n23584__;
  assign new_new_n23586__ = ~new_new_n22898__ & ~new_new_n22899__;
  assign new_new_n23587__ = new_new_n22903__ & new_new_n23586__;
  assign new_new_n23588__ = ~new_new_n22903__ & ~new_new_n23586__;
  assign new_new_n23589__ = ~new_new_n23587__ & ~new_new_n23588__;
  assign new_new_n23590__ = ~new_new_n23585__ & ~new_new_n23589__;
  assign new_new_n23591__ = new_new_n23585__ & new_new_n23589__;
  assign new_new_n23592__ = new_new_n8474__ & new_new_n15572__;
  assign new_new_n23593__ = ~new_new_n8479__ & new_new_n15564__;
  assign new_new_n23594__ = new_new_n8470__ & new_new_n18944__;
  assign new_new_n23595__ = ~new_new_n23592__ & ~new_new_n23593__;
  assign new_new_n23596__ = ~new_new_n23594__ & new_new_n23595__;
  assign new_new_n23597__ = new_new_n8469__ & new_new_n15560__;
  assign new_new_n23598__ = pi11 & ~new_new_n23597__;
  assign new_new_n23599__ = new_new_n11368__ & new_new_n15560__;
  assign new_new_n23600__ = ~new_new_n23598__ & ~new_new_n23599__;
  assign new_new_n23601__ = new_new_n23596__ & ~new_new_n23600__;
  assign new_new_n23602__ = ~pi11 & ~new_new_n23596__;
  assign new_new_n23603__ = ~new_new_n23601__ & ~new_new_n23602__;
  assign new_new_n23604__ = ~new_new_n23591__ & new_new_n23603__;
  assign new_new_n23605__ = ~new_new_n23590__ & ~new_new_n23604__;
  assign new_new_n23606__ = ~new_new_n22905__ & ~new_new_n22928__;
  assign new_new_n23607__ = ~new_new_n22929__ & ~new_new_n23606__;
  assign new_new_n23608__ = new_new_n8474__ & new_new_n15560__;
  assign new_new_n23609__ = ~new_new_n8479__ & new_new_n15572__;
  assign new_new_n23610__ = new_new_n8470__ & ~new_new_n18454__;
  assign new_new_n23611__ = ~new_new_n23608__ & ~new_new_n23609__;
  assign new_new_n23612__ = ~new_new_n23610__ & new_new_n23611__;
  assign new_new_n23613__ = new_new_n8469__ & new_new_n15767__;
  assign new_new_n23614__ = pi11 & ~new_new_n23613__;
  assign new_new_n23615__ = new_new_n11368__ & new_new_n15767__;
  assign new_new_n23616__ = ~new_new_n23614__ & ~new_new_n23615__;
  assign new_new_n23617__ = new_new_n23612__ & ~new_new_n23616__;
  assign new_new_n23618__ = ~pi11 & ~new_new_n23612__;
  assign new_new_n23619__ = ~new_new_n23617__ & ~new_new_n23618__;
  assign new_new_n23620__ = new_new_n23607__ & new_new_n23619__;
  assign new_new_n23621__ = new_new_n23605__ & ~new_new_n23620__;
  assign new_new_n23622__ = ~new_new_n23607__ & ~new_new_n23619__;
  assign new_new_n23623__ = ~new_new_n23621__ & ~new_new_n23622__;
  assign new_new_n23624__ = ~new_new_n23365__ & new_new_n23623__;
  assign new_new_n23625__ = new_new_n23365__ & ~new_new_n23623__;
  assign new_new_n23626__ = ~new_new_n22936__ & ~new_new_n22937__;
  assign new_new_n23627__ = new_new_n22952__ & ~new_new_n23626__;
  assign new_new_n23628__ = ~new_new_n22952__ & new_new_n23626__;
  assign new_new_n23629__ = ~new_new_n23627__ & ~new_new_n23628__;
  assign new_new_n23630__ = ~new_new_n23625__ & ~new_new_n23629__;
  assign new_new_n23631__ = ~new_new_n23624__ & ~new_new_n23630__;
  assign new_new_n23632__ = new_new_n23355__ & new_new_n23631__;
  assign new_new_n23633__ = ~new_new_n23355__ & ~new_new_n23631__;
  assign new_new_n23634__ = ~new_new_n22959__ & ~new_new_n22960__;
  assign new_new_n23635__ = new_new_n22977__ & new_new_n23634__;
  assign new_new_n23636__ = ~new_new_n22977__ & ~new_new_n23634__;
  assign new_new_n23637__ = ~new_new_n23635__ & ~new_new_n23636__;
  assign new_new_n23638__ = ~new_new_n23633__ & ~new_new_n23637__;
  assign new_new_n23639__ = ~new_new_n23632__ & ~new_new_n23638__;
  assign new_new_n23640__ = ~new_new_n23343__ & ~new_new_n23639__;
  assign new_new_n23641__ = new_new_n23343__ & new_new_n23639__;
  assign new_new_n23642__ = new_new_n8474__ & new_new_n15520__;
  assign new_new_n23643__ = ~new_new_n8479__ & ~new_new_n15533__;
  assign new_new_n23644__ = ~new_new_n23642__ & ~new_new_n23643__;
  assign new_new_n23645__ = new_new_n8469__ & new_new_n18923__;
  assign new_new_n23646__ = new_new_n23644__ & ~new_new_n23645__;
  assign new_new_n23647__ = pi11 & ~new_new_n23646__;
  assign new_new_n23648__ = new_new_n8469__ & ~new_new_n18914__;
  assign new_new_n23649__ = ~pi11 & ~new_new_n23648__;
  assign new_new_n23650__ = ~pi10 & new_new_n15524__;
  assign new_new_n23651__ = pi10 & ~new_new_n15524__;
  assign new_new_n23652__ = new_new_n8469__ & ~new_new_n23650__;
  assign new_new_n23653__ = ~new_new_n23651__ & new_new_n23652__;
  assign new_new_n23654__ = new_new_n18913__ & new_new_n23653__;
  assign new_new_n23655__ = ~new_new_n23649__ & ~new_new_n23654__;
  assign new_new_n23656__ = new_new_n23644__ & ~new_new_n23655__;
  assign new_new_n23657__ = ~new_new_n23647__ & ~new_new_n23656__;
  assign new_new_n23658__ = ~new_new_n23641__ & new_new_n23657__;
  assign new_new_n23659__ = ~new_new_n23640__ & ~new_new_n23658__;
  assign new_new_n23660__ = ~new_new_n23339__ & ~new_new_n23659__;
  assign new_new_n23661__ = ~new_new_n23338__ & ~new_new_n23660__;
  assign new_new_n23662__ = ~new_new_n22990__ & ~new_new_n22991__;
  assign new_new_n23663__ = ~new_new_n22995__ & new_new_n23662__;
  assign new_new_n23664__ = new_new_n22995__ & ~new_new_n23662__;
  assign new_new_n23665__ = ~new_new_n23663__ & ~new_new_n23664__;
  assign new_new_n23666__ = new_new_n23661__ & ~new_new_n23665__;
  assign new_new_n23667__ = ~new_new_n23661__ & new_new_n23665__;
  assign new_new_n23668__ = new_new_n8858__ & ~new_new_n15809__;
  assign new_new_n23669__ = ~new_new_n8479__ & new_new_n15524__;
  assign new_new_n23670__ = new_new_n8474__ & ~new_new_n15487__;
  assign new_new_n23671__ = new_new_n8470__ & new_new_n18020__;
  assign new_new_n23672__ = ~new_new_n23669__ & ~new_new_n23670__;
  assign new_new_n23673__ = ~new_new_n23668__ & new_new_n23672__;
  assign new_new_n23674__ = ~new_new_n23671__ & new_new_n23673__;
  assign new_new_n23675__ = pi11 & ~new_new_n23674__;
  assign new_new_n23676__ = ~pi11 & new_new_n23674__;
  assign new_new_n23677__ = ~new_new_n23675__ & ~new_new_n23676__;
  assign new_new_n23678__ = ~new_new_n23667__ & ~new_new_n23677__;
  assign new_new_n23679__ = ~new_new_n23666__ & ~new_new_n23678__;
  assign new_new_n23680__ = new_new_n23321__ & ~new_new_n23679__;
  assign new_new_n23681__ = ~new_new_n23321__ & new_new_n23679__;
  assign new_new_n23682__ = new_new_n8470__ & ~new_new_n18633__;
  assign new_new_n23683__ = new_new_n8474__ & ~new_new_n15809__;
  assign new_new_n23684__ = ~new_new_n8479__ & ~new_new_n15487__;
  assign new_new_n23685__ = new_new_n8858__ & ~new_new_n15471__;
  assign new_new_n23686__ = ~new_new_n23683__ & ~new_new_n23684__;
  assign new_new_n23687__ = ~new_new_n23685__ & new_new_n23686__;
  assign new_new_n23688__ = ~new_new_n23682__ & new_new_n23687__;
  assign new_new_n23689__ = ~pi11 & new_new_n23688__;
  assign new_new_n23690__ = pi11 & ~new_new_n23688__;
  assign new_new_n23691__ = ~new_new_n23689__ & ~new_new_n23690__;
  assign new_new_n23692__ = ~new_new_n23681__ & ~new_new_n23691__;
  assign new_new_n23693__ = ~new_new_n23680__ & ~new_new_n23692__;
  assign new_new_n23694__ = ~new_new_n23317__ & new_new_n23693__;
  assign new_new_n23695__ = ~new_new_n23316__ & ~new_new_n23694__;
  assign new_new_n23696__ = ~new_new_n23299__ & ~new_new_n23695__;
  assign new_new_n23697__ = new_new_n23299__ & new_new_n23695__;
  assign new_new_n23698__ = new_new_n8858__ & ~new_new_n15439__;
  assign new_new_n23699__ = ~new_new_n8479__ & ~new_new_n15471__;
  assign new_new_n23700__ = new_new_n8474__ & new_new_n15464__;
  assign new_new_n23701__ = ~new_new_n23698__ & ~new_new_n23699__;
  assign new_new_n23702__ = ~new_new_n23700__ & new_new_n23701__;
  assign new_new_n23703__ = new_new_n8469__ & ~new_new_n17240__;
  assign new_new_n23704__ = pi11 & ~new_new_n23703__;
  assign new_new_n23705__ = new_new_n11530__ & ~new_new_n17240__;
  assign new_new_n23706__ = ~new_new_n23704__ & ~new_new_n23705__;
  assign new_new_n23707__ = new_new_n23702__ & ~new_new_n23706__;
  assign new_new_n23708__ = ~pi11 & ~new_new_n23702__;
  assign new_new_n23709__ = ~new_new_n23707__ & ~new_new_n23708__;
  assign new_new_n23710__ = ~new_new_n23697__ & ~new_new_n23709__;
  assign new_new_n23711__ = ~new_new_n23696__ & ~new_new_n23710__;
  assign new_new_n23712__ = new_new_n23295__ & ~new_new_n23711__;
  assign new_new_n23713__ = ~new_new_n23295__ & new_new_n23711__;
  assign new_new_n23714__ = ~new_new_n23037__ & ~new_new_n23038__;
  assign new_new_n23715__ = new_new_n23055__ & new_new_n23714__;
  assign new_new_n23716__ = ~new_new_n23055__ & ~new_new_n23714__;
  assign new_new_n23717__ = ~new_new_n23715__ & ~new_new_n23716__;
  assign new_new_n23718__ = ~new_new_n23713__ & ~new_new_n23717__;
  assign new_new_n23719__ = ~new_new_n23712__ & ~new_new_n23718__;
  assign new_new_n23720__ = ~new_new_n23283__ & ~new_new_n23719__;
  assign new_new_n23721__ = new_new_n23283__ & new_new_n23719__;
  assign new_new_n23722__ = ~new_new_n22304__ & ~new_new_n22583__;
  assign new_new_n23723__ = new_new_n22304__ & new_new_n22583__;
  assign new_new_n23724__ = ~new_new_n23722__ & ~new_new_n23723__;
  assign new_new_n23725__ = ~new_new_n21985__ & ~new_new_n23057__;
  assign new_new_n23726__ = new_new_n21985__ & new_new_n23057__;
  assign new_new_n23727__ = ~new_new_n23725__ & ~new_new_n23726__;
  assign new_new_n23728__ = new_new_n23724__ & new_new_n23727__;
  assign new_new_n23729__ = ~new_new_n23724__ & ~new_new_n23727__;
  assign new_new_n23730__ = ~new_new_n23728__ & ~new_new_n23729__;
  assign new_new_n23731__ = ~new_new_n23721__ & ~new_new_n23730__;
  assign new_new_n23732__ = ~new_new_n23720__ & ~new_new_n23731__;
  assign new_new_n23733__ = ~new_new_n23271__ & ~new_new_n23732__;
  assign new_new_n23734__ = ~new_new_n23270__ & ~new_new_n23733__;
  assign new_new_n23735__ = new_new_n23249__ & new_new_n23734__;
  assign new_new_n23736__ = ~new_new_n23249__ & ~new_new_n23734__;
  assign new_new_n23737__ = ~new_new_n23066__ & ~new_new_n23067__;
  assign new_new_n23738__ = new_new_n23084__ & ~new_new_n23737__;
  assign new_new_n23739__ = ~new_new_n23084__ & new_new_n23737__;
  assign new_new_n23740__ = ~new_new_n23738__ & ~new_new_n23739__;
  assign new_new_n23741__ = ~new_new_n23736__ & new_new_n23740__;
  assign new_new_n23742__ = ~new_new_n23735__ & ~new_new_n23741__;
  assign new_new_n23743__ = ~new_new_n23233__ & ~new_new_n23742__;
  assign new_new_n23744__ = new_new_n23233__ & new_new_n23742__;
  assign new_new_n23745__ = new_new_n8858__ & ~new_new_n15349__;
  assign new_new_n23746__ = ~new_new_n8479__ & new_new_n15390__;
  assign new_new_n23747__ = new_new_n8474__ & ~new_new_n15398__;
  assign new_new_n23748__ = new_new_n8470__ & ~new_new_n17180__;
  assign new_new_n23749__ = ~new_new_n23746__ & ~new_new_n23747__;
  assign new_new_n23750__ = ~new_new_n23745__ & new_new_n23749__;
  assign new_new_n23751__ = ~new_new_n23748__ & new_new_n23750__;
  assign new_new_n23752__ = pi11 & ~new_new_n23751__;
  assign new_new_n23753__ = ~pi11 & new_new_n23751__;
  assign new_new_n23754__ = ~new_new_n23752__ & ~new_new_n23753__;
  assign new_new_n23755__ = ~new_new_n23744__ & ~new_new_n23754__;
  assign new_new_n23756__ = ~new_new_n23743__ & ~new_new_n23755__;
  assign new_new_n23757__ = ~new_new_n23229__ & ~new_new_n23756__;
  assign new_new_n23758__ = ~new_new_n23228__ & ~new_new_n23757__;
  assign new_new_n23759__ = new_new_n23213__ & ~new_new_n23758__;
  assign new_new_n23760__ = ~new_new_n23213__ & new_new_n23758__;
  assign new_new_n23761__ = new_new_n8474__ & ~new_new_n15321__;
  assign new_new_n23762__ = ~new_new_n8479__ & ~new_new_n15349__;
  assign new_new_n23763__ = new_new_n8858__ & ~new_new_n15273__;
  assign new_new_n23764__ = ~new_new_n23761__ & ~new_new_n23762__;
  assign new_new_n23765__ = ~new_new_n23763__ & new_new_n23764__;
  assign new_new_n23766__ = new_new_n8469__ & ~new_new_n17103__;
  assign new_new_n23767__ = pi11 & ~new_new_n23766__;
  assign new_new_n23768__ = new_new_n11530__ & ~new_new_n17103__;
  assign new_new_n23769__ = ~new_new_n23767__ & ~new_new_n23768__;
  assign new_new_n23770__ = new_new_n23765__ & ~new_new_n23769__;
  assign new_new_n23771__ = ~pi11 & ~new_new_n23765__;
  assign new_new_n23772__ = ~new_new_n23770__ & ~new_new_n23771__;
  assign new_new_n23773__ = ~new_new_n23760__ & new_new_n23772__;
  assign new_new_n23774__ = ~new_new_n23759__ & ~new_new_n23773__;
  assign new_new_n23775__ = ~new_new_n23209__ & ~new_new_n23774__;
  assign new_new_n23776__ = new_new_n23209__ & new_new_n23774__;
  assign new_new_n23777__ = new_new_n8858__ & new_new_n15285__;
  assign new_new_n23778__ = ~new_new_n8479__ & ~new_new_n15321__;
  assign new_new_n23779__ = new_new_n8474__ & ~new_new_n15273__;
  assign new_new_n23780__ = new_new_n8470__ & new_new_n16078__;
  assign new_new_n23781__ = ~new_new_n23778__ & ~new_new_n23779__;
  assign new_new_n23782__ = ~new_new_n23777__ & new_new_n23781__;
  assign new_new_n23783__ = ~new_new_n23780__ & new_new_n23782__;
  assign new_new_n23784__ = ~pi11 & ~new_new_n23783__;
  assign new_new_n23785__ = pi11 & new_new_n23783__;
  assign new_new_n23786__ = ~new_new_n23784__ & ~new_new_n23785__;
  assign new_new_n23787__ = ~new_new_n23776__ & new_new_n23786__;
  assign new_new_n23788__ = ~new_new_n23775__ & ~new_new_n23787__;
  assign new_new_n23789__ = ~new_new_n23205__ & new_new_n23788__;
  assign new_new_n23790__ = new_new_n23205__ & ~new_new_n23788__;
  assign new_new_n23791__ = ~new_new_n22374__ & new_new_n23130__;
  assign new_new_n23792__ = new_new_n22374__ & ~new_new_n23130__;
  assign new_new_n23793__ = ~new_new_n23791__ & ~new_new_n23792__;
  assign new_new_n23794__ = new_new_n22474__ & ~new_new_n23793__;
  assign new_new_n23795__ = ~new_new_n22474__ & new_new_n23793__;
  assign new_new_n23796__ = ~new_new_n23794__ & ~new_new_n23795__;
  assign new_new_n23797__ = new_new_n22397__ & new_new_n23796__;
  assign new_new_n23798__ = ~new_new_n22397__ & ~new_new_n23796__;
  assign new_new_n23799__ = ~new_new_n23797__ & ~new_new_n23798__;
  assign new_new_n23800__ = ~new_new_n23790__ & ~new_new_n23799__;
  assign new_new_n23801__ = ~new_new_n23789__ & ~new_new_n23800__;
  assign new_new_n23802__ = ~new_new_n23193__ & ~new_new_n23801__;
  assign new_new_n23803__ = new_new_n23193__ & new_new_n23801__;
  assign new_new_n23804__ = ~new_new_n23153__ & ~new_new_n23155__;
  assign new_new_n23805__ = ~new_new_n23156__ & ~new_new_n23804__;
  assign new_new_n23806__ = ~new_new_n23803__ & ~new_new_n23805__;
  assign new_new_n23807__ = ~new_new_n23802__ & ~new_new_n23806__;
  assign new_new_n23808__ = ~new_new_n23162__ & ~new_new_n23163__;
  assign new_new_n23809__ = ~new_new_n23173__ & new_new_n23808__;
  assign new_new_n23810__ = new_new_n23173__ & ~new_new_n23808__;
  assign new_new_n23811__ = ~new_new_n23809__ & ~new_new_n23810__;
  assign new_new_n23812__ = new_new_n23807__ & new_new_n23811__;
  assign new_new_n23813__ = ~new_new_n23176__ & ~new_new_n23177__;
  assign new_new_n23814__ = ~new_new_n23179__ & ~new_new_n23813__;
  assign new_new_n23815__ = new_new_n23179__ & new_new_n23813__;
  assign new_new_n23816__ = ~new_new_n23814__ & ~new_new_n23815__;
  assign new_new_n23817__ = new_new_n23812__ & new_new_n23816__;
  assign new_new_n23818__ = ~new_new_n23789__ & ~new_new_n23790__;
  assign new_new_n23819__ = ~new_new_n22474__ & ~new_new_n23134__;
  assign new_new_n23820__ = new_new_n22474__ & new_new_n23134__;
  assign new_new_n23821__ = ~new_new_n23819__ & ~new_new_n23820__;
  assign new_new_n23822__ = ~new_new_n23130__ & new_new_n23821__;
  assign new_new_n23823__ = new_new_n23130__ & ~new_new_n23821__;
  assign new_new_n23824__ = ~new_new_n23822__ & ~new_new_n23823__;
  assign new_new_n23825__ = new_new_n23818__ & ~new_new_n23824__;
  assign new_new_n23826__ = ~new_new_n23818__ & new_new_n23824__;
  assign new_new_n23827__ = ~new_new_n23825__ & ~new_new_n23826__;
  assign new_new_n23828__ = new_new_n10702__ & ~new_new_n15314__;
  assign new_new_n23829__ = ~new_new_n11409__ & new_new_n15285__;
  assign new_new_n23830__ = new_new_n10698__ & ~new_new_n15248__;
  assign new_new_n23831__ = ~new_new_n23828__ & ~new_new_n23829__;
  assign new_new_n23832__ = ~new_new_n23830__ & new_new_n23831__;
  assign new_new_n23833__ = new_new_n10694__ & new_new_n16725__;
  assign new_new_n23834__ = pi08 & ~new_new_n23833__;
  assign new_new_n23835__ = new_new_n11498__ & new_new_n16725__;
  assign new_new_n23836__ = ~new_new_n23834__ & ~new_new_n23835__;
  assign new_new_n23837__ = new_new_n23832__ & ~new_new_n23836__;
  assign new_new_n23838__ = ~pi08 & ~new_new_n23832__;
  assign new_new_n23839__ = ~new_new_n23837__ & ~new_new_n23838__;
  assign new_new_n23840__ = new_new_n11378__ & new_new_n17140__;
  assign new_new_n23841__ = ~new_new_n11409__ & ~new_new_n15273__;
  assign new_new_n23842__ = new_new_n10702__ & new_new_n15285__;
  assign new_new_n23843__ = ~new_new_n23841__ & ~new_new_n23842__;
  assign new_new_n23844__ = ~new_new_n23840__ & new_new_n23843__;
  assign new_new_n23845__ = new_new_n10694__ & ~new_new_n15314__;
  assign new_new_n23846__ = ~pi08 & ~new_new_n23845__;
  assign new_new_n23847__ = new_new_n11498__ & ~new_new_n15314__;
  assign new_new_n23848__ = ~new_new_n23846__ & ~new_new_n23847__;
  assign new_new_n23849__ = new_new_n23844__ & ~new_new_n23848__;
  assign new_new_n23850__ = pi08 & ~new_new_n23844__;
  assign new_new_n23851__ = ~new_new_n23849__ & ~new_new_n23850__;
  assign new_new_n23852__ = ~new_new_n23743__ & ~new_new_n23744__;
  assign new_new_n23853__ = ~new_new_n23754__ & new_new_n23852__;
  assign new_new_n23854__ = new_new_n23754__ & ~new_new_n23852__;
  assign new_new_n23855__ = ~new_new_n23853__ & ~new_new_n23854__;
  assign new_new_n23856__ = ~new_new_n23735__ & ~new_new_n23736__;
  assign new_new_n23857__ = ~new_new_n23740__ & new_new_n23856__;
  assign new_new_n23858__ = new_new_n23740__ & ~new_new_n23856__;
  assign new_new_n23859__ = ~new_new_n23857__ & ~new_new_n23858__;
  assign new_new_n23860__ = new_new_n11378__ & new_new_n16458__;
  assign new_new_n23861__ = ~new_new_n11409__ & ~new_new_n15398__;
  assign new_new_n23862__ = new_new_n10702__ & ~new_new_n15349__;
  assign new_new_n23863__ = new_new_n10698__ & ~new_new_n15321__;
  assign new_new_n23864__ = ~new_new_n23861__ & ~new_new_n23862__;
  assign new_new_n23865__ = ~new_new_n23863__ & new_new_n23864__;
  assign new_new_n23866__ = ~new_new_n23860__ & new_new_n23865__;
  assign new_new_n23867__ = pi08 & ~new_new_n23866__;
  assign new_new_n23868__ = ~pi08 & new_new_n23866__;
  assign new_new_n23869__ = ~new_new_n23867__ & ~new_new_n23868__;
  assign new_new_n23870__ = new_new_n10698__ & ~new_new_n15349__;
  assign new_new_n23871__ = new_new_n10702__ & ~new_new_n15398__;
  assign new_new_n23872__ = ~new_new_n11409__ & new_new_n15390__;
  assign new_new_n23873__ = new_new_n11378__ & ~new_new_n17180__;
  assign new_new_n23874__ = ~new_new_n23871__ & ~new_new_n23872__;
  assign new_new_n23875__ = ~new_new_n23870__ & new_new_n23874__;
  assign new_new_n23876__ = ~new_new_n23873__ & new_new_n23875__;
  assign new_new_n23877__ = pi08 & ~new_new_n23876__;
  assign new_new_n23878__ = ~pi08 & new_new_n23876__;
  assign new_new_n23879__ = ~new_new_n23877__ & ~new_new_n23878__;
  assign new_new_n23880__ = ~new_new_n23057__ & new_new_n23719__;
  assign new_new_n23881__ = new_new_n23057__ & ~new_new_n23719__;
  assign new_new_n23882__ = ~new_new_n23880__ & ~new_new_n23881__;
  assign new_new_n23883__ = new_new_n21985__ & new_new_n23882__;
  assign new_new_n23884__ = ~new_new_n21985__ & ~new_new_n23882__;
  assign new_new_n23885__ = ~new_new_n23883__ & ~new_new_n23884__;
  assign new_new_n23886__ = new_new_n23724__ & ~new_new_n23885__;
  assign new_new_n23887__ = ~new_new_n23724__ & new_new_n23885__;
  assign new_new_n23888__ = ~new_new_n23886__ & ~new_new_n23887__;
  assign new_new_n23889__ = new_new_n23283__ & new_new_n23888__;
  assign new_new_n23890__ = ~new_new_n23283__ & ~new_new_n23888__;
  assign new_new_n23891__ = ~new_new_n23889__ & ~new_new_n23890__;
  assign new_new_n23892__ = new_new_n23879__ & ~new_new_n23891__;
  assign new_new_n23893__ = ~new_new_n23879__ & new_new_n23891__;
  assign new_new_n23894__ = new_new_n10702__ & new_new_n15390__;
  assign new_new_n23895__ = ~new_new_n11409__ & ~new_new_n15362__;
  assign new_new_n23896__ = ~new_new_n23894__ & ~new_new_n23895__;
  assign new_new_n23897__ = new_new_n10694__ & ~new_new_n17364__;
  assign new_new_n23898__ = pi08 & ~new_new_n23897__;
  assign new_new_n23899__ = ~pi07 & new_new_n15398__;
  assign new_new_n23900__ = pi07 & ~new_new_n15398__;
  assign new_new_n23901__ = new_new_n10694__ & ~new_new_n23899__;
  assign new_new_n23902__ = ~new_new_n23900__ & new_new_n23901__;
  assign new_new_n23903__ = new_new_n16956__ & new_new_n23902__;
  assign new_new_n23904__ = ~new_new_n23898__ & ~new_new_n23903__;
  assign new_new_n23905__ = new_new_n23896__ & ~new_new_n23904__;
  assign new_new_n23906__ = new_new_n10694__ & new_new_n17360__;
  assign new_new_n23907__ = new_new_n23896__ & ~new_new_n23906__;
  assign new_new_n23908__ = ~pi08 & ~new_new_n23907__;
  assign new_new_n23909__ = ~new_new_n23905__ & ~new_new_n23908__;
  assign new_new_n23910__ = ~new_new_n23712__ & ~new_new_n23713__;
  assign new_new_n23911__ = ~new_new_n23717__ & new_new_n23910__;
  assign new_new_n23912__ = new_new_n23717__ & ~new_new_n23910__;
  assign new_new_n23913__ = ~new_new_n23911__ & ~new_new_n23912__;
  assign new_new_n23914__ = ~new_new_n23909__ & new_new_n23913__;
  assign new_new_n23915__ = ~new_new_n11409__ & ~new_new_n15432__;
  assign new_new_n23916__ = new_new_n10702__ & ~new_new_n15362__;
  assign new_new_n23917__ = ~new_new_n23915__ & ~new_new_n23916__;
  assign new_new_n23918__ = new_new_n10694__ & new_new_n17914__;
  assign new_new_n23919__ = new_new_n23917__ & ~new_new_n23918__;
  assign new_new_n23920__ = pi08 & ~new_new_n23919__;
  assign new_new_n23921__ = new_new_n10694__ & ~new_new_n17918__;
  assign new_new_n23922__ = ~pi08 & ~new_new_n23921__;
  assign new_new_n23923__ = ~pi07 & new_new_n15390__;
  assign new_new_n23924__ = pi07 & ~new_new_n15390__;
  assign new_new_n23925__ = new_new_n10694__ & new_new_n15829__;
  assign new_new_n23926__ = ~new_new_n23923__ & ~new_new_n23924__;
  assign new_new_n23927__ = new_new_n23925__ & new_new_n23926__;
  assign new_new_n23928__ = ~new_new_n23922__ & ~new_new_n23927__;
  assign new_new_n23929__ = new_new_n23917__ & ~new_new_n23928__;
  assign new_new_n23930__ = ~new_new_n23920__ & ~new_new_n23929__;
  assign new_new_n23931__ = ~new_new_n23316__ & ~new_new_n23317__;
  assign new_new_n23932__ = new_new_n23693__ & new_new_n23931__;
  assign new_new_n23933__ = ~new_new_n23693__ & ~new_new_n23931__;
  assign new_new_n23934__ = ~new_new_n23932__ & ~new_new_n23933__;
  assign new_new_n23935__ = new_new_n11378__ & new_new_n17204__;
  assign new_new_n23936__ = ~new_new_n11409__ & new_new_n15464__;
  assign new_new_n23937__ = new_new_n10702__ & ~new_new_n15439__;
  assign new_new_n23938__ = ~new_new_n23936__ & ~new_new_n23937__;
  assign new_new_n23939__ = ~new_new_n23935__ & new_new_n23938__;
  assign new_new_n23940__ = new_new_n10694__ & ~new_new_n15432__;
  assign new_new_n23941__ = ~pi08 & ~new_new_n23940__;
  assign new_new_n23942__ = new_new_n11498__ & ~new_new_n15432__;
  assign new_new_n23943__ = ~new_new_n23941__ & ~new_new_n23942__;
  assign new_new_n23944__ = new_new_n23939__ & ~new_new_n23943__;
  assign new_new_n23945__ = pi08 & ~new_new_n23939__;
  assign new_new_n23946__ = ~new_new_n23944__ & ~new_new_n23945__;
  assign new_new_n23947__ = new_new_n11378__ & ~new_new_n17240__;
  assign new_new_n23948__ = ~new_new_n11409__ & ~new_new_n15471__;
  assign new_new_n23949__ = new_new_n10702__ & new_new_n15464__;
  assign new_new_n23950__ = ~new_new_n23948__ & ~new_new_n23949__;
  assign new_new_n23951__ = ~new_new_n23947__ & new_new_n23950__;
  assign new_new_n23952__ = new_new_n10694__ & ~new_new_n15439__;
  assign new_new_n23953__ = ~pi08 & ~new_new_n23952__;
  assign new_new_n23954__ = new_new_n11498__ & ~new_new_n15439__;
  assign new_new_n23955__ = ~new_new_n23953__ & ~new_new_n23954__;
  assign new_new_n23956__ = new_new_n23951__ & ~new_new_n23955__;
  assign new_new_n23957__ = pi08 & ~new_new_n23951__;
  assign new_new_n23958__ = ~new_new_n23956__ & ~new_new_n23957__;
  assign new_new_n23959__ = new_new_n11378__ & ~new_new_n18633__;
  assign new_new_n23960__ = ~new_new_n11409__ & ~new_new_n15487__;
  assign new_new_n23961__ = new_new_n10702__ & ~new_new_n15809__;
  assign new_new_n23962__ = ~new_new_n23960__ & ~new_new_n23961__;
  assign new_new_n23963__ = ~new_new_n23959__ & new_new_n23962__;
  assign new_new_n23964__ = new_new_n10694__ & ~new_new_n15471__;
  assign new_new_n23965__ = ~pi08 & ~new_new_n23964__;
  assign new_new_n23966__ = new_new_n11498__ & ~new_new_n15471__;
  assign new_new_n23967__ = ~new_new_n23965__ & ~new_new_n23966__;
  assign new_new_n23968__ = new_new_n23963__ & ~new_new_n23967__;
  assign new_new_n23969__ = pi08 & ~new_new_n23963__;
  assign new_new_n23970__ = ~new_new_n23968__ & ~new_new_n23969__;
  assign new_new_n23971__ = new_new_n10702__ & ~new_new_n15487__;
  assign new_new_n23972__ = ~new_new_n11409__ & new_new_n15524__;
  assign new_new_n23973__ = ~new_new_n23971__ & ~new_new_n23972__;
  assign new_new_n23974__ = new_new_n10694__ & ~new_new_n15809__;
  assign new_new_n23975__ = new_new_n18020__ & new_new_n23974__;
  assign new_new_n23976__ = new_new_n23973__ & ~new_new_n23975__;
  assign new_new_n23977__ = ~pi08 & ~new_new_n23976__;
  assign new_new_n23978__ = new_new_n10694__ & ~new_new_n18019__;
  assign new_new_n23979__ = pi08 & ~new_new_n23978__;
  assign new_new_n23980__ = ~pi07 & ~new_new_n18018__;
  assign new_new_n23981__ = pi07 & ~new_new_n20943__;
  assign new_new_n23982__ = new_new_n10694__ & ~new_new_n23980__;
  assign new_new_n23983__ = ~new_new_n23981__ & new_new_n23982__;
  assign new_new_n23984__ = ~new_new_n23979__ & ~new_new_n23983__;
  assign new_new_n23985__ = new_new_n23973__ & ~new_new_n23984__;
  assign new_new_n23986__ = ~new_new_n23977__ & ~new_new_n23985__;
  assign new_new_n23987__ = ~new_new_n23632__ & ~new_new_n23633__;
  assign new_new_n23988__ = ~new_new_n23637__ & new_new_n23987__;
  assign new_new_n23989__ = new_new_n23637__ & ~new_new_n23987__;
  assign new_new_n23990__ = ~new_new_n23988__ & ~new_new_n23989__;
  assign new_new_n23991__ = ~new_new_n23986__ & new_new_n23990__;
  assign new_new_n23992__ = new_new_n23986__ & ~new_new_n23990__;
  assign new_new_n23993__ = new_new_n10702__ & new_new_n15520__;
  assign new_new_n23994__ = ~new_new_n11409__ & ~new_new_n15533__;
  assign new_new_n23995__ = ~new_new_n23993__ & ~new_new_n23994__;
  assign new_new_n23996__ = new_new_n10694__ & ~new_new_n18914__;
  assign new_new_n23997__ = pi08 & ~new_new_n23996__;
  assign new_new_n23998__ = pi07 & ~new_new_n15524__;
  assign new_new_n23999__ = ~pi07 & new_new_n15524__;
  assign new_new_n24000__ = ~new_new_n23998__ & ~new_new_n23999__;
  assign new_new_n24001__ = new_new_n10694__ & ~new_new_n24000__;
  assign new_new_n24002__ = new_new_n18913__ & new_new_n24001__;
  assign new_new_n24003__ = ~new_new_n23997__ & ~new_new_n24002__;
  assign new_new_n24004__ = new_new_n23995__ & ~new_new_n24003__;
  assign new_new_n24005__ = new_new_n10694__ & new_new_n18923__;
  assign new_new_n24006__ = new_new_n23995__ & ~new_new_n24005__;
  assign new_new_n24007__ = ~pi08 & ~new_new_n24006__;
  assign new_new_n24008__ = ~new_new_n24004__ & ~new_new_n24007__;
  assign new_new_n24009__ = ~new_new_n23382__ & ~new_new_n23383__;
  assign new_new_n24010__ = ~new_new_n23583__ & new_new_n24009__;
  assign new_new_n24011__ = new_new_n23583__ & ~new_new_n24009__;
  assign new_new_n24012__ = ~new_new_n24010__ & ~new_new_n24011__;
  assign new_new_n24013__ = ~new_new_n11409__ & new_new_n15572__;
  assign new_new_n24014__ = new_new_n10702__ & new_new_n15560__;
  assign new_new_n24015__ = ~new_new_n10697__ & new_new_n18454__;
  assign new_new_n24016__ = new_new_n10697__ & ~new_new_n15767__;
  assign new_new_n24017__ = new_new_n10694__ & ~new_new_n24016__;
  assign new_new_n24018__ = ~new_new_n24015__ & new_new_n24017__;
  assign new_new_n24019__ = ~new_new_n24013__ & ~new_new_n24014__;
  assign new_new_n24020__ = ~new_new_n24018__ & new_new_n24019__;
  assign new_new_n24021__ = ~new_new_n24012__ & ~new_new_n24020__;
  assign new_new_n24022__ = ~new_new_n23545__ & ~new_new_n23546__;
  assign new_new_n24023__ = ~new_new_n23557__ & new_new_n24022__;
  assign new_new_n24024__ = new_new_n23557__ & ~new_new_n24022__;
  assign new_new_n24025__ = ~new_new_n24023__ & ~new_new_n24024__;
  assign new_new_n24026__ = ~new_new_n23531__ & ~new_new_n23532__;
  assign new_new_n24027__ = ~new_new_n23542__ & new_new_n24026__;
  assign new_new_n24028__ = new_new_n23542__ & ~new_new_n24026__;
  assign new_new_n24029__ = ~new_new_n24027__ & ~new_new_n24028__;
  assign new_new_n24030__ = ~new_new_n23517__ & ~new_new_n23518__;
  assign new_new_n24031__ = new_new_n23528__ & new_new_n24030__;
  assign new_new_n24032__ = ~new_new_n23528__ & ~new_new_n24030__;
  assign new_new_n24033__ = ~new_new_n24031__ & ~new_new_n24032__;
  assign new_new_n24034__ = ~new_new_n23508__ & ~new_new_n23509__;
  assign new_new_n24035__ = new_new_n23514__ & ~new_new_n24034__;
  assign new_new_n24036__ = ~new_new_n23514__ & new_new_n24034__;
  assign new_new_n24037__ = ~new_new_n24035__ & ~new_new_n24036__;
  assign new_new_n24038__ = ~new_new_n23494__ & ~new_new_n23495__;
  assign new_new_n24039__ = new_new_n23505__ & ~new_new_n24038__;
  assign new_new_n24040__ = ~new_new_n23505__ & new_new_n24038__;
  assign new_new_n24041__ = ~new_new_n24039__ & ~new_new_n24040__;
  assign new_new_n24042__ = pi11 & ~new_new_n8469__;
  assign new_new_n24043__ = new_new_n15674__ & new_new_n24042__;
  assign new_new_n24044__ = new_new_n8474__ & new_new_n15668__;
  assign new_new_n24045__ = ~pi11 & ~new_new_n24044__;
  assign new_new_n24046__ = new_new_n23471__ & ~new_new_n24043__;
  assign new_new_n24047__ = ~new_new_n24045__ & new_new_n24046__;
  assign new_new_n24048__ = new_new_n23480__ & ~new_new_n24047__;
  assign new_new_n24049__ = new_new_n8474__ & ~new_new_n15674__;
  assign new_new_n24050__ = new_new_n20003__ & ~new_new_n20628__;
  assign new_new_n24051__ = ~new_new_n24049__ & new_new_n24050__;
  assign new_new_n24052__ = ~new_new_n23480__ & new_new_n24051__;
  assign new_new_n24053__ = ~new_new_n24048__ & ~new_new_n24052__;
  assign new_new_n24054__ = ~new_new_n11409__ & new_new_n15668__;
  assign new_new_n24055__ = new_new_n10702__ & ~new_new_n15661__;
  assign new_new_n24056__ = ~new_new_n24054__ & ~new_new_n24055__;
  assign new_new_n24057__ = new_new_n10694__ & ~new_new_n20177__;
  assign new_new_n24058__ = pi08 & ~new_new_n24057__;
  assign new_new_n24059__ = pi07 & ~new_new_n15643__;
  assign new_new_n24060__ = ~pi07 & new_new_n15643__;
  assign new_new_n24061__ = ~new_new_n24059__ & ~new_new_n24060__;
  assign new_new_n24062__ = new_new_n10694__ & new_new_n20176__;
  assign new_new_n24063__ = ~new_new_n24061__ & new_new_n24062__;
  assign new_new_n24064__ = ~new_new_n24058__ & ~new_new_n24063__;
  assign new_new_n24065__ = new_new_n24056__ & ~new_new_n24064__;
  assign new_new_n24066__ = new_new_n10694__ & new_new_n20187__;
  assign new_new_n24067__ = new_new_n24056__ & ~new_new_n24066__;
  assign new_new_n24068__ = ~pi08 & ~new_new_n24067__;
  assign new_new_n24069__ = ~new_new_n24065__ & ~new_new_n24068__;
  assign new_new_n24070__ = new_new_n8469__ & ~new_new_n15673__;
  assign new_new_n24071__ = ~new_new_n12276__ & ~new_new_n20628__;
  assign new_new_n24072__ = new_new_n10694__ & ~new_new_n15661__;
  assign new_new_n24073__ = new_new_n11409__ & ~new_new_n24072__;
  assign new_new_n24074__ = ~new_new_n15673__ & ~new_new_n24073__;
  assign new_new_n24075__ = ~new_new_n10697__ & new_new_n15668__;
  assign new_new_n24076__ = ~new_new_n15679__ & new_new_n24075__;
  assign new_new_n24077__ = new_new_n15661__ & ~new_new_n24075__;
  assign new_new_n24078__ = new_new_n10694__ & ~new_new_n24077__;
  assign new_new_n24079__ = ~new_new_n24076__ & new_new_n24078__;
  assign new_new_n24080__ = ~new_new_n24074__ & ~new_new_n24079__;
  assign new_new_n24081__ = pi08 & ~new_new_n24071__;
  assign new_new_n24082__ = new_new_n24080__ & new_new_n24081__;
  assign new_new_n24083__ = ~new_new_n24070__ & ~new_new_n24082__;
  assign new_new_n24084__ = ~new_new_n24069__ & ~new_new_n24083__;
  assign new_new_n24085__ = new_new_n8472__ & new_new_n15674__;
  assign new_new_n24086__ = ~new_new_n8469__ & new_new_n20195__;
  assign new_new_n24087__ = ~new_new_n8301__ & new_new_n15668__;
  assign new_new_n24088__ = new_new_n8473__ & ~new_new_n24087__;
  assign new_new_n24089__ = ~new_new_n8855__ & ~new_new_n20628__;
  assign new_new_n24090__ = ~new_new_n24085__ & new_new_n24089__;
  assign new_new_n24091__ = ~new_new_n24086__ & ~new_new_n24088__;
  assign new_new_n24092__ = new_new_n24090__ & new_new_n24091__;
  assign new_new_n24093__ = new_new_n24084__ & new_new_n24092__;
  assign new_new_n24094__ = ~new_new_n24084__ & ~new_new_n24092__;
  assign new_new_n24095__ = new_new_n10698__ & new_new_n15656__;
  assign new_new_n24096__ = new_new_n10702__ & new_new_n15643__;
  assign new_new_n24097__ = ~new_new_n11409__ & ~new_new_n15661__;
  assign new_new_n24098__ = new_new_n11378__ & new_new_n15687__;
  assign new_new_n24099__ = ~new_new_n24096__ & ~new_new_n24097__;
  assign new_new_n24100__ = ~new_new_n24095__ & new_new_n24099__;
  assign new_new_n24101__ = ~new_new_n24098__ & new_new_n24100__;
  assign new_new_n24102__ = pi08 & ~new_new_n24101__;
  assign new_new_n24103__ = ~pi08 & new_new_n24101__;
  assign new_new_n24104__ = ~new_new_n24102__ & ~new_new_n24103__;
  assign new_new_n24105__ = ~new_new_n24094__ & new_new_n24104__;
  assign new_new_n24106__ = ~new_new_n24093__ & ~new_new_n24105__;
  assign new_new_n24107__ = new_new_n24053__ & ~new_new_n24106__;
  assign new_new_n24108__ = ~new_new_n24053__ & new_new_n24106__;
  assign new_new_n24109__ = new_new_n10698__ & ~new_new_n15710__;
  assign new_new_n24110__ = new_new_n10702__ & new_new_n15656__;
  assign new_new_n24111__ = ~new_new_n11409__ & new_new_n15643__;
  assign new_new_n24112__ = new_new_n11378__ & ~new_new_n19466__;
  assign new_new_n24113__ = ~new_new_n24110__ & ~new_new_n24111__;
  assign new_new_n24114__ = ~new_new_n24109__ & new_new_n24113__;
  assign new_new_n24115__ = ~new_new_n24112__ & new_new_n24114__;
  assign new_new_n24116__ = pi08 & ~new_new_n24115__;
  assign new_new_n24117__ = ~pi08 & new_new_n24115__;
  assign new_new_n24118__ = ~new_new_n24116__ & ~new_new_n24117__;
  assign new_new_n24119__ = ~new_new_n24108__ & new_new_n24118__;
  assign new_new_n24120__ = ~new_new_n24107__ & ~new_new_n24119__;
  assign new_new_n24121__ = ~new_new_n23468__ & ~new_new_n23469__;
  assign new_new_n24122__ = new_new_n23482__ & ~new_new_n24121__;
  assign new_new_n24123__ = new_new_n23468__ & ~new_new_n23469__;
  assign new_new_n24124__ = ~new_new_n23484__ & ~new_new_n24123__;
  assign new_new_n24125__ = ~new_new_n24122__ & ~new_new_n24124__;
  assign new_new_n24126__ = new_new_n10702__ & ~new_new_n15710__;
  assign new_new_n24127__ = ~new_new_n11409__ & new_new_n15656__;
  assign new_new_n24128__ = new_new_n10698__ & ~new_new_n15647__;
  assign new_new_n24129__ = ~new_new_n24126__ & ~new_new_n24127__;
  assign new_new_n24130__ = ~new_new_n24128__ & new_new_n24129__;
  assign new_new_n24131__ = new_new_n10694__ & ~new_new_n19118__;
  assign new_new_n24132__ = pi08 & ~new_new_n24131__;
  assign new_new_n24133__ = new_new_n11498__ & ~new_new_n19118__;
  assign new_new_n24134__ = ~new_new_n24132__ & ~new_new_n24133__;
  assign new_new_n24135__ = new_new_n24130__ & ~new_new_n24134__;
  assign new_new_n24136__ = ~pi08 & ~new_new_n24130__;
  assign new_new_n24137__ = ~new_new_n24135__ & ~new_new_n24136__;
  assign new_new_n24138__ = ~new_new_n24125__ & ~new_new_n24137__;
  assign new_new_n24139__ = new_new_n24120__ & ~new_new_n24138__;
  assign new_new_n24140__ = ~new_new_n24124__ & new_new_n24137__;
  assign new_new_n24141__ = ~new_new_n24139__ & ~new_new_n24140__;
  assign new_new_n24142__ = new_new_n24041__ & ~new_new_n24141__;
  assign new_new_n24143__ = ~new_new_n24041__ & new_new_n24141__;
  assign new_new_n24144__ = new_new_n10698__ & ~new_new_n15582__;
  assign new_new_n24145__ = new_new_n10702__ & ~new_new_n15647__;
  assign new_new_n24146__ = ~new_new_n11409__ & ~new_new_n15710__;
  assign new_new_n24147__ = new_new_n11378__ & ~new_new_n15736__;
  assign new_new_n24148__ = ~new_new_n24145__ & ~new_new_n24146__;
  assign new_new_n24149__ = ~new_new_n24144__ & new_new_n24148__;
  assign new_new_n24150__ = ~new_new_n24147__ & new_new_n24149__;
  assign new_new_n24151__ = pi08 & ~new_new_n24150__;
  assign new_new_n24152__ = ~pi08 & new_new_n24150__;
  assign new_new_n24153__ = ~new_new_n24151__ & ~new_new_n24152__;
  assign new_new_n24154__ = ~new_new_n24143__ & ~new_new_n24153__;
  assign new_new_n24155__ = ~new_new_n24142__ & ~new_new_n24154__;
  assign new_new_n24156__ = ~new_new_n24037__ & new_new_n24155__;
  assign new_new_n24157__ = new_new_n24037__ & ~new_new_n24155__;
  assign new_new_n24158__ = new_new_n10698__ & ~new_new_n15638__;
  assign new_new_n24159__ = new_new_n10702__ & ~new_new_n15582__;
  assign new_new_n24160__ = ~new_new_n11409__ & ~new_new_n15647__;
  assign new_new_n24161__ = new_new_n11378__ & new_new_n19487__;
  assign new_new_n24162__ = ~new_new_n24159__ & ~new_new_n24160__;
  assign new_new_n24163__ = ~new_new_n24158__ & new_new_n24162__;
  assign new_new_n24164__ = ~new_new_n24161__ & new_new_n24163__;
  assign new_new_n24165__ = ~pi08 & ~new_new_n24164__;
  assign new_new_n24166__ = pi08 & new_new_n24164__;
  assign new_new_n24167__ = ~new_new_n24165__ & ~new_new_n24166__;
  assign new_new_n24168__ = ~new_new_n24157__ & ~new_new_n24167__;
  assign new_new_n24169__ = ~new_new_n24156__ & ~new_new_n24168__;
  assign new_new_n24170__ = ~new_new_n24033__ & new_new_n24169__;
  assign new_new_n24171__ = new_new_n24033__ & ~new_new_n24169__;
  assign new_new_n24172__ = new_new_n11378__ & new_new_n19494__;
  assign new_new_n24173__ = new_new_n10702__ & ~new_new_n15638__;
  assign new_new_n24174__ = ~new_new_n11409__ & ~new_new_n15582__;
  assign new_new_n24175__ = new_new_n10698__ & new_new_n15743__;
  assign new_new_n24176__ = ~new_new_n24173__ & ~new_new_n24174__;
  assign new_new_n24177__ = ~new_new_n24175__ & new_new_n24176__;
  assign new_new_n24178__ = ~new_new_n24172__ & new_new_n24177__;
  assign new_new_n24179__ = pi08 & ~new_new_n24178__;
  assign new_new_n24180__ = ~pi08 & new_new_n24178__;
  assign new_new_n24181__ = ~new_new_n24179__ & ~new_new_n24180__;
  assign new_new_n24182__ = ~new_new_n24171__ & ~new_new_n24181__;
  assign new_new_n24183__ = ~new_new_n24170__ & ~new_new_n24182__;
  assign new_new_n24184__ = ~new_new_n24029__ & ~new_new_n24183__;
  assign new_new_n24185__ = new_new_n24029__ & new_new_n24183__;
  assign new_new_n24186__ = new_new_n10698__ & ~new_new_n15615__;
  assign new_new_n24187__ = ~new_new_n11409__ & ~new_new_n15638__;
  assign new_new_n24188__ = new_new_n10702__ & new_new_n15743__;
  assign new_new_n24189__ = ~new_new_n24187__ & ~new_new_n24188__;
  assign new_new_n24190__ = ~new_new_n24186__ & new_new_n24189__;
  assign new_new_n24191__ = new_new_n10694__ & new_new_n19005__;
  assign new_new_n24192__ = pi08 & ~new_new_n24191__;
  assign new_new_n24193__ = new_new_n11498__ & new_new_n19005__;
  assign new_new_n24194__ = ~new_new_n24192__ & ~new_new_n24193__;
  assign new_new_n24195__ = new_new_n24190__ & ~new_new_n24194__;
  assign new_new_n24196__ = ~pi08 & ~new_new_n24190__;
  assign new_new_n24197__ = ~new_new_n24195__ & ~new_new_n24196__;
  assign new_new_n24198__ = ~new_new_n24185__ & new_new_n24197__;
  assign new_new_n24199__ = ~new_new_n24184__ & ~new_new_n24198__;
  assign new_new_n24200__ = ~new_new_n24025__ & new_new_n24199__;
  assign new_new_n24201__ = new_new_n24025__ & ~new_new_n24199__;
  assign new_new_n24202__ = ~new_new_n24200__ & ~new_new_n24201__;
  assign new_new_n24203__ = new_new_n10698__ & new_new_n15564__;
  assign new_new_n24204__ = ~new_new_n11409__ & new_new_n15743__;
  assign new_new_n24205__ = new_new_n10702__ & ~new_new_n15615__;
  assign new_new_n24206__ = new_new_n11378__ & new_new_n18512__;
  assign new_new_n24207__ = ~new_new_n24204__ & ~new_new_n24205__;
  assign new_new_n24208__ = ~new_new_n24203__ & new_new_n24207__;
  assign new_new_n24209__ = ~new_new_n24206__ & new_new_n24208__;
  assign new_new_n24210__ = pi08 & ~new_new_n24209__;
  assign new_new_n24211__ = ~pi08 & new_new_n24209__;
  assign new_new_n24212__ = ~new_new_n24210__ & ~new_new_n24211__;
  assign new_new_n24213__ = new_new_n24202__ & new_new_n24212__;
  assign new_new_n24214__ = ~new_new_n24200__ & ~new_new_n24213__;
  assign new_new_n24215__ = ~new_new_n23416__ & ~new_new_n23417__;
  assign new_new_n24216__ = new_new_n23559__ & ~new_new_n24215__;
  assign new_new_n24217__ = ~new_new_n23559__ & new_new_n24215__;
  assign new_new_n24218__ = ~new_new_n24216__ & ~new_new_n24217__;
  assign new_new_n24219__ = ~new_new_n24214__ & new_new_n24218__;
  assign new_new_n24220__ = new_new_n24214__ & ~new_new_n24218__;
  assign new_new_n24221__ = new_new_n10698__ & new_new_n15572__;
  assign new_new_n24222__ = new_new_n10702__ & new_new_n15564__;
  assign new_new_n24223__ = ~new_new_n11409__ & ~new_new_n15615__;
  assign new_new_n24224__ = new_new_n11378__ & ~new_new_n20114__;
  assign new_new_n24225__ = ~new_new_n24222__ & ~new_new_n24223__;
  assign new_new_n24226__ = ~new_new_n24221__ & new_new_n24225__;
  assign new_new_n24227__ = ~new_new_n24224__ & new_new_n24226__;
  assign new_new_n24228__ = ~pi08 & ~new_new_n24227__;
  assign new_new_n24229__ = pi08 & new_new_n24227__;
  assign new_new_n24230__ = ~new_new_n24228__ & ~new_new_n24229__;
  assign new_new_n24231__ = ~new_new_n24220__ & ~new_new_n24230__;
  assign new_new_n24232__ = ~new_new_n24219__ & ~new_new_n24231__;
  assign new_new_n24233__ = ~new_new_n23562__ & ~new_new_n23563__;
  assign new_new_n24234__ = ~new_new_n23573__ & new_new_n24233__;
  assign new_new_n24235__ = new_new_n23573__ & ~new_new_n24233__;
  assign new_new_n24236__ = ~new_new_n24234__ & ~new_new_n24235__;
  assign new_new_n24237__ = ~new_new_n24232__ & ~new_new_n24236__;
  assign new_new_n24238__ = new_new_n24232__ & new_new_n24236__;
  assign new_new_n24239__ = new_new_n10698__ & new_new_n15560__;
  assign new_new_n24240__ = new_new_n10702__ & new_new_n15572__;
  assign new_new_n24241__ = ~new_new_n11409__ & new_new_n15564__;
  assign new_new_n24242__ = new_new_n11378__ & new_new_n18944__;
  assign new_new_n24243__ = ~new_new_n24240__ & ~new_new_n24241__;
  assign new_new_n24244__ = ~new_new_n24239__ & new_new_n24243__;
  assign new_new_n24245__ = ~new_new_n24242__ & new_new_n24244__;
  assign new_new_n24246__ = pi08 & ~new_new_n24245__;
  assign new_new_n24247__ = ~pi08 & new_new_n24245__;
  assign new_new_n24248__ = ~new_new_n24246__ & ~new_new_n24247__;
  assign new_new_n24249__ = ~new_new_n24238__ & new_new_n24248__;
  assign new_new_n24250__ = ~new_new_n24237__ & ~new_new_n24249__;
  assign new_new_n24251__ = ~new_new_n24020__ & new_new_n24250__;
  assign new_new_n24252__ = pi08 & ~new_new_n24251__;
  assign new_new_n24253__ = ~new_new_n24021__ & ~new_new_n24252__;
  assign new_new_n24254__ = new_new_n10698__ & ~new_new_n15533__;
  assign new_new_n24255__ = new_new_n10702__ & new_new_n15767__;
  assign new_new_n24256__ = ~new_new_n11409__ & new_new_n15560__;
  assign new_new_n24257__ = new_new_n11378__ & new_new_n19893__;
  assign new_new_n24258__ = ~new_new_n24255__ & ~new_new_n24256__;
  assign new_new_n24259__ = ~new_new_n24254__ & new_new_n24258__;
  assign new_new_n24260__ = ~new_new_n24257__ & new_new_n24259__;
  assign new_new_n24261__ = ~new_new_n24253__ & new_new_n24260__;
  assign new_new_n24262__ = ~pi08 & ~new_new_n24020__;
  assign new_new_n24263__ = ~new_new_n24012__ & new_new_n24020__;
  assign new_new_n24264__ = ~new_new_n24262__ & ~new_new_n24263__;
  assign new_new_n24265__ = ~new_new_n24260__ & ~new_new_n24264__;
  assign new_new_n24266__ = ~pi08 & ~new_new_n24260__;
  assign new_new_n24267__ = new_new_n24012__ & ~new_new_n24266__;
  assign new_new_n24268__ = ~new_new_n24250__ & ~new_new_n24267__;
  assign new_new_n24269__ = ~new_new_n24265__ & ~new_new_n24268__;
  assign new_new_n24270__ = ~new_new_n24261__ & new_new_n24269__;
  assign new_new_n24271__ = ~new_new_n23576__ & ~new_new_n23577__;
  assign new_new_n24272__ = new_new_n23581__ & new_new_n24271__;
  assign new_new_n24273__ = ~new_new_n23581__ & ~new_new_n24271__;
  assign new_new_n24274__ = ~new_new_n24272__ & ~new_new_n24273__;
  assign new_new_n24275__ = ~new_new_n24270__ & ~new_new_n24274__;
  assign new_new_n24276__ = pi08 & ~new_new_n24012__;
  assign new_new_n24277__ = pi08 & new_new_n24020__;
  assign new_new_n24278__ = ~new_new_n24021__ & ~new_new_n24277__;
  assign new_new_n24279__ = ~new_new_n24250__ & ~new_new_n24278__;
  assign new_new_n24280__ = ~new_new_n24276__ & ~new_new_n24279__;
  assign new_new_n24281__ = new_new_n24260__ & ~new_new_n24280__;
  assign new_new_n24282__ = ~pi08 & ~new_new_n24012__;
  assign new_new_n24283__ = ~new_new_n24250__ & ~new_new_n24264__;
  assign new_new_n24284__ = ~new_new_n24282__ & ~new_new_n24283__;
  assign new_new_n24285__ = ~new_new_n24260__ & ~new_new_n24284__;
  assign new_new_n24286__ = ~new_new_n24281__ & ~new_new_n24285__;
  assign new_new_n24287__ = ~new_new_n24275__ & new_new_n24286__;
  assign new_new_n24288__ = new_new_n11378__ & new_new_n19731__;
  assign new_new_n24289__ = ~new_new_n11409__ & new_new_n15767__;
  assign new_new_n24290__ = new_new_n10702__ & ~new_new_n15533__;
  assign new_new_n24291__ = ~new_new_n24289__ & ~new_new_n24290__;
  assign new_new_n24292__ = ~new_new_n24288__ & new_new_n24291__;
  assign new_new_n24293__ = new_new_n10694__ & new_new_n15520__;
  assign new_new_n24294__ = pi08 & ~new_new_n24293__;
  assign new_new_n24295__ = new_new_n12121__ & new_new_n15520__;
  assign new_new_n24296__ = ~new_new_n24294__ & ~new_new_n24295__;
  assign new_new_n24297__ = new_new_n24292__ & ~new_new_n24296__;
  assign new_new_n24298__ = ~pi08 & ~new_new_n24292__;
  assign new_new_n24299__ = ~new_new_n24297__ & ~new_new_n24298__;
  assign new_new_n24300__ = new_new_n24287__ & new_new_n24299__;
  assign new_new_n24301__ = ~new_new_n24287__ & ~new_new_n24299__;
  assign new_new_n24302__ = ~new_new_n23590__ & ~new_new_n23591__;
  assign new_new_n24303__ = ~new_new_n23603__ & new_new_n24302__;
  assign new_new_n24304__ = new_new_n23603__ & ~new_new_n24302__;
  assign new_new_n24305__ = ~new_new_n24303__ & ~new_new_n24304__;
  assign new_new_n24306__ = ~new_new_n24301__ & ~new_new_n24305__;
  assign new_new_n24307__ = ~new_new_n24300__ & ~new_new_n24306__;
  assign new_new_n24308__ = new_new_n22905__ & ~new_new_n22928__;
  assign new_new_n24309__ = ~new_new_n22905__ & new_new_n22928__;
  assign new_new_n24310__ = ~new_new_n24308__ & ~new_new_n24309__;
  assign new_new_n24311__ = ~new_new_n23605__ & new_new_n23619__;
  assign new_new_n24312__ = new_new_n23605__ & ~new_new_n23619__;
  assign new_new_n24313__ = ~new_new_n24311__ & ~new_new_n24312__;
  assign new_new_n24314__ = new_new_n24310__ & new_new_n24313__;
  assign new_new_n24315__ = ~new_new_n24310__ & ~new_new_n24313__;
  assign new_new_n24316__ = ~new_new_n24314__ & ~new_new_n24315__;
  assign new_new_n24317__ = new_new_n24307__ & new_new_n24316__;
  assign new_new_n24318__ = new_new_n24008__ & ~new_new_n24317__;
  assign new_new_n24319__ = ~new_new_n24307__ & ~new_new_n24316__;
  assign new_new_n24320__ = ~new_new_n24318__ & ~new_new_n24319__;
  assign new_new_n24321__ = ~new_new_n11409__ & new_new_n15520__;
  assign new_new_n24322__ = new_new_n10702__ & new_new_n15524__;
  assign new_new_n24323__ = new_new_n11378__ & new_new_n17587__;
  assign new_new_n24324__ = ~new_new_n24321__ & ~new_new_n24322__;
  assign new_new_n24325__ = ~new_new_n24323__ & new_new_n24324__;
  assign new_new_n24326__ = new_new_n10694__ & ~new_new_n15487__;
  assign new_new_n24327__ = pi08 & ~new_new_n24326__;
  assign new_new_n24328__ = new_new_n12121__ & ~new_new_n15487__;
  assign new_new_n24329__ = ~new_new_n24327__ & ~new_new_n24328__;
  assign new_new_n24330__ = new_new_n24325__ & ~new_new_n24329__;
  assign new_new_n24331__ = ~pi08 & ~new_new_n24325__;
  assign new_new_n24332__ = ~new_new_n24330__ & ~new_new_n24331__;
  assign new_new_n24333__ = new_new_n24320__ & ~new_new_n24332__;
  assign new_new_n24334__ = ~new_new_n24320__ & new_new_n24332__;
  assign new_new_n24335__ = ~new_new_n23624__ & ~new_new_n23625__;
  assign new_new_n24336__ = new_new_n23629__ & new_new_n24335__;
  assign new_new_n24337__ = ~new_new_n23629__ & ~new_new_n24335__;
  assign new_new_n24338__ = ~new_new_n24336__ & ~new_new_n24337__;
  assign new_new_n24339__ = ~new_new_n24334__ & new_new_n24338__;
  assign new_new_n24340__ = ~new_new_n24333__ & ~new_new_n24339__;
  assign new_new_n24341__ = ~new_new_n23992__ & ~new_new_n24340__;
  assign new_new_n24342__ = ~new_new_n23991__ & ~new_new_n24341__;
  assign new_new_n24343__ = new_new_n23970__ & ~new_new_n24342__;
  assign new_new_n24344__ = ~new_new_n23970__ & new_new_n24342__;
  assign new_new_n24345__ = ~new_new_n23640__ & ~new_new_n23641__;
  assign new_new_n24346__ = ~new_new_n23657__ & new_new_n24345__;
  assign new_new_n24347__ = new_new_n23657__ & ~new_new_n24345__;
  assign new_new_n24348__ = ~new_new_n24346__ & ~new_new_n24347__;
  assign new_new_n24349__ = ~new_new_n24344__ & ~new_new_n24348__;
  assign new_new_n24350__ = ~new_new_n24343__ & ~new_new_n24349__;
  assign new_new_n24351__ = ~new_new_n23338__ & ~new_new_n23339__;
  assign new_new_n24352__ = new_new_n23659__ & ~new_new_n24351__;
  assign new_new_n24353__ = ~new_new_n23659__ & new_new_n24351__;
  assign new_new_n24354__ = ~new_new_n24352__ & ~new_new_n24353__;
  assign new_new_n24355__ = ~new_new_n24350__ & new_new_n24354__;
  assign new_new_n24356__ = new_new_n24350__ & ~new_new_n24354__;
  assign new_new_n24357__ = new_new_n10698__ & new_new_n15464__;
  assign new_new_n24358__ = new_new_n10702__ & ~new_new_n15471__;
  assign new_new_n24359__ = ~new_new_n11409__ & ~new_new_n15809__;
  assign new_new_n24360__ = new_new_n11378__ & new_new_n15819__;
  assign new_new_n24361__ = ~new_new_n24358__ & ~new_new_n24359__;
  assign new_new_n24362__ = ~new_new_n24357__ & new_new_n24361__;
  assign new_new_n24363__ = ~new_new_n24360__ & new_new_n24362__;
  assign new_new_n24364__ = pi08 & ~new_new_n24363__;
  assign new_new_n24365__ = ~pi08 & new_new_n24363__;
  assign new_new_n24366__ = ~new_new_n24364__ & ~new_new_n24365__;
  assign new_new_n24367__ = ~new_new_n24356__ & new_new_n24366__;
  assign new_new_n24368__ = ~new_new_n24355__ & ~new_new_n24367__;
  assign new_new_n24369__ = new_new_n23958__ & ~new_new_n24368__;
  assign new_new_n24370__ = ~new_new_n23958__ & new_new_n24368__;
  assign new_new_n24371__ = ~new_new_n23666__ & ~new_new_n23667__;
  assign new_new_n24372__ = ~new_new_n23677__ & new_new_n24371__;
  assign new_new_n24373__ = new_new_n23677__ & ~new_new_n24371__;
  assign new_new_n24374__ = ~new_new_n24372__ & ~new_new_n24373__;
  assign new_new_n24375__ = ~new_new_n24370__ & ~new_new_n24374__;
  assign new_new_n24376__ = ~new_new_n24369__ & ~new_new_n24375__;
  assign new_new_n24377__ = new_new_n23946__ & ~new_new_n24376__;
  assign new_new_n24378__ = ~new_new_n23946__ & new_new_n24376__;
  assign new_new_n24379__ = ~new_new_n23680__ & ~new_new_n23681__;
  assign new_new_n24380__ = ~new_new_n23691__ & new_new_n24379__;
  assign new_new_n24381__ = new_new_n23691__ & ~new_new_n24379__;
  assign new_new_n24382__ = ~new_new_n24380__ & ~new_new_n24381__;
  assign new_new_n24383__ = ~new_new_n24378__ & ~new_new_n24382__;
  assign new_new_n24384__ = ~new_new_n24377__ & ~new_new_n24383__;
  assign new_new_n24385__ = new_new_n23934__ & ~new_new_n24384__;
  assign new_new_n24386__ = ~new_new_n23934__ & new_new_n24384__;
  assign new_new_n24387__ = new_new_n11378__ & new_new_n16771__;
  assign new_new_n24388__ = ~new_new_n11409__ & ~new_new_n15439__;
  assign new_new_n24389__ = new_new_n10702__ & ~new_new_n15432__;
  assign new_new_n24390__ = new_new_n10698__ & ~new_new_n15362__;
  assign new_new_n24391__ = ~new_new_n24388__ & ~new_new_n24389__;
  assign new_new_n24392__ = ~new_new_n24390__ & new_new_n24391__;
  assign new_new_n24393__ = ~new_new_n24387__ & new_new_n24392__;
  assign new_new_n24394__ = ~pi08 & ~new_new_n24393__;
  assign new_new_n24395__ = pi08 & new_new_n24393__;
  assign new_new_n24396__ = ~new_new_n24394__ & ~new_new_n24395__;
  assign new_new_n24397__ = ~new_new_n24386__ & ~new_new_n24396__;
  assign new_new_n24398__ = ~new_new_n24385__ & ~new_new_n24397__;
  assign new_new_n24399__ = new_new_n23930__ & ~new_new_n24398__;
  assign new_new_n24400__ = ~new_new_n23930__ & new_new_n24398__;
  assign new_new_n24401__ = ~new_new_n23696__ & ~new_new_n23697__;
  assign new_new_n24402__ = new_new_n23709__ & ~new_new_n24401__;
  assign new_new_n24403__ = ~new_new_n23709__ & new_new_n24401__;
  assign new_new_n24404__ = ~new_new_n24402__ & ~new_new_n24403__;
  assign new_new_n24405__ = ~new_new_n24400__ & new_new_n24404__;
  assign new_new_n24406__ = ~new_new_n24399__ & ~new_new_n24405__;
  assign new_new_n24407__ = new_new_n23909__ & ~new_new_n23913__;
  assign new_new_n24408__ = ~new_new_n24406__ & ~new_new_n24407__;
  assign new_new_n24409__ = ~new_new_n23914__ & ~new_new_n24408__;
  assign new_new_n24410__ = ~new_new_n23893__ & ~new_new_n24409__;
  assign new_new_n24411__ = ~new_new_n23892__ & ~new_new_n24410__;
  assign new_new_n24412__ = new_new_n23869__ & ~new_new_n24411__;
  assign new_new_n24413__ = ~new_new_n23869__ & new_new_n24411__;
  assign new_new_n24414__ = ~new_new_n23270__ & ~new_new_n23271__;
  assign new_new_n24415__ = ~new_new_n23732__ & ~new_new_n24414__;
  assign new_new_n24416__ = new_new_n23732__ & new_new_n24414__;
  assign new_new_n24417__ = ~new_new_n24415__ & ~new_new_n24416__;
  assign new_new_n24418__ = ~new_new_n24413__ & ~new_new_n24417__;
  assign new_new_n24419__ = ~new_new_n24412__ & ~new_new_n24418__;
  assign new_new_n24420__ = ~new_new_n23859__ & new_new_n24419__;
  assign new_new_n24421__ = new_new_n23859__ & ~new_new_n24419__;
  assign new_new_n24422__ = new_new_n10698__ & ~new_new_n15273__;
  assign new_new_n24423__ = new_new_n10702__ & ~new_new_n15321__;
  assign new_new_n24424__ = ~new_new_n11409__ & ~new_new_n15349__;
  assign new_new_n24425__ = new_new_n11378__ & ~new_new_n17103__;
  assign new_new_n24426__ = ~new_new_n24423__ & ~new_new_n24424__;
  assign new_new_n24427__ = ~new_new_n24422__ & new_new_n24426__;
  assign new_new_n24428__ = ~new_new_n24425__ & new_new_n24427__;
  assign new_new_n24429__ = pi08 & ~new_new_n24428__;
  assign new_new_n24430__ = ~pi08 & new_new_n24428__;
  assign new_new_n24431__ = ~new_new_n24429__ & ~new_new_n24430__;
  assign new_new_n24432__ = ~new_new_n24421__ & ~new_new_n24431__;
  assign new_new_n24433__ = ~new_new_n24420__ & ~new_new_n24432__;
  assign new_new_n24434__ = ~new_new_n23855__ & new_new_n24433__;
  assign new_new_n24435__ = new_new_n23855__ & ~new_new_n24433__;
  assign new_new_n24436__ = new_new_n11378__ & new_new_n16078__;
  assign new_new_n24437__ = ~new_new_n11409__ & ~new_new_n15321__;
  assign new_new_n24438__ = new_new_n10702__ & ~new_new_n15273__;
  assign new_new_n24439__ = new_new_n10698__ & new_new_n15285__;
  assign new_new_n24440__ = ~new_new_n24437__ & ~new_new_n24438__;
  assign new_new_n24441__ = ~new_new_n24439__ & new_new_n24440__;
  assign new_new_n24442__ = ~new_new_n24436__ & new_new_n24441__;
  assign new_new_n24443__ = ~pi08 & ~new_new_n24442__;
  assign new_new_n24444__ = pi08 & new_new_n24442__;
  assign new_new_n24445__ = ~new_new_n24443__ & ~new_new_n24444__;
  assign new_new_n24446__ = ~new_new_n24435__ & ~new_new_n24445__;
  assign new_new_n24447__ = ~new_new_n24434__ & ~new_new_n24446__;
  assign new_new_n24448__ = new_new_n23851__ & ~new_new_n24447__;
  assign new_new_n24449__ = ~new_new_n23851__ & new_new_n24447__;
  assign new_new_n24450__ = ~new_new_n22507__ & new_new_n23227__;
  assign new_new_n24451__ = new_new_n22507__ & ~new_new_n23227__;
  assign new_new_n24452__ = ~new_new_n24450__ & ~new_new_n24451__;
  assign new_new_n24453__ = new_new_n23094__ & new_new_n23756__;
  assign new_new_n24454__ = ~new_new_n23094__ & ~new_new_n23756__;
  assign new_new_n24455__ = ~new_new_n24453__ & ~new_new_n24454__;
  assign new_new_n24456__ = new_new_n24452__ & new_new_n24455__;
  assign new_new_n24457__ = ~new_new_n24452__ & ~new_new_n24455__;
  assign new_new_n24458__ = ~new_new_n24456__ & ~new_new_n24457__;
  assign new_new_n24459__ = ~new_new_n24449__ & new_new_n24458__;
  assign new_new_n24460__ = ~new_new_n24448__ & ~new_new_n24459__;
  assign new_new_n24461__ = new_new_n23839__ & new_new_n24460__;
  assign new_new_n24462__ = ~new_new_n23839__ & ~new_new_n24460__;
  assign new_new_n24463__ = ~new_new_n23759__ & ~new_new_n23760__;
  assign new_new_n24464__ = new_new_n23772__ & new_new_n24463__;
  assign new_new_n24465__ = ~new_new_n23772__ & ~new_new_n24463__;
  assign new_new_n24466__ = ~new_new_n24464__ & ~new_new_n24465__;
  assign new_new_n24467__ = ~new_new_n24462__ & new_new_n24466__;
  assign new_new_n24468__ = ~new_new_n24461__ & ~new_new_n24467__;
  assign new_new_n24469__ = ~pi11 & new_new_n23774__;
  assign new_new_n24470__ = pi11 & ~new_new_n23774__;
  assign new_new_n24471__ = ~new_new_n24469__ & ~new_new_n24470__;
  assign new_new_n24472__ = ~new_new_n23783__ & new_new_n24471__;
  assign new_new_n24473__ = new_new_n23783__ & ~new_new_n24471__;
  assign new_new_n24474__ = ~new_new_n24472__ & ~new_new_n24473__;
  assign new_new_n24475__ = new_new_n23209__ & new_new_n24474__;
  assign new_new_n24476__ = ~new_new_n23209__ & ~new_new_n24474__;
  assign new_new_n24477__ = ~new_new_n24475__ & ~new_new_n24476__;
  assign new_new_n24478__ = ~new_new_n24468__ & new_new_n24477__;
  assign new_new_n24479__ = new_new_n24468__ & ~new_new_n24477__;
  assign new_new_n24480__ = new_new_n10698__ & new_new_n15244__;
  assign new_new_n24481__ = new_new_n10702__ & ~new_new_n15248__;
  assign new_new_n24482__ = ~new_new_n11409__ & ~new_new_n15314__;
  assign new_new_n24483__ = new_new_n11378__ & new_new_n16378__;
  assign new_new_n24484__ = ~new_new_n24481__ & ~new_new_n24482__;
  assign new_new_n24485__ = ~new_new_n24480__ & new_new_n24484__;
  assign new_new_n24486__ = ~new_new_n24483__ & new_new_n24485__;
  assign new_new_n24487__ = pi08 & ~new_new_n24486__;
  assign new_new_n24488__ = ~pi08 & new_new_n24486__;
  assign new_new_n24489__ = ~new_new_n24487__ & ~new_new_n24488__;
  assign new_new_n24490__ = ~new_new_n24479__ & ~new_new_n24489__;
  assign new_new_n24491__ = ~new_new_n24478__ & ~new_new_n24490__;
  assign new_new_n24492__ = ~new_new_n23827__ & ~new_new_n24491__;
  assign new_new_n24493__ = new_new_n23827__ & new_new_n24491__;
  assign new_new_n24494__ = new_new_n10698__ & new_new_n15237__;
  assign new_new_n24495__ = new_new_n10702__ & new_new_n15244__;
  assign new_new_n24496__ = ~new_new_n11409__ & ~new_new_n15248__;
  assign new_new_n24497__ = new_new_n11378__ & ~new_new_n16603__;
  assign new_new_n24498__ = ~new_new_n24495__ & ~new_new_n24496__;
  assign new_new_n24499__ = ~new_new_n24494__ & new_new_n24498__;
  assign new_new_n24500__ = ~new_new_n24497__ & new_new_n24499__;
  assign new_new_n24501__ = pi08 & ~new_new_n24500__;
  assign new_new_n24502__ = ~pi08 & new_new_n24500__;
  assign new_new_n24503__ = ~new_new_n24501__ & ~new_new_n24502__;
  assign new_new_n24504__ = ~new_new_n24493__ & ~new_new_n24503__;
  assign new_new_n24505__ = ~new_new_n24492__ & ~new_new_n24504__;
  assign new_new_n24506__ = ~new_new_n23802__ & ~new_new_n23803__;
  assign new_new_n24507__ = ~new_new_n23805__ & new_new_n24506__;
  assign new_new_n24508__ = new_new_n23805__ & ~new_new_n24506__;
  assign new_new_n24509__ = ~new_new_n24507__ & ~new_new_n24508__;
  assign new_new_n24510__ = new_new_n24505__ & new_new_n24509__;
  assign new_new_n24511__ = ~new_new_n24505__ & ~new_new_n24509__;
  assign new_new_n24512__ = new_new_n12832__ & ~new_new_n15998__;
  assign new_new_n24513__ = new_new_n13069__ & new_new_n16630__;
  assign new_new_n24514__ = new_new_n11475__ & ~new_new_n16056__;
  assign new_new_n24515__ = ~new_new_n12850__ & ~new_new_n24514__;
  assign new_new_n24516__ = ~new_new_n24512__ & new_new_n24515__;
  assign new_new_n24517__ = ~new_new_n24513__ & new_new_n24516__;
  assign new_new_n24518__ = pi05 & ~new_new_n24517__;
  assign new_new_n24519__ = ~pi05 & new_new_n24517__;
  assign new_new_n24520__ = ~new_new_n24518__ & ~new_new_n24519__;
  assign new_new_n24521__ = ~new_new_n24511__ & new_new_n24520__;
  assign new_new_n24522__ = ~new_new_n24510__ & ~new_new_n24521__;
  assign new_new_n24523__ = new_new_n12850__ & ~new_new_n15998__;
  assign new_new_n24524__ = new_new_n11475__ & new_new_n15905__;
  assign new_new_n24525__ = new_new_n11471__ & new_new_n15237__;
  assign new_new_n24526__ = new_new_n13069__ & new_new_n16025__;
  assign new_new_n24527__ = ~new_new_n24524__ & ~new_new_n24525__;
  assign new_new_n24528__ = ~new_new_n24523__ & new_new_n24527__;
  assign new_new_n24529__ = ~new_new_n24526__ & new_new_n24528__;
  assign new_new_n24530__ = ~pi05 & ~new_new_n24529__;
  assign new_new_n24531__ = pi05 & new_new_n24529__;
  assign new_new_n24532__ = ~new_new_n24530__ & ~new_new_n24531__;
  assign new_new_n24533__ = ~new_new_n24448__ & ~new_new_n24449__;
  assign new_new_n24534__ = new_new_n24452__ & ~new_new_n24455__;
  assign new_new_n24535__ = ~new_new_n24452__ & new_new_n24455__;
  assign new_new_n24536__ = ~new_new_n24534__ & ~new_new_n24535__;
  assign new_new_n24537__ = new_new_n24533__ & new_new_n24536__;
  assign new_new_n24538__ = ~new_new_n24533__ & ~new_new_n24536__;
  assign new_new_n24539__ = ~new_new_n24537__ & ~new_new_n24538__;
  assign new_new_n24540__ = ~new_new_n24434__ & ~new_new_n24435__;
  assign new_new_n24541__ = ~new_new_n24445__ & new_new_n24540__;
  assign new_new_n24542__ = new_new_n24445__ & ~new_new_n24540__;
  assign new_new_n24543__ = ~new_new_n24541__ & ~new_new_n24542__;
  assign new_new_n24544__ = new_new_n11475__ & ~new_new_n15273__;
  assign new_new_n24545__ = new_new_n11471__ & ~new_new_n15321__;
  assign new_new_n24546__ = new_new_n12850__ & new_new_n15285__;
  assign new_new_n24547__ = ~new_new_n24544__ & ~new_new_n24545__;
  assign new_new_n24548__ = ~new_new_n24546__ & new_new_n24547__;
  assign new_new_n24549__ = pi05 & ~new_new_n24548__;
  assign new_new_n24550__ = new_new_n12856__ & new_new_n16078__;
  assign new_new_n24551__ = new_new_n11469__ & new_new_n16078__;
  assign new_new_n24552__ = ~pi05 & ~new_new_n24551__;
  assign new_new_n24553__ = ~new_new_n24550__ & ~new_new_n24552__;
  assign new_new_n24554__ = new_new_n24548__ & ~new_new_n24553__;
  assign new_new_n24555__ = ~new_new_n24549__ & ~new_new_n24554__;
  assign new_new_n24556__ = ~new_new_n23892__ & ~new_new_n23893__;
  assign new_new_n24557__ = new_new_n24409__ & new_new_n24556__;
  assign new_new_n24558__ = ~new_new_n24409__ & ~new_new_n24556__;
  assign new_new_n24559__ = ~new_new_n24557__ & ~new_new_n24558__;
  assign new_new_n24560__ = ~new_new_n24555__ & new_new_n24559__;
  assign new_new_n24561__ = new_new_n24555__ & ~new_new_n24559__;
  assign new_new_n24562__ = new_new_n11471__ & ~new_new_n15362__;
  assign new_new_n24563__ = new_new_n11475__ & new_new_n15390__;
  assign new_new_n24564__ = new_new_n11478__ & new_new_n16956__;
  assign new_new_n24565__ = new_new_n15398__ & ~new_new_n24564__;
  assign new_new_n24566__ = ~new_new_n15398__ & new_new_n24564__;
  assign new_new_n24567__ = new_new_n11469__ & ~new_new_n24565__;
  assign new_new_n24568__ = ~new_new_n24566__ & new_new_n24567__;
  assign new_new_n24569__ = ~new_new_n24562__ & ~new_new_n24563__;
  assign new_new_n24570__ = ~new_new_n24568__ & new_new_n24569__;
  assign new_new_n24571__ = ~new_new_n24385__ & ~new_new_n24386__;
  assign new_new_n24572__ = ~new_new_n24396__ & new_new_n24571__;
  assign new_new_n24573__ = new_new_n24396__ & ~new_new_n24571__;
  assign new_new_n24574__ = ~new_new_n24572__ & ~new_new_n24573__;
  assign new_new_n24575__ = ~new_new_n24570__ & new_new_n24574__;
  assign new_new_n24576__ = new_new_n12832__ & ~new_new_n15439__;
  assign new_new_n24577__ = new_new_n11475__ & ~new_new_n15432__;
  assign new_new_n24578__ = ~new_new_n11478__ & new_new_n15362__;
  assign new_new_n24579__ = new_new_n11478__ & ~new_new_n16771__;
  assign new_new_n24580__ = ~new_new_n11482__ & ~new_new_n24578__;
  assign new_new_n24581__ = ~new_new_n24579__ & new_new_n24580__;
  assign new_new_n24582__ = ~new_new_n24576__ & ~new_new_n24577__;
  assign new_new_n24583__ = ~new_new_n24581__ & new_new_n24582__;
  assign new_new_n24584__ = ~pi05 & new_new_n24583__;
  assign new_new_n24585__ = pi05 & ~new_new_n24583__;
  assign new_new_n24586__ = ~new_new_n24584__ & ~new_new_n24585__;
  assign new_new_n24587__ = ~new_new_n24355__ & ~new_new_n24356__;
  assign new_new_n24588__ = new_new_n24366__ & new_new_n24587__;
  assign new_new_n24589__ = ~new_new_n24366__ & ~new_new_n24587__;
  assign new_new_n24590__ = ~new_new_n24588__ & ~new_new_n24589__;
  assign new_new_n24591__ = ~new_new_n24586__ & ~new_new_n24590__;
  assign new_new_n24592__ = new_new_n24586__ & new_new_n24590__;
  assign new_new_n24593__ = ~new_new_n24343__ & ~new_new_n24344__;
  assign new_new_n24594__ = ~new_new_n24348__ & new_new_n24593__;
  assign new_new_n24595__ = new_new_n24348__ & ~new_new_n24593__;
  assign new_new_n24596__ = ~new_new_n24594__ & ~new_new_n24595__;
  assign new_new_n24597__ = new_new_n13111__ & ~new_new_n15809__;
  assign new_new_n24598__ = new_new_n11469__ & new_new_n15819__;
  assign new_new_n24599__ = ~new_new_n24597__ & ~new_new_n24598__;
  assign new_new_n24600__ = new_new_n11478__ & ~new_new_n24599__;
  assign new_new_n24601__ = new_new_n11475__ & ~new_new_n15471__;
  assign new_new_n24602__ = ~new_new_n24600__ & ~new_new_n24601__;
  assign new_new_n24603__ = ~pi05 & ~new_new_n24602__;
  assign new_new_n24604__ = new_new_n12856__ & new_new_n15464__;
  assign new_new_n24605__ = new_new_n11469__ & new_new_n15464__;
  assign new_new_n24606__ = pi05 & ~new_new_n24605__;
  assign new_new_n24607__ = ~new_new_n24604__ & ~new_new_n24606__;
  assign new_new_n24608__ = new_new_n24602__ & ~new_new_n24607__;
  assign new_new_n24609__ = ~new_new_n24603__ & ~new_new_n24608__;
  assign new_new_n24610__ = new_new_n11475__ & ~new_new_n15809__;
  assign new_new_n24611__ = new_new_n11471__ & ~new_new_n15487__;
  assign new_new_n24612__ = new_new_n12850__ & ~new_new_n15471__;
  assign new_new_n24613__ = ~new_new_n24610__ & ~new_new_n24611__;
  assign new_new_n24614__ = ~new_new_n24612__ & new_new_n24613__;
  assign new_new_n24615__ = pi05 & ~new_new_n24614__;
  assign new_new_n24616__ = new_new_n12856__ & ~new_new_n18633__;
  assign new_new_n24617__ = new_new_n11469__ & ~new_new_n18633__;
  assign new_new_n24618__ = ~pi05 & ~new_new_n24617__;
  assign new_new_n24619__ = ~new_new_n24616__ & ~new_new_n24618__;
  assign new_new_n24620__ = new_new_n24614__ & ~new_new_n24619__;
  assign new_new_n24621__ = ~new_new_n24615__ & ~new_new_n24620__;
  assign new_new_n24622__ = new_new_n12850__ & ~new_new_n15809__;
  assign new_new_n24623__ = new_new_n11471__ & new_new_n15524__;
  assign new_new_n24624__ = new_new_n11475__ & ~new_new_n15487__;
  assign new_new_n24625__ = ~new_new_n24623__ & ~new_new_n24624__;
  assign new_new_n24626__ = ~new_new_n24622__ & new_new_n24625__;
  assign new_new_n24627__ = pi05 & ~new_new_n24626__;
  assign new_new_n24628__ = new_new_n12856__ & new_new_n18020__;
  assign new_new_n24629__ = new_new_n11469__ & new_new_n18020__;
  assign new_new_n24630__ = ~pi05 & ~new_new_n24629__;
  assign new_new_n24631__ = ~new_new_n24628__ & ~new_new_n24630__;
  assign new_new_n24632__ = new_new_n24626__ & ~new_new_n24631__;
  assign new_new_n24633__ = ~new_new_n24627__ & ~new_new_n24632__;
  assign new_new_n24634__ = ~new_new_n24300__ & ~new_new_n24301__;
  assign new_new_n24635__ = ~new_new_n24305__ & new_new_n24634__;
  assign new_new_n24636__ = new_new_n24305__ & ~new_new_n24634__;
  assign new_new_n24637__ = ~new_new_n24635__ & ~new_new_n24636__;
  assign new_new_n24638__ = new_new_n24633__ & ~new_new_n24637__;
  assign new_new_n24639__ = ~new_new_n24633__ & new_new_n24637__;
  assign new_new_n24640__ = new_new_n24250__ & new_new_n24274__;
  assign new_new_n24641__ = ~pi08 & new_new_n24012__;
  assign new_new_n24642__ = ~new_new_n24276__ & ~new_new_n24641__;
  assign new_new_n24643__ = ~new_new_n24260__ & new_new_n24642__;
  assign new_new_n24644__ = new_new_n24260__ & ~new_new_n24642__;
  assign new_new_n24645__ = ~new_new_n24643__ & ~new_new_n24644__;
  assign new_new_n24646__ = new_new_n24640__ & ~new_new_n24645__;
  assign new_new_n24647__ = ~new_new_n24250__ & ~new_new_n24274__;
  assign new_new_n24648__ = ~new_new_n24640__ & ~new_new_n24647__;
  assign new_new_n24649__ = new_new_n24012__ & ~new_new_n24020__;
  assign new_new_n24650__ = ~new_new_n24263__ & ~new_new_n24649__;
  assign new_new_n24651__ = new_new_n24260__ & ~new_new_n24650__;
  assign new_new_n24652__ = ~new_new_n24260__ & new_new_n24650__;
  assign new_new_n24653__ = ~new_new_n24651__ & ~new_new_n24652__;
  assign new_new_n24654__ = new_new_n24648__ & new_new_n24653__;
  assign new_new_n24655__ = new_new_n24645__ & new_new_n24647__;
  assign new_new_n24656__ = ~new_new_n24646__ & ~new_new_n24655__;
  assign new_new_n24657__ = ~new_new_n24654__ & new_new_n24656__;
  assign new_new_n24658__ = new_new_n12832__ & ~new_new_n15533__;
  assign new_new_n24659__ = new_new_n11475__ & new_new_n15520__;
  assign new_new_n24660__ = ~new_new_n24658__ & ~new_new_n24659__;
  assign new_new_n24661__ = new_new_n11469__ & new_new_n18923__;
  assign new_new_n24662__ = new_new_n24660__ & ~new_new_n24661__;
  assign new_new_n24663__ = pi05 & ~new_new_n24662__;
  assign new_new_n24664__ = ~pi04 & new_new_n15524__;
  assign new_new_n24665__ = pi04 & ~new_new_n15524__;
  assign new_new_n24666__ = ~new_new_n11482__ & ~new_new_n24664__;
  assign new_new_n24667__ = ~new_new_n24665__ & new_new_n24666__;
  assign new_new_n24668__ = new_new_n18913__ & new_new_n24667__;
  assign new_new_n24669__ = new_new_n11469__ & ~new_new_n18914__;
  assign new_new_n24670__ = ~pi05 & ~new_new_n24669__;
  assign new_new_n24671__ = ~new_new_n24668__ & ~new_new_n24670__;
  assign new_new_n24672__ = new_new_n24660__ & ~new_new_n24671__;
  assign new_new_n24673__ = ~new_new_n24663__ & ~new_new_n24672__;
  assign new_new_n24674__ = ~new_new_n24237__ & ~new_new_n24238__;
  assign new_new_n24675__ = ~new_new_n24248__ & new_new_n24674__;
  assign new_new_n24676__ = new_new_n24248__ & ~new_new_n24674__;
  assign new_new_n24677__ = ~new_new_n24675__ & ~new_new_n24676__;
  assign new_new_n24678__ = new_new_n11475__ & new_new_n15560__;
  assign new_new_n24679__ = new_new_n11471__ & new_new_n15572__;
  assign new_new_n24680__ = new_new_n12850__ & new_new_n15767__;
  assign new_new_n24681__ = ~new_new_n24679__ & ~new_new_n24680__;
  assign new_new_n24682__ = ~new_new_n24678__ & new_new_n24681__;
  assign new_new_n24683__ = pi05 & ~new_new_n24682__;
  assign new_new_n24684__ = new_new_n12856__ & ~new_new_n18454__;
  assign new_new_n24685__ = new_new_n11469__ & ~new_new_n18454__;
  assign new_new_n24686__ = ~pi05 & ~new_new_n24685__;
  assign new_new_n24687__ = ~new_new_n24684__ & ~new_new_n24686__;
  assign new_new_n24688__ = new_new_n24682__ & ~new_new_n24687__;
  assign new_new_n24689__ = ~new_new_n24683__ & ~new_new_n24688__;
  assign new_new_n24690__ = new_new_n11475__ & new_new_n15572__;
  assign new_new_n24691__ = ~new_new_n11478__ & ~new_new_n15560__;
  assign new_new_n24692__ = new_new_n11478__ & ~new_new_n18944__;
  assign new_new_n24693__ = ~new_new_n11482__ & ~new_new_n24691__;
  assign new_new_n24694__ = ~new_new_n24692__ & new_new_n24693__;
  assign new_new_n24695__ = ~new_new_n24690__ & ~new_new_n24694__;
  assign new_new_n24696__ = new_new_n11466__ & new_new_n15564__;
  assign new_new_n24697__ = pi05 & ~new_new_n24696__;
  assign new_new_n24698__ = new_new_n11467__ & new_new_n15564__;
  assign new_new_n24699__ = ~pi05 & ~new_new_n24698__;
  assign new_new_n24700__ = pi02 & ~new_new_n24699__;
  assign new_new_n24701__ = ~new_new_n24697__ & ~new_new_n24700__;
  assign new_new_n24702__ = new_new_n24695__ & ~new_new_n24701__;
  assign new_new_n24703__ = ~pi05 & ~new_new_n24695__;
  assign new_new_n24704__ = ~new_new_n24702__ & ~new_new_n24703__;
  assign new_new_n24705__ = ~new_new_n24156__ & ~new_new_n24157__;
  assign new_new_n24706__ = new_new_n24167__ & new_new_n24705__;
  assign new_new_n24707__ = ~new_new_n24167__ & ~new_new_n24705__;
  assign new_new_n24708__ = ~new_new_n24706__ & ~new_new_n24707__;
  assign new_new_n24709__ = ~new_new_n24142__ & ~new_new_n24143__;
  assign new_new_n24710__ = ~new_new_n24153__ & new_new_n24709__;
  assign new_new_n24711__ = new_new_n24153__ & ~new_new_n24709__;
  assign new_new_n24712__ = ~new_new_n24710__ & ~new_new_n24711__;
  assign new_new_n24713__ = ~new_new_n24120__ & new_new_n24137__;
  assign new_new_n24714__ = new_new_n24120__ & ~new_new_n24137__;
  assign new_new_n24715__ = ~new_new_n24713__ & ~new_new_n24714__;
  assign new_new_n24716__ = new_new_n24125__ & new_new_n24715__;
  assign new_new_n24717__ = new_new_n24121__ & ~new_new_n24715__;
  assign new_new_n24718__ = new_new_n23468__ & new_new_n23469__;
  assign new_new_n24719__ = new_new_n24713__ & new_new_n24718__;
  assign new_new_n24720__ = ~new_new_n24717__ & ~new_new_n24719__;
  assign new_new_n24721__ = ~new_new_n23482__ & ~new_new_n24720__;
  assign new_new_n24722__ = ~new_new_n24122__ & ~new_new_n24718__;
  assign new_new_n24723__ = new_new_n24714__ & ~new_new_n24722__;
  assign new_new_n24724__ = ~new_new_n24716__ & ~new_new_n24723__;
  assign new_new_n24725__ = ~new_new_n24721__ & new_new_n24724__;
  assign new_new_n24726__ = new_new_n13069__ & new_new_n19494__;
  assign new_new_n24727__ = new_new_n11475__ & ~new_new_n15638__;
  assign new_new_n24728__ = new_new_n11471__ & ~new_new_n15582__;
  assign new_new_n24729__ = new_new_n12850__ & new_new_n15743__;
  assign new_new_n24730__ = ~new_new_n24727__ & ~new_new_n24728__;
  assign new_new_n24731__ = ~new_new_n24729__ & new_new_n24730__;
  assign new_new_n24732__ = ~new_new_n24726__ & new_new_n24731__;
  assign new_new_n24733__ = new_new_n12850__ & ~new_new_n15638__;
  assign new_new_n24734__ = new_new_n11475__ & ~new_new_n15582__;
  assign new_new_n24735__ = new_new_n11471__ & ~new_new_n15647__;
  assign new_new_n24736__ = new_new_n13069__ & new_new_n19487__;
  assign new_new_n24737__ = ~new_new_n24734__ & ~new_new_n24735__;
  assign new_new_n24738__ = ~new_new_n24733__ & new_new_n24737__;
  assign new_new_n24739__ = ~new_new_n24736__ & new_new_n24738__;
  assign new_new_n24740__ = ~new_new_n24732__ & new_new_n24739__;
  assign new_new_n24741__ = new_new_n24732__ & ~new_new_n24739__;
  assign new_new_n24742__ = ~new_new_n24740__ & ~new_new_n24741__;
  assign new_new_n24743__ = new_new_n24725__ & ~new_new_n24742__;
  assign new_new_n24744__ = ~new_new_n24107__ & ~new_new_n24108__;
  assign new_new_n24745__ = new_new_n24118__ & new_new_n24744__;
  assign new_new_n24746__ = ~new_new_n24118__ & ~new_new_n24744__;
  assign new_new_n24747__ = ~new_new_n24745__ & ~new_new_n24746__;
  assign new_new_n24748__ = ~new_new_n24093__ & ~new_new_n24094__;
  assign new_new_n24749__ = new_new_n24104__ & new_new_n24748__;
  assign new_new_n24750__ = ~new_new_n24104__ & ~new_new_n24748__;
  assign new_new_n24751__ = ~new_new_n24749__ & ~new_new_n24750__;
  assign new_new_n24752__ = new_new_n11471__ & new_new_n15656__;
  assign new_new_n24753__ = new_new_n11475__ & ~new_new_n15710__;
  assign new_new_n24754__ = new_new_n11478__ & new_new_n19118__;
  assign new_new_n24755__ = ~new_new_n11478__ & new_new_n15647__;
  assign new_new_n24756__ = ~new_new_n11482__ & ~new_new_n24755__;
  assign new_new_n24757__ = ~new_new_n24754__ & new_new_n24756__;
  assign new_new_n24758__ = ~new_new_n24752__ & ~new_new_n24753__;
  assign new_new_n24759__ = ~new_new_n24757__ & new_new_n24758__;
  assign new_new_n24760__ = ~pi05 & ~new_new_n24759__;
  assign new_new_n24761__ = pi05 & new_new_n24759__;
  assign new_new_n24762__ = ~new_new_n24760__ & ~new_new_n24761__;
  assign new_new_n24763__ = new_new_n10694__ & ~new_new_n20628__;
  assign new_new_n24764__ = new_new_n24080__ & new_new_n24763__;
  assign new_new_n24765__ = new_new_n10702__ & ~new_new_n15673__;
  assign new_new_n24766__ = ~new_new_n15668__ & new_new_n24765__;
  assign new_new_n24767__ = ~new_new_n24764__ & ~new_new_n24766__;
  assign new_new_n24768__ = pi08 & ~new_new_n24767__;
  assign new_new_n24769__ = pi08 & new_new_n24763__;
  assign new_new_n24770__ = ~new_new_n24080__ & ~new_new_n24769__;
  assign new_new_n24771__ = pi08 & ~new_new_n15673__;
  assign new_new_n24772__ = new_new_n10702__ & ~new_new_n24771__;
  assign new_new_n24773__ = new_new_n15668__ & new_new_n24772__;
  assign new_new_n24774__ = ~new_new_n24770__ & ~new_new_n24773__;
  assign new_new_n24775__ = ~new_new_n24768__ & new_new_n24774__;
  assign new_new_n24776__ = new_new_n12850__ & new_new_n15656__;
  assign new_new_n24777__ = new_new_n11471__ & ~new_new_n15661__;
  assign new_new_n24778__ = new_new_n11475__ & new_new_n15643__;
  assign new_new_n24779__ = ~new_new_n24777__ & ~new_new_n24778__;
  assign new_new_n24780__ = ~new_new_n24776__ & new_new_n24779__;
  assign new_new_n24781__ = pi05 & ~new_new_n24780__;
  assign new_new_n24782__ = new_new_n12856__ & new_new_n15687__;
  assign new_new_n24783__ = new_new_n11469__ & new_new_n15687__;
  assign new_new_n24784__ = ~pi05 & ~new_new_n24783__;
  assign new_new_n24785__ = ~new_new_n24782__ & ~new_new_n24784__;
  assign new_new_n24786__ = new_new_n24780__ & ~new_new_n24785__;
  assign new_new_n24787__ = ~new_new_n24781__ & ~new_new_n24786__;
  assign new_new_n24788__ = new_new_n11468__ & ~new_new_n15673__;
  assign new_new_n24789__ = new_new_n11469__ & ~new_new_n20628__;
  assign new_new_n24790__ = ~new_new_n24788__ & ~new_new_n24789__;
  assign new_new_n24791__ = new_new_n12832__ & new_new_n15668__;
  assign new_new_n24792__ = new_new_n11475__ & ~new_new_n15661__;
  assign new_new_n24793__ = new_new_n11478__ & new_new_n20176__;
  assign new_new_n24794__ = ~new_new_n15643__ & ~new_new_n24793__;
  assign new_new_n24795__ = new_new_n11478__ & new_new_n21085__;
  assign new_new_n24796__ = ~new_new_n11482__ & ~new_new_n24794__;
  assign new_new_n24797__ = ~new_new_n24795__ & new_new_n24796__;
  assign new_new_n24798__ = ~new_new_n24791__ & ~new_new_n24792__;
  assign new_new_n24799__ = ~new_new_n24797__ & new_new_n24798__;
  assign new_new_n24800__ = pi05 & new_new_n24799__;
  assign new_new_n24801__ = new_new_n11471__ & ~new_new_n15673__;
  assign new_new_n24802__ = new_new_n13069__ & new_new_n15679__;
  assign new_new_n24803__ = new_new_n13082__ & ~new_new_n24802__;
  assign new_new_n24804__ = new_new_n15668__ & ~new_new_n24803__;
  assign new_new_n24805__ = new_new_n11478__ & new_new_n20195__;
  assign new_new_n24806__ = ~new_new_n11482__ & ~new_new_n15661__;
  assign new_new_n24807__ = ~new_new_n24805__ & new_new_n24806__;
  assign new_new_n24808__ = ~new_new_n24801__ & ~new_new_n24807__;
  assign new_new_n24809__ = ~new_new_n24804__ & new_new_n24808__;
  assign new_new_n24810__ = new_new_n24790__ & new_new_n24809__;
  assign new_new_n24811__ = new_new_n24800__ & new_new_n24810__;
  assign new_new_n24812__ = pi06 & ~new_new_n24799__;
  assign new_new_n24813__ = ~new_new_n24800__ & ~new_new_n24812__;
  assign new_new_n24814__ = ~new_new_n9701__ & ~new_new_n15673__;
  assign new_new_n24815__ = ~new_new_n24813__ & new_new_n24814__;
  assign new_new_n24816__ = ~new_new_n24811__ & ~new_new_n24815__;
  assign new_new_n24817__ = new_new_n24787__ & ~new_new_n24816__;
  assign new_new_n24818__ = ~new_new_n24787__ & new_new_n24816__;
  assign new_new_n24819__ = new_new_n10694__ & new_new_n15668__;
  assign new_new_n24820__ = new_new_n15673__ & ~new_new_n24819__;
  assign new_new_n24821__ = new_new_n10700__ & new_new_n15674__;
  assign new_new_n24822__ = ~new_new_n9697__ & new_new_n15668__;
  assign new_new_n24823__ = new_new_n10701__ & ~new_new_n24822__;
  assign new_new_n24824__ = ~new_new_n17566__ & ~new_new_n24820__;
  assign new_new_n24825__ = ~new_new_n24821__ & ~new_new_n24823__;
  assign new_new_n24826__ = new_new_n24824__ & new_new_n24825__;
  assign new_new_n24827__ = ~new_new_n24818__ & new_new_n24826__;
  assign new_new_n24828__ = ~new_new_n24817__ & ~new_new_n24827__;
  assign new_new_n24829__ = new_new_n24775__ & new_new_n24828__;
  assign new_new_n24830__ = new_new_n12850__ & ~new_new_n15710__;
  assign new_new_n24831__ = new_new_n11471__ & new_new_n15643__;
  assign new_new_n24832__ = new_new_n11475__ & new_new_n15656__;
  assign new_new_n24833__ = ~new_new_n24831__ & ~new_new_n24832__;
  assign new_new_n24834__ = ~new_new_n24830__ & new_new_n24833__;
  assign new_new_n24835__ = ~pi05 & ~new_new_n24834__;
  assign new_new_n24836__ = new_new_n12873__ & ~new_new_n19466__;
  assign new_new_n24837__ = new_new_n11469__ & ~new_new_n19466__;
  assign new_new_n24838__ = pi05 & ~new_new_n24837__;
  assign new_new_n24839__ = ~new_new_n24836__ & ~new_new_n24838__;
  assign new_new_n24840__ = new_new_n24834__ & ~new_new_n24839__;
  assign new_new_n24841__ = ~new_new_n24835__ & ~new_new_n24840__;
  assign new_new_n24842__ = ~new_new_n24775__ & ~new_new_n24828__;
  assign new_new_n24843__ = new_new_n24841__ & ~new_new_n24842__;
  assign new_new_n24844__ = ~new_new_n24829__ & ~new_new_n24843__;
  assign new_new_n24845__ = ~new_new_n24762__ & new_new_n24844__;
  assign new_new_n24846__ = new_new_n24762__ & ~new_new_n24844__;
  assign new_new_n24847__ = new_new_n24070__ & new_new_n24082__;
  assign new_new_n24848__ = ~new_new_n24069__ & ~new_new_n24847__;
  assign new_new_n24849__ = new_new_n24083__ & ~new_new_n24848__;
  assign new_new_n24850__ = ~new_new_n24083__ & new_new_n24848__;
  assign new_new_n24851__ = ~new_new_n24849__ & ~new_new_n24850__;
  assign new_new_n24852__ = ~new_new_n24846__ & new_new_n24851__;
  assign new_new_n24853__ = ~new_new_n24845__ & ~new_new_n24852__;
  assign new_new_n24854__ = ~new_new_n24751__ & new_new_n24853__;
  assign new_new_n24855__ = new_new_n24751__ & ~new_new_n24853__;
  assign new_new_n24856__ = new_new_n12850__ & ~new_new_n15582__;
  assign new_new_n24857__ = new_new_n11475__ & ~new_new_n15647__;
  assign new_new_n24858__ = new_new_n12832__ & ~new_new_n15710__;
  assign new_new_n24859__ = new_new_n13069__ & ~new_new_n15736__;
  assign new_new_n24860__ = ~new_new_n24857__ & ~new_new_n24858__;
  assign new_new_n24861__ = ~new_new_n24856__ & new_new_n24860__;
  assign new_new_n24862__ = ~new_new_n24859__ & new_new_n24861__;
  assign new_new_n24863__ = ~pi05 & ~new_new_n24862__;
  assign new_new_n24864__ = pi05 & new_new_n24862__;
  assign new_new_n24865__ = ~new_new_n24863__ & ~new_new_n24864__;
  assign new_new_n24866__ = ~new_new_n24855__ & new_new_n24865__;
  assign new_new_n24867__ = ~new_new_n24854__ & ~new_new_n24866__;
  assign new_new_n24868__ = new_new_n24747__ & new_new_n24867__;
  assign new_new_n24869__ = ~pi05 & new_new_n24732__;
  assign new_new_n24870__ = pi05 & ~new_new_n24732__;
  assign new_new_n24871__ = ~new_new_n24869__ & ~new_new_n24870__;
  assign new_new_n24872__ = new_new_n24742__ & new_new_n24871__;
  assign new_new_n24873__ = ~new_new_n24743__ & ~new_new_n24868__;
  assign new_new_n24874__ = ~new_new_n24872__ & new_new_n24873__;
  assign new_new_n24875__ = new_new_n24725__ & new_new_n24871__;
  assign new_new_n24876__ = ~new_new_n24747__ & ~new_new_n24867__;
  assign new_new_n24877__ = ~new_new_n24725__ & ~new_new_n24871__;
  assign new_new_n24878__ = ~new_new_n24876__ & ~new_new_n24877__;
  assign new_new_n24879__ = ~new_new_n24875__ & ~new_new_n24878__;
  assign new_new_n24880__ = ~new_new_n24874__ & ~new_new_n24879__;
  assign new_new_n24881__ = ~new_new_n24712__ & new_new_n24880__;
  assign new_new_n24882__ = new_new_n24712__ & ~new_new_n24880__;
  assign new_new_n24883__ = new_new_n12850__ & ~new_new_n15615__;
  assign new_new_n24884__ = new_new_n11475__ & new_new_n15743__;
  assign new_new_n24885__ = new_new_n11471__ & ~new_new_n15638__;
  assign new_new_n24886__ = new_new_n13069__ & new_new_n19005__;
  assign new_new_n24887__ = ~new_new_n24884__ & ~new_new_n24885__;
  assign new_new_n24888__ = ~new_new_n24883__ & new_new_n24887__;
  assign new_new_n24889__ = ~new_new_n24886__ & new_new_n24888__;
  assign new_new_n24890__ = pi05 & ~new_new_n24889__;
  assign new_new_n24891__ = ~pi05 & new_new_n24889__;
  assign new_new_n24892__ = ~new_new_n24890__ & ~new_new_n24891__;
  assign new_new_n24893__ = ~new_new_n24882__ & new_new_n24892__;
  assign new_new_n24894__ = ~new_new_n24881__ & ~new_new_n24893__;
  assign new_new_n24895__ = ~new_new_n24708__ & ~new_new_n24894__;
  assign new_new_n24896__ = new_new_n24708__ & new_new_n24894__;
  assign new_new_n24897__ = new_new_n11471__ & new_new_n15743__;
  assign new_new_n24898__ = new_new_n11475__ & ~new_new_n15615__;
  assign new_new_n24899__ = ~new_new_n11478__ & ~new_new_n15564__;
  assign new_new_n24900__ = new_new_n11478__ & ~new_new_n18512__;
  assign new_new_n24901__ = ~new_new_n11482__ & ~new_new_n24899__;
  assign new_new_n24902__ = ~new_new_n24900__ & new_new_n24901__;
  assign new_new_n24903__ = ~new_new_n24897__ & ~new_new_n24898__;
  assign new_new_n24904__ = ~new_new_n24902__ & new_new_n24903__;
  assign new_new_n24905__ = pi05 & ~new_new_n24904__;
  assign new_new_n24906__ = ~pi05 & new_new_n24904__;
  assign new_new_n24907__ = ~new_new_n24905__ & ~new_new_n24906__;
  assign new_new_n24908__ = ~new_new_n24896__ & new_new_n24907__;
  assign new_new_n24909__ = ~new_new_n24895__ & ~new_new_n24908__;
  assign new_new_n24910__ = ~new_new_n24170__ & ~new_new_n24171__;
  assign new_new_n24911__ = ~new_new_n24181__ & new_new_n24910__;
  assign new_new_n24912__ = new_new_n24181__ & ~new_new_n24910__;
  assign new_new_n24913__ = ~new_new_n24911__ & ~new_new_n24912__;
  assign new_new_n24914__ = new_new_n24909__ & new_new_n24913__;
  assign new_new_n24915__ = ~new_new_n24909__ & ~new_new_n24913__;
  assign new_new_n24916__ = new_new_n12850__ & new_new_n15572__;
  assign new_new_n24917__ = new_new_n11475__ & new_new_n15564__;
  assign new_new_n24918__ = new_new_n11471__ & ~new_new_n15615__;
  assign new_new_n24919__ = new_new_n13069__ & ~new_new_n20114__;
  assign new_new_n24920__ = ~new_new_n24917__ & ~new_new_n24918__;
  assign new_new_n24921__ = ~new_new_n24916__ & new_new_n24920__;
  assign new_new_n24922__ = ~new_new_n24919__ & new_new_n24921__;
  assign new_new_n24923__ = pi05 & ~new_new_n24922__;
  assign new_new_n24924__ = ~pi05 & new_new_n24922__;
  assign new_new_n24925__ = ~new_new_n24923__ & ~new_new_n24924__;
  assign new_new_n24926__ = ~new_new_n24915__ & ~new_new_n24925__;
  assign new_new_n24927__ = ~new_new_n24914__ & ~new_new_n24926__;
  assign new_new_n24928__ = ~new_new_n24704__ & new_new_n24927__;
  assign new_new_n24929__ = new_new_n24704__ & ~new_new_n24927__;
  assign new_new_n24930__ = ~new_new_n24184__ & ~new_new_n24185__;
  assign new_new_n24931__ = ~new_new_n24197__ & new_new_n24930__;
  assign new_new_n24932__ = new_new_n24197__ & ~new_new_n24930__;
  assign new_new_n24933__ = ~new_new_n24931__ & ~new_new_n24932__;
  assign new_new_n24934__ = ~new_new_n24929__ & new_new_n24933__;
  assign new_new_n24935__ = ~new_new_n24928__ & ~new_new_n24934__;
  assign new_new_n24936__ = ~new_new_n24689__ & new_new_n24935__;
  assign new_new_n24937__ = new_new_n24689__ & ~new_new_n24935__;
  assign new_new_n24938__ = ~new_new_n24202__ & ~new_new_n24212__;
  assign new_new_n24939__ = ~new_new_n24213__ & ~new_new_n24938__;
  assign new_new_n24940__ = ~new_new_n24937__ & ~new_new_n24939__;
  assign new_new_n24941__ = ~new_new_n24936__ & ~new_new_n24940__;
  assign new_new_n24942__ = ~new_new_n24219__ & ~new_new_n24220__;
  assign new_new_n24943__ = ~new_new_n24230__ & new_new_n24942__;
  assign new_new_n24944__ = new_new_n24230__ & ~new_new_n24942__;
  assign new_new_n24945__ = ~new_new_n24943__ & ~new_new_n24944__;
  assign new_new_n24946__ = ~new_new_n24941__ & ~new_new_n24945__;
  assign new_new_n24947__ = new_new_n24941__ & new_new_n24945__;
  assign new_new_n24948__ = new_new_n12850__ & ~new_new_n15533__;
  assign new_new_n24949__ = new_new_n11475__ & new_new_n15767__;
  assign new_new_n24950__ = new_new_n11471__ & new_new_n15560__;
  assign new_new_n24951__ = new_new_n13069__ & new_new_n19893__;
  assign new_new_n24952__ = ~new_new_n24949__ & ~new_new_n24950__;
  assign new_new_n24953__ = ~new_new_n24948__ & new_new_n24952__;
  assign new_new_n24954__ = ~new_new_n24951__ & new_new_n24953__;
  assign new_new_n24955__ = pi05 & new_new_n24954__;
  assign new_new_n24956__ = ~pi05 & ~new_new_n24954__;
  assign new_new_n24957__ = ~new_new_n24955__ & ~new_new_n24956__;
  assign new_new_n24958__ = ~new_new_n24947__ & new_new_n24957__;
  assign new_new_n24959__ = ~new_new_n24946__ & ~new_new_n24958__;
  assign new_new_n24960__ = ~new_new_n24677__ & new_new_n24959__;
  assign new_new_n24961__ = new_new_n24677__ & ~new_new_n24959__;
  assign new_new_n24962__ = new_new_n12850__ & new_new_n15520__;
  assign new_new_n24963__ = new_new_n11475__ & ~new_new_n15533__;
  assign new_new_n24964__ = new_new_n11471__ & new_new_n15767__;
  assign new_new_n24965__ = new_new_n13069__ & new_new_n19731__;
  assign new_new_n24966__ = ~new_new_n24963__ & ~new_new_n24964__;
  assign new_new_n24967__ = ~new_new_n24962__ & new_new_n24966__;
  assign new_new_n24968__ = ~new_new_n24965__ & new_new_n24967__;
  assign new_new_n24969__ = ~pi05 & ~new_new_n24968__;
  assign new_new_n24970__ = pi05 & new_new_n24968__;
  assign new_new_n24971__ = ~new_new_n24969__ & ~new_new_n24970__;
  assign new_new_n24972__ = ~new_new_n24961__ & ~new_new_n24971__;
  assign new_new_n24973__ = ~new_new_n24960__ & ~new_new_n24972__;
  assign new_new_n24974__ = new_new_n24673__ & ~new_new_n24973__;
  assign new_new_n24975__ = ~new_new_n24673__ & new_new_n24973__;
  assign new_new_n24976__ = ~new_new_n24262__ & ~new_new_n24277__;
  assign new_new_n24977__ = new_new_n24648__ & ~new_new_n24976__;
  assign new_new_n24978__ = ~new_new_n24648__ & new_new_n24976__;
  assign new_new_n24979__ = ~new_new_n24977__ & ~new_new_n24978__;
  assign new_new_n24980__ = ~new_new_n24975__ & new_new_n24979__;
  assign new_new_n24981__ = ~new_new_n24974__ & ~new_new_n24980__;
  assign new_new_n24982__ = new_new_n24657__ & ~new_new_n24981__;
  assign new_new_n24983__ = ~new_new_n24657__ & new_new_n24981__;
  assign new_new_n24984__ = new_new_n11471__ & new_new_n15520__;
  assign new_new_n24985__ = new_new_n11475__ & new_new_n15524__;
  assign new_new_n24986__ = new_new_n12850__ & ~new_new_n15487__;
  assign new_new_n24987__ = ~new_new_n24984__ & ~new_new_n24985__;
  assign new_new_n24988__ = ~new_new_n24986__ & new_new_n24987__;
  assign new_new_n24989__ = ~pi05 & ~new_new_n24988__;
  assign new_new_n24990__ = new_new_n12873__ & new_new_n17587__;
  assign new_new_n24991__ = new_new_n11469__ & new_new_n17587__;
  assign new_new_n24992__ = pi05 & ~new_new_n24991__;
  assign new_new_n24993__ = ~new_new_n24990__ & ~new_new_n24992__;
  assign new_new_n24994__ = new_new_n24988__ & ~new_new_n24993__;
  assign new_new_n24995__ = ~new_new_n24989__ & ~new_new_n24994__;
  assign new_new_n24996__ = ~new_new_n24983__ & ~new_new_n24995__;
  assign new_new_n24997__ = ~new_new_n24982__ & ~new_new_n24996__;
  assign new_new_n24998__ = ~new_new_n24639__ & ~new_new_n24997__;
  assign new_new_n24999__ = ~new_new_n24638__ & ~new_new_n24998__;
  assign new_new_n25000__ = new_new_n24621__ & ~new_new_n24999__;
  assign new_new_n25001__ = ~new_new_n24621__ & new_new_n24999__;
  assign new_new_n25002__ = ~new_new_n24317__ & ~new_new_n24319__;
  assign new_new_n25003__ = new_new_n24008__ & ~new_new_n25002__;
  assign new_new_n25004__ = ~new_new_n24008__ & new_new_n25002__;
  assign new_new_n25005__ = ~new_new_n25003__ & ~new_new_n25004__;
  assign new_new_n25006__ = ~new_new_n25001__ & new_new_n25005__;
  assign new_new_n25007__ = ~new_new_n25000__ & ~new_new_n25006__;
  assign new_new_n25008__ = ~new_new_n24609__ & ~new_new_n25007__;
  assign new_new_n25009__ = new_new_n24609__ & new_new_n25007__;
  assign new_new_n25010__ = ~new_new_n24333__ & ~new_new_n24334__;
  assign new_new_n25011__ = ~new_new_n24338__ & new_new_n25010__;
  assign new_new_n25012__ = new_new_n24338__ & ~new_new_n25010__;
  assign new_new_n25013__ = ~new_new_n25011__ & ~new_new_n25012__;
  assign new_new_n25014__ = ~new_new_n25009__ & ~new_new_n25013__;
  assign new_new_n25015__ = ~new_new_n25008__ & ~new_new_n25014__;
  assign new_new_n25016__ = ~new_new_n23991__ & ~new_new_n23992__;
  assign new_new_n25017__ = ~new_new_n24340__ & new_new_n25016__;
  assign new_new_n25018__ = new_new_n24340__ & ~new_new_n25016__;
  assign new_new_n25019__ = ~new_new_n25017__ & ~new_new_n25018__;
  assign new_new_n25020__ = new_new_n25015__ & ~new_new_n25019__;
  assign new_new_n25021__ = ~new_new_n25015__ & new_new_n25019__;
  assign new_new_n25022__ = new_new_n12850__ & ~new_new_n15439__;
  assign new_new_n25023__ = new_new_n13111__ & ~new_new_n15471__;
  assign new_new_n25024__ = new_new_n11469__ & ~new_new_n17240__;
  assign new_new_n25025__ = ~new_new_n25023__ & ~new_new_n25024__;
  assign new_new_n25026__ = new_new_n11478__ & ~new_new_n25025__;
  assign new_new_n25027__ = new_new_n11475__ & new_new_n15464__;
  assign new_new_n25028__ = ~new_new_n25022__ & ~new_new_n25027__;
  assign new_new_n25029__ = ~new_new_n25026__ & new_new_n25028__;
  assign new_new_n25030__ = pi05 & ~new_new_n25029__;
  assign new_new_n25031__ = ~pi05 & new_new_n25029__;
  assign new_new_n25032__ = ~new_new_n25030__ & ~new_new_n25031__;
  assign new_new_n25033__ = ~new_new_n25021__ & ~new_new_n25032__;
  assign new_new_n25034__ = ~new_new_n25020__ & ~new_new_n25033__;
  assign new_new_n25035__ = ~new_new_n24596__ & ~new_new_n25034__;
  assign new_new_n25036__ = new_new_n24596__ & new_new_n25034__;
  assign new_new_n25037__ = new_new_n12850__ & ~new_new_n15432__;
  assign new_new_n25038__ = new_new_n11471__ & new_new_n15464__;
  assign new_new_n25039__ = new_new_n11475__ & ~new_new_n15439__;
  assign new_new_n25040__ = ~new_new_n25038__ & ~new_new_n25039__;
  assign new_new_n25041__ = ~new_new_n25037__ & new_new_n25040__;
  assign new_new_n25042__ = pi05 & ~new_new_n25041__;
  assign new_new_n25043__ = new_new_n12856__ & new_new_n17204__;
  assign new_new_n25044__ = new_new_n11469__ & new_new_n17204__;
  assign new_new_n25045__ = ~pi05 & ~new_new_n25044__;
  assign new_new_n25046__ = ~new_new_n25043__ & ~new_new_n25045__;
  assign new_new_n25047__ = new_new_n25041__ & ~new_new_n25046__;
  assign new_new_n25048__ = ~new_new_n25042__ & ~new_new_n25047__;
  assign new_new_n25049__ = ~new_new_n25036__ & ~new_new_n25048__;
  assign new_new_n25050__ = ~new_new_n25035__ & ~new_new_n25049__;
  assign new_new_n25051__ = ~new_new_n24592__ & ~new_new_n25050__;
  assign new_new_n25052__ = ~new_new_n24591__ & ~new_new_n25051__;
  assign new_new_n25053__ = ~new_new_n24369__ & ~new_new_n24370__;
  assign new_new_n25054__ = ~new_new_n24374__ & new_new_n25053__;
  assign new_new_n25055__ = new_new_n24374__ & ~new_new_n25053__;
  assign new_new_n25056__ = ~new_new_n25054__ & ~new_new_n25055__;
  assign new_new_n25057__ = ~new_new_n25052__ & ~new_new_n25056__;
  assign new_new_n25058__ = new_new_n25052__ & new_new_n25056__;
  assign new_new_n25059__ = new_new_n11475__ & ~new_new_n15362__;
  assign new_new_n25060__ = new_new_n11471__ & ~new_new_n15432__;
  assign new_new_n25061__ = ~new_new_n11478__ & ~new_new_n15390__;
  assign new_new_n25062__ = new_new_n11478__ & new_new_n22497__;
  assign new_new_n25063__ = new_new_n11469__ & ~new_new_n25061__;
  assign new_new_n25064__ = ~new_new_n17918__ & new_new_n25063__;
  assign new_new_n25065__ = ~new_new_n25062__ & new_new_n25064__;
  assign new_new_n25066__ = ~new_new_n25059__ & ~new_new_n25060__;
  assign new_new_n25067__ = ~new_new_n25065__ & new_new_n25066__;
  assign new_new_n25068__ = pi05 & ~new_new_n25067__;
  assign new_new_n25069__ = ~pi05 & new_new_n25067__;
  assign new_new_n25070__ = ~new_new_n25068__ & ~new_new_n25069__;
  assign new_new_n25071__ = ~new_new_n25058__ & ~new_new_n25070__;
  assign new_new_n25072__ = ~new_new_n25057__ & ~new_new_n25071__;
  assign new_new_n25073__ = ~new_new_n24570__ & ~new_new_n25072__;
  assign new_new_n25074__ = pi05 & ~new_new_n25073__;
  assign new_new_n25075__ = ~new_new_n24575__ & ~new_new_n25074__;
  assign new_new_n25076__ = new_new_n12850__ & ~new_new_n15349__;
  assign new_new_n25077__ = new_new_n11475__ & ~new_new_n15398__;
  assign new_new_n25078__ = new_new_n11471__ & new_new_n15390__;
  assign new_new_n25079__ = new_new_n13069__ & ~new_new_n17180__;
  assign new_new_n25080__ = ~new_new_n25077__ & ~new_new_n25078__;
  assign new_new_n25081__ = ~new_new_n25076__ & new_new_n25080__;
  assign new_new_n25082__ = ~new_new_n25079__ & new_new_n25081__;
  assign new_new_n25083__ = ~new_new_n25075__ & new_new_n25082__;
  assign new_new_n25084__ = pi05 & ~new_new_n24570__;
  assign new_new_n25085__ = new_new_n24570__ & ~new_new_n24574__;
  assign new_new_n25086__ = ~new_new_n25084__ & ~new_new_n25085__;
  assign new_new_n25087__ = ~new_new_n25082__ & new_new_n25086__;
  assign new_new_n25088__ = ~pi05 & ~new_new_n25082__;
  assign new_new_n25089__ = ~new_new_n24574__ & ~new_new_n25088__;
  assign new_new_n25090__ = new_new_n25072__ & ~new_new_n25089__;
  assign new_new_n25091__ = ~new_new_n25087__ & ~new_new_n25090__;
  assign new_new_n25092__ = ~new_new_n25083__ & new_new_n25091__;
  assign new_new_n25093__ = ~new_new_n24377__ & ~new_new_n24378__;
  assign new_new_n25094__ = ~new_new_n24382__ & new_new_n25093__;
  assign new_new_n25095__ = new_new_n24382__ & ~new_new_n25093__;
  assign new_new_n25096__ = ~new_new_n25094__ & ~new_new_n25095__;
  assign new_new_n25097__ = ~new_new_n25092__ & new_new_n25096__;
  assign new_new_n25098__ = pi05 & new_new_n24574__;
  assign new_new_n25099__ = pi05 & new_new_n24570__;
  assign new_new_n25100__ = ~new_new_n24575__ & ~new_new_n25099__;
  assign new_new_n25101__ = new_new_n25072__ & ~new_new_n25100__;
  assign new_new_n25102__ = ~new_new_n25098__ & ~new_new_n25101__;
  assign new_new_n25103__ = new_new_n25082__ & ~new_new_n25102__;
  assign new_new_n25104__ = ~pi05 & new_new_n24574__;
  assign new_new_n25105__ = new_new_n25072__ & new_new_n25086__;
  assign new_new_n25106__ = ~new_new_n25104__ & ~new_new_n25105__;
  assign new_new_n25107__ = ~new_new_n25082__ & ~new_new_n25106__;
  assign new_new_n25108__ = ~new_new_n25103__ & ~new_new_n25107__;
  assign new_new_n25109__ = ~new_new_n25097__ & new_new_n25108__;
  assign new_new_n25110__ = ~new_new_n24399__ & ~new_new_n24400__;
  assign new_new_n25111__ = new_new_n24404__ & new_new_n25110__;
  assign new_new_n25112__ = ~new_new_n24404__ & ~new_new_n25110__;
  assign new_new_n25113__ = ~new_new_n25111__ & ~new_new_n25112__;
  assign new_new_n25114__ = new_new_n25109__ & ~new_new_n25113__;
  assign new_new_n25115__ = ~new_new_n25109__ & new_new_n25113__;
  assign new_new_n25116__ = new_new_n13069__ & new_new_n16458__;
  assign new_new_n25117__ = new_new_n11471__ & ~new_new_n15398__;
  assign new_new_n25118__ = new_new_n11475__ & ~new_new_n15349__;
  assign new_new_n25119__ = new_new_n12850__ & ~new_new_n15321__;
  assign new_new_n25120__ = ~new_new_n25117__ & ~new_new_n25118__;
  assign new_new_n25121__ = ~new_new_n25119__ & new_new_n25120__;
  assign new_new_n25122__ = ~new_new_n25116__ & new_new_n25121__;
  assign new_new_n25123__ = pi05 & ~new_new_n25122__;
  assign new_new_n25124__ = ~pi05 & new_new_n25122__;
  assign new_new_n25125__ = ~new_new_n25123__ & ~new_new_n25124__;
  assign new_new_n25126__ = ~new_new_n25115__ & ~new_new_n25125__;
  assign new_new_n25127__ = ~new_new_n25114__ & ~new_new_n25126__;
  assign new_new_n25128__ = new_new_n12850__ & ~new_new_n15273__;
  assign new_new_n25129__ = new_new_n11471__ & ~new_new_n15349__;
  assign new_new_n25130__ = new_new_n11475__ & ~new_new_n15321__;
  assign new_new_n25131__ = ~new_new_n25129__ & ~new_new_n25130__;
  assign new_new_n25132__ = ~new_new_n25128__ & new_new_n25131__;
  assign new_new_n25133__ = pi05 & ~new_new_n25132__;
  assign new_new_n25134__ = new_new_n12856__ & ~new_new_n17103__;
  assign new_new_n25135__ = new_new_n11469__ & ~new_new_n17103__;
  assign new_new_n25136__ = ~pi05 & ~new_new_n25135__;
  assign new_new_n25137__ = ~new_new_n25134__ & ~new_new_n25136__;
  assign new_new_n25138__ = new_new_n25132__ & ~new_new_n25137__;
  assign new_new_n25139__ = ~new_new_n25133__ & ~new_new_n25138__;
  assign new_new_n25140__ = ~new_new_n23914__ & ~new_new_n24407__;
  assign new_new_n25141__ = new_new_n24406__ & ~new_new_n25140__;
  assign new_new_n25142__ = ~new_new_n24406__ & new_new_n25140__;
  assign new_new_n25143__ = ~new_new_n25141__ & ~new_new_n25142__;
  assign new_new_n25144__ = new_new_n25139__ & new_new_n25143__;
  assign new_new_n25145__ = ~new_new_n25127__ & ~new_new_n25144__;
  assign new_new_n25146__ = ~new_new_n25139__ & ~new_new_n25143__;
  assign new_new_n25147__ = ~new_new_n25145__ & ~new_new_n25146__;
  assign new_new_n25148__ = ~new_new_n24561__ & ~new_new_n25147__;
  assign new_new_n25149__ = ~new_new_n24560__ & ~new_new_n25148__;
  assign new_new_n25150__ = ~new_new_n24412__ & ~new_new_n24413__;
  assign new_new_n25151__ = ~new_new_n23732__ & new_new_n24414__;
  assign new_new_n25152__ = new_new_n23732__ & ~new_new_n24414__;
  assign new_new_n25153__ = ~new_new_n25151__ & ~new_new_n25152__;
  assign new_new_n25154__ = new_new_n25150__ & new_new_n25153__;
  assign new_new_n25155__ = ~new_new_n25150__ & ~new_new_n25153__;
  assign new_new_n25156__ = ~new_new_n25154__ & ~new_new_n25155__;
  assign new_new_n25157__ = ~new_new_n25149__ & ~new_new_n25156__;
  assign new_new_n25158__ = new_new_n12850__ & ~new_new_n15314__;
  assign new_new_n25159__ = new_new_n11471__ & ~new_new_n15273__;
  assign new_new_n25160__ = new_new_n11475__ & new_new_n15285__;
  assign new_new_n25161__ = ~new_new_n25159__ & ~new_new_n25160__;
  assign new_new_n25162__ = ~new_new_n25158__ & new_new_n25161__;
  assign new_new_n25163__ = pi05 & ~new_new_n25162__;
  assign new_new_n25164__ = new_new_n12856__ & new_new_n17140__;
  assign new_new_n25165__ = new_new_n11469__ & new_new_n17140__;
  assign new_new_n25166__ = ~pi05 & ~new_new_n25165__;
  assign new_new_n25167__ = ~new_new_n25164__ & ~new_new_n25166__;
  assign new_new_n25168__ = new_new_n25162__ & ~new_new_n25167__;
  assign new_new_n25169__ = ~new_new_n25163__ & ~new_new_n25168__;
  assign new_new_n25170__ = ~new_new_n25157__ & new_new_n25169__;
  assign new_new_n25171__ = new_new_n11475__ & ~new_new_n15314__;
  assign new_new_n25172__ = new_new_n11471__ & new_new_n15285__;
  assign new_new_n25173__ = new_new_n12850__ & ~new_new_n15248__;
  assign new_new_n25174__ = ~new_new_n25171__ & ~new_new_n25172__;
  assign new_new_n25175__ = ~new_new_n25173__ & new_new_n25174__;
  assign new_new_n25176__ = ~new_new_n11482__ & new_new_n16725__;
  assign new_new_n25177__ = ~new_new_n24420__ & ~new_new_n24421__;
  assign new_new_n25178__ = new_new_n24431__ & new_new_n25177__;
  assign new_new_n25179__ = ~new_new_n24431__ & ~new_new_n25177__;
  assign new_new_n25180__ = ~new_new_n25178__ & ~new_new_n25179__;
  assign new_new_n25181__ = pi04 & ~new_new_n25180__;
  assign new_new_n25182__ = ~pi04 & new_new_n25180__;
  assign new_new_n25183__ = ~new_new_n25181__ & ~new_new_n25182__;
  assign new_new_n25184__ = new_new_n25176__ & ~new_new_n25183__;
  assign new_new_n25185__ = pi05 & new_new_n25180__;
  assign new_new_n25186__ = ~pi05 & ~new_new_n25180__;
  assign new_new_n25187__ = ~new_new_n25185__ & ~new_new_n25186__;
  assign new_new_n25188__ = ~new_new_n25176__ & new_new_n25187__;
  assign new_new_n25189__ = ~new_new_n25184__ & ~new_new_n25188__;
  assign new_new_n25190__ = new_new_n25175__ & ~new_new_n25189__;
  assign new_new_n25191__ = ~new_new_n25175__ & ~new_new_n25187__;
  assign new_new_n25192__ = ~new_new_n25190__ & ~new_new_n25191__;
  assign new_new_n25193__ = new_new_n25170__ & ~new_new_n25192__;
  assign new_new_n25194__ = new_new_n25180__ & new_new_n25192__;
  assign new_new_n25195__ = new_new_n25149__ & new_new_n25156__;
  assign new_new_n25196__ = ~new_new_n25192__ & new_new_n25195__;
  assign new_new_n25197__ = ~new_new_n25193__ & ~new_new_n25194__;
  assign new_new_n25198__ = ~new_new_n25196__ & new_new_n25197__;
  assign new_new_n25199__ = ~new_new_n24543__ & new_new_n25198__;
  assign new_new_n25200__ = new_new_n24543__ & ~new_new_n25198__;
  assign new_new_n25201__ = new_new_n12850__ & new_new_n15244__;
  assign new_new_n25202__ = new_new_n13111__ & ~new_new_n15314__;
  assign new_new_n25203__ = new_new_n11469__ & new_new_n16378__;
  assign new_new_n25204__ = ~new_new_n25202__ & ~new_new_n25203__;
  assign new_new_n25205__ = new_new_n11478__ & ~new_new_n25204__;
  assign new_new_n25206__ = new_new_n11475__ & ~new_new_n15248__;
  assign new_new_n25207__ = ~new_new_n25201__ & ~new_new_n25206__;
  assign new_new_n25208__ = ~new_new_n25205__ & new_new_n25207__;
  assign new_new_n25209__ = pi05 & ~new_new_n25208__;
  assign new_new_n25210__ = ~pi05 & new_new_n25208__;
  assign new_new_n25211__ = ~new_new_n25209__ & ~new_new_n25210__;
  assign new_new_n25212__ = ~new_new_n25200__ & ~new_new_n25211__;
  assign new_new_n25213__ = ~new_new_n25199__ & ~new_new_n25212__;
  assign new_new_n25214__ = ~new_new_n24539__ & new_new_n25213__;
  assign new_new_n25215__ = new_new_n24539__ & ~new_new_n25213__;
  assign new_new_n25216__ = new_new_n13069__ & ~new_new_n16603__;
  assign new_new_n25217__ = new_new_n12832__ & ~new_new_n15248__;
  assign new_new_n25218__ = ~new_new_n25216__ & ~new_new_n25217__;
  assign new_new_n25219__ = new_new_n12850__ & new_new_n15237__;
  assign new_new_n25220__ = new_new_n11475__ & new_new_n15244__;
  assign new_new_n25221__ = ~new_new_n25219__ & ~new_new_n25220__;
  assign new_new_n25222__ = new_new_n25218__ & new_new_n25221__;
  assign new_new_n25223__ = pi05 & ~new_new_n25222__;
  assign new_new_n25224__ = new_new_n13082__ & ~new_new_n15237__;
  assign new_new_n25225__ = new_new_n12850__ & ~new_new_n25224__;
  assign new_new_n25226__ = ~pi05 & ~new_new_n25220__;
  assign new_new_n25227__ = ~new_new_n25225__ & new_new_n25226__;
  assign new_new_n25228__ = new_new_n25218__ & new_new_n25227__;
  assign new_new_n25229__ = ~new_new_n25223__ & ~new_new_n25228__;
  assign new_new_n25230__ = ~new_new_n25215__ & new_new_n25229__;
  assign new_new_n25231__ = ~new_new_n25214__ & ~new_new_n25230__;
  assign new_new_n25232__ = ~new_new_n24461__ & ~new_new_n24462__;
  assign new_new_n25233__ = new_new_n24466__ & new_new_n25232__;
  assign new_new_n25234__ = ~new_new_n24466__ & ~new_new_n25232__;
  assign new_new_n25235__ = ~new_new_n25233__ & ~new_new_n25234__;
  assign new_new_n25236__ = ~new_new_n25231__ & ~new_new_n25235__;
  assign new_new_n25237__ = new_new_n25231__ & new_new_n25235__;
  assign new_new_n25238__ = new_new_n13111__ & new_new_n15244__;
  assign new_new_n25239__ = new_new_n11469__ & ~new_new_n15917__;
  assign new_new_n25240__ = ~new_new_n25238__ & ~new_new_n25239__;
  assign new_new_n25241__ = new_new_n11478__ & ~new_new_n25240__;
  assign new_new_n25242__ = new_new_n11475__ & new_new_n15237__;
  assign new_new_n25243__ = ~new_new_n25241__ & ~new_new_n25242__;
  assign new_new_n25244__ = pi05 & ~new_new_n25243__;
  assign new_new_n25245__ = new_new_n12873__ & new_new_n15905__;
  assign new_new_n25246__ = new_new_n11469__ & new_new_n15905__;
  assign new_new_n25247__ = ~pi05 & ~new_new_n25246__;
  assign new_new_n25248__ = ~new_new_n25245__ & ~new_new_n25247__;
  assign new_new_n25249__ = new_new_n25243__ & ~new_new_n25248__;
  assign new_new_n25250__ = ~new_new_n25244__ & ~new_new_n25249__;
  assign new_new_n25251__ = ~new_new_n25237__ & new_new_n25250__;
  assign new_new_n25252__ = ~new_new_n25236__ & ~new_new_n25251__;
  assign new_new_n25253__ = new_new_n24532__ & new_new_n25252__;
  assign new_new_n25254__ = ~new_new_n24532__ & ~new_new_n25252__;
  assign new_new_n25255__ = ~new_new_n25253__ & ~new_new_n25254__;
  assign new_new_n25256__ = ~new_new_n24478__ & ~new_new_n24479__;
  assign new_new_n25257__ = ~new_new_n24489__ & new_new_n25256__;
  assign new_new_n25258__ = new_new_n24489__ & ~new_new_n25256__;
  assign new_new_n25259__ = ~new_new_n25257__ & ~new_new_n25258__;
  assign new_new_n25260__ = ~new_new_n25255__ & new_new_n25259__;
  assign new_new_n25261__ = new_new_n25255__ & ~new_new_n25259__;
  assign new_new_n25262__ = ~new_new_n25260__ & ~new_new_n25261__;
  assign new_new_n25263__ = pi02 & new_new_n25262__;
  assign new_new_n25264__ = ~pi01 & ~new_new_n16630__;
  assign new_new_n25265__ = ~pi02 & ~new_new_n16056__;
  assign new_new_n25266__ = ~new_new_n16048__ & new_new_n25265__;
  assign new_new_n25267__ = ~new_new_n25264__ & ~new_new_n25266__;
  assign new_new_n25268__ = pi00 & ~new_new_n25267__;
  assign new_new_n25269__ = pi02 & new_new_n15998__;
  assign new_new_n25270__ = ~pi01 & ~new_new_n25269__;
  assign new_new_n25271__ = pi02 & new_new_n16056__;
  assign new_new_n25272__ = pi01 & ~new_new_n25265__;
  assign new_new_n25273__ = ~new_new_n25271__ & new_new_n25272__;
  assign new_new_n25274__ = ~pi00 & ~new_new_n25273__;
  assign new_new_n25275__ = ~new_new_n25270__ & new_new_n25274__;
  assign new_new_n25276__ = ~new_new_n25268__ & ~new_new_n25275__;
  assign new_new_n25277__ = ~pi02 & ~new_new_n15998__;
  assign new_new_n25278__ = ~new_new_n25269__ & ~new_new_n25277__;
  assign new_new_n25279__ = pi01 & ~new_new_n25278__;
  assign new_new_n25280__ = new_new_n12798__ & ~new_new_n15905__;
  assign new_new_n25281__ = ~new_new_n25279__ & ~new_new_n25280__;
  assign new_new_n25282__ = ~pi00 & ~new_new_n25281__;
  assign new_new_n25283__ = pi02 & ~new_new_n16051__;
  assign new_new_n25284__ = pi01 & new_new_n16051__;
  assign new_new_n25285__ = ~new_new_n16056__ & ~new_new_n25283__;
  assign new_new_n25286__ = ~new_new_n25284__ & new_new_n25285__;
  assign new_new_n25287__ = ~new_new_n25271__ & ~new_new_n25286__;
  assign new_new_n25288__ = pi00 & ~new_new_n25287__;
  assign new_new_n25289__ = ~new_new_n25282__ & ~new_new_n25288__;
  assign new_new_n25290__ = ~pi01 & ~pi02;
  assign new_new_n25291__ = pi02 & new_new_n14441__;
  assign new_new_n25292__ = ~new_new_n25290__ & ~new_new_n25291__;
  assign new_new_n25293__ = new_new_n15998__ & ~new_new_n25292__;
  assign new_new_n25294__ = ~new_new_n12798__ & ~new_new_n13508__;
  assign new_new_n25295__ = pi00 & ~new_new_n25294__;
  assign new_new_n25296__ = ~new_new_n16025__ & new_new_n25295__;
  assign new_new_n25297__ = new_new_n12798__ & new_new_n15237__;
  assign new_new_n25298__ = pi01 & new_new_n15905__;
  assign new_new_n25299__ = ~pi00 & ~new_new_n25297__;
  assign new_new_n25300__ = ~new_new_n25298__ & new_new_n25299__;
  assign new_new_n25301__ = ~new_new_n25293__ & ~new_new_n25300__;
  assign new_new_n25302__ = ~new_new_n25296__ & new_new_n25301__;
  assign new_new_n25303__ = ~pi02 & new_new_n25302__;
  assign new_new_n25304__ = pi02 & ~new_new_n25302__;
  assign new_new_n25305__ = ~new_new_n25303__ & ~new_new_n25304__;
  assign new_new_n25306__ = ~new_new_n25199__ & ~new_new_n25200__;
  assign new_new_n25307__ = ~new_new_n25211__ & new_new_n25306__;
  assign new_new_n25308__ = new_new_n25211__ & ~new_new_n25306__;
  assign new_new_n25309__ = ~new_new_n25307__ & ~new_new_n25308__;
  assign new_new_n25310__ = new_new_n25305__ & new_new_n25309__;
  assign new_new_n25311__ = new_new_n25192__ & ~new_new_n25195__;
  assign new_new_n25312__ = ~new_new_n25170__ & new_new_n25311__;
  assign new_new_n25313__ = pi02 & ~new_new_n15851__;
  assign new_new_n25314__ = pi01 & new_new_n15851__;
  assign new_new_n25315__ = ~new_new_n25313__ & ~new_new_n25314__;
  assign new_new_n25316__ = new_new_n15237__ & new_new_n25315__;
  assign new_new_n25317__ = ~new_new_n15237__ & ~new_new_n25315__;
  assign new_new_n25318__ = pi00 & ~new_new_n25316__;
  assign new_new_n25319__ = ~new_new_n25317__ & new_new_n25318__;
  assign new_new_n25320__ = ~pi02 & new_new_n15244__;
  assign new_new_n25321__ = pi01 & new_new_n25320__;
  assign new_new_n25322__ = pi01 & ~new_new_n15244__;
  assign new_new_n25323__ = ~pi01 & new_new_n15248__;
  assign new_new_n25324__ = ~new_new_n25322__ & ~new_new_n25323__;
  assign new_new_n25325__ = pi02 & ~new_new_n25324__;
  assign new_new_n25326__ = ~pi00 & ~new_new_n25321__;
  assign new_new_n25327__ = ~new_new_n25325__ & new_new_n25326__;
  assign new_new_n25328__ = ~new_new_n25319__ & ~new_new_n25327__;
  assign new_new_n25329__ = pi01 & ~new_new_n15248__;
  assign new_new_n25330__ = ~pi01 & ~new_new_n15314__;
  assign new_new_n25331__ = pi02 & ~new_new_n25330__;
  assign new_new_n25332__ = ~new_new_n25329__ & new_new_n25331__;
  assign new_new_n25333__ = new_new_n13508__ & ~new_new_n15248__;
  assign new_new_n25334__ = ~new_new_n25332__ & ~new_new_n25333__;
  assign new_new_n25335__ = ~pi00 & ~new_new_n25334__;
  assign new_new_n25336__ = ~new_new_n25320__ & ~new_new_n25322__;
  assign new_new_n25337__ = new_new_n16378__ & ~new_new_n25336__;
  assign new_new_n25338__ = ~pi02 & ~new_new_n15244__;
  assign new_new_n25339__ = pi01 & new_new_n15244__;
  assign new_new_n25340__ = ~new_new_n25338__ & ~new_new_n25339__;
  assign new_new_n25341__ = ~new_new_n16378__ & new_new_n25340__;
  assign new_new_n25342__ = ~new_new_n25337__ & ~new_new_n25341__;
  assign new_new_n25343__ = pi00 & ~new_new_n25342__;
  assign new_new_n25344__ = ~new_new_n25335__ & ~new_new_n25343__;
  assign new_new_n25345__ = ~new_new_n24560__ & ~new_new_n24561__;
  assign new_new_n25346__ = ~new_new_n25147__ & new_new_n25345__;
  assign new_new_n25347__ = new_new_n25147__ & ~new_new_n25345__;
  assign new_new_n25348__ = ~new_new_n25346__ & ~new_new_n25347__;
  assign new_new_n25349__ = ~new_new_n25344__ & ~new_new_n25348__;
  assign new_new_n25350__ = new_new_n25344__ & new_new_n25348__;
  assign new_new_n25351__ = new_new_n13508__ & new_new_n15285__;
  assign new_new_n25352__ = ~pi01 & ~new_new_n15273__;
  assign new_new_n25353__ = pi01 & new_new_n15285__;
  assign new_new_n25354__ = pi02 & ~new_new_n25352__;
  assign new_new_n25355__ = ~new_new_n25353__ & new_new_n25354__;
  assign new_new_n25356__ = ~pi00 & ~new_new_n25351__;
  assign new_new_n25357__ = ~new_new_n25355__ & new_new_n25356__;
  assign new_new_n25358__ = ~pi01 & new_new_n16082__;
  assign new_new_n25359__ = ~pi02 & ~new_new_n16082__;
  assign new_new_n25360__ = ~new_new_n25358__ & ~new_new_n25359__;
  assign new_new_n25361__ = ~new_new_n15314__ & ~new_new_n25360__;
  assign new_new_n25362__ = new_new_n15314__ & new_new_n25360__;
  assign new_new_n25363__ = pi00 & ~new_new_n25361__;
  assign new_new_n25364__ = ~new_new_n25362__ & new_new_n25363__;
  assign new_new_n25365__ = ~new_new_n25357__ & ~new_new_n25364__;
  assign new_new_n25366__ = ~new_new_n25114__ & ~new_new_n25115__;
  assign new_new_n25367__ = new_new_n25125__ & new_new_n25366__;
  assign new_new_n25368__ = ~new_new_n25125__ & ~new_new_n25366__;
  assign new_new_n25369__ = ~new_new_n25367__ & ~new_new_n25368__;
  assign new_new_n25370__ = ~new_new_n25365__ & ~new_new_n25369__;
  assign new_new_n25371__ = new_new_n25365__ & new_new_n25369__;
  assign new_new_n25372__ = ~pi01 & ~new_new_n17103__;
  assign new_new_n25373__ = ~pi02 & new_new_n17103__;
  assign new_new_n25374__ = new_new_n15273__ & ~new_new_n25372__;
  assign new_new_n25375__ = ~new_new_n25373__ & new_new_n25374__;
  assign new_new_n25376__ = pi01 & new_new_n17103__;
  assign new_new_n25377__ = pi02 & ~new_new_n17103__;
  assign new_new_n25378__ = ~new_new_n15273__ & ~new_new_n25376__;
  assign new_new_n25379__ = ~new_new_n25377__ & new_new_n25378__;
  assign new_new_n25380__ = ~new_new_n25375__ & ~new_new_n25379__;
  assign new_new_n25381__ = pi00 & ~new_new_n25380__;
  assign new_new_n25382__ = ~pi02 & ~new_new_n15321__;
  assign new_new_n25383__ = pi02 & new_new_n15321__;
  assign new_new_n25384__ = ~new_new_n25382__ & ~new_new_n25383__;
  assign new_new_n25385__ = pi01 & ~new_new_n25384__;
  assign new_new_n25386__ = new_new_n12798__ & new_new_n15349__;
  assign new_new_n25387__ = ~new_new_n25385__ & ~new_new_n25386__;
  assign new_new_n25388__ = ~pi00 & ~new_new_n25387__;
  assign new_new_n25389__ = ~new_new_n25381__ & ~new_new_n25388__;
  assign new_new_n25390__ = pi01 & ~new_new_n15349__;
  assign new_new_n25391__ = ~pi01 & ~new_new_n15398__;
  assign new_new_n25392__ = ~new_new_n25390__ & ~new_new_n25391__;
  assign new_new_n25393__ = pi02 & ~new_new_n25392__;
  assign new_new_n25394__ = ~pi02 & ~new_new_n25390__;
  assign new_new_n25395__ = ~pi00 & ~new_new_n25394__;
  assign new_new_n25396__ = ~new_new_n25393__ & new_new_n25395__;
  assign new_new_n25397__ = ~pi01 & ~new_new_n15321__;
  assign new_new_n25398__ = ~new_new_n25383__ & ~new_new_n25397__;
  assign new_new_n25399__ = ~new_new_n16458__ & new_new_n25398__;
  assign new_new_n25400__ = pi01 & new_new_n15321__;
  assign new_new_n25401__ = ~new_new_n25382__ & ~new_new_n25400__;
  assign new_new_n25402__ = new_new_n16458__ & new_new_n25401__;
  assign new_new_n25403__ = pi00 & ~new_new_n25399__;
  assign new_new_n25404__ = ~new_new_n25402__ & new_new_n25403__;
  assign new_new_n25405__ = ~new_new_n25396__ & ~new_new_n25404__;
  assign new_new_n25406__ = ~new_new_n25057__ & ~new_new_n25058__;
  assign new_new_n25407__ = new_new_n25070__ & new_new_n25406__;
  assign new_new_n25408__ = ~new_new_n25070__ & ~new_new_n25406__;
  assign new_new_n25409__ = ~new_new_n25407__ & ~new_new_n25408__;
  assign new_new_n25410__ = ~new_new_n25405__ & new_new_n25409__;
  assign new_new_n25411__ = new_new_n25405__ & ~new_new_n25409__;
  assign new_new_n25412__ = new_new_n24586__ & ~new_new_n24590__;
  assign new_new_n25413__ = ~new_new_n24586__ & new_new_n24590__;
  assign new_new_n25414__ = ~new_new_n25412__ & ~new_new_n25413__;
  assign new_new_n25415__ = new_new_n25050__ & new_new_n25414__;
  assign new_new_n25416__ = ~new_new_n25050__ & ~new_new_n25414__;
  assign new_new_n25417__ = ~new_new_n25415__ & ~new_new_n25416__;
  assign new_new_n25418__ = new_new_n13508__ & new_new_n15390__;
  assign new_new_n25419__ = pi01 & new_new_n15390__;
  assign new_new_n25420__ = ~pi01 & ~new_new_n15362__;
  assign new_new_n25421__ = pi02 & ~new_new_n25420__;
  assign new_new_n25422__ = ~new_new_n25419__ & new_new_n25421__;
  assign new_new_n25423__ = ~pi00 & ~new_new_n25418__;
  assign new_new_n25424__ = ~new_new_n25422__ & new_new_n25423__;
  assign new_new_n25425__ = pi02 & ~new_new_n16956__;
  assign new_new_n25426__ = pi01 & new_new_n16956__;
  assign new_new_n25427__ = ~new_new_n25425__ & ~new_new_n25426__;
  assign new_new_n25428__ = new_new_n15398__ & ~new_new_n25427__;
  assign new_new_n25429__ = ~new_new_n15398__ & new_new_n25427__;
  assign new_new_n25430__ = pi00 & ~new_new_n25428__;
  assign new_new_n25431__ = ~new_new_n25429__ & new_new_n25430__;
  assign new_new_n25432__ = ~new_new_n25424__ & ~new_new_n25431__;
  assign new_new_n25433__ = new_new_n13508__ & ~new_new_n15362__;
  assign new_new_n25434__ = ~pi01 & ~new_new_n15432__;
  assign new_new_n25435__ = pi01 & ~new_new_n15362__;
  assign new_new_n25436__ = pi02 & ~new_new_n25434__;
  assign new_new_n25437__ = ~new_new_n25435__ & new_new_n25436__;
  assign new_new_n25438__ = ~pi00 & ~new_new_n25433__;
  assign new_new_n25439__ = ~new_new_n25437__ & new_new_n25438__;
  assign new_new_n25440__ = pi02 & ~new_new_n15829__;
  assign new_new_n25441__ = pi01 & new_new_n15829__;
  assign new_new_n25442__ = ~new_new_n25440__ & ~new_new_n25441__;
  assign new_new_n25443__ = new_new_n15390__ & new_new_n25442__;
  assign new_new_n25444__ = ~new_new_n15390__ & ~new_new_n25442__;
  assign new_new_n25445__ = pi00 & ~new_new_n25443__;
  assign new_new_n25446__ = ~new_new_n25444__ & new_new_n25445__;
  assign new_new_n25447__ = ~new_new_n25439__ & ~new_new_n25446__;
  assign new_new_n25448__ = ~new_new_n25020__ & ~new_new_n25021__;
  assign new_new_n25449__ = new_new_n25032__ & new_new_n25448__;
  assign new_new_n25450__ = ~new_new_n25032__ & ~new_new_n25448__;
  assign new_new_n25451__ = ~new_new_n25449__ & ~new_new_n25450__;
  assign new_new_n25452__ = ~new_new_n25447__ & ~new_new_n25451__;
  assign new_new_n25453__ = new_new_n25447__ & new_new_n25451__;
  assign new_new_n25454__ = ~new_new_n25008__ & ~new_new_n25009__;
  assign new_new_n25455__ = ~new_new_n25013__ & new_new_n25454__;
  assign new_new_n25456__ = new_new_n25013__ & ~new_new_n25454__;
  assign new_new_n25457__ = ~new_new_n25455__ & ~new_new_n25456__;
  assign new_new_n25458__ = ~new_new_n25000__ & ~new_new_n25001__;
  assign new_new_n25459__ = new_new_n25005__ & new_new_n25458__;
  assign new_new_n25460__ = ~new_new_n25005__ & ~new_new_n25458__;
  assign new_new_n25461__ = ~pi02 & ~new_new_n17204__;
  assign new_new_n25462__ = ~pi01 & new_new_n17204__;
  assign new_new_n25463__ = new_new_n15432__ & ~new_new_n25461__;
  assign new_new_n25464__ = ~new_new_n25462__ & new_new_n25463__;
  assign new_new_n25465__ = pi02 & new_new_n17204__;
  assign new_new_n25466__ = pi01 & ~new_new_n17204__;
  assign new_new_n25467__ = ~new_new_n15432__ & ~new_new_n25465__;
  assign new_new_n25468__ = ~new_new_n25466__ & new_new_n25467__;
  assign new_new_n25469__ = ~new_new_n25464__ & ~new_new_n25468__;
  assign new_new_n25470__ = pi00 & ~new_new_n25469__;
  assign new_new_n25471__ = pi02 & new_new_n15439__;
  assign new_new_n25472__ = ~pi02 & ~new_new_n15439__;
  assign new_new_n25473__ = pi01 & ~new_new_n25471__;
  assign new_new_n25474__ = ~new_new_n25472__ & new_new_n25473__;
  assign new_new_n25475__ = pi02 & ~new_new_n15464__;
  assign new_new_n25476__ = ~pi01 & ~new_new_n25475__;
  assign new_new_n25477__ = ~pi00 & ~new_new_n25476__;
  assign new_new_n25478__ = ~new_new_n25474__ & new_new_n25477__;
  assign new_new_n25479__ = ~new_new_n25470__ & ~new_new_n25478__;
  assign new_new_n25480__ = ~pi01 & new_new_n15471__;
  assign new_new_n25481__ = pi01 & ~new_new_n15464__;
  assign new_new_n25482__ = ~new_new_n25480__ & ~new_new_n25481__;
  assign new_new_n25483__ = pi02 & ~new_new_n25482__;
  assign new_new_n25484__ = new_new_n13508__ & new_new_n15464__;
  assign new_new_n25485__ = ~new_new_n25483__ & ~new_new_n25484__;
  assign new_new_n25486__ = ~pi00 & ~new_new_n25485__;
  assign new_new_n25487__ = pi01 & new_new_n15439__;
  assign new_new_n25488__ = ~new_new_n25472__ & ~new_new_n25487__;
  assign new_new_n25489__ = ~new_new_n17240__ & new_new_n25488__;
  assign new_new_n25490__ = ~pi01 & ~new_new_n15439__;
  assign new_new_n25491__ = ~new_new_n25471__ & ~new_new_n25490__;
  assign new_new_n25492__ = new_new_n17240__ & new_new_n25491__;
  assign new_new_n25493__ = pi00 & ~new_new_n25489__;
  assign new_new_n25494__ = ~new_new_n25492__ & new_new_n25493__;
  assign new_new_n25495__ = ~new_new_n25486__ & ~new_new_n25494__;
  assign new_new_n25496__ = ~new_new_n24638__ & ~new_new_n24639__;
  assign new_new_n25497__ = ~new_new_n24997__ & new_new_n25496__;
  assign new_new_n25498__ = new_new_n24997__ & ~new_new_n25496__;
  assign new_new_n25499__ = ~new_new_n25497__ & ~new_new_n25498__;
  assign new_new_n25500__ = pi02 & new_new_n15471__;
  assign new_new_n25501__ = ~pi02 & ~new_new_n15471__;
  assign new_new_n25502__ = ~new_new_n25500__ & ~new_new_n25501__;
  assign new_new_n25503__ = pi01 & ~new_new_n25502__;
  assign new_new_n25504__ = new_new_n12798__ & new_new_n15809__;
  assign new_new_n25505__ = ~new_new_n25503__ & ~new_new_n25504__;
  assign new_new_n25506__ = ~pi00 & ~new_new_n25505__;
  assign new_new_n25507__ = ~pi01 & new_new_n15464__;
  assign new_new_n25508__ = ~new_new_n25475__ & ~new_new_n25507__;
  assign new_new_n25509__ = ~new_new_n15819__ & new_new_n25508__;
  assign new_new_n25510__ = ~pi02 & new_new_n15464__;
  assign new_new_n25511__ = ~new_new_n25481__ & ~new_new_n25510__;
  assign new_new_n25512__ = new_new_n15819__ & new_new_n25511__;
  assign new_new_n25513__ = pi00 & ~new_new_n25509__;
  assign new_new_n25514__ = ~new_new_n25512__ & new_new_n25513__;
  assign new_new_n25515__ = ~new_new_n25506__ & ~new_new_n25514__;
  assign new_new_n25516__ = pi01 & new_new_n15809__;
  assign new_new_n25517__ = ~pi01 & new_new_n15487__;
  assign new_new_n25518__ = ~new_new_n25516__ & ~new_new_n25517__;
  assign new_new_n25519__ = pi02 & ~new_new_n25518__;
  assign new_new_n25520__ = new_new_n13508__ & ~new_new_n15809__;
  assign new_new_n25521__ = ~new_new_n25519__ & ~new_new_n25520__;
  assign new_new_n25522__ = ~pi00 & ~new_new_n25521__;
  assign new_new_n25523__ = ~new_new_n18630__ & new_new_n25502__;
  assign new_new_n25524__ = pi01 & ~new_new_n15471__;
  assign new_new_n25525__ = ~new_new_n25480__ & ~new_new_n25524__;
  assign new_new_n25526__ = new_new_n18630__ & ~new_new_n25525__;
  assign new_new_n25527__ = pi00 & ~new_new_n25523__;
  assign new_new_n25528__ = ~new_new_n25526__ & new_new_n25527__;
  assign new_new_n25529__ = ~new_new_n25522__ & ~new_new_n25528__;
  assign new_new_n25530__ = ~new_new_n24974__ & ~new_new_n24975__;
  assign new_new_n25531__ = new_new_n24979__ & new_new_n25530__;
  assign new_new_n25532__ = ~new_new_n24979__ & ~new_new_n25530__;
  assign new_new_n25533__ = ~new_new_n25531__ & ~new_new_n25532__;
  assign new_new_n25534__ = new_new_n25529__ & ~new_new_n25533__;
  assign new_new_n25535__ = ~new_new_n25529__ & new_new_n25533__;
  assign new_new_n25536__ = ~new_new_n24960__ & ~new_new_n24961__;
  assign new_new_n25537__ = ~new_new_n24971__ & new_new_n25536__;
  assign new_new_n25538__ = new_new_n24971__ & ~new_new_n25536__;
  assign new_new_n25539__ = ~new_new_n25537__ & ~new_new_n25538__;
  assign new_new_n25540__ = pi02 & new_new_n17587__;
  assign new_new_n25541__ = pi01 & ~new_new_n17587__;
  assign new_new_n25542__ = ~new_new_n15487__ & ~new_new_n25540__;
  assign new_new_n25543__ = ~new_new_n25541__ & new_new_n25542__;
  assign new_new_n25544__ = ~pi02 & ~new_new_n17587__;
  assign new_new_n25545__ = ~pi01 & new_new_n17587__;
  assign new_new_n25546__ = new_new_n15487__ & ~new_new_n25544__;
  assign new_new_n25547__ = ~new_new_n25545__ & new_new_n25546__;
  assign new_new_n25548__ = ~new_new_n25543__ & ~new_new_n25547__;
  assign new_new_n25549__ = pi00 & ~new_new_n25548__;
  assign new_new_n25550__ = pi02 & ~new_new_n15520__;
  assign new_new_n25551__ = ~pi01 & ~new_new_n25550__;
  assign new_new_n25552__ = pi02 & new_new_n15524__;
  assign new_new_n25553__ = ~pi02 & ~new_new_n15524__;
  assign new_new_n25554__ = ~new_new_n25552__ & ~new_new_n25553__;
  assign new_new_n25555__ = pi01 & ~new_new_n25554__;
  assign new_new_n25556__ = ~pi00 & ~new_new_n25551__;
  assign new_new_n25557__ = ~new_new_n25555__ & new_new_n25556__;
  assign new_new_n25558__ = ~new_new_n25549__ & ~new_new_n25557__;
  assign new_new_n25559__ = ~new_new_n18913__ & ~new_new_n25554__;
  assign new_new_n25560__ = ~pi01 & ~new_new_n15524__;
  assign new_new_n25561__ = pi01 & new_new_n15524__;
  assign new_new_n25562__ = ~new_new_n25560__ & ~new_new_n25561__;
  assign new_new_n25563__ = new_new_n18913__ & ~new_new_n25562__;
  assign new_new_n25564__ = pi00 & ~new_new_n25559__;
  assign new_new_n25565__ = ~new_new_n25563__ & new_new_n25564__;
  assign new_new_n25566__ = ~pi00 & ~new_new_n25290__;
  assign new_new_n25567__ = ~pi02 & ~new_new_n15520__;
  assign new_new_n25568__ = pi01 & ~new_new_n15520__;
  assign new_new_n25569__ = ~pi01 & new_new_n15533__;
  assign new_new_n25570__ = pi02 & ~new_new_n25569__;
  assign new_new_n25571__ = ~new_new_n25568__ & new_new_n25570__;
  assign new_new_n25572__ = new_new_n25566__ & ~new_new_n25567__;
  assign new_new_n25573__ = ~new_new_n25571__ & new_new_n25572__;
  assign new_new_n25574__ = ~new_new_n25565__ & ~new_new_n25573__;
  assign new_new_n25575__ = ~new_new_n24936__ & ~new_new_n24937__;
  assign new_new_n25576__ = ~new_new_n24939__ & new_new_n25575__;
  assign new_new_n25577__ = new_new_n24939__ & ~new_new_n25575__;
  assign new_new_n25578__ = ~new_new_n25576__ & ~new_new_n25577__;
  assign new_new_n25579__ = new_new_n25574__ & new_new_n25578__;
  assign new_new_n25580__ = ~new_new_n25574__ & ~new_new_n25578__;
  assign new_new_n25581__ = pi02 & new_new_n14393__;
  assign new_new_n25582__ = ~new_new_n15767__ & new_new_n25581__;
  assign new_new_n25583__ = ~pi00 & pi01;
  assign new_new_n25584__ = ~pi02 & ~new_new_n15533__;
  assign new_new_n25585__ = pi02 & new_new_n15533__;
  assign new_new_n25586__ = ~new_new_n25584__ & ~new_new_n25585__;
  assign new_new_n25587__ = new_new_n25583__ & ~new_new_n25586__;
  assign new_new_n25588__ = pi01 & new_new_n18124__;
  assign new_new_n25589__ = new_new_n15520__ & new_new_n25584__;
  assign new_new_n25590__ = ~new_new_n25588__ & ~new_new_n25589__;
  assign new_new_n25591__ = ~new_new_n15771__ & ~new_new_n25590__;
  assign new_new_n25592__ = ~pi01 & ~new_new_n19731__;
  assign new_new_n25593__ = ~new_new_n25568__ & ~new_new_n25592__;
  assign new_new_n25594__ = ~new_new_n25567__ & ~new_new_n25593__;
  assign new_new_n25595__ = pi01 & ~new_new_n15533__;
  assign new_new_n25596__ = ~pi02 & new_new_n15520__;
  assign new_new_n25597__ = ~new_new_n25595__ & ~new_new_n25596__;
  assign new_new_n25598__ = ~new_new_n15534__ & new_new_n15771__;
  assign new_new_n25599__ = ~new_new_n25597__ & new_new_n25598__;
  assign new_new_n25600__ = ~new_new_n25591__ & ~new_new_n25599__;
  assign new_new_n25601__ = ~new_new_n25594__ & new_new_n25600__;
  assign new_new_n25602__ = pi00 & ~new_new_n25601__;
  assign new_new_n25603__ = ~new_new_n24928__ & ~new_new_n24929__;
  assign new_new_n25604__ = new_new_n24933__ & new_new_n25603__;
  assign new_new_n25605__ = ~new_new_n24933__ & ~new_new_n25603__;
  assign new_new_n25606__ = ~new_new_n25604__ & ~new_new_n25605__;
  assign new_new_n25607__ = ~pi01 & new_new_n15572__;
  assign new_new_n25608__ = pi01 & new_new_n15560__;
  assign new_new_n25609__ = pi02 & ~new_new_n25607__;
  assign new_new_n25610__ = ~new_new_n25608__ & new_new_n25609__;
  assign new_new_n25611__ = new_new_n13508__ & new_new_n15560__;
  assign new_new_n25612__ = ~new_new_n25610__ & ~new_new_n25611__;
  assign new_new_n25613__ = ~pi00 & ~new_new_n25612__;
  assign new_new_n25614__ = pi01 & ~new_new_n15767__;
  assign new_new_n25615__ = ~pi02 & new_new_n15767__;
  assign new_new_n25616__ = ~new_new_n25614__ & ~new_new_n25615__;
  assign new_new_n25617__ = ~new_new_n18454__ & ~new_new_n25616__;
  assign new_new_n25618__ = ~pi02 & ~new_new_n15767__;
  assign new_new_n25619__ = pi01 & new_new_n15767__;
  assign new_new_n25620__ = ~new_new_n25618__ & ~new_new_n25619__;
  assign new_new_n25621__ = new_new_n18454__ & new_new_n25620__;
  assign new_new_n25622__ = ~new_new_n25617__ & ~new_new_n25621__;
  assign new_new_n25623__ = pi00 & ~new_new_n25622__;
  assign new_new_n25624__ = ~new_new_n25613__ & ~new_new_n25623__;
  assign new_new_n25625__ = new_new_n13508__ & new_new_n15572__;
  assign new_new_n25626__ = ~pi01 & new_new_n15564__;
  assign new_new_n25627__ = pi01 & new_new_n15572__;
  assign new_new_n25628__ = pi02 & ~new_new_n25626__;
  assign new_new_n25629__ = ~new_new_n25627__ & new_new_n25628__;
  assign new_new_n25630__ = ~pi00 & ~new_new_n25625__;
  assign new_new_n25631__ = ~new_new_n25629__ & new_new_n25630__;
  assign new_new_n25632__ = ~pi01 & ~new_new_n15560__;
  assign new_new_n25633__ = pi02 & new_new_n15560__;
  assign new_new_n25634__ = ~new_new_n25632__ & ~new_new_n25633__;
  assign new_new_n25635__ = new_new_n18944__ & new_new_n25634__;
  assign new_new_n25636__ = ~pi02 & ~new_new_n15560__;
  assign new_new_n25637__ = ~new_new_n25608__ & ~new_new_n25636__;
  assign new_new_n25638__ = ~new_new_n18944__ & new_new_n25637__;
  assign new_new_n25639__ = pi00 & ~new_new_n25635__;
  assign new_new_n25640__ = ~new_new_n25638__ & new_new_n25639__;
  assign new_new_n25641__ = ~new_new_n25631__ & ~new_new_n25640__;
  assign new_new_n25642__ = ~new_new_n24881__ & ~new_new_n24882__;
  assign new_new_n25643__ = new_new_n24892__ & new_new_n25642__;
  assign new_new_n25644__ = ~new_new_n24892__ & ~new_new_n25642__;
  assign new_new_n25645__ = ~new_new_n25643__ & ~new_new_n25644__;
  assign new_new_n25646__ = ~new_new_n25641__ & ~new_new_n25645__;
  assign new_new_n25647__ = new_new_n25641__ & new_new_n25645__;
  assign new_new_n25648__ = new_new_n13508__ & new_new_n15564__;
  assign new_new_n25649__ = pi01 & ~new_new_n15564__;
  assign new_new_n25650__ = ~pi01 & new_new_n15615__;
  assign new_new_n25651__ = ~new_new_n25649__ & ~new_new_n25650__;
  assign new_new_n25652__ = pi02 & ~new_new_n25651__;
  assign new_new_n25653__ = ~pi00 & ~new_new_n25648__;
  assign new_new_n25654__ = ~new_new_n25652__ & new_new_n25653__;
  assign new_new_n25655__ = pi02 & ~new_new_n19534__;
  assign new_new_n25656__ = pi01 & new_new_n19534__;
  assign new_new_n25657__ = ~new_new_n25655__ & ~new_new_n25656__;
  assign new_new_n25658__ = ~new_new_n15572__ & ~new_new_n25657__;
  assign new_new_n25659__ = new_new_n15572__ & new_new_n25657__;
  assign new_new_n25660__ = pi00 & ~new_new_n25658__;
  assign new_new_n25661__ = ~new_new_n25659__ & new_new_n25660__;
  assign new_new_n25662__ = ~new_new_n25654__ & ~new_new_n25661__;
  assign new_new_n25663__ = pi01 & ~new_new_n15615__;
  assign new_new_n25664__ = ~pi01 & new_new_n15743__;
  assign new_new_n25665__ = pi02 & ~new_new_n25664__;
  assign new_new_n25666__ = ~new_new_n25663__ & ~new_new_n25665__;
  assign new_new_n25667__ = pi02 & new_new_n25663__;
  assign new_new_n25668__ = ~pi00 & ~new_new_n25666__;
  assign new_new_n25669__ = ~new_new_n25667__ & new_new_n25668__;
  assign new_new_n25670__ = pi02 & ~new_new_n15564__;
  assign new_new_n25671__ = ~new_new_n25626__ & ~new_new_n25670__;
  assign new_new_n25672__ = ~new_new_n18512__ & new_new_n25671__;
  assign new_new_n25673__ = ~pi02 & new_new_n15564__;
  assign new_new_n25674__ = ~new_new_n25649__ & ~new_new_n25673__;
  assign new_new_n25675__ = new_new_n18512__ & new_new_n25674__;
  assign new_new_n25676__ = pi00 & ~new_new_n25672__;
  assign new_new_n25677__ = ~new_new_n25675__ & new_new_n25676__;
  assign new_new_n25678__ = ~new_new_n25669__ & ~new_new_n25677__;
  assign new_new_n25679__ = ~pi01 & ~new_new_n15638__;
  assign new_new_n25680__ = pi01 & new_new_n15743__;
  assign new_new_n25681__ = pi02 & ~new_new_n25679__;
  assign new_new_n25682__ = ~new_new_n25680__ & new_new_n25681__;
  assign new_new_n25683__ = new_new_n13508__ & new_new_n15743__;
  assign new_new_n25684__ = ~new_new_n25682__ & ~new_new_n25683__;
  assign new_new_n25685__ = ~pi00 & ~new_new_n25684__;
  assign new_new_n25686__ = ~pi02 & ~new_new_n19005__;
  assign new_new_n25687__ = ~pi01 & new_new_n19005__;
  assign new_new_n25688__ = new_new_n15615__ & ~new_new_n25686__;
  assign new_new_n25689__ = ~new_new_n25687__ & new_new_n25688__;
  assign new_new_n25690__ = pi02 & new_new_n19005__;
  assign new_new_n25691__ = pi01 & ~new_new_n19005__;
  assign new_new_n25692__ = ~new_new_n15615__ & ~new_new_n25690__;
  assign new_new_n25693__ = ~new_new_n25691__ & new_new_n25692__;
  assign new_new_n25694__ = ~new_new_n25689__ & ~new_new_n25693__;
  assign new_new_n25695__ = pi00 & ~new_new_n25694__;
  assign new_new_n25696__ = ~new_new_n25685__ & ~new_new_n25695__;
  assign new_new_n25697__ = pi02 & ~new_new_n19491__;
  assign new_new_n25698__ = pi01 & new_new_n19491__;
  assign new_new_n25699__ = ~new_new_n25697__ & ~new_new_n25698__;
  assign new_new_n25700__ = new_new_n15743__ & ~new_new_n25699__;
  assign new_new_n25701__ = ~new_new_n15743__ & new_new_n25699__;
  assign new_new_n25702__ = pi00 & ~new_new_n25700__;
  assign new_new_n25703__ = ~new_new_n25701__ & new_new_n25702__;
  assign new_new_n25704__ = pi02 & new_new_n15582__;
  assign new_new_n25705__ = ~pi01 & ~new_new_n25704__;
  assign new_new_n25706__ = ~pi02 & new_new_n15638__;
  assign new_new_n25707__ = pi02 & ~new_new_n15638__;
  assign new_new_n25708__ = ~new_new_n25706__ & ~new_new_n25707__;
  assign new_new_n25709__ = pi01 & ~new_new_n25708__;
  assign new_new_n25710__ = ~pi00 & ~new_new_n25705__;
  assign new_new_n25711__ = ~new_new_n25709__ & new_new_n25710__;
  assign new_new_n25712__ = ~new_new_n25703__ & ~new_new_n25711__;
  assign new_new_n25713__ = new_new_n13508__ & ~new_new_n15582__;
  assign new_new_n25714__ = pi01 & new_new_n15582__;
  assign new_new_n25715__ = ~pi01 & new_new_n15647__;
  assign new_new_n25716__ = ~new_new_n25714__ & ~new_new_n25715__;
  assign new_new_n25717__ = pi02 & ~new_new_n25716__;
  assign new_new_n25718__ = ~new_new_n25713__ & ~new_new_n25717__;
  assign new_new_n25719__ = ~pi00 & ~new_new_n25718__;
  assign new_new_n25720__ = pi01 & new_new_n15638__;
  assign new_new_n25721__ = new_new_n15716__ & ~new_new_n15736__;
  assign new_new_n25722__ = new_new_n15718__ & new_new_n15736__;
  assign new_new_n25723__ = ~new_new_n25721__ & ~new_new_n25722__;
  assign new_new_n25724__ = ~new_new_n25679__ & ~new_new_n25720__;
  assign new_new_n25725__ = ~new_new_n25723__ & new_new_n25724__;
  assign new_new_n25726__ = ~new_new_n25708__ & new_new_n25723__;
  assign new_new_n25727__ = pi00 & ~new_new_n25725__;
  assign new_new_n25728__ = ~new_new_n25726__ & new_new_n25727__;
  assign new_new_n25729__ = ~new_new_n25719__ & ~new_new_n25728__;
  assign new_new_n25730__ = ~pi01 & ~new_new_n15710__;
  assign new_new_n25731__ = pi01 & ~new_new_n15647__;
  assign new_new_n25732__ = pi02 & ~new_new_n25730__;
  assign new_new_n25733__ = ~new_new_n25731__ & new_new_n25732__;
  assign new_new_n25734__ = new_new_n13508__ & ~new_new_n15647__;
  assign new_new_n25735__ = ~new_new_n25733__ & ~new_new_n25734__;
  assign new_new_n25736__ = ~pi00 & ~new_new_n25735__;
  assign new_new_n25737__ = ~pi01 & ~new_new_n15736__;
  assign new_new_n25738__ = ~pi02 & new_new_n15736__;
  assign new_new_n25739__ = new_new_n15582__ & ~new_new_n25737__;
  assign new_new_n25740__ = ~new_new_n25738__ & new_new_n25739__;
  assign new_new_n25741__ = pi01 & new_new_n15736__;
  assign new_new_n25742__ = pi02 & ~new_new_n15736__;
  assign new_new_n25743__ = ~new_new_n15582__ & ~new_new_n25741__;
  assign new_new_n25744__ = ~new_new_n25742__ & new_new_n25743__;
  assign new_new_n25745__ = ~new_new_n25740__ & ~new_new_n25744__;
  assign new_new_n25746__ = pi00 & ~new_new_n25745__;
  assign new_new_n25747__ = ~new_new_n25736__ & ~new_new_n25746__;
  assign new_new_n25748__ = ~new_new_n15673__ & ~new_new_n24799__;
  assign new_new_n25749__ = ~new_new_n24811__ & ~new_new_n25748__;
  assign new_new_n25750__ = pi06 & ~new_new_n25749__;
  assign new_new_n25751__ = pi05 & ~new_new_n24790__;
  assign new_new_n25752__ = new_new_n24809__ & ~new_new_n25751__;
  assign new_new_n25753__ = pi05 & ~new_new_n25752__;
  assign new_new_n25754__ = new_new_n15673__ & ~new_new_n25753__;
  assign new_new_n25755__ = pi05 & new_new_n25752__;
  assign new_new_n25756__ = ~pi06 & ~new_new_n15673__;
  assign new_new_n25757__ = ~new_new_n25755__ & new_new_n25756__;
  assign new_new_n25758__ = ~new_new_n25754__ & ~new_new_n25757__;
  assign new_new_n25759__ = new_new_n24799__ & ~new_new_n25758__;
  assign new_new_n25760__ = new_new_n15673__ & new_new_n25753__;
  assign new_new_n25761__ = ~new_new_n24799__ & new_new_n25760__;
  assign new_new_n25762__ = ~new_new_n25759__ & ~new_new_n25761__;
  assign new_new_n25763__ = ~new_new_n25750__ & new_new_n25762__;
  assign new_new_n25764__ = pi01 & new_new_n15710__;
  assign new_new_n25765__ = ~pi01 & ~new_new_n15656__;
  assign new_new_n25766__ = ~new_new_n25764__ & ~new_new_n25765__;
  assign new_new_n25767__ = pi02 & ~new_new_n25766__;
  assign new_new_n25768__ = new_new_n13508__ & ~new_new_n15710__;
  assign new_new_n25769__ = ~new_new_n25767__ & ~new_new_n25768__;
  assign new_new_n25770__ = ~pi00 & ~new_new_n25769__;
  assign new_new_n25771__ = pi02 & ~new_new_n15647__;
  assign new_new_n25772__ = ~new_new_n25715__ & ~new_new_n25771__;
  assign new_new_n25773__ = ~new_new_n19118__ & ~new_new_n25772__;
  assign new_new_n25774__ = ~pi02 & new_new_n15647__;
  assign new_new_n25775__ = ~new_new_n25731__ & ~new_new_n25774__;
  assign new_new_n25776__ = new_new_n19118__ & ~new_new_n25775__;
  assign new_new_n25777__ = pi00 & ~new_new_n25773__;
  assign new_new_n25778__ = ~new_new_n25776__ & new_new_n25777__;
  assign new_new_n25779__ = ~new_new_n25770__ & ~new_new_n25778__;
  assign new_new_n25780__ = new_new_n25763__ & ~new_new_n25779__;
  assign new_new_n25781__ = ~new_new_n25763__ & new_new_n25779__;
  assign new_new_n25782__ = ~new_new_n24809__ & new_new_n25751__;
  assign new_new_n25783__ = ~new_new_n25752__ & ~new_new_n25782__;
  assign new_new_n25784__ = ~pi02 & ~new_new_n15710__;
  assign new_new_n25785__ = ~new_new_n25764__ & ~new_new_n25784__;
  assign new_new_n25786__ = ~new_new_n19466__ & new_new_n25785__;
  assign new_new_n25787__ = pi02 & new_new_n15710__;
  assign new_new_n25788__ = ~new_new_n25730__ & ~new_new_n25787__;
  assign new_new_n25789__ = new_new_n19466__ & new_new_n25788__;
  assign new_new_n25790__ = pi00 & ~new_new_n25786__;
  assign new_new_n25791__ = ~new_new_n25789__ & new_new_n25790__;
  assign new_new_n25792__ = pi02 & ~new_new_n15643__;
  assign new_new_n25793__ = ~pi01 & ~new_new_n25792__;
  assign new_new_n25794__ = pi02 & new_new_n15656__;
  assign new_new_n25795__ = ~pi02 & ~new_new_n15656__;
  assign new_new_n25796__ = ~new_new_n25794__ & ~new_new_n25795__;
  assign new_new_n25797__ = pi01 & ~new_new_n25796__;
  assign new_new_n25798__ = ~pi00 & ~new_new_n25793__;
  assign new_new_n25799__ = ~new_new_n25797__ & new_new_n25798__;
  assign new_new_n25800__ = ~new_new_n25791__ & ~new_new_n25799__;
  assign new_new_n25801__ = new_new_n25783__ & ~new_new_n25800__;
  assign new_new_n25802__ = ~new_new_n25783__ & new_new_n25800__;
  assign new_new_n25803__ = ~new_new_n15677__ & ~new_new_n25796__;
  assign new_new_n25804__ = pi01 & new_new_n15656__;
  assign new_new_n25805__ = ~new_new_n25765__ & ~new_new_n25804__;
  assign new_new_n25806__ = new_new_n15677__ & ~new_new_n25805__;
  assign new_new_n25807__ = pi00 & ~new_new_n25803__;
  assign new_new_n25808__ = ~new_new_n25806__ & new_new_n25807__;
  assign new_new_n25809__ = pi02 & new_new_n15661__;
  assign new_new_n25810__ = ~pi01 & ~new_new_n25809__;
  assign new_new_n25811__ = ~pi02 & new_new_n15643__;
  assign new_new_n25812__ = ~new_new_n25792__ & ~new_new_n25811__;
  assign new_new_n25813__ = pi01 & new_new_n25812__;
  assign new_new_n25814__ = ~pi00 & ~new_new_n25810__;
  assign new_new_n25815__ = ~new_new_n25813__ & new_new_n25814__;
  assign new_new_n25816__ = ~new_new_n25808__ & ~new_new_n25815__;
  assign new_new_n25817__ = pi01 & ~new_new_n15661__;
  assign new_new_n25818__ = ~pi02 & ~new_new_n25817__;
  assign new_new_n25819__ = ~pi01 & new_new_n15668__;
  assign new_new_n25820__ = ~new_new_n25817__ & ~new_new_n25819__;
  assign new_new_n25821__ = pi02 & ~new_new_n25820__;
  assign new_new_n25822__ = ~pi00 & ~new_new_n25818__;
  assign new_new_n25823__ = ~new_new_n25821__ & new_new_n25822__;
  assign new_new_n25824__ = ~pi01 & ~new_new_n15643__;
  assign new_new_n25825__ = pi01 & new_new_n15643__;
  assign new_new_n25826__ = ~new_new_n25824__ & ~new_new_n25825__;
  assign new_new_n25827__ = new_new_n20176__ & ~new_new_n25826__;
  assign new_new_n25828__ = ~new_new_n20176__ & new_new_n25812__;
  assign new_new_n25829__ = pi00 & ~new_new_n25827__;
  assign new_new_n25830__ = ~new_new_n25828__ & new_new_n25829__;
  assign new_new_n25831__ = ~new_new_n25823__ & ~new_new_n25830__;
  assign new_new_n25832__ = ~new_new_n11482__ & ~new_new_n15673__;
  assign new_new_n25833__ = ~new_new_n25831__ & new_new_n25832__;
  assign new_new_n25834__ = new_new_n25816__ & ~new_new_n25833__;
  assign new_new_n25835__ = new_new_n11474__ & new_new_n15674__;
  assign new_new_n25836__ = ~new_new_n10726__ & new_new_n15668__;
  assign new_new_n25837__ = new_new_n11473__ & ~new_new_n25836__;
  assign new_new_n25838__ = new_new_n11482__ & new_new_n20195__;
  assign new_new_n25839__ = ~new_new_n12828__ & ~new_new_n20628__;
  assign new_new_n25840__ = ~new_new_n25835__ & new_new_n25839__;
  assign new_new_n25841__ = ~new_new_n25837__ & ~new_new_n25838__;
  assign new_new_n25842__ = new_new_n25840__ & new_new_n25841__;
  assign new_new_n25843__ = ~new_new_n25834__ & new_new_n25842__;
  assign new_new_n25844__ = new_new_n20628__ & new_new_n25809__;
  assign new_new_n25845__ = ~new_new_n25832__ & ~new_new_n25844__;
  assign new_new_n25846__ = ~new_new_n25831__ & ~new_new_n25845__;
  assign new_new_n25847__ = ~new_new_n25816__ & new_new_n25846__;
  assign new_new_n25848__ = ~new_new_n25843__ & ~new_new_n25847__;
  assign new_new_n25849__ = ~new_new_n25802__ & ~new_new_n25848__;
  assign new_new_n25850__ = ~new_new_n25801__ & ~new_new_n25849__;
  assign new_new_n25851__ = ~new_new_n25781__ & ~new_new_n25850__;
  assign new_new_n25852__ = ~new_new_n25780__ & ~new_new_n25851__;
  assign new_new_n25853__ = ~new_new_n25747__ & ~new_new_n25852__;
  assign new_new_n25854__ = new_new_n25747__ & new_new_n25852__;
  assign new_new_n25855__ = ~new_new_n24817__ & ~new_new_n24818__;
  assign new_new_n25856__ = new_new_n24826__ & ~new_new_n25855__;
  assign new_new_n25857__ = ~new_new_n24826__ & new_new_n25855__;
  assign new_new_n25858__ = ~new_new_n25856__ & ~new_new_n25857__;
  assign new_new_n25859__ = ~new_new_n25854__ & ~new_new_n25858__;
  assign new_new_n25860__ = ~new_new_n25853__ & ~new_new_n25859__;
  assign new_new_n25861__ = ~new_new_n25729__ & ~new_new_n25860__;
  assign new_new_n25862__ = new_new_n25729__ & new_new_n25860__;
  assign new_new_n25863__ = ~new_new_n24829__ & ~new_new_n24842__;
  assign new_new_n25864__ = new_new_n24841__ & ~new_new_n25863__;
  assign new_new_n25865__ = ~new_new_n24841__ & new_new_n25863__;
  assign new_new_n25866__ = ~new_new_n25864__ & ~new_new_n25865__;
  assign new_new_n25867__ = ~new_new_n25862__ & new_new_n25866__;
  assign new_new_n25868__ = ~new_new_n25861__ & ~new_new_n25867__;
  assign new_new_n25869__ = new_new_n25712__ & new_new_n25868__;
  assign new_new_n25870__ = ~new_new_n25712__ & ~new_new_n25868__;
  assign new_new_n25871__ = ~new_new_n24845__ & ~new_new_n24846__;
  assign new_new_n25872__ = ~new_new_n24851__ & new_new_n25871__;
  assign new_new_n25873__ = new_new_n24851__ & ~new_new_n25871__;
  assign new_new_n25874__ = ~new_new_n25872__ & ~new_new_n25873__;
  assign new_new_n25875__ = ~new_new_n25870__ & new_new_n25874__;
  assign new_new_n25876__ = ~new_new_n25869__ & ~new_new_n25875__;
  assign new_new_n25877__ = ~new_new_n25696__ & new_new_n25876__;
  assign new_new_n25878__ = new_new_n25696__ & ~new_new_n25876__;
  assign new_new_n25879__ = ~new_new_n24854__ & ~new_new_n24855__;
  assign new_new_n25880__ = new_new_n24865__ & new_new_n25879__;
  assign new_new_n25881__ = ~new_new_n24865__ & ~new_new_n25879__;
  assign new_new_n25882__ = ~new_new_n25880__ & ~new_new_n25881__;
  assign new_new_n25883__ = ~new_new_n25878__ & ~new_new_n25882__;
  assign new_new_n25884__ = ~new_new_n25877__ & ~new_new_n25883__;
  assign new_new_n25885__ = new_new_n25678__ & new_new_n25884__;
  assign new_new_n25886__ = ~new_new_n25678__ & ~new_new_n25884__;
  assign new_new_n25887__ = pi05 & new_new_n24747__;
  assign new_new_n25888__ = ~pi05 & ~new_new_n24747__;
  assign new_new_n25889__ = ~new_new_n25887__ & ~new_new_n25888__;
  assign new_new_n25890__ = new_new_n24739__ & ~new_new_n25889__;
  assign new_new_n25891__ = ~new_new_n24739__ & new_new_n25889__;
  assign new_new_n25892__ = ~new_new_n25890__ & ~new_new_n25891__;
  assign new_new_n25893__ = new_new_n24867__ & new_new_n25892__;
  assign new_new_n25894__ = ~new_new_n24867__ & ~new_new_n25892__;
  assign new_new_n25895__ = ~new_new_n25893__ & ~new_new_n25894__;
  assign new_new_n25896__ = ~new_new_n25886__ & ~new_new_n25895__;
  assign new_new_n25897__ = ~new_new_n25885__ & ~new_new_n25896__;
  assign new_new_n25898__ = ~new_new_n25662__ & ~new_new_n25897__;
  assign new_new_n25899__ = new_new_n25662__ & new_new_n25897__;
  assign new_new_n25900__ = ~new_new_n24868__ & ~new_new_n24876__;
  assign new_new_n25901__ = ~new_new_n24739__ & new_new_n25900__;
  assign new_new_n25902__ = new_new_n25889__ & ~new_new_n25900__;
  assign new_new_n25903__ = ~new_new_n25901__ & ~new_new_n25902__;
  assign new_new_n25904__ = ~new_new_n24732__ & ~new_new_n25903__;
  assign new_new_n25905__ = new_new_n24732__ & new_new_n25903__;
  assign new_new_n25906__ = ~new_new_n25904__ & ~new_new_n25905__;
  assign new_new_n25907__ = new_new_n24725__ & new_new_n25906__;
  assign new_new_n25908__ = ~new_new_n24725__ & ~new_new_n25906__;
  assign new_new_n25909__ = ~new_new_n25907__ & ~new_new_n25908__;
  assign new_new_n25910__ = ~new_new_n25899__ & ~new_new_n25909__;
  assign new_new_n25911__ = ~new_new_n25898__ & ~new_new_n25910__;
  assign new_new_n25912__ = ~new_new_n25647__ & ~new_new_n25911__;
  assign new_new_n25913__ = ~new_new_n25646__ & ~new_new_n25912__;
  assign new_new_n25914__ = ~new_new_n25624__ & new_new_n25913__;
  assign new_new_n25915__ = new_new_n25624__ & ~new_new_n25913__;
  assign new_new_n25916__ = ~new_new_n24895__ & ~new_new_n24896__;
  assign new_new_n25917__ = new_new_n24907__ & ~new_new_n25916__;
  assign new_new_n25918__ = ~new_new_n24907__ & new_new_n25916__;
  assign new_new_n25919__ = ~new_new_n25917__ & ~new_new_n25918__;
  assign new_new_n25920__ = ~new_new_n25915__ & ~new_new_n25919__;
  assign new_new_n25921__ = ~new_new_n25914__ & ~new_new_n25920__;
  assign new_new_n25922__ = ~new_new_n25614__ & ~new_new_n25632__;
  assign new_new_n25923__ = pi02 & ~new_new_n25922__;
  assign new_new_n25924__ = pi01 & new_new_n25615__;
  assign new_new_n25925__ = ~new_new_n25923__ & ~new_new_n25924__;
  assign new_new_n25926__ = ~pi00 & ~new_new_n25925__;
  assign new_new_n25927__ = ~new_new_n25569__ & ~new_new_n25595__;
  assign new_new_n25928__ = new_new_n19890__ & ~new_new_n25927__;
  assign new_new_n25929__ = ~new_new_n19890__ & new_new_n25586__;
  assign new_new_n25930__ = pi00 & ~new_new_n25928__;
  assign new_new_n25931__ = ~new_new_n25929__ & new_new_n25930__;
  assign new_new_n25932__ = ~new_new_n25926__ & ~new_new_n25931__;
  assign new_new_n25933__ = ~new_new_n24914__ & ~new_new_n24915__;
  assign new_new_n25934__ = ~new_new_n24925__ & ~new_new_n25933__;
  assign new_new_n25935__ = new_new_n24925__ & new_new_n25933__;
  assign new_new_n25936__ = ~new_new_n25934__ & ~new_new_n25935__;
  assign new_new_n25937__ = new_new_n25932__ & ~new_new_n25936__;
  assign new_new_n25938__ = ~new_new_n25921__ & ~new_new_n25937__;
  assign new_new_n25939__ = ~new_new_n25932__ & new_new_n25936__;
  assign new_new_n25940__ = ~new_new_n25938__ & ~new_new_n25939__;
  assign new_new_n25941__ = new_new_n25606__ & ~new_new_n25940__;
  assign new_new_n25942__ = ~new_new_n25582__ & ~new_new_n25587__;
  assign new_new_n25943__ = ~new_new_n25602__ & new_new_n25942__;
  assign new_new_n25944__ = ~new_new_n25941__ & new_new_n25943__;
  assign new_new_n25945__ = ~new_new_n25606__ & new_new_n25940__;
  assign new_new_n25946__ = ~new_new_n25944__ & ~new_new_n25945__;
  assign new_new_n25947__ = ~new_new_n25580__ & ~new_new_n25946__;
  assign new_new_n25948__ = ~new_new_n25579__ & ~new_new_n25947__;
  assign new_new_n25949__ = ~new_new_n25558__ & new_new_n25948__;
  assign new_new_n25950__ = new_new_n25558__ & ~new_new_n25948__;
  assign new_new_n25951__ = ~new_new_n24946__ & ~new_new_n24947__;
  assign new_new_n25952__ = ~new_new_n24957__ & ~new_new_n25951__;
  assign new_new_n25953__ = new_new_n24957__ & new_new_n25951__;
  assign new_new_n25954__ = ~new_new_n25952__ & ~new_new_n25953__;
  assign new_new_n25955__ = ~new_new_n25950__ & ~new_new_n25954__;
  assign new_new_n25956__ = ~new_new_n25949__ & ~new_new_n25955__;
  assign new_new_n25957__ = ~new_new_n25539__ & new_new_n25956__;
  assign new_new_n25958__ = new_new_n25539__ & ~new_new_n25956__;
  assign new_new_n25959__ = ~pi02 & ~new_new_n18017__;
  assign new_new_n25960__ = ~pi01 & new_new_n18017__;
  assign new_new_n25961__ = ~new_new_n25959__ & ~new_new_n25960__;
  assign new_new_n25962__ = ~new_new_n15809__ & ~new_new_n25961__;
  assign new_new_n25963__ = new_new_n15809__ & new_new_n25961__;
  assign new_new_n25964__ = pi00 & ~new_new_n25962__;
  assign new_new_n25965__ = ~new_new_n25963__ & new_new_n25964__;
  assign new_new_n25966__ = new_new_n13508__ & ~new_new_n15487__;
  assign new_new_n25967__ = pi01 & new_new_n15487__;
  assign new_new_n25968__ = ~new_new_n25560__ & ~new_new_n25967__;
  assign new_new_n25969__ = pi02 & ~new_new_n25968__;
  assign new_new_n25970__ = ~pi00 & ~new_new_n25966__;
  assign new_new_n25971__ = ~new_new_n25969__ & new_new_n25970__;
  assign new_new_n25972__ = ~new_new_n25965__ & ~new_new_n25971__;
  assign new_new_n25973__ = ~new_new_n25958__ & ~new_new_n25972__;
  assign new_new_n25974__ = ~new_new_n25957__ & ~new_new_n25973__;
  assign new_new_n25975__ = ~new_new_n25535__ & ~new_new_n25974__;
  assign new_new_n25976__ = ~new_new_n25534__ & ~new_new_n25975__;
  assign new_new_n25977__ = ~new_new_n25515__ & new_new_n25976__;
  assign new_new_n25978__ = new_new_n25515__ & ~new_new_n25976__;
  assign new_new_n25979__ = ~new_new_n24982__ & ~new_new_n24983__;
  assign new_new_n25980__ = ~new_new_n24995__ & new_new_n25979__;
  assign new_new_n25981__ = new_new_n24995__ & ~new_new_n25979__;
  assign new_new_n25982__ = ~new_new_n25980__ & ~new_new_n25981__;
  assign new_new_n25983__ = ~new_new_n25978__ & new_new_n25982__;
  assign new_new_n25984__ = ~new_new_n25977__ & ~new_new_n25983__;
  assign new_new_n25985__ = ~new_new_n25499__ & new_new_n25984__;
  assign new_new_n25986__ = ~new_new_n25495__ & ~new_new_n25985__;
  assign new_new_n25987__ = new_new_n25499__ & ~new_new_n25984__;
  assign new_new_n25988__ = ~new_new_n25986__ & ~new_new_n25987__;
  assign new_new_n25989__ = new_new_n25479__ & new_new_n25988__;
  assign new_new_n25990__ = ~new_new_n25459__ & ~new_new_n25460__;
  assign new_new_n25991__ = ~new_new_n25989__ & new_new_n25990__;
  assign new_new_n25992__ = ~new_new_n25479__ & ~new_new_n25988__;
  assign new_new_n25993__ = ~new_new_n25991__ & ~new_new_n25992__;
  assign new_new_n25994__ = ~new_new_n25457__ & new_new_n25993__;
  assign new_new_n25995__ = pi02 & ~new_new_n16768__;
  assign new_new_n25996__ = pi01 & new_new_n16768__;
  assign new_new_n25997__ = ~new_new_n25995__ & ~new_new_n25996__;
  assign new_new_n25998__ = ~new_new_n15362__ & new_new_n25997__;
  assign new_new_n25999__ = new_new_n15362__ & ~new_new_n25997__;
  assign new_new_n26000__ = pi00 & ~new_new_n25998__;
  assign new_new_n26001__ = ~new_new_n25999__ & new_new_n26000__;
  assign new_new_n26002__ = new_new_n13508__ & ~new_new_n15432__;
  assign new_new_n26003__ = pi01 & ~new_new_n15432__;
  assign new_new_n26004__ = pi02 & ~new_new_n25490__;
  assign new_new_n26005__ = ~new_new_n26003__ & new_new_n26004__;
  assign new_new_n26006__ = ~pi00 & ~new_new_n26002__;
  assign new_new_n26007__ = ~new_new_n26005__ & new_new_n26006__;
  assign new_new_n26008__ = ~new_new_n26001__ & ~new_new_n26007__;
  assign new_new_n26009__ = new_new_n25457__ & ~new_new_n25993__;
  assign new_new_n26010__ = ~new_new_n26008__ & ~new_new_n26009__;
  assign new_new_n26011__ = ~new_new_n25994__ & ~new_new_n26010__;
  assign new_new_n26012__ = ~new_new_n25453__ & ~new_new_n26011__;
  assign new_new_n26013__ = ~new_new_n25452__ & ~new_new_n26012__;
  assign new_new_n26014__ = ~new_new_n25432__ & ~new_new_n26013__;
  assign new_new_n26015__ = new_new_n25432__ & new_new_n26013__;
  assign new_new_n26016__ = ~new_new_n25035__ & ~new_new_n25036__;
  assign new_new_n26017__ = ~new_new_n25048__ & ~new_new_n26016__;
  assign new_new_n26018__ = new_new_n25048__ & new_new_n26016__;
  assign new_new_n26019__ = ~new_new_n26017__ & ~new_new_n26018__;
  assign new_new_n26020__ = ~new_new_n26015__ & ~new_new_n26019__;
  assign new_new_n26021__ = ~new_new_n26014__ & ~new_new_n26020__;
  assign new_new_n26022__ = ~new_new_n25417__ & new_new_n26021__;
  assign new_new_n26023__ = pi01 & new_new_n17180__;
  assign new_new_n26024__ = pi02 & ~new_new_n17180__;
  assign new_new_n26025__ = ~new_new_n15349__ & ~new_new_n26023__;
  assign new_new_n26026__ = ~new_new_n26024__ & new_new_n26025__;
  assign new_new_n26027__ = ~pi01 & ~new_new_n17180__;
  assign new_new_n26028__ = ~pi02 & new_new_n17180__;
  assign new_new_n26029__ = new_new_n15349__ & ~new_new_n26027__;
  assign new_new_n26030__ = ~new_new_n26028__ & new_new_n26029__;
  assign new_new_n26031__ = ~new_new_n26026__ & ~new_new_n26030__;
  assign new_new_n26032__ = pi00 & ~new_new_n26031__;
  assign new_new_n26033__ = pi01 & ~new_new_n15398__;
  assign new_new_n26034__ = ~pi01 & new_new_n15390__;
  assign new_new_n26035__ = ~new_new_n26033__ & ~new_new_n26034__;
  assign new_new_n26036__ = pi02 & ~new_new_n26035__;
  assign new_new_n26037__ = ~pi02 & ~new_new_n26033__;
  assign new_new_n26038__ = ~pi00 & ~new_new_n26037__;
  assign new_new_n26039__ = ~new_new_n26036__ & new_new_n26038__;
  assign new_new_n26040__ = ~new_new_n26032__ & ~new_new_n26039__;
  assign new_new_n26041__ = new_new_n25417__ & ~new_new_n26021__;
  assign new_new_n26042__ = ~new_new_n26040__ & ~new_new_n26041__;
  assign new_new_n26043__ = ~new_new_n26022__ & ~new_new_n26042__;
  assign new_new_n26044__ = ~new_new_n25411__ & ~new_new_n26043__;
  assign new_new_n26045__ = ~new_new_n25410__ & ~new_new_n26044__;
  assign new_new_n26046__ = ~new_new_n25389__ & ~new_new_n26045__;
  assign new_new_n26047__ = new_new_n25389__ & new_new_n26045__;
  assign new_new_n26048__ = ~new_new_n25072__ & ~new_new_n25096__;
  assign new_new_n26049__ = new_new_n25072__ & new_new_n25096__;
  assign new_new_n26050__ = ~new_new_n26048__ & ~new_new_n26049__;
  assign new_new_n26051__ = ~pi05 & new_new_n24570__;
  assign new_new_n26052__ = ~new_new_n25084__ & ~new_new_n26051__;
  assign new_new_n26053__ = new_new_n26050__ & ~new_new_n26052__;
  assign new_new_n26054__ = ~new_new_n26050__ & new_new_n26052__;
  assign new_new_n26055__ = ~new_new_n26053__ & ~new_new_n26054__;
  assign new_new_n26056__ = ~new_new_n26047__ & ~new_new_n26055__;
  assign new_new_n26057__ = pi01 & ~new_new_n15273__;
  assign new_new_n26058__ = ~pi02 & new_new_n26057__;
  assign new_new_n26059__ = pi02 & ~new_new_n25397__;
  assign new_new_n26060__ = ~new_new_n26057__ & new_new_n26059__;
  assign new_new_n26061__ = ~pi00 & ~new_new_n26058__;
  assign new_new_n26062__ = ~new_new_n26060__ & new_new_n26061__;
  assign new_new_n26063__ = ~pi02 & ~new_new_n15285__;
  assign new_new_n26064__ = ~new_new_n25353__ & ~new_new_n26063__;
  assign new_new_n26065__ = ~new_new_n16078__ & new_new_n26064__;
  assign new_new_n26066__ = ~pi01 & ~new_new_n15285__;
  assign new_new_n26067__ = pi02 & new_new_n15285__;
  assign new_new_n26068__ = ~new_new_n26066__ & ~new_new_n26067__;
  assign new_new_n26069__ = new_new_n16078__ & new_new_n26068__;
  assign new_new_n26070__ = pi00 & ~new_new_n26065__;
  assign new_new_n26071__ = ~new_new_n26069__ & new_new_n26070__;
  assign new_new_n26072__ = ~new_new_n26062__ & ~new_new_n26071__;
  assign new_new_n26073__ = pi05 & ~new_new_n24574__;
  assign new_new_n26074__ = ~new_new_n25104__ & ~new_new_n26073__;
  assign new_new_n26075__ = new_new_n25082__ & ~new_new_n26074__;
  assign new_new_n26076__ = ~new_new_n25082__ & new_new_n26074__;
  assign new_new_n26077__ = ~new_new_n26075__ & ~new_new_n26076__;
  assign new_new_n26078__ = new_new_n26048__ & ~new_new_n26077__;
  assign new_new_n26079__ = ~new_new_n24575__ & ~new_new_n25085__;
  assign new_new_n26080__ = new_new_n25082__ & ~new_new_n26079__;
  assign new_new_n26081__ = ~new_new_n25082__ & new_new_n26079__;
  assign new_new_n26082__ = new_new_n26050__ & ~new_new_n26080__;
  assign new_new_n26083__ = ~new_new_n26081__ & new_new_n26082__;
  assign new_new_n26084__ = new_new_n26049__ & new_new_n26077__;
  assign new_new_n26085__ = ~new_new_n26078__ & ~new_new_n26083__;
  assign new_new_n26086__ = ~new_new_n26084__ & new_new_n26085__;
  assign new_new_n26087__ = new_new_n26072__ & ~new_new_n26086__;
  assign new_new_n26088__ = ~new_new_n26046__ & ~new_new_n26056__;
  assign new_new_n26089__ = ~new_new_n26087__ & new_new_n26088__;
  assign new_new_n26090__ = ~new_new_n26072__ & new_new_n26086__;
  assign new_new_n26091__ = ~new_new_n26089__ & ~new_new_n26090__;
  assign new_new_n26092__ = ~new_new_n25371__ & ~new_new_n26091__;
  assign new_new_n26093__ = ~new_new_n25370__ & ~new_new_n26092__;
  assign new_new_n26094__ = new_new_n25127__ & ~new_new_n26093__;
  assign new_new_n26095__ = ~new_new_n25127__ & new_new_n26093__;
  assign new_new_n26096__ = ~new_new_n26094__ & ~new_new_n26095__;
  assign new_new_n26097__ = new_new_n13508__ & ~new_new_n15314__;
  assign new_new_n26098__ = pi01 & new_new_n15314__;
  assign new_new_n26099__ = ~new_new_n26066__ & ~new_new_n26098__;
  assign new_new_n26100__ = pi02 & ~new_new_n26099__;
  assign new_new_n26101__ = ~pi00 & ~new_new_n26097__;
  assign new_new_n26102__ = ~new_new_n26100__ & new_new_n26101__;
  assign new_new_n26103__ = ~pi02 & new_new_n15248__;
  assign new_new_n26104__ = ~new_new_n25329__ & ~new_new_n26103__;
  assign new_new_n26105__ = ~new_new_n16725__ & new_new_n26104__;
  assign new_new_n26106__ = pi02 & ~new_new_n15248__;
  assign new_new_n26107__ = ~new_new_n25323__ & ~new_new_n26106__;
  assign new_new_n26108__ = new_new_n16725__ & new_new_n26107__;
  assign new_new_n26109__ = pi00 & ~new_new_n26105__;
  assign new_new_n26110__ = ~new_new_n26108__ & new_new_n26109__;
  assign new_new_n26111__ = ~new_new_n26102__ & ~new_new_n26110__;
  assign new_new_n26112__ = ~new_new_n25144__ & ~new_new_n25146__;
  assign new_new_n26113__ = new_new_n26111__ & ~new_new_n26112__;
  assign new_new_n26114__ = ~new_new_n26111__ & new_new_n26112__;
  assign new_new_n26115__ = ~new_new_n26113__ & ~new_new_n26114__;
  assign new_new_n26116__ = new_new_n26096__ & new_new_n26115__;
  assign new_new_n26117__ = ~new_new_n26096__ & ~new_new_n26115__;
  assign new_new_n26118__ = ~new_new_n26116__ & ~new_new_n26117__;
  assign new_new_n26119__ = ~new_new_n26093__ & new_new_n26118__;
  assign new_new_n26120__ = new_new_n26093__ & ~new_new_n26118__;
  assign new_new_n26121__ = ~new_new_n26111__ & ~new_new_n26120__;
  assign new_new_n26122__ = ~new_new_n26119__ & ~new_new_n26121__;
  assign new_new_n26123__ = ~new_new_n25350__ & new_new_n26122__;
  assign new_new_n26124__ = ~new_new_n25349__ & ~new_new_n26123__;
  assign new_new_n26125__ = new_new_n25328__ & ~new_new_n26124__;
  assign new_new_n26126__ = ~new_new_n25157__ & ~new_new_n25192__;
  assign new_new_n26127__ = ~new_new_n25312__ & ~new_new_n26126__;
  assign new_new_n26128__ = new_new_n26125__ & new_new_n26127__;
  assign new_new_n26129__ = ~new_new_n25157__ & ~new_new_n25195__;
  assign new_new_n26130__ = ~new_new_n25169__ & ~new_new_n26129__;
  assign new_new_n26131__ = ~new_new_n25328__ & new_new_n26124__;
  assign new_new_n26132__ = ~new_new_n25193__ & ~new_new_n26130__;
  assign new_new_n26133__ = ~new_new_n25311__ & new_new_n26132__;
  assign new_new_n26134__ = ~new_new_n26131__ & new_new_n26133__;
  assign new_new_n26135__ = ~new_new_n26128__ & ~new_new_n26134__;
  assign new_new_n26136__ = new_new_n25157__ & new_new_n25192__;
  assign new_new_n26137__ = ~new_new_n25196__ & ~new_new_n26136__;
  assign new_new_n26138__ = ~new_new_n25169__ & ~new_new_n26137__;
  assign new_new_n26139__ = new_new_n25193__ & ~new_new_n25195__;
  assign new_new_n26140__ = ~new_new_n26138__ & ~new_new_n26139__;
  assign new_new_n26141__ = ~new_new_n26125__ & ~new_new_n26140__;
  assign new_new_n26142__ = ~new_new_n25196__ & ~new_new_n25312__;
  assign new_new_n26143__ = new_new_n26131__ & ~new_new_n26142__;
  assign new_new_n26144__ = ~new_new_n26141__ & ~new_new_n26143__;
  assign new_new_n26145__ = ~new_new_n25305__ & ~new_new_n25309__;
  assign new_new_n26146__ = ~new_new_n26144__ & ~new_new_n26145__;
  assign new_new_n26147__ = ~new_new_n25302__ & ~new_new_n25309__;
  assign new_new_n26148__ = ~new_new_n15905__ & ~new_new_n25292__;
  assign new_new_n26149__ = new_new_n15917__ & new_new_n25295__;
  assign new_new_n26150__ = new_new_n12798__ & new_new_n15244__;
  assign new_new_n26151__ = pi01 & new_new_n15237__;
  assign new_new_n26152__ = ~pi00 & ~new_new_n26150__;
  assign new_new_n26153__ = ~new_new_n26151__ & new_new_n26152__;
  assign new_new_n26154__ = ~new_new_n26148__ & ~new_new_n26153__;
  assign new_new_n26155__ = ~new_new_n26149__ & new_new_n26154__;
  assign new_new_n26156__ = ~new_new_n25303__ & new_new_n26155__;
  assign new_new_n26157__ = ~new_new_n26147__ & new_new_n26156__;
  assign new_new_n26158__ = new_new_n25302__ & ~new_new_n25309__;
  assign new_new_n26159__ = ~new_new_n25304__ & ~new_new_n26155__;
  assign new_new_n26160__ = ~new_new_n26158__ & new_new_n26159__;
  assign new_new_n26161__ = ~new_new_n26146__ & ~new_new_n26157__;
  assign new_new_n26162__ = ~new_new_n26160__ & new_new_n26161__;
  assign new_new_n26163__ = new_new_n26135__ & ~new_new_n26162__;
  assign new_new_n26164__ = ~new_new_n25310__ & ~new_new_n26163__;
  assign new_new_n26165__ = new_new_n25289__ & ~new_new_n26164__;
  assign new_new_n26166__ = ~new_new_n25289__ & new_new_n26164__;
  assign new_new_n26167__ = ~new_new_n25214__ & ~new_new_n25215__;
  assign new_new_n26168__ = new_new_n25229__ & new_new_n26167__;
  assign new_new_n26169__ = ~new_new_n25229__ & ~new_new_n26167__;
  assign new_new_n26170__ = ~new_new_n26168__ & ~new_new_n26169__;
  assign new_new_n26171__ = ~new_new_n26166__ & ~new_new_n26170__;
  assign new_new_n26172__ = ~new_new_n26165__ & ~new_new_n26171__;
  assign new_new_n26173__ = new_new_n25276__ & ~new_new_n26172__;
  assign new_new_n26174__ = ~new_new_n25276__ & new_new_n26172__;
  assign new_new_n26175__ = ~new_new_n25236__ & ~new_new_n25237__;
  assign new_new_n26176__ = new_new_n25250__ & ~new_new_n26175__;
  assign new_new_n26177__ = ~new_new_n25250__ & new_new_n26175__;
  assign new_new_n26178__ = ~new_new_n26176__ & ~new_new_n26177__;
  assign new_new_n26179__ = ~new_new_n26174__ & new_new_n26178__;
  assign new_new_n26180__ = ~new_new_n26173__ & ~new_new_n26179__;
  assign new_new_n26181__ = ~new_new_n25263__ & ~new_new_n26180__;
  assign new_new_n26182__ = new_new_n14393__ & new_new_n16056__;
  assign new_new_n26183__ = ~new_new_n26181__ & new_new_n26182__;
  assign new_new_n26184__ = pi02 & ~new_new_n25262__;
  assign new_new_n26185__ = new_new_n26180__ & ~new_new_n26184__;
  assign new_new_n26186__ = new_new_n18146__ & new_new_n25262__;
  assign new_new_n26187__ = ~new_new_n26185__ & ~new_new_n26186__;
  assign new_new_n26188__ = ~new_new_n26183__ & new_new_n26187__;
  assign new_new_n26189__ = ~new_new_n25253__ & ~new_new_n25259__;
  assign new_new_n26190__ = ~new_new_n25254__ & ~new_new_n26189__;
  assign new_new_n26191__ = ~new_new_n26188__ & ~new_new_n26190__;
  assign new_new_n26192__ = new_new_n11471__ & new_new_n15905__;
  assign new_new_n26193__ = new_new_n11475__ & ~new_new_n15998__;
  assign new_new_n26194__ = new_new_n11478__ & new_new_n16051__;
  assign new_new_n26195__ = ~new_new_n11482__ & ~new_new_n16056__;
  assign new_new_n26196__ = ~new_new_n26194__ & new_new_n26195__;
  assign new_new_n26197__ = ~new_new_n26192__ & ~new_new_n26193__;
  assign new_new_n26198__ = ~new_new_n26196__ & new_new_n26197__;
  assign new_new_n26199__ = pi05 & ~new_new_n26198__;
  assign new_new_n26200__ = ~pi05 & new_new_n26198__;
  assign new_new_n26201__ = ~new_new_n26199__ & ~new_new_n26200__;
  assign new_new_n26202__ = ~new_new_n24492__ & ~new_new_n24493__;
  assign new_new_n26203__ = new_new_n24503__ & new_new_n26202__;
  assign new_new_n26204__ = ~new_new_n24503__ & ~new_new_n26202__;
  assign new_new_n26205__ = ~new_new_n26203__ & ~new_new_n26204__;
  assign new_new_n26206__ = ~new_new_n26201__ & ~new_new_n26205__;
  assign new_new_n26207__ = new_new_n26201__ & new_new_n26205__;
  assign new_new_n26208__ = ~new_new_n18146__ & ~new_new_n26207__;
  assign new_new_n26209__ = ~new_new_n26206__ & ~new_new_n26208__;
  assign new_new_n26210__ = ~new_new_n26191__ & ~new_new_n26209__;
  assign new_new_n26211__ = ~new_new_n24510__ & ~new_new_n24511__;
  assign new_new_n26212__ = new_new_n24520__ & new_new_n26211__;
  assign new_new_n26213__ = ~new_new_n24520__ & ~new_new_n26211__;
  assign new_new_n26214__ = ~new_new_n26212__ & ~new_new_n26213__;
  assign new_new_n26215__ = ~new_new_n26210__ & new_new_n26214__;
  assign new_new_n26216__ = new_new_n26188__ & new_new_n26190__;
  assign new_new_n26217__ = new_new_n18146__ & new_new_n26207__;
  assign new_new_n26218__ = ~new_new_n18146__ & new_new_n26206__;
  assign new_new_n26219__ = new_new_n26214__ & ~new_new_n26218__;
  assign new_new_n26220__ = ~new_new_n26217__ & ~new_new_n26219__;
  assign new_new_n26221__ = ~new_new_n26216__ & ~new_new_n26220__;
  assign new_new_n26222__ = new_new_n26191__ & new_new_n26209__;
  assign new_new_n26223__ = ~new_new_n26221__ & ~new_new_n26222__;
  assign new_new_n26224__ = ~new_new_n26215__ & new_new_n26223__;
  assign new_new_n26225__ = ~new_new_n24522__ & ~new_new_n26224__;
  assign new_new_n26226__ = new_new_n23816__ & ~new_new_n26225__;
  assign new_new_n26227__ = pi05 & new_new_n16056__;
  assign new_new_n26228__ = pi03 & ~new_new_n16056__;
  assign new_new_n26229__ = new_new_n11470__ & ~new_new_n26227__;
  assign new_new_n26230__ = ~new_new_n26228__ & new_new_n26229__;
  assign new_new_n26231__ = ~new_new_n14117__ & ~new_new_n26230__;
  assign new_new_n26232__ = ~new_new_n26226__ & new_new_n26231__;
  assign new_new_n26233__ = ~new_new_n23807__ & ~new_new_n23811__;
  assign new_new_n26234__ = new_new_n24522__ & new_new_n26224__;
  assign new_new_n26235__ = ~new_new_n23816__ & ~new_new_n26234__;
  assign new_new_n26236__ = ~new_new_n26233__ & ~new_new_n26235__;
  assign new_new_n26237__ = ~new_new_n26232__ & new_new_n26236__;
  assign new_new_n26238__ = ~new_new_n23812__ & ~new_new_n23816__;
  assign new_new_n26239__ = ~new_new_n26225__ & ~new_new_n26231__;
  assign new_new_n26240__ = ~new_new_n26234__ & ~new_new_n26239__;
  assign new_new_n26241__ = ~new_new_n26238__ & ~new_new_n26240__;
  assign new_new_n26242__ = ~new_new_n23817__ & ~new_new_n26237__;
  assign new_new_n26243__ = ~new_new_n26241__ & new_new_n26242__;
  assign new_new_n26244__ = ~new_new_n23181__ & ~new_new_n26243__;
  assign new_new_n26245__ = ~new_new_n22429__ & new_new_n22454__;
  assign new_new_n26246__ = ~new_new_n22428__ & ~new_new_n26245__;
  assign new_new_n26247__ = new_new_n8474__ & new_new_n15237__;
  assign new_new_n26248__ = ~new_new_n8479__ & new_new_n15244__;
  assign new_new_n26249__ = ~new_new_n26247__ & ~new_new_n26248__;
  assign new_new_n26250__ = new_new_n8469__ & new_new_n17974__;
  assign new_new_n26251__ = new_new_n26249__ & ~new_new_n26250__;
  assign new_new_n26252__ = pi11 & ~new_new_n26251__;
  assign new_new_n26253__ = new_new_n8469__ & ~new_new_n17978__;
  assign new_new_n26254__ = ~pi11 & ~new_new_n26253__;
  assign new_new_n26255__ = ~pi10 & ~new_new_n17981__;
  assign new_new_n26256__ = pi10 & ~new_new_n17983__;
  assign new_new_n26257__ = new_new_n8469__ & ~new_new_n26255__;
  assign new_new_n26258__ = ~new_new_n26256__ & new_new_n26257__;
  assign new_new_n26259__ = ~new_new_n26254__ & ~new_new_n26258__;
  assign new_new_n26260__ = new_new_n26249__ & ~new_new_n26259__;
  assign new_new_n26261__ = ~new_new_n26252__ & ~new_new_n26260__;
  assign new_new_n26262__ = ~new_new_n21353__ & ~new_new_n21354__;
  assign new_new_n26263__ = ~new_new_n21358__ & new_new_n26262__;
  assign new_new_n26264__ = new_new_n21358__ & ~new_new_n26262__;
  assign new_new_n26265__ = ~new_new_n26263__ & ~new_new_n26264__;
  assign new_new_n26266__ = new_new_n26261__ & new_new_n26265__;
  assign new_new_n26267__ = ~new_new_n26261__ & ~new_new_n26265__;
  assign new_new_n26268__ = ~new_new_n26266__ & ~new_new_n26267__;
  assign new_new_n26269__ = ~new_new_n22438__ & ~new_new_n22451__;
  assign new_new_n26270__ = ~new_new_n22437__ & ~new_new_n26269__;
  assign new_new_n26271__ = new_new_n26268__ & ~new_new_n26270__;
  assign new_new_n26272__ = ~new_new_n26268__ & new_new_n26270__;
  assign new_new_n26273__ = ~new_new_n26271__ & ~new_new_n26272__;
  assign new_new_n26274__ = new_new_n26246__ & ~new_new_n26273__;
  assign new_new_n26275__ = ~new_new_n26246__ & new_new_n26273__;
  assign new_new_n26276__ = ~new_new_n11409__ & ~new_new_n15998__;
  assign new_new_n26277__ = new_new_n10702__ & ~new_new_n16056__;
  assign new_new_n26278__ = ~new_new_n10698__ & ~new_new_n26277__;
  assign new_new_n26279__ = ~new_new_n26276__ & new_new_n26278__;
  assign new_new_n26280__ = new_new_n10694__ & new_new_n16630__;
  assign new_new_n26281__ = ~pi08 & ~new_new_n26280__;
  assign new_new_n26282__ = new_new_n12121__ & new_new_n16630__;
  assign new_new_n26283__ = ~new_new_n26281__ & ~new_new_n26282__;
  assign new_new_n26284__ = new_new_n26279__ & ~new_new_n26283__;
  assign new_new_n26285__ = pi08 & ~new_new_n26279__;
  assign new_new_n26286__ = ~new_new_n26284__ & ~new_new_n26285__;
  assign new_new_n26287__ = ~new_new_n26275__ & ~new_new_n26286__;
  assign new_new_n26288__ = ~new_new_n26274__ & ~new_new_n26287__;
  assign new_new_n26289__ = ~new_new_n26244__ & new_new_n26288__;
  assign new_new_n26290__ = ~new_new_n26267__ & ~new_new_n26270__;
  assign new_new_n26291__ = ~new_new_n26266__ & ~new_new_n26290__;
  assign new_new_n26292__ = ~new_new_n21365__ & ~new_new_n21366__;
  assign new_new_n26293__ = new_new_n21378__ & ~new_new_n26292__;
  assign new_new_n26294__ = ~new_new_n21378__ & new_new_n26292__;
  assign new_new_n26295__ = ~new_new_n26293__ & ~new_new_n26294__;
  assign new_new_n26296__ = ~new_new_n26291__ & new_new_n26295__;
  assign new_new_n26297__ = new_new_n26291__ & ~new_new_n26295__;
  assign new_new_n26298__ = ~new_new_n26296__ & ~new_new_n26297__;
  assign new_new_n26299__ = new_new_n10712__ & new_new_n16056__;
  assign new_new_n26300__ = ~new_new_n10709__ & ~new_new_n26299__;
  assign new_new_n26301__ = pi08 & new_new_n16056__;
  assign new_new_n26302__ = ~new_new_n10694__ & ~new_new_n26301__;
  assign new_new_n26303__ = ~new_new_n26300__ & new_new_n26302__;
  assign new_new_n26304__ = ~new_new_n13064__ & ~new_new_n26303__;
  assign new_new_n26305__ = new_new_n26298__ & ~new_new_n26304__;
  assign new_new_n26306__ = ~new_new_n26298__ & new_new_n26304__;
  assign new_new_n26307__ = ~new_new_n26305__ & ~new_new_n26306__;
  assign new_new_n26308__ = ~new_new_n26289__ & new_new_n26307__;
  assign new_new_n26309__ = new_new_n26275__ & new_new_n26286__;
  assign new_new_n26310__ = new_new_n23181__ & new_new_n26243__;
  assign new_new_n26311__ = new_new_n26274__ & ~new_new_n26286__;
  assign new_new_n26312__ = ~new_new_n26307__ & ~new_new_n26311__;
  assign new_new_n26313__ = ~new_new_n26309__ & ~new_new_n26312__;
  assign new_new_n26314__ = ~new_new_n26310__ & new_new_n26313__;
  assign new_new_n26315__ = new_new_n26244__ & ~new_new_n26288__;
  assign new_new_n26316__ = ~new_new_n26314__ & ~new_new_n26315__;
  assign new_new_n26317__ = ~new_new_n26308__ & new_new_n26316__;
  assign new_new_n26318__ = ~new_new_n21383__ & ~new_new_n26317__;
  assign new_new_n26319__ = new_new_n21383__ & new_new_n26317__;
  assign new_new_n26320__ = ~new_new_n26296__ & ~new_new_n26304__;
  assign new_new_n26321__ = ~new_new_n26297__ & ~new_new_n26320__;
  assign new_new_n26322__ = ~new_new_n26319__ & ~new_new_n26321__;
  assign new_new_n26323__ = ~new_new_n26318__ & ~new_new_n26322__;
  assign new_new_n26324__ = ~new_new_n20881__ & ~new_new_n21380__;
  assign new_new_n26325__ = ~new_new_n20882__ & ~new_new_n26324__;
  assign new_new_n26326__ = new_new_n26323__ & ~new_new_n26325__;
  assign new_new_n26327__ = ~new_new_n20871__ & ~new_new_n20877__;
  assign new_new_n26328__ = ~new_new_n20878__ & ~new_new_n26327__;
  assign new_new_n26329__ = ~new_new_n20413__ & ~new_new_n20414__;
  assign new_new_n26330__ = new_new_n20429__ & new_new_n26329__;
  assign new_new_n26331__ = ~new_new_n20429__ & ~new_new_n26329__;
  assign new_new_n26332__ = ~new_new_n26330__ & ~new_new_n26331__;
  assign new_new_n26333__ = new_new_n26328__ & ~new_new_n26332__;
  assign new_new_n26334__ = ~new_new_n26328__ & new_new_n26332__;
  assign new_new_n26335__ = ~new_new_n8479__ & ~new_new_n15998__;
  assign new_new_n26336__ = new_new_n8474__ & ~new_new_n16056__;
  assign new_new_n26337__ = ~new_new_n8858__ & ~new_new_n26336__;
  assign new_new_n26338__ = ~new_new_n26335__ & new_new_n26337__;
  assign new_new_n26339__ = new_new_n8469__ & new_new_n16630__;
  assign new_new_n26340__ = pi11 & ~new_new_n26339__;
  assign new_new_n26341__ = new_new_n11530__ & new_new_n16630__;
  assign new_new_n26342__ = ~new_new_n26340__ & ~new_new_n26341__;
  assign new_new_n26343__ = new_new_n26338__ & ~new_new_n26342__;
  assign new_new_n26344__ = ~pi11 & ~new_new_n26338__;
  assign new_new_n26345__ = ~new_new_n26343__ & ~new_new_n26344__;
  assign new_new_n26346__ = ~new_new_n26334__ & ~new_new_n26345__;
  assign new_new_n26347__ = ~new_new_n26333__ & ~new_new_n26346__;
  assign new_new_n26348__ = ~new_new_n26326__ & new_new_n26347__;
  assign new_new_n26349__ = ~new_new_n20006__ & ~new_new_n20007__;
  assign new_new_n26350__ = new_new_n20431__ & new_new_n26349__;
  assign new_new_n26351__ = ~new_new_n20431__ & ~new_new_n26349__;
  assign new_new_n26352__ = ~new_new_n26350__ & ~new_new_n26351__;
  assign new_new_n26353__ = ~new_new_n26348__ & ~new_new_n26352__;
  assign new_new_n26354__ = ~new_new_n26334__ & ~new_new_n26352__;
  assign new_new_n26355__ = new_new_n26345__ & ~new_new_n26354__;
  assign new_new_n26356__ = ~new_new_n26323__ & new_new_n26325__;
  assign new_new_n26357__ = ~new_new_n26333__ & new_new_n26352__;
  assign new_new_n26358__ = ~new_new_n26355__ & ~new_new_n26357__;
  assign new_new_n26359__ = ~new_new_n26356__ & new_new_n26358__;
  assign new_new_n26360__ = new_new_n26326__ & ~new_new_n26347__;
  assign new_new_n26361__ = ~new_new_n26359__ & ~new_new_n26360__;
  assign new_new_n26362__ = ~new_new_n26353__ & new_new_n26361__;
  assign new_new_n26363__ = ~new_new_n20433__ & ~new_new_n26362__;
  assign new_new_n26364__ = new_new_n20433__ & new_new_n26362__;
  assign new_new_n26365__ = ~new_new_n19981__ & ~new_new_n19982__;
  assign new_new_n26366__ = new_new_n17447__ & ~new_new_n26365__;
  assign new_new_n26367__ = ~new_new_n17447__ & new_new_n26365__;
  assign new_new_n26368__ = ~new_new_n26366__ & ~new_new_n26367__;
  assign new_new_n26369__ = ~new_new_n26364__ & new_new_n26368__;
  assign new_new_n26370__ = ~new_new_n26363__ & ~new_new_n26369__;
  assign new_new_n26371__ = new_new_n19666__ & ~new_new_n19818__;
  assign new_new_n26372__ = ~new_new_n19817__ & ~new_new_n26371__;
  assign new_new_n26373__ = ~new_new_n26370__ & new_new_n26372__;
  assign new_new_n26374__ = ~new_new_n18860__ & ~new_new_n18861__;
  assign new_new_n26375__ = ~new_new_n19649__ & new_new_n26374__;
  assign new_new_n26376__ = new_new_n19649__ & ~new_new_n26374__;
  assign new_new_n26377__ = ~new_new_n26375__ & ~new_new_n26376__;
  assign new_new_n26378__ = ~new_new_n26373__ & new_new_n26377__;
  assign new_new_n26379__ = ~new_new_n19989__ & ~new_new_n26378__;
  assign new_new_n26380__ = ~new_new_n19662__ & new_new_n26379__;
  assign new_new_n26381__ = new_new_n26370__ & ~new_new_n26372__;
  assign new_new_n26382__ = ~new_new_n19989__ & ~new_new_n26377__;
  assign new_new_n26383__ = new_new_n19662__ & ~new_new_n26382__;
  assign new_new_n26384__ = ~new_new_n26381__ & ~new_new_n26383__;
  assign new_new_n26385__ = ~new_new_n26373__ & ~new_new_n26384__;
  assign new_new_n26386__ = ~new_new_n26377__ & ~new_new_n26385__;
  assign new_new_n26387__ = ~new_new_n26379__ & ~new_new_n26384__;
  assign new_new_n26388__ = ~new_new_n19984__ & ~new_new_n19988__;
  assign new_new_n26389__ = ~new_new_n26387__ & new_new_n26388__;
  assign new_new_n26390__ = ~new_new_n26380__ & ~new_new_n26386__;
  assign new_new_n26391__ = ~new_new_n26389__ & new_new_n26390__;
  assign new_new_n26392__ = new_new_n19651__ & ~new_new_n26391__;
  assign new_new_n26393__ = ~new_new_n18851__ & new_new_n18856__;
  assign new_new_n26394__ = ~new_new_n18850__ & ~new_new_n26393__;
  assign new_new_n26395__ = new_new_n18358__ & ~new_new_n18661__;
  assign new_new_n26396__ = ~new_new_n18358__ & new_new_n18661__;
  assign new_new_n26397__ = ~new_new_n26395__ & ~new_new_n26396__;
  assign new_new_n26398__ = new_new_n18316__ & ~new_new_n18335__;
  assign new_new_n26399__ = ~new_new_n18316__ & new_new_n18335__;
  assign new_new_n26400__ = ~new_new_n26398__ & ~new_new_n26399__;
  assign new_new_n26401__ = new_new_n26397__ & new_new_n26400__;
  assign new_new_n26402__ = ~new_new_n26397__ & ~new_new_n26400__;
  assign new_new_n26403__ = ~new_new_n26401__ & ~new_new_n26402__;
  assign new_new_n26404__ = ~new_new_n26394__ & new_new_n26403__;
  assign new_new_n26405__ = new_new_n26394__ & ~new_new_n26403__;
  assign new_new_n26406__ = new_new_n16844__ & ~new_new_n26405__;
  assign new_new_n26407__ = ~new_new_n26404__ & ~new_new_n26406__;
  assign new_new_n26408__ = ~new_new_n26392__ & ~new_new_n26407__;
  assign new_new_n26409__ = ~new_new_n18666__ & ~new_new_n18667__;
  assign new_new_n26410__ = ~new_new_n18676__ & new_new_n26409__;
  assign new_new_n26411__ = new_new_n18676__ & ~new_new_n26409__;
  assign new_new_n26412__ = ~new_new_n26410__ & ~new_new_n26411__;
  assign new_new_n26413__ = ~new_new_n26408__ & ~new_new_n26412__;
  assign new_new_n26414__ = new_new_n16844__ & new_new_n26404__;
  assign new_new_n26415__ = ~new_new_n19651__ & new_new_n26391__;
  assign new_new_n26416__ = ~new_new_n16844__ & new_new_n26405__;
  assign new_new_n26417__ = new_new_n26412__ & ~new_new_n26416__;
  assign new_new_n26418__ = ~new_new_n26414__ & ~new_new_n26417__;
  assign new_new_n26419__ = ~new_new_n26415__ & new_new_n26418__;
  assign new_new_n26420__ = new_new_n26392__ & new_new_n26407__;
  assign new_new_n26421__ = ~new_new_n26419__ & ~new_new_n26420__;
  assign new_new_n26422__ = ~new_new_n26413__ & new_new_n26421__;
  assign new_new_n26423__ = ~new_new_n18716__ & ~new_new_n26422__;
  assign new_new_n26424__ = new_new_n18711__ & ~new_new_n26423__;
  assign new_new_n26425__ = pi17 & new_new_n16056__;
  assign new_new_n26426__ = new_new_n10340__ & new_new_n16056__;
  assign new_new_n26427__ = ~new_new_n10337__ & ~new_new_n26426__;
  assign new_new_n26428__ = ~new_new_n6958__ & ~new_new_n26425__;
  assign new_new_n26429__ = ~new_new_n26427__ & new_new_n26428__;
  assign new_new_n26430__ = pi17 & new_new_n6963__;
  assign new_new_n26431__ = ~new_new_n26429__ & ~new_new_n26430__;
  assign new_new_n26432__ = ~new_new_n26424__ & new_new_n26431__;
  assign new_new_n26433__ = ~new_new_n18340__ & new_new_n18678__;
  assign new_new_n26434__ = new_new_n18716__ & new_new_n26422__;
  assign new_new_n26435__ = ~new_new_n18711__ & ~new_new_n26434__;
  assign new_new_n26436__ = ~new_new_n26433__ & ~new_new_n26435__;
  assign new_new_n26437__ = ~new_new_n26432__ & new_new_n26436__;
  assign new_new_n26438__ = ~new_new_n18679__ & ~new_new_n18711__;
  assign new_new_n26439__ = ~new_new_n26423__ & ~new_new_n26431__;
  assign new_new_n26440__ = ~new_new_n26434__ & ~new_new_n26439__;
  assign new_new_n26441__ = ~new_new_n26438__ & ~new_new_n26440__;
  assign new_new_n26442__ = ~new_new_n18712__ & ~new_new_n26437__;
  assign new_new_n26443__ = ~new_new_n26441__ & new_new_n26442__;
  assign new_new_n26444__ = ~new_new_n17970__ & ~new_new_n26443__;
  assign new_new_n26445__ = ~new_new_n17343__ & ~new_new_n17344__;
  assign new_new_n26446__ = new_new_n17736__ & new_new_n26445__;
  assign new_new_n26447__ = ~new_new_n17736__ & ~new_new_n26445__;
  assign new_new_n26448__ = ~new_new_n26446__ & ~new_new_n26447__;
  assign new_new_n26449__ = new_new_n26444__ & ~new_new_n26448__;
  assign new_new_n26450__ = ~new_new_n17719__ & ~new_new_n17720__;
  assign new_new_n26451__ = new_new_n17734__ & ~new_new_n26450__;
  assign new_new_n26452__ = ~new_new_n17734__ & new_new_n26450__;
  assign new_new_n26453__ = ~new_new_n26451__ & ~new_new_n26452__;
  assign new_new_n26454__ = ~new_new_n18702__ & ~new_new_n18708__;
  assign new_new_n26455__ = ~new_new_n18703__ & ~new_new_n26454__;
  assign new_new_n26456__ = new_new_n26453__ & ~new_new_n26455__;
  assign new_new_n26457__ = new_new_n6629__ & ~new_new_n16056__;
  assign new_new_n26458__ = ~new_new_n6633__ & ~new_new_n16630__;
  assign new_new_n26459__ = new_new_n6631__ & ~new_new_n26458__;
  assign new_new_n26460__ = ~new_new_n26457__ & ~new_new_n26459__;
  assign new_new_n26461__ = new_new_n9797__ & ~new_new_n15998__;
  assign new_new_n26462__ = pi20 & ~new_new_n26461__;
  assign new_new_n26463__ = ~pi17 & ~new_new_n26462__;
  assign new_new_n26464__ = new_new_n9800__ & ~new_new_n15998__;
  assign new_new_n26465__ = ~pi20 & ~new_new_n26464__;
  assign new_new_n26466__ = ~new_new_n26463__ & ~new_new_n26465__;
  assign new_new_n26467__ = new_new_n26460__ & ~new_new_n26466__;
  assign new_new_n26468__ = pi20 & ~new_new_n26460__;
  assign new_new_n26469__ = ~new_new_n26467__ & ~new_new_n26468__;
  assign new_new_n26470__ = ~new_new_n26456__ & new_new_n26469__;
  assign new_new_n26471__ = ~new_new_n26444__ & new_new_n26448__;
  assign new_new_n26472__ = ~new_new_n26453__ & new_new_n26455__;
  assign new_new_n26473__ = ~new_new_n26470__ & ~new_new_n26472__;
  assign new_new_n26474__ = ~new_new_n26471__ & new_new_n26473__;
  assign new_new_n26475__ = new_new_n26469__ & new_new_n26472__;
  assign new_new_n26476__ = new_new_n26456__ & ~new_new_n26469__;
  assign new_new_n26477__ = new_new_n26448__ & ~new_new_n26476__;
  assign new_new_n26478__ = new_new_n17970__ & new_new_n26443__;
  assign new_new_n26479__ = ~new_new_n26475__ & ~new_new_n26477__;
  assign new_new_n26480__ = ~new_new_n26478__ & new_new_n26479__;
  assign new_new_n26481__ = ~new_new_n26449__ & ~new_new_n26480__;
  assign new_new_n26482__ = ~new_new_n26474__ & new_new_n26481__;
  assign new_new_n26483__ = new_new_n17868__ & ~new_new_n26482__;
  assign new_new_n26484__ = new_new_n17864__ & ~new_new_n26483__;
  assign new_new_n26485__ = new_new_n16185__ & ~new_new_n26484__;
  assign new_new_n26486__ = ~new_new_n17868__ & new_new_n26482__;
  assign new_new_n26487__ = ~new_new_n17864__ & ~new_new_n26486__;
  assign new_new_n26488__ = ~new_new_n17866__ & ~new_new_n26487__;
  assign new_new_n26489__ = ~new_new_n26485__ & new_new_n26488__;
  assign new_new_n26490__ = ~new_new_n17820__ & ~new_new_n17864__;
  assign new_new_n26491__ = ~new_new_n16185__ & ~new_new_n26483__;
  assign new_new_n26492__ = ~new_new_n26486__ & ~new_new_n26491__;
  assign new_new_n26493__ = ~new_new_n26490__ & ~new_new_n26492__;
  assign new_new_n26494__ = ~new_new_n17865__ & ~new_new_n26489__;
  assign new_new_n26495__ = ~new_new_n26493__ & new_new_n26494__;
  assign new_new_n26496__ = ~new_new_n17851__ & ~new_new_n17861__;
  assign new_new_n26497__ = ~new_new_n17850__ & ~new_new_n26496__;
  assign new_new_n26498__ = ~new_new_n26495__ & new_new_n26497__;
  assign new_new_n26499__ = ~new_new_n16695__ & ~new_new_n16696__;
  assign new_new_n26500__ = new_new_n16993__ & ~new_new_n26499__;
  assign new_new_n26501__ = ~new_new_n16993__ & new_new_n26499__;
  assign new_new_n26502__ = ~new_new_n26500__ & ~new_new_n26501__;
  assign new_new_n26503__ = ~new_new_n17840__ & ~new_new_n17846__;
  assign new_new_n26504__ = ~new_new_n17841__ & ~new_new_n26503__;
  assign new_new_n26505__ = ~new_new_n26502__ & ~new_new_n26504__;
  assign new_new_n26506__ = new_new_n26502__ & new_new_n26504__;
  assign new_new_n26507__ = ~new_new_n5195__ & ~new_new_n21064__;
  assign new_new_n26508__ = pi23 & ~new_new_n26507__;
  assign new_new_n26509__ = pi21 & ~new_new_n16056__;
  assign new_new_n26510__ = pi23 & new_new_n16056__;
  assign new_new_n26511__ = new_new_n26507__ & ~new_new_n26509__;
  assign new_new_n26512__ = ~new_new_n26510__ & new_new_n26511__;
  assign new_new_n26513__ = ~new_new_n26508__ & ~new_new_n26512__;
  assign new_new_n26514__ = ~new_new_n26506__ & ~new_new_n26513__;
  assign new_new_n26515__ = ~new_new_n26505__ & ~new_new_n26514__;
  assign new_new_n26516__ = ~new_new_n26498__ & ~new_new_n26515__;
  assign new_new_n26517__ = ~new_new_n16996__ & ~new_new_n16997__;
  assign new_new_n26518__ = ~new_new_n16999__ & ~new_new_n26517__;
  assign new_new_n26519__ = new_new_n16999__ & new_new_n26517__;
  assign new_new_n26520__ = ~new_new_n26518__ & ~new_new_n26519__;
  assign new_new_n26521__ = ~new_new_n26516__ & ~new_new_n26520__;
  assign new_new_n26522__ = new_new_n26495__ & ~new_new_n26497__;
  assign new_new_n26523__ = new_new_n26506__ & new_new_n26513__;
  assign new_new_n26524__ = new_new_n26505__ & ~new_new_n26513__;
  assign new_new_n26525__ = ~new_new_n26520__ & ~new_new_n26524__;
  assign new_new_n26526__ = ~new_new_n26523__ & ~new_new_n26525__;
  assign new_new_n26527__ = ~new_new_n26522__ & ~new_new_n26526__;
  assign new_new_n26528__ = new_new_n26498__ & new_new_n26515__;
  assign new_new_n26529__ = ~new_new_n26527__ & ~new_new_n26528__;
  assign new_new_n26530__ = ~new_new_n26521__ & new_new_n26529__;
  assign new_new_n26531__ = ~new_new_n17003__ & new_new_n26530__;
  assign new_new_n26532__ = ~new_new_n17002__ & ~new_new_n26531__;
  assign new_new_n26533__ = new_new_n16624__ & new_new_n16661__;
  assign new_new_n26534__ = new_new_n16667__ & ~new_new_n26533__;
  assign new_new_n26535__ = ~new_new_n16624__ & ~new_new_n16661__;
  assign new_new_n26536__ = ~new_new_n26534__ & ~new_new_n26535__;
  assign new_new_n26537__ = new_new_n26532__ & ~new_new_n26536__;
  assign new_new_n26538__ = ~new_new_n16654__ & ~new_new_n16658__;
  assign new_new_n26539__ = ~new_new_n16655__ & ~new_new_n26538__;
  assign new_new_n26540__ = ~new_new_n16384__ & ~new_new_n16388__;
  assign new_new_n26541__ = ~new_new_n15960__ & new_new_n16397__;
  assign new_new_n26542__ = new_new_n15960__ & ~new_new_n16397__;
  assign new_new_n26543__ = ~new_new_n26541__ & ~new_new_n26542__;
  assign new_new_n26544__ = new_new_n26540__ & new_new_n26543__;
  assign new_new_n26545__ = ~new_new_n26540__ & ~new_new_n26543__;
  assign new_new_n26546__ = ~new_new_n26544__ & ~new_new_n26545__;
  assign new_new_n26547__ = new_new_n26539__ & ~new_new_n26546__;
  assign new_new_n26548__ = ~new_new_n26539__ & new_new_n26546__;
  assign new_new_n26549__ = ~pi26 & ~new_new_n16056__;
  assign new_new_n26550__ = ~new_new_n272__ & ~new_new_n26549__;
  assign new_new_n26551__ = pi23 & ~new_new_n26550__;
  assign new_new_n26552__ = new_new_n145__ & new_new_n16056__;
  assign new_new_n26553__ = new_new_n15928__ & ~new_new_n26552__;
  assign new_new_n26554__ = ~new_new_n429__ & ~new_new_n19220__;
  assign new_new_n26555__ = new_new_n16056__ & new_new_n26554__;
  assign new_new_n26556__ = ~new_new_n26553__ & ~new_new_n26555__;
  assign new_new_n26557__ = ~new_new_n26551__ & new_new_n26556__;
  assign new_new_n26558__ = ~new_new_n26548__ & new_new_n26557__;
  assign new_new_n26559__ = ~new_new_n26547__ & ~new_new_n26558__;
  assign new_new_n26560__ = ~new_new_n26537__ & ~new_new_n26559__;
  assign new_new_n26561__ = new_new_n15929__ & ~new_new_n16408__;
  assign new_new_n26562__ = ~new_new_n15929__ & new_new_n16408__;
  assign new_new_n26563__ = ~new_new_n26561__ & ~new_new_n26562__;
  assign new_new_n26564__ = ~new_new_n4818__ & new_new_n15905__;
  assign new_new_n26565__ = pi29 & new_new_n26564__;
  assign new_new_n26566__ = ~new_new_n16413__ & ~new_new_n26564__;
  assign new_new_n26567__ = ~new_new_n26565__ & ~new_new_n26566__;
  assign new_new_n26568__ = new_new_n26563__ & new_new_n26567__;
  assign new_new_n26569__ = new_new_n16414__ & ~new_new_n26563__;
  assign new_new_n26570__ = new_new_n16061__ & new_new_n26561__;
  assign new_new_n26571__ = new_new_n26562__ & new_new_n26565__;
  assign new_new_n26572__ = ~new_new_n26570__ & ~new_new_n26571__;
  assign new_new_n26573__ = ~new_new_n26568__ & new_new_n26572__;
  assign new_new_n26574__ = ~new_new_n26569__ & new_new_n26573__;
  assign new_new_n26575__ = ~new_new_n26560__ & ~new_new_n26574__;
  assign new_new_n26576__ = new_new_n26547__ & new_new_n26557__;
  assign new_new_n26577__ = ~new_new_n26532__ & new_new_n26536__;
  assign new_new_n26578__ = new_new_n26548__ & ~new_new_n26557__;
  assign new_new_n26579__ = new_new_n26574__ & ~new_new_n26578__;
  assign new_new_n26580__ = ~new_new_n26576__ & ~new_new_n26579__;
  assign new_new_n26581__ = ~new_new_n26577__ & new_new_n26580__;
  assign new_new_n26582__ = new_new_n26537__ & new_new_n26559__;
  assign new_new_n26583__ = ~new_new_n26581__ & ~new_new_n26582__;
  assign new_new_n26584__ = ~new_new_n26575__ & new_new_n26583__;
  assign new_new_n26585__ = new_new_n16419__ & ~new_new_n26584__;
  assign new_new_n26586__ = new_new_n15960__ & ~new_new_n16366__;
  assign new_new_n26587__ = new_new_n16383__ & new_new_n26586__;
  assign new_new_n26588__ = ~new_new_n15960__ & new_new_n16366__;
  assign new_new_n26589__ = ~new_new_n16383__ & new_new_n26588__;
  assign new_new_n26590__ = new_new_n16356__ & ~new_new_n26589__;
  assign new_new_n26591__ = ~new_new_n16383__ & ~new_new_n26586__;
  assign new_new_n26592__ = ~new_new_n26588__ & ~new_new_n26591__;
  assign new_new_n26593__ = ~new_new_n26590__ & ~new_new_n26592__;
  assign new_new_n26594__ = ~new_new_n16369__ & ~new_new_n26593__;
  assign new_new_n26595__ = new_new_n16356__ & new_new_n26592__;
  assign new_new_n26596__ = ~new_new_n26587__ & ~new_new_n26595__;
  assign new_new_n26597__ = ~new_new_n26594__ & new_new_n26596__;
  assign new_new_n26598__ = new_new_n16392__ & ~new_new_n26597__;
  assign new_new_n26599__ = new_new_n16356__ & new_new_n16388__;
  assign new_new_n26600__ = ~new_new_n16366__ & new_new_n26599__;
  assign new_new_n26601__ = ~new_new_n16356__ & new_new_n16384__;
  assign new_new_n26602__ = new_new_n16366__ & new_new_n26601__;
  assign new_new_n26603__ = ~new_new_n15960__ & ~new_new_n16392__;
  assign new_new_n26604__ = ~new_new_n26602__ & new_new_n26603__;
  assign new_new_n26605__ = ~new_new_n26600__ & ~new_new_n26604__;
  assign new_new_n26606__ = ~new_new_n26598__ & new_new_n26605__;
  assign new_new_n26607__ = new_new_n15923__ & new_new_n15941__;
  assign new_new_n26608__ = ~new_new_n15923__ & ~new_new_n15941__;
  assign new_new_n26609__ = ~new_new_n26607__ & ~new_new_n26608__;
  assign new_new_n26610__ = ~new_new_n15874__ & new_new_n15960__;
  assign new_new_n26611__ = ~new_new_n15925__ & ~new_new_n15960__;
  assign new_new_n26612__ = ~new_new_n26610__ & ~new_new_n26611__;
  assign new_new_n26613__ = new_new_n26609__ & ~new_new_n26612__;
  assign new_new_n26614__ = ~new_new_n26609__ & new_new_n26612__;
  assign new_new_n26615__ = ~new_new_n26613__ & ~new_new_n26614__;
  assign new_new_n26616__ = new_new_n26606__ & ~new_new_n26615__;
  assign new_new_n26617__ = ~new_new_n26606__ & new_new_n26615__;
  assign new_new_n26618__ = ~pi26 & pi29;
  assign new_new_n26619__ = pi26 & ~new_new_n16630__;
  assign new_new_n26620__ = ~pi29 & ~new_new_n26619__;
  assign new_new_n26621__ = ~pi27 & ~new_new_n26620__;
  assign new_new_n26622__ = ~pi26 & new_new_n16630__;
  assign new_new_n26623__ = pi27 & ~pi29;
  assign new_new_n26624__ = new_new_n15998__ & new_new_n26623__;
  assign new_new_n26625__ = ~new_new_n26622__ & new_new_n26624__;
  assign new_new_n26626__ = ~new_new_n26618__ & ~new_new_n26625__;
  assign new_new_n26627__ = ~new_new_n26621__ & new_new_n26626__;
  assign new_new_n26628__ = pi28 & ~new_new_n26627__;
  assign new_new_n26629__ = ~pi29 & new_new_n4221__;
  assign new_new_n26630__ = ~new_new_n3889__ & ~new_new_n16630__;
  assign new_new_n26631__ = ~pi28 & ~new_new_n26630__;
  assign new_new_n26632__ = ~new_new_n4209__ & ~new_new_n26631__;
  assign new_new_n26633__ = new_new_n4209__ & new_new_n15998__;
  assign new_new_n26634__ = pi29 & ~new_new_n26633__;
  assign new_new_n26635__ = ~new_new_n26632__ & new_new_n26634__;
  assign new_new_n26636__ = ~new_new_n26629__ & ~new_new_n26635__;
  assign new_new_n26637__ = ~new_new_n26628__ & new_new_n26636__;
  assign new_new_n26638__ = ~new_new_n26617__ & new_new_n26637__;
  assign new_new_n26639__ = ~new_new_n26616__ & ~new_new_n26638__;
  assign new_new_n26640__ = new_new_n26585__ & new_new_n26639__;
  assign new_new_n26641__ = new_new_n26617__ & ~new_new_n26637__;
  assign new_new_n26642__ = ~new_new_n16419__ & new_new_n26584__;
  assign new_new_n26643__ = ~new_new_n26585__ & ~new_new_n26642__;
  assign new_new_n26644__ = new_new_n26616__ & new_new_n26637__;
  assign new_new_n26645__ = ~new_new_n26641__ & ~new_new_n26644__;
  assign new_new_n26646__ = new_new_n26643__ & new_new_n26645__;
  assign new_new_n26647__ = ~new_new_n26639__ & new_new_n26642__;
  assign new_new_n26648__ = new_new_n16044__ & ~new_new_n26640__;
  assign new_new_n26649__ = ~new_new_n26647__ & new_new_n26648__;
  assign new_new_n26650__ = ~new_new_n26646__ & new_new_n26649__;
  assign new_new_n26651__ = new_new_n26585__ & new_new_n26606__;
  assign new_new_n26652__ = ~new_new_n26615__ & new_new_n26651__;
  assign new_new_n26653__ = ~new_new_n26585__ & ~new_new_n26606__;
  assign new_new_n26654__ = ~new_new_n26615__ & ~new_new_n26642__;
  assign new_new_n26655__ = ~new_new_n26653__ & new_new_n26654__;
  assign new_new_n26656__ = ~new_new_n26651__ & ~new_new_n26655__;
  assign new_new_n26657__ = new_new_n26637__ & ~new_new_n26656__;
  assign new_new_n26658__ = new_new_n26617__ & new_new_n26642__;
  assign new_new_n26659__ = ~new_new_n26616__ & new_new_n26642__;
  assign new_new_n26660__ = new_new_n26615__ & new_new_n26653__;
  assign new_new_n26661__ = ~new_new_n26659__ & ~new_new_n26660__;
  assign new_new_n26662__ = ~new_new_n26637__ & ~new_new_n26661__;
  assign new_new_n26663__ = ~new_new_n16044__ & ~new_new_n26658__;
  assign new_new_n26664__ = ~new_new_n26652__ & new_new_n26663__;
  assign new_new_n26665__ = ~new_new_n26657__ & new_new_n26664__;
  assign new_new_n26666__ = ~new_new_n26662__ & new_new_n26665__;
  assign new_new_n26667__ = ~new_new_n26650__ & ~new_new_n26666__;
  assign new_new_n26668__ = ~new_new_n26616__ & ~new_new_n26617__;
  assign new_new_n26669__ = ~new_new_n26637__ & new_new_n26643__;
  assign new_new_n26670__ = new_new_n26637__ & ~new_new_n26643__;
  assign new_new_n26671__ = ~new_new_n26669__ & ~new_new_n26670__;
  assign new_new_n26672__ = new_new_n26668__ & new_new_n26671__;
  assign new_new_n26673__ = ~new_new_n26668__ & ~new_new_n26671__;
  assign new_new_n26674__ = ~new_new_n26672__ & ~new_new_n26673__;
  assign new_new_n26675__ = new_new_n26559__ & ~new_new_n26577__;
  assign new_new_n26676__ = ~new_new_n26560__ & ~new_new_n26675__;
  assign new_new_n26677__ = ~new_new_n26537__ & ~new_new_n26577__;
  assign new_new_n26678__ = ~new_new_n26576__ & ~new_new_n26578__;
  assign new_new_n26679__ = new_new_n26677__ & new_new_n26678__;
  assign new_new_n26680__ = ~new_new_n26676__ & ~new_new_n26679__;
  assign new_new_n26681__ = ~new_new_n26574__ & ~new_new_n26680__;
  assign new_new_n26682__ = new_new_n26537__ & new_new_n26546__;
  assign new_new_n26683__ = ~new_new_n26539__ & new_new_n26682__;
  assign new_new_n26684__ = ~new_new_n26537__ & ~new_new_n26546__;
  assign new_new_n26685__ = ~new_new_n26539__ & ~new_new_n26577__;
  assign new_new_n26686__ = ~new_new_n26684__ & new_new_n26685__;
  assign new_new_n26687__ = ~new_new_n26682__ & ~new_new_n26686__;
  assign new_new_n26688__ = ~new_new_n26557__ & ~new_new_n26687__;
  assign new_new_n26689__ = new_new_n26547__ & new_new_n26577__;
  assign new_new_n26690__ = ~new_new_n26548__ & new_new_n26577__;
  assign new_new_n26691__ = new_new_n26539__ & new_new_n26684__;
  assign new_new_n26692__ = ~new_new_n26690__ & ~new_new_n26691__;
  assign new_new_n26693__ = new_new_n26557__ & ~new_new_n26692__;
  assign new_new_n26694__ = ~new_new_n26683__ & ~new_new_n26689__;
  assign new_new_n26695__ = ~new_new_n26688__ & new_new_n26694__;
  assign new_new_n26696__ = ~new_new_n26693__ & new_new_n26695__;
  assign new_new_n26697__ = new_new_n26574__ & ~new_new_n26696__;
  assign new_new_n26698__ = ~new_new_n26681__ & ~new_new_n26697__;
  assign new_new_n26699__ = new_new_n26515__ & ~new_new_n26522__;
  assign new_new_n26700__ = ~new_new_n26516__ & ~new_new_n26699__;
  assign new_new_n26701__ = ~new_new_n26498__ & ~new_new_n26522__;
  assign new_new_n26702__ = ~new_new_n26523__ & ~new_new_n26524__;
  assign new_new_n26703__ = new_new_n26701__ & new_new_n26702__;
  assign new_new_n26704__ = ~new_new_n26700__ & ~new_new_n26703__;
  assign new_new_n26705__ = ~new_new_n26520__ & ~new_new_n26704__;
  assign new_new_n26706__ = new_new_n26498__ & new_new_n26506__;
  assign new_new_n26707__ = new_new_n26498__ & new_new_n26504__;
  assign new_new_n26708__ = ~new_new_n26498__ & ~new_new_n26504__;
  assign new_new_n26709__ = new_new_n26502__ & ~new_new_n26522__;
  assign new_new_n26710__ = ~new_new_n26708__ & new_new_n26709__;
  assign new_new_n26711__ = ~new_new_n26707__ & ~new_new_n26710__;
  assign new_new_n26712__ = new_new_n26513__ & ~new_new_n26711__;
  assign new_new_n26713__ = ~new_new_n26506__ & new_new_n26522__;
  assign new_new_n26714__ = ~new_new_n26502__ & new_new_n26708__;
  assign new_new_n26715__ = ~new_new_n26713__ & ~new_new_n26714__;
  assign new_new_n26716__ = ~new_new_n26513__ & ~new_new_n26715__;
  assign new_new_n26717__ = new_new_n26505__ & new_new_n26522__;
  assign new_new_n26718__ = ~new_new_n26706__ & ~new_new_n26717__;
  assign new_new_n26719__ = ~new_new_n26712__ & new_new_n26718__;
  assign new_new_n26720__ = ~new_new_n26716__ & new_new_n26719__;
  assign new_new_n26721__ = new_new_n26520__ & ~new_new_n26720__;
  assign new_new_n26722__ = ~new_new_n26705__ & ~new_new_n26721__;
  assign new_new_n26723__ = ~new_new_n26505__ & ~new_new_n26506__;
  assign new_new_n26724__ = ~new_new_n26513__ & new_new_n26723__;
  assign new_new_n26725__ = new_new_n26513__ & ~new_new_n26723__;
  assign new_new_n26726__ = ~new_new_n26724__ & ~new_new_n26725__;
  assign new_new_n26727__ = ~new_new_n26701__ & new_new_n26726__;
  assign new_new_n26728__ = new_new_n26701__ & ~new_new_n26726__;
  assign new_new_n26729__ = ~new_new_n26727__ & ~new_new_n26728__;
  assign new_new_n26730__ = ~new_new_n17970__ & new_new_n26453__;
  assign new_new_n26731__ = new_new_n17970__ & ~new_new_n26453__;
  assign new_new_n26732__ = ~new_new_n26730__ & ~new_new_n26731__;
  assign new_new_n26733__ = ~new_new_n26443__ & ~new_new_n26455__;
  assign new_new_n26734__ = new_new_n26443__ & new_new_n26455__;
  assign new_new_n26735__ = ~new_new_n26733__ & ~new_new_n26734__;
  assign new_new_n26736__ = ~new_new_n26469__ & new_new_n26735__;
  assign new_new_n26737__ = new_new_n26469__ & ~new_new_n26735__;
  assign new_new_n26738__ = ~new_new_n26736__ & ~new_new_n26737__;
  assign new_new_n26739__ = new_new_n26732__ & new_new_n26738__;
  assign new_new_n26740__ = ~new_new_n26732__ & ~new_new_n26738__;
  assign new_new_n26741__ = ~new_new_n26739__ & ~new_new_n26740__;
  assign new_new_n26742__ = ~new_new_n17819__ & new_new_n17868__;
  assign new_new_n26743__ = new_new_n16185__ & new_new_n26742__;
  assign new_new_n26744__ = new_new_n17738__ & ~new_new_n26482__;
  assign new_new_n26745__ = ~new_new_n17738__ & new_new_n26482__;
  assign new_new_n26746__ = ~new_new_n26744__ & ~new_new_n26745__;
  assign new_new_n26747__ = new_new_n17819__ & ~new_new_n17868__;
  assign new_new_n26748__ = ~new_new_n16185__ & new_new_n26747__;
  assign new_new_n26749__ = ~new_new_n26743__ & ~new_new_n26748__;
  assign new_new_n26750__ = new_new_n26746__ & new_new_n26749__;
  assign new_new_n26751__ = new_new_n16185__ & ~new_new_n26747__;
  assign new_new_n26752__ = ~new_new_n26742__ & ~new_new_n26751__;
  assign new_new_n26753__ = new_new_n26745__ & ~new_new_n26752__;
  assign new_new_n26754__ = new_new_n26744__ & new_new_n26752__;
  assign new_new_n26755__ = ~new_new_n26753__ & ~new_new_n26754__;
  assign new_new_n26756__ = ~new_new_n26750__ & new_new_n26755__;
  assign new_new_n26757__ = new_new_n17864__ & ~new_new_n26756__;
  assign new_new_n26758__ = new_new_n17820__ & new_new_n26482__;
  assign new_new_n26759__ = ~new_new_n17868__ & new_new_n26758__;
  assign new_new_n26760__ = ~new_new_n17819__ & ~new_new_n26745__;
  assign new_new_n26761__ = ~new_new_n26744__ & ~new_new_n26760__;
  assign new_new_n26762__ = ~new_new_n17868__ & new_new_n26761__;
  assign new_new_n26763__ = ~new_new_n26758__ & ~new_new_n26762__;
  assign new_new_n26764__ = ~new_new_n16185__ & ~new_new_n26763__;
  assign new_new_n26765__ = new_new_n17868__ & ~new_new_n26761__;
  assign new_new_n26766__ = new_new_n17866__ & ~new_new_n26482__;
  assign new_new_n26767__ = ~new_new_n26765__ & ~new_new_n26766__;
  assign new_new_n26768__ = new_new_n16185__ & ~new_new_n26767__;
  assign new_new_n26769__ = new_new_n17866__ & new_new_n26483__;
  assign new_new_n26770__ = ~new_new_n26759__ & ~new_new_n26769__;
  assign new_new_n26771__ = ~new_new_n26764__ & new_new_n26770__;
  assign new_new_n26772__ = ~new_new_n26768__ & new_new_n26771__;
  assign new_new_n26773__ = ~new_new_n17864__ & ~new_new_n26772__;
  assign new_new_n26774__ = ~new_new_n26757__ & ~new_new_n26773__;
  assign new_new_n26775__ = new_new_n26469__ & new_new_n26731__;
  assign new_new_n26776__ = ~new_new_n26469__ & new_new_n26730__;
  assign new_new_n26777__ = ~new_new_n26775__ & ~new_new_n26776__;
  assign new_new_n26778__ = new_new_n26735__ & new_new_n26777__;
  assign new_new_n26779__ = ~new_new_n26469__ & ~new_new_n26731__;
  assign new_new_n26780__ = ~new_new_n26730__ & ~new_new_n26779__;
  assign new_new_n26781__ = new_new_n26734__ & ~new_new_n26780__;
  assign new_new_n26782__ = new_new_n26733__ & new_new_n26780__;
  assign new_new_n26783__ = ~new_new_n26781__ & ~new_new_n26782__;
  assign new_new_n26784__ = ~new_new_n26778__ & new_new_n26783__;
  assign new_new_n26785__ = ~new_new_n26448__ & ~new_new_n26784__;
  assign new_new_n26786__ = ~new_new_n26443__ & new_new_n26456__;
  assign new_new_n26787__ = ~new_new_n17970__ & new_new_n26786__;
  assign new_new_n26788__ = ~new_new_n26443__ & ~new_new_n26472__;
  assign new_new_n26789__ = ~new_new_n26456__ & ~new_new_n26788__;
  assign new_new_n26790__ = new_new_n17970__ & new_new_n26789__;
  assign new_new_n26791__ = new_new_n26443__ & new_new_n26472__;
  assign new_new_n26792__ = ~new_new_n26790__ & ~new_new_n26791__;
  assign new_new_n26793__ = new_new_n26469__ & ~new_new_n26792__;
  assign new_new_n26794__ = new_new_n17970__ & ~new_new_n26786__;
  assign new_new_n26795__ = ~new_new_n26469__ & ~new_new_n26789__;
  assign new_new_n26796__ = ~new_new_n26794__ & new_new_n26795__;
  assign new_new_n26797__ = new_new_n26472__ & new_new_n26478__;
  assign new_new_n26798__ = ~new_new_n26787__ & ~new_new_n26797__;
  assign new_new_n26799__ = ~new_new_n26796__ & new_new_n26798__;
  assign new_new_n26800__ = ~new_new_n26793__ & new_new_n26799__;
  assign new_new_n26801__ = new_new_n26448__ & ~new_new_n26800__;
  assign new_new_n26802__ = ~new_new_n26785__ & ~new_new_n26801__;
  assign new_new_n26803__ = ~new_new_n26774__ & new_new_n26802__;
  assign new_new_n26804__ = ~new_new_n26742__ & ~new_new_n26747__;
  assign new_new_n26805__ = new_new_n26746__ & ~new_new_n26804__;
  assign new_new_n26806__ = ~new_new_n26746__ & new_new_n26804__;
  assign new_new_n26807__ = ~new_new_n26805__ & ~new_new_n26806__;
  assign new_new_n26808__ = new_new_n16185__ & new_new_n26807__;
  assign new_new_n26809__ = ~new_new_n16185__ & ~new_new_n26807__;
  assign new_new_n26810__ = ~new_new_n26808__ & ~new_new_n26809__;
  assign new_new_n26811__ = ~new_new_n26729__ & ~new_new_n26810__;
  assign new_new_n26812__ = ~new_new_n18340__ & ~new_new_n18716__;
  assign new_new_n26813__ = new_new_n18340__ & new_new_n18716__;
  assign new_new_n26814__ = ~new_new_n26812__ & ~new_new_n26813__;
  assign new_new_n26815__ = new_new_n18678__ & ~new_new_n26422__;
  assign new_new_n26816__ = ~new_new_n18678__ & new_new_n26422__;
  assign new_new_n26817__ = ~new_new_n26815__ & ~new_new_n26816__;
  assign new_new_n26818__ = new_new_n26814__ & ~new_new_n26817__;
  assign new_new_n26819__ = ~new_new_n26814__ & new_new_n26817__;
  assign new_new_n26820__ = ~new_new_n26818__ & ~new_new_n26819__;
  assign new_new_n26821__ = new_new_n26431__ & new_new_n26820__;
  assign new_new_n26822__ = ~new_new_n26431__ & ~new_new_n26820__;
  assign new_new_n26823__ = ~new_new_n26821__ & ~new_new_n26822__;
  assign new_new_n26824__ = new_new_n26407__ & ~new_new_n26415__;
  assign new_new_n26825__ = ~new_new_n26408__ & ~new_new_n26824__;
  assign new_new_n26826__ = ~new_new_n26392__ & ~new_new_n26415__;
  assign new_new_n26827__ = ~new_new_n26414__ & ~new_new_n26416__;
  assign new_new_n26828__ = new_new_n26826__ & new_new_n26827__;
  assign new_new_n26829__ = new_new_n26412__ & ~new_new_n26825__;
  assign new_new_n26830__ = ~new_new_n26828__ & new_new_n26829__;
  assign new_new_n26831__ = new_new_n26404__ & new_new_n26415__;
  assign new_new_n26832__ = new_new_n26403__ & new_new_n26415__;
  assign new_new_n26833__ = ~new_new_n26403__ & ~new_new_n26415__;
  assign new_new_n26834__ = ~new_new_n26392__ & ~new_new_n26394__;
  assign new_new_n26835__ = ~new_new_n26833__ & new_new_n26834__;
  assign new_new_n26836__ = ~new_new_n26832__ & ~new_new_n26835__;
  assign new_new_n26837__ = new_new_n16844__ & ~new_new_n26836__;
  assign new_new_n26838__ = new_new_n26392__ & new_new_n26405__;
  assign new_new_n26839__ = new_new_n26392__ & ~new_new_n26404__;
  assign new_new_n26840__ = new_new_n26405__ & ~new_new_n26415__;
  assign new_new_n26841__ = ~new_new_n26839__ & ~new_new_n26840__;
  assign new_new_n26842__ = ~new_new_n16844__ & ~new_new_n26841__;
  assign new_new_n26843__ = ~new_new_n26412__ & ~new_new_n26831__;
  assign new_new_n26844__ = ~new_new_n26838__ & new_new_n26843__;
  assign new_new_n26845__ = ~new_new_n26842__ & new_new_n26844__;
  assign new_new_n26846__ = ~new_new_n26837__ & new_new_n26845__;
  assign new_new_n26847__ = ~new_new_n26830__ & ~new_new_n26846__;
  assign new_new_n26848__ = ~new_new_n26404__ & ~new_new_n26405__;
  assign new_new_n26849__ = ~new_new_n16844__ & new_new_n26848__;
  assign new_new_n26850__ = new_new_n16844__ & ~new_new_n26848__;
  assign new_new_n26851__ = ~new_new_n26849__ & ~new_new_n26850__;
  assign new_new_n26852__ = new_new_n26826__ & ~new_new_n26851__;
  assign new_new_n26853__ = ~new_new_n26826__ & new_new_n26851__;
  assign new_new_n26854__ = ~new_new_n26852__ & ~new_new_n26853__;
  assign new_new_n26855__ = new_new_n26847__ & ~new_new_n26854__;
  assign new_new_n26856__ = ~new_new_n19984__ & ~new_new_n26370__;
  assign new_new_n26857__ = ~new_new_n19988__ & new_new_n26372__;
  assign new_new_n26858__ = new_new_n19988__ & ~new_new_n26372__;
  assign new_new_n26859__ = ~new_new_n19662__ & ~new_new_n26858__;
  assign new_new_n26860__ = ~new_new_n26857__ & ~new_new_n26859__;
  assign new_new_n26861__ = new_new_n26856__ & new_new_n26860__;
  assign new_new_n26862__ = new_new_n19984__ & new_new_n26370__;
  assign new_new_n26863__ = ~new_new_n26856__ & ~new_new_n26862__;
  assign new_new_n26864__ = ~new_new_n19662__ & new_new_n26857__;
  assign new_new_n26865__ = new_new_n19662__ & new_new_n26858__;
  assign new_new_n26866__ = ~new_new_n26864__ & ~new_new_n26865__;
  assign new_new_n26867__ = new_new_n26863__ & new_new_n26866__;
  assign new_new_n26868__ = ~new_new_n26860__ & new_new_n26862__;
  assign new_new_n26869__ = ~new_new_n26377__ & ~new_new_n26861__;
  assign new_new_n26870__ = ~new_new_n26868__ & new_new_n26869__;
  assign new_new_n26871__ = ~new_new_n26867__ & new_new_n26870__;
  assign new_new_n26872__ = new_new_n19984__ & new_new_n26381__;
  assign new_new_n26873__ = new_new_n19988__ & new_new_n26872__;
  assign new_new_n26874__ = new_new_n19984__ & ~new_new_n26373__;
  assign new_new_n26875__ = ~new_new_n26381__ & ~new_new_n26874__;
  assign new_new_n26876__ = ~new_new_n19988__ & new_new_n26875__;
  assign new_new_n26877__ = ~new_new_n19984__ & new_new_n26373__;
  assign new_new_n26878__ = ~new_new_n26876__ & ~new_new_n26877__;
  assign new_new_n26879__ = ~new_new_n19662__ & ~new_new_n26878__;
  assign new_new_n26880__ = ~new_new_n19988__ & ~new_new_n26872__;
  assign new_new_n26881__ = new_new_n19662__ & ~new_new_n26875__;
  assign new_new_n26882__ = ~new_new_n26880__ & new_new_n26881__;
  assign new_new_n26883__ = new_new_n26856__ & new_new_n26857__;
  assign new_new_n26884__ = new_new_n26377__ & ~new_new_n26883__;
  assign new_new_n26885__ = ~new_new_n26873__ & new_new_n26884__;
  assign new_new_n26886__ = ~new_new_n26882__ & new_new_n26885__;
  assign new_new_n26887__ = ~new_new_n26879__ & new_new_n26886__;
  assign new_new_n26888__ = ~new_new_n26871__ & ~new_new_n26887__;
  assign new_new_n26889__ = new_new_n26847__ & ~new_new_n26888__;
  assign new_new_n26890__ = ~new_new_n26326__ & ~new_new_n26356__;
  assign new_new_n26891__ = new_new_n26328__ & ~new_new_n26345__;
  assign new_new_n26892__ = ~new_new_n26328__ & new_new_n26345__;
  assign new_new_n26893__ = ~new_new_n26891__ & ~new_new_n26892__;
  assign new_new_n26894__ = ~new_new_n26333__ & ~new_new_n26334__;
  assign new_new_n26895__ = ~new_new_n26893__ & ~new_new_n26894__;
  assign new_new_n26896__ = new_new_n26890__ & ~new_new_n26895__;
  assign new_new_n26897__ = ~new_new_n26347__ & ~new_new_n26356__;
  assign new_new_n26898__ = ~new_new_n26348__ & ~new_new_n26897__;
  assign new_new_n26899__ = ~new_new_n26896__ & ~new_new_n26898__;
  assign new_new_n26900__ = ~new_new_n26352__ & ~new_new_n26899__;
  assign new_new_n26901__ = new_new_n26326__ & ~new_new_n26332__;
  assign new_new_n26902__ = new_new_n26328__ & new_new_n26901__;
  assign new_new_n26903__ = ~new_new_n26326__ & new_new_n26332__;
  assign new_new_n26904__ = new_new_n26328__ & ~new_new_n26356__;
  assign new_new_n26905__ = ~new_new_n26903__ & new_new_n26904__;
  assign new_new_n26906__ = ~new_new_n26901__ & ~new_new_n26905__;
  assign new_new_n26907__ = ~new_new_n26345__ & ~new_new_n26906__;
  assign new_new_n26908__ = new_new_n26334__ & new_new_n26356__;
  assign new_new_n26909__ = ~new_new_n26333__ & new_new_n26356__;
  assign new_new_n26910__ = ~new_new_n26328__ & new_new_n26903__;
  assign new_new_n26911__ = ~new_new_n26909__ & ~new_new_n26910__;
  assign new_new_n26912__ = new_new_n26345__ & ~new_new_n26911__;
  assign new_new_n26913__ = ~new_new_n26902__ & ~new_new_n26908__;
  assign new_new_n26914__ = ~new_new_n26907__ & new_new_n26913__;
  assign new_new_n26915__ = ~new_new_n26912__ & new_new_n26914__;
  assign new_new_n26916__ = new_new_n26352__ & ~new_new_n26915__;
  assign new_new_n26917__ = ~new_new_n26900__ & ~new_new_n26916__;
  assign new_new_n26918__ = new_new_n26860__ & ~new_new_n26865__;
  assign new_new_n26919__ = ~new_new_n26864__ & ~new_new_n26918__;
  assign new_new_n26920__ = new_new_n26863__ & ~new_new_n26919__;
  assign new_new_n26921__ = ~new_new_n26863__ & new_new_n26919__;
  assign new_new_n26922__ = ~new_new_n26920__ & ~new_new_n26921__;
  assign new_new_n26923__ = ~new_new_n26332__ & new_new_n26890__;
  assign new_new_n26924__ = new_new_n26332__ & ~new_new_n26890__;
  assign new_new_n26925__ = ~new_new_n26923__ & ~new_new_n26924__;
  assign new_new_n26926__ = new_new_n26893__ & new_new_n26925__;
  assign new_new_n26927__ = ~new_new_n26893__ & ~new_new_n26925__;
  assign new_new_n26928__ = ~new_new_n26926__ & ~new_new_n26927__;
  assign new_new_n26929__ = ~new_new_n26917__ & ~new_new_n26928__;
  assign new_new_n26930__ = ~new_new_n26274__ & ~new_new_n26275__;
  assign new_new_n26931__ = ~new_new_n26244__ & ~new_new_n26310__;
  assign new_new_n26932__ = new_new_n26930__ & ~new_new_n26931__;
  assign new_new_n26933__ = ~new_new_n26930__ & new_new_n26931__;
  assign new_new_n26934__ = ~new_new_n26932__ & ~new_new_n26933__;
  assign new_new_n26935__ = new_new_n26286__ & new_new_n26934__;
  assign new_new_n26936__ = ~new_new_n26286__ & ~new_new_n26934__;
  assign new_new_n26937__ = ~new_new_n26935__ & ~new_new_n26936__;
  assign new_new_n26938__ = ~new_new_n26318__ & ~new_new_n26319__;
  assign new_new_n26939__ = ~new_new_n26321__ & new_new_n26938__;
  assign new_new_n26940__ = new_new_n26321__ & ~new_new_n26938__;
  assign new_new_n26941__ = ~new_new_n26939__ & ~new_new_n26940__;
  assign new_new_n26942__ = ~new_new_n26917__ & new_new_n26941__;
  assign new_new_n26943__ = new_new_n26231__ & new_new_n26233__;
  assign new_new_n26944__ = ~new_new_n26225__ & ~new_new_n26234__;
  assign new_new_n26945__ = new_new_n23812__ & ~new_new_n26231__;
  assign new_new_n26946__ = ~new_new_n26943__ & ~new_new_n26945__;
  assign new_new_n26947__ = new_new_n26944__ & new_new_n26946__;
  assign new_new_n26948__ = ~new_new_n23812__ & new_new_n26231__;
  assign new_new_n26949__ = ~new_new_n26233__ & ~new_new_n26948__;
  assign new_new_n26950__ = new_new_n26234__ & ~new_new_n26949__;
  assign new_new_n26951__ = new_new_n26225__ & new_new_n26949__;
  assign new_new_n26952__ = ~new_new_n26950__ & ~new_new_n26951__;
  assign new_new_n26953__ = ~new_new_n26947__ & new_new_n26952__;
  assign new_new_n26954__ = ~new_new_n23816__ & ~new_new_n26953__;
  assign new_new_n26955__ = new_new_n26225__ & new_new_n26233__;
  assign new_new_n26956__ = ~new_new_n23807__ & new_new_n26225__;
  assign new_new_n26957__ = new_new_n23807__ & ~new_new_n26225__;
  assign new_new_n26958__ = ~new_new_n23811__ & ~new_new_n26234__;
  assign new_new_n26959__ = ~new_new_n26957__ & new_new_n26958__;
  assign new_new_n26960__ = ~new_new_n26956__ & ~new_new_n26959__;
  assign new_new_n26961__ = new_new_n26231__ & ~new_new_n26960__;
  assign new_new_n26962__ = ~new_new_n26233__ & new_new_n26234__;
  assign new_new_n26963__ = new_new_n23811__ & new_new_n26957__;
  assign new_new_n26964__ = ~new_new_n26962__ & ~new_new_n26963__;
  assign new_new_n26965__ = ~new_new_n26231__ & ~new_new_n26964__;
  assign new_new_n26966__ = new_new_n23812__ & new_new_n26234__;
  assign new_new_n26967__ = ~new_new_n26955__ & ~new_new_n26966__;
  assign new_new_n26968__ = ~new_new_n26961__ & new_new_n26967__;
  assign new_new_n26969__ = ~new_new_n26965__ & new_new_n26968__;
  assign new_new_n26970__ = new_new_n23816__ & ~new_new_n26969__;
  assign new_new_n26971__ = ~new_new_n26954__ & ~new_new_n26970__;
  assign new_new_n26972__ = ~new_new_n23812__ & ~new_new_n26233__;
  assign new_new_n26973__ = new_new_n26944__ & ~new_new_n26972__;
  assign new_new_n26974__ = ~new_new_n26944__ & new_new_n26972__;
  assign new_new_n26975__ = ~new_new_n26973__ & ~new_new_n26974__;
  assign new_new_n26976__ = new_new_n26231__ & new_new_n26975__;
  assign new_new_n26977__ = ~new_new_n26231__ & ~new_new_n26975__;
  assign new_new_n26978__ = ~new_new_n26976__ & ~new_new_n26977__;
  assign new_new_n26979__ = ~new_new_n26937__ & ~new_new_n26978__;
  assign new_new_n26980__ = ~new_new_n26205__ & new_new_n26216__;
  assign new_new_n26981__ = new_new_n26205__ & ~new_new_n26216__;
  assign new_new_n26982__ = ~new_new_n26191__ & ~new_new_n26201__;
  assign new_new_n26983__ = ~new_new_n26981__ & new_new_n26982__;
  assign new_new_n26984__ = ~new_new_n26980__ & ~new_new_n26983__;
  assign new_new_n26985__ = ~new_new_n18146__ & ~new_new_n26984__;
  assign new_new_n26986__ = new_new_n26206__ & new_new_n26216__;
  assign new_new_n26987__ = new_new_n26191__ & ~new_new_n26206__;
  assign new_new_n26988__ = new_new_n26207__ & ~new_new_n26216__;
  assign new_new_n26989__ = ~new_new_n26987__ & ~new_new_n26988__;
  assign new_new_n26990__ = new_new_n18146__ & ~new_new_n26989__;
  assign new_new_n26991__ = new_new_n26191__ & new_new_n26207__;
  assign new_new_n26992__ = ~new_new_n26214__ & ~new_new_n26986__;
  assign new_new_n26993__ = ~new_new_n26991__ & new_new_n26992__;
  assign new_new_n26994__ = ~new_new_n26990__ & new_new_n26993__;
  assign new_new_n26995__ = ~new_new_n26985__ & new_new_n26994__;
  assign new_new_n26996__ = new_new_n26209__ & ~new_new_n26216__;
  assign new_new_n26997__ = ~new_new_n26210__ & ~new_new_n26996__;
  assign new_new_n26998__ = ~new_new_n26191__ & ~new_new_n26216__;
  assign new_new_n26999__ = ~new_new_n26217__ & ~new_new_n26218__;
  assign new_new_n27000__ = new_new_n26998__ & new_new_n26999__;
  assign new_new_n27001__ = new_new_n26214__ & ~new_new_n26997__;
  assign new_new_n27002__ = ~new_new_n27000__ & new_new_n27001__;
  assign new_new_n27003__ = ~new_new_n26995__ & ~new_new_n27002__;
  assign new_new_n27004__ = ~pi02 & new_new_n25262__;
  assign new_new_n27005__ = new_new_n25262__ & new_new_n26180__;
  assign new_new_n27006__ = ~new_new_n26180__ & new_new_n26184__;
  assign new_new_n27007__ = ~new_new_n27005__ & ~new_new_n27006__;
  assign new_new_n27008__ = new_new_n16056__ & ~new_new_n27007__;
  assign new_new_n27009__ = ~new_new_n27004__ & ~new_new_n27008__;
  assign new_new_n27010__ = new_new_n14393__ & ~new_new_n27009__;
  assign new_new_n27011__ = new_new_n26180__ & new_new_n27004__;
  assign new_new_n27012__ = ~new_new_n14393__ & ~new_new_n27004__;
  assign new_new_n27013__ = ~new_new_n26185__ & new_new_n27012__;
  assign new_new_n27014__ = ~new_new_n27006__ & new_new_n27013__;
  assign new_new_n27015__ = new_new_n14393__ & new_new_n25262__;
  assign new_new_n27016__ = ~new_new_n26180__ & ~new_new_n27015__;
  assign new_new_n27017__ = ~new_new_n16056__ & ~new_new_n26185__;
  assign new_new_n27018__ = ~new_new_n27016__ & new_new_n27017__;
  assign new_new_n27019__ = ~new_new_n27011__ & ~new_new_n27014__;
  assign new_new_n27020__ = ~new_new_n27018__ & new_new_n27019__;
  assign new_new_n27021__ = ~new_new_n27010__ & new_new_n27020__;
  assign new_new_n27022__ = ~new_new_n27003__ & ~new_new_n27021__;
  assign new_new_n27023__ = ~new_new_n26206__ & ~new_new_n26207__;
  assign new_new_n27024__ = new_new_n18146__ & ~new_new_n27023__;
  assign new_new_n27025__ = ~new_new_n18146__ & new_new_n27023__;
  assign new_new_n27026__ = ~new_new_n27024__ & ~new_new_n27025__;
  assign new_new_n27027__ = new_new_n26998__ & new_new_n27026__;
  assign new_new_n27028__ = ~new_new_n26998__ & ~new_new_n27026__;
  assign new_new_n27029__ = ~new_new_n27027__ & ~new_new_n27028__;
  assign new_new_n27030__ = ~new_new_n26165__ & ~new_new_n26166__;
  assign new_new_n27031__ = new_new_n26170__ & ~new_new_n27030__;
  assign new_new_n27032__ = ~new_new_n26170__ & new_new_n27030__;
  assign new_new_n27033__ = ~new_new_n27031__ & ~new_new_n27032__;
  assign new_new_n27034__ = new_new_n26135__ & new_new_n26144__;
  assign new_new_n27035__ = new_new_n26155__ & ~new_new_n27034__;
  assign new_new_n27036__ = new_new_n26144__ & ~new_new_n26155__;
  assign new_new_n27037__ = new_new_n26135__ & new_new_n27036__;
  assign new_new_n27038__ = ~new_new_n27035__ & ~new_new_n27037__;
  assign new_new_n27039__ = pi02 & ~new_new_n27038__;
  assign new_new_n27040__ = ~pi02 & new_new_n27038__;
  assign new_new_n27041__ = ~new_new_n27039__ & ~new_new_n27040__;
  assign new_new_n27042__ = new_new_n25302__ & new_new_n25309__;
  assign new_new_n27043__ = ~new_new_n26147__ & ~new_new_n27042__;
  assign new_new_n27044__ = pi02 & ~new_new_n26135__;
  assign new_new_n27045__ = new_new_n26144__ & new_new_n27044__;
  assign new_new_n27046__ = ~pi02 & ~new_new_n26144__;
  assign new_new_n27047__ = ~new_new_n27036__ & ~new_new_n27046__;
  assign new_new_n27048__ = new_new_n26135__ & ~new_new_n27047__;
  assign new_new_n27049__ = ~new_new_n27045__ & ~new_new_n27048__;
  assign new_new_n27050__ = ~new_new_n27043__ & ~new_new_n27049__;
  assign new_new_n27051__ = ~new_new_n27044__ & ~new_new_n27046__;
  assign new_new_n27052__ = ~new_new_n27037__ & new_new_n27051__;
  assign new_new_n27053__ = new_new_n27043__ & new_new_n27052__;
  assign new_new_n27054__ = ~new_new_n27050__ & ~new_new_n27053__;
  assign new_new_n27055__ = new_new_n27041__ & ~new_new_n27054__;
  assign new_new_n27056__ = ~new_new_n25349__ & ~new_new_n25350__;
  assign new_new_n27057__ = new_new_n26122__ & new_new_n27056__;
  assign new_new_n27058__ = ~new_new_n26122__ & ~new_new_n27056__;
  assign new_new_n27059__ = ~new_new_n27057__ & ~new_new_n27058__;
  assign new_new_n27060__ = new_new_n27055__ & new_new_n27059__;
  assign new_new_n27061__ = ~new_new_n27041__ & new_new_n27054__;
  assign new_new_n27062__ = ~new_new_n26125__ & ~new_new_n26131__;
  assign new_new_n27063__ = new_new_n25149__ & new_new_n27062__;
  assign new_new_n27064__ = ~new_new_n25149__ & ~new_new_n27062__;
  assign new_new_n27065__ = ~new_new_n27063__ & ~new_new_n27064__;
  assign new_new_n27066__ = new_new_n25169__ & ~new_new_n27065__;
  assign new_new_n27067__ = ~new_new_n25169__ & new_new_n27065__;
  assign new_new_n27068__ = ~new_new_n27066__ & ~new_new_n27067__;
  assign new_new_n27069__ = new_new_n25156__ & new_new_n27068__;
  assign new_new_n27070__ = ~new_new_n25156__ & ~new_new_n27068__;
  assign new_new_n27071__ = ~new_new_n27069__ & ~new_new_n27070__;
  assign new_new_n27072__ = ~new_new_n25370__ & ~new_new_n25371__;
  assign new_new_n27073__ = new_new_n26091__ & ~new_new_n27072__;
  assign new_new_n27074__ = ~new_new_n26091__ & new_new_n27072__;
  assign new_new_n27075__ = ~new_new_n27073__ & ~new_new_n27074__;
  assign new_new_n27076__ = ~new_new_n27071__ & ~new_new_n27075__;
  assign new_new_n27077__ = new_new_n27061__ & new_new_n27076__;
  assign new_new_n27078__ = ~new_new_n27060__ & ~new_new_n27077__;
  assign new_new_n27079__ = new_new_n26118__ & ~new_new_n27078__;
  assign new_new_n27080__ = new_new_n27059__ & new_new_n27061__;
  assign new_new_n27081__ = ~new_new_n27055__ & ~new_new_n27080__;
  assign new_new_n27082__ = ~new_new_n27071__ & ~new_new_n27081__;
  assign new_new_n27083__ = ~new_new_n27041__ & new_new_n27071__;
  assign new_new_n27084__ = new_new_n26118__ & new_new_n27059__;
  assign new_new_n27085__ = new_new_n27071__ & ~new_new_n27084__;
  assign new_new_n27086__ = new_new_n27054__ & new_new_n27085__;
  assign new_new_n27087__ = new_new_n26118__ & ~new_new_n27075__;
  assign new_new_n27088__ = ~new_new_n27059__ & ~new_new_n27087__;
  assign new_new_n27089__ = ~new_new_n27041__ & new_new_n27088__;
  assign new_new_n27090__ = ~new_new_n27083__ & ~new_new_n27089__;
  assign new_new_n27091__ = ~new_new_n27086__ & new_new_n27090__;
  assign new_new_n27092__ = ~new_new_n27061__ & ~new_new_n27091__;
  assign new_new_n27093__ = ~new_new_n27079__ & ~new_new_n27092__;
  assign new_new_n27094__ = ~new_new_n27082__ & new_new_n27093__;
  assign new_new_n27095__ = new_new_n27041__ & new_new_n27084__;
  assign new_new_n27096__ = new_new_n27071__ & ~new_new_n27095__;
  assign new_new_n27097__ = ~new_new_n27089__ & ~new_new_n27096__;
  assign new_new_n27098__ = ~new_new_n27041__ & ~new_new_n27097__;
  assign new_new_n27099__ = ~new_new_n27094__ & new_new_n27098__;
  assign new_new_n27100__ = new_new_n27041__ & ~new_new_n27085__;
  assign new_new_n27101__ = new_new_n27094__ & new_new_n27100__;
  assign new_new_n27102__ = ~new_new_n27099__ & ~new_new_n27101__;
  assign new_new_n27103__ = new_new_n27033__ & ~new_new_n27102__;
  assign new_new_n27104__ = new_new_n27054__ & new_new_n27102__;
  assign new_new_n27105__ = ~new_new_n27103__ & ~new_new_n27104__;
  assign new_new_n27106__ = ~new_new_n27029__ & new_new_n27105__;
  assign new_new_n27107__ = ~new_new_n27022__ & ~new_new_n27106__;
  assign new_new_n27108__ = ~new_new_n26173__ & ~new_new_n26174__;
  assign new_new_n27109__ = ~new_new_n26178__ & new_new_n27108__;
  assign new_new_n27110__ = new_new_n26178__ & ~new_new_n27108__;
  assign new_new_n27111__ = ~new_new_n27109__ & ~new_new_n27110__;
  assign new_new_n27112__ = ~new_new_n27107__ & new_new_n27111__;
  assign new_new_n27113__ = ~new_new_n27003__ & ~new_new_n27029__;
  assign new_new_n27114__ = ~new_new_n27029__ & new_new_n27111__;
  assign new_new_n27115__ = new_new_n27022__ & new_new_n27105__;
  assign new_new_n27116__ = ~new_new_n27114__ & ~new_new_n27115__;
  assign new_new_n27117__ = ~new_new_n27033__ & ~new_new_n27116__;
  assign new_new_n27118__ = ~new_new_n27021__ & ~new_new_n27029__;
  assign new_new_n27119__ = ~new_new_n27113__ & ~new_new_n27118__;
  assign new_new_n27120__ = ~new_new_n27112__ & new_new_n27119__;
  assign new_new_n27121__ = ~new_new_n27117__ & new_new_n27120__;
  assign new_new_n27122__ = new_new_n27003__ & new_new_n27121__;
  assign new_new_n27123__ = new_new_n26979__ & ~new_new_n27122__;
  assign new_new_n27124__ = ~new_new_n26971__ & ~new_new_n27123__;
  assign new_new_n27125__ = new_new_n26937__ & new_new_n26978__;
  assign new_new_n27126__ = ~new_new_n27003__ & ~new_new_n27121__;
  assign new_new_n27127__ = new_new_n27125__ & ~new_new_n27126__;
  assign new_new_n27128__ = ~new_new_n27124__ & ~new_new_n27127__;
  assign new_new_n27129__ = new_new_n26942__ & ~new_new_n27128__;
  assign new_new_n27130__ = ~new_new_n26288__ & ~new_new_n26310__;
  assign new_new_n27131__ = ~new_new_n26289__ & ~new_new_n27130__;
  assign new_new_n27132__ = ~new_new_n26309__ & ~new_new_n26311__;
  assign new_new_n27133__ = new_new_n26931__ & new_new_n27132__;
  assign new_new_n27134__ = ~new_new_n27131__ & ~new_new_n27133__;
  assign new_new_n27135__ = ~new_new_n26307__ & ~new_new_n27134__;
  assign new_new_n27136__ = new_new_n26244__ & new_new_n26274__;
  assign new_new_n27137__ = new_new_n26244__ & new_new_n26246__;
  assign new_new_n27138__ = ~new_new_n26244__ & ~new_new_n26246__;
  assign new_new_n27139__ = ~new_new_n26273__ & ~new_new_n26310__;
  assign new_new_n27140__ = ~new_new_n27138__ & new_new_n27139__;
  assign new_new_n27141__ = ~new_new_n27137__ & ~new_new_n27140__;
  assign new_new_n27142__ = ~new_new_n26286__ & ~new_new_n27141__;
  assign new_new_n27143__ = ~new_new_n26274__ & new_new_n26310__;
  assign new_new_n27144__ = new_new_n26273__ & new_new_n27138__;
  assign new_new_n27145__ = ~new_new_n27143__ & ~new_new_n27144__;
  assign new_new_n27146__ = new_new_n26286__ & ~new_new_n27145__;
  assign new_new_n27147__ = new_new_n26275__ & new_new_n26310__;
  assign new_new_n27148__ = ~new_new_n27136__ & ~new_new_n27147__;
  assign new_new_n27149__ = ~new_new_n27142__ & new_new_n27148__;
  assign new_new_n27150__ = ~new_new_n27146__ & new_new_n27149__;
  assign new_new_n27151__ = new_new_n26307__ & ~new_new_n27150__;
  assign new_new_n27152__ = ~new_new_n27135__ & ~new_new_n27151__;
  assign new_new_n27153__ = ~new_new_n26928__ & ~new_new_n27152__;
  assign new_new_n27154__ = ~new_new_n27129__ & ~new_new_n27153__;
  assign new_new_n27155__ = new_new_n26937__ & ~new_new_n27154__;
  assign new_new_n27156__ = ~new_new_n26928__ & ~new_new_n27128__;
  assign new_new_n27157__ = ~new_new_n26942__ & ~new_new_n27156__;
  assign new_new_n27158__ = ~new_new_n27152__ & ~new_new_n27157__;
  assign new_new_n27159__ = ~new_new_n26928__ & new_new_n26941__;
  assign new_new_n27160__ = ~new_new_n26929__ & ~new_new_n27159__;
  assign new_new_n27161__ = ~new_new_n27158__ & new_new_n27160__;
  assign new_new_n27162__ = ~new_new_n27155__ & new_new_n27161__;
  assign new_new_n27163__ = ~new_new_n26922__ & ~new_new_n27162__;
  assign new_new_n27164__ = ~new_new_n26917__ & new_new_n27163__;
  assign new_new_n27165__ = ~new_new_n26363__ & ~new_new_n26364__;
  assign new_new_n27166__ = ~new_new_n26368__ & new_new_n27165__;
  assign new_new_n27167__ = new_new_n26368__ & ~new_new_n27165__;
  assign new_new_n27168__ = ~new_new_n27166__ & ~new_new_n27167__;
  assign new_new_n27169__ = ~new_new_n27164__ & ~new_new_n27168__;
  assign new_new_n27170__ = new_new_n26922__ & new_new_n27162__;
  assign new_new_n27171__ = new_new_n26917__ & new_new_n27170__;
  assign new_new_n27172__ = ~new_new_n27169__ & ~new_new_n27171__;
  assign new_new_n27173__ = ~new_new_n26854__ & ~new_new_n27172__;
  assign new_new_n27174__ = ~new_new_n26889__ & ~new_new_n27173__;
  assign new_new_n27175__ = new_new_n26922__ & ~new_new_n27172__;
  assign new_new_n27176__ = ~new_new_n26922__ & ~new_new_n27169__;
  assign new_new_n27177__ = ~new_new_n27175__ & ~new_new_n27176__;
  assign new_new_n27178__ = new_new_n26888__ & ~new_new_n27177__;
  assign new_new_n27179__ = ~new_new_n26888__ & new_new_n27177__;
  assign new_new_n27180__ = ~new_new_n27178__ & ~new_new_n27179__;
  assign new_new_n27181__ = ~new_new_n27174__ & ~new_new_n27180__;
  assign new_new_n27182__ = new_new_n26847__ & new_new_n26922__;
  assign new_new_n27183__ = new_new_n26854__ & ~new_new_n27182__;
  assign new_new_n27184__ = ~new_new_n26888__ & ~new_new_n27183__;
  assign new_new_n27185__ = ~new_new_n27181__ & ~new_new_n27184__;
  assign new_new_n27186__ = ~new_new_n26855__ & new_new_n27185__;
  assign new_new_n27187__ = ~new_new_n26823__ & new_new_n27186__;
  assign new_new_n27188__ = ~new_new_n26847__ & new_new_n27187__;
  assign new_new_n27189__ = new_new_n26823__ & ~new_new_n27186__;
  assign new_new_n27190__ = new_new_n26847__ & new_new_n27189__;
  assign new_new_n27191__ = ~new_new_n27188__ & ~new_new_n27190__;
  assign new_new_n27192__ = new_new_n26741__ & new_new_n27191__;
  assign new_new_n27193__ = new_new_n26823__ & new_new_n27192__;
  assign new_new_n27194__ = new_new_n18340__ & new_new_n26816__;
  assign new_new_n27195__ = ~new_new_n18340__ & ~new_new_n26816__;
  assign new_new_n27196__ = ~new_new_n26815__ & ~new_new_n27195__;
  assign new_new_n27197__ = new_new_n18716__ & new_new_n27196__;
  assign new_new_n27198__ = ~new_new_n26431__ & ~new_new_n27194__;
  assign new_new_n27199__ = ~new_new_n27197__ & new_new_n27198__;
  assign new_new_n27200__ = ~new_new_n18340__ & new_new_n26815__;
  assign new_new_n27201__ = ~new_new_n18716__ & ~new_new_n27196__;
  assign new_new_n27202__ = new_new_n26431__ & ~new_new_n27200__;
  assign new_new_n27203__ = ~new_new_n27201__ & new_new_n27202__;
  assign new_new_n27204__ = ~new_new_n27199__ & ~new_new_n27203__;
  assign new_new_n27205__ = ~new_new_n26423__ & ~new_new_n26816__;
  assign new_new_n27206__ = ~new_new_n26433__ & ~new_new_n26813__;
  assign new_new_n27207__ = ~new_new_n27205__ & ~new_new_n27206__;
  assign new_new_n27208__ = new_new_n18711__ & ~new_new_n27207__;
  assign new_new_n27209__ = ~new_new_n27204__ & new_new_n27208__;
  assign new_new_n27210__ = new_new_n26431__ & ~new_new_n26813__;
  assign new_new_n27211__ = ~new_new_n26812__ & ~new_new_n27210__;
  assign new_new_n27212__ = new_new_n26815__ & new_new_n27211__;
  assign new_new_n27213__ = new_new_n26431__ & new_new_n26812__;
  assign new_new_n27214__ = ~new_new_n26431__ & new_new_n26813__;
  assign new_new_n27215__ = ~new_new_n27213__ & ~new_new_n27214__;
  assign new_new_n27216__ = new_new_n26817__ & new_new_n27215__;
  assign new_new_n27217__ = new_new_n26816__ & ~new_new_n27211__;
  assign new_new_n27218__ = ~new_new_n18711__ & ~new_new_n27212__;
  assign new_new_n27219__ = ~new_new_n27217__ & new_new_n27218__;
  assign new_new_n27220__ = ~new_new_n27216__ & new_new_n27219__;
  assign new_new_n27221__ = ~new_new_n27209__ & ~new_new_n27220__;
  assign new_new_n27222__ = ~new_new_n26847__ & new_new_n27185__;
  assign new_new_n27223__ = ~new_new_n26823__ & ~new_new_n27222__;
  assign new_new_n27224__ = ~new_new_n27192__ & new_new_n27223__;
  assign new_new_n27225__ = new_new_n27221__ & ~new_new_n27224__;
  assign new_new_n27226__ = ~new_new_n27193__ & ~new_new_n27225__;
  assign new_new_n27227__ = new_new_n26811__ & ~new_new_n27226__;
  assign new_new_n27228__ = ~new_new_n26803__ & ~new_new_n27227__;
  assign new_new_n27229__ = new_new_n26741__ & ~new_new_n27228__;
  assign new_new_n27230__ = new_new_n26729__ & new_new_n26810__;
  assign new_new_n27231__ = ~new_new_n26774__ & ~new_new_n27230__;
  assign new_new_n27232__ = ~new_new_n26774__ & ~new_new_n27226__;
  assign new_new_n27233__ = ~new_new_n26811__ & ~new_new_n27232__;
  assign new_new_n27234__ = new_new_n26802__ & ~new_new_n27233__;
  assign new_new_n27235__ = ~new_new_n27231__ & ~new_new_n27234__;
  assign new_new_n27236__ = ~new_new_n27229__ & new_new_n27235__;
  assign new_new_n27237__ = ~new_new_n26729__ & ~new_new_n27236__;
  assign new_new_n27238__ = new_new_n26722__ & ~new_new_n27237__;
  assign new_new_n27239__ = ~new_new_n17002__ & ~new_new_n17003__;
  assign new_new_n27240__ = new_new_n26530__ & new_new_n27239__;
  assign new_new_n27241__ = ~new_new_n26530__ & ~new_new_n27239__;
  assign new_new_n27242__ = ~new_new_n27240__ & ~new_new_n27241__;
  assign new_new_n27243__ = ~new_new_n27238__ & new_new_n27242__;
  assign new_new_n27244__ = ~new_new_n26547__ & ~new_new_n26548__;
  assign new_new_n27245__ = new_new_n26557__ & ~new_new_n27244__;
  assign new_new_n27246__ = ~new_new_n26557__ & new_new_n27244__;
  assign new_new_n27247__ = ~new_new_n27245__ & ~new_new_n27246__;
  assign new_new_n27248__ = new_new_n26677__ & new_new_n27247__;
  assign new_new_n27249__ = ~new_new_n26677__ & ~new_new_n27247__;
  assign new_new_n27250__ = ~new_new_n27248__ & ~new_new_n27249__;
  assign new_new_n27251__ = new_new_n27242__ & new_new_n27250__;
  assign new_new_n27252__ = ~new_new_n27242__ & ~new_new_n27250__;
  assign new_new_n27253__ = ~new_new_n27236__ & new_new_n27252__;
  assign new_new_n27254__ = ~new_new_n27251__ & ~new_new_n27253__;
  assign new_new_n27255__ = ~new_new_n26722__ & ~new_new_n27254__;
  assign new_new_n27256__ = ~new_new_n27242__ & new_new_n27250__;
  assign new_new_n27257__ = new_new_n27242__ & ~new_new_n27250__;
  assign new_new_n27258__ = new_new_n27236__ & new_new_n27257__;
  assign new_new_n27259__ = ~new_new_n27256__ & ~new_new_n27258__;
  assign new_new_n27260__ = new_new_n26722__ & ~new_new_n27259__;
  assign new_new_n27261__ = new_new_n27236__ & new_new_n27256__;
  assign new_new_n27262__ = new_new_n26722__ & new_new_n27257__;
  assign new_new_n27263__ = new_new_n26729__ & ~new_new_n27261__;
  assign new_new_n27264__ = ~new_new_n27262__ & new_new_n27263__;
  assign new_new_n27265__ = ~new_new_n26722__ & new_new_n27252__;
  assign new_new_n27266__ = ~new_new_n27236__ & new_new_n27251__;
  assign new_new_n27267__ = ~new_new_n26729__ & ~new_new_n27265__;
  assign new_new_n27268__ = ~new_new_n27266__ & new_new_n27267__;
  assign new_new_n27269__ = ~new_new_n27264__ & ~new_new_n27268__;
  assign new_new_n27270__ = ~new_new_n27255__ & ~new_new_n27260__;
  assign new_new_n27271__ = ~new_new_n27269__ & new_new_n27270__;
  assign new_new_n27272__ = ~new_new_n27250__ & ~new_new_n27271__;
  assign new_new_n27273__ = ~new_new_n27243__ & ~new_new_n27272__;
  assign new_new_n27274__ = new_new_n26674__ & new_new_n27273__;
  assign new_new_n27275__ = ~new_new_n26674__ & ~new_new_n27273__;
  assign new_new_n27276__ = ~new_new_n27274__ & ~new_new_n27275__;
  assign new_new_n27277__ = new_new_n27243__ & new_new_n27250__;
  assign new_new_n27278__ = ~new_new_n27250__ & new_new_n27271__;
  assign new_new_n27279__ = ~new_new_n27243__ & new_new_n27278__;
  assign new_new_n27280__ = ~new_new_n26698__ & ~new_new_n27279__;
  assign new_new_n27281__ = ~new_new_n27277__ & ~new_new_n27280__;
  assign new_new_n27282__ = new_new_n27276__ & ~new_new_n27281__;
  assign new_new_n27283__ = ~new_new_n27276__ & new_new_n27281__;
  assign new_new_n27284__ = ~new_new_n27282__ & ~new_new_n27283__;
  assign new_new_n27285__ = new_new_n26698__ & ~new_new_n27284__;
  assign new_new_n27286__ = new_new_n26674__ & ~new_new_n27285__;
  assign new_new_n27287__ = ~new_new_n26674__ & new_new_n26698__;
  assign new_new_n27288__ = ~new_new_n26674__ & ~new_new_n27284__;
  assign new_new_n27289__ = ~new_new_n27287__ & ~new_new_n27288__;
  assign new_new_n27290__ = ~new_new_n27286__ & new_new_n27289__;
  assign new_new_n27291__ = pi02 & ~new_new_n27290__;
  assign new_new_n27292__ = pi01 & new_new_n27290__;
  assign new_new_n27293__ = ~new_new_n27291__ & ~new_new_n27292__;
  assign new_new_n27294__ = ~new_new_n26667__ & new_new_n27293__;
  assign new_new_n27295__ = new_new_n26667__ & ~new_new_n27293__;
  assign new_new_n27296__ = pi00 & ~new_new_n27294__;
  assign new_new_n27297__ = ~new_new_n27295__ & new_new_n27296__;
  assign new_new_n27298__ = new_new_n13508__ & ~new_new_n26674__;
  assign new_new_n27299__ = ~pi01 & ~new_new_n26698__;
  assign new_new_n27300__ = pi01 & new_new_n26674__;
  assign new_new_n27301__ = ~new_new_n27299__ & ~new_new_n27300__;
  assign new_new_n27302__ = pi02 & ~new_new_n27301__;
  assign new_new_n27303__ = ~pi00 & ~new_new_n27298__;
  assign new_new_n27304__ = ~new_new_n27302__ & new_new_n27303__;
  assign new_new_n27305__ = ~new_new_n27297__ & ~new_new_n27304__;
  assign new_new_n27306__ = new_new_n11471__ & new_new_n26722__;
  assign new_new_n27307__ = new_new_n11475__ & ~new_new_n27242__;
  assign new_new_n27308__ = new_new_n12850__ & new_new_n27250__;
  assign new_new_n27309__ = ~new_new_n27306__ & ~new_new_n27307__;
  assign new_new_n27310__ = ~new_new_n27308__ & new_new_n27309__;
  assign new_new_n27311__ = pi05 & ~new_new_n27310__;
  assign new_new_n27312__ = new_new_n12856__ & ~new_new_n27271__;
  assign new_new_n27313__ = new_new_n11469__ & ~new_new_n27271__;
  assign new_new_n27314__ = ~pi05 & ~new_new_n27313__;
  assign new_new_n27315__ = ~new_new_n27312__ & ~new_new_n27314__;
  assign new_new_n27316__ = new_new_n27310__ & ~new_new_n27315__;
  assign new_new_n27317__ = ~new_new_n27311__ & ~new_new_n27316__;
  assign new_new_n27318__ = new_new_n12832__ & new_new_n26729__;
  assign new_new_n27319__ = new_new_n11475__ & new_new_n26722__;
  assign new_new_n27320__ = ~new_new_n27318__ & ~new_new_n27319__;
  assign new_new_n27321__ = new_new_n26722__ & ~new_new_n26729__;
  assign new_new_n27322__ = ~new_new_n26722__ & new_new_n26729__;
  assign new_new_n27323__ = ~new_new_n27321__ & ~new_new_n27322__;
  assign new_new_n27324__ = ~new_new_n26774__ & new_new_n27322__;
  assign new_new_n27325__ = ~new_new_n26741__ & ~new_new_n27225__;
  assign new_new_n27326__ = new_new_n26810__ & new_new_n27325__;
  assign new_new_n27327__ = ~new_new_n26810__ & ~new_new_n27226__;
  assign new_new_n27328__ = new_new_n26741__ & new_new_n27327__;
  assign new_new_n27329__ = ~new_new_n26802__ & ~new_new_n27328__;
  assign new_new_n27330__ = ~new_new_n27326__ & ~new_new_n27329__;
  assign new_new_n27331__ = new_new_n27321__ & new_new_n27330__;
  assign new_new_n27332__ = ~new_new_n27324__ & ~new_new_n27331__;
  assign new_new_n27333__ = ~new_new_n26810__ & ~new_new_n27332__;
  assign new_new_n27334__ = ~new_new_n26722__ & ~new_new_n26729__;
  assign new_new_n27335__ = new_new_n26774__ & new_new_n27334__;
  assign new_new_n27336__ = new_new_n26722__ & new_new_n26729__;
  assign new_new_n27337__ = ~new_new_n27330__ & new_new_n27336__;
  assign new_new_n27338__ = ~new_new_n27335__ & ~new_new_n27337__;
  assign new_new_n27339__ = new_new_n26810__ & ~new_new_n27338__;
  assign new_new_n27340__ = new_new_n27322__ & new_new_n27330__;
  assign new_new_n27341__ = ~new_new_n27321__ & ~new_new_n27340__;
  assign new_new_n27342__ = ~new_new_n26774__ & ~new_new_n27341__;
  assign new_new_n27343__ = ~new_new_n27330__ & new_new_n27334__;
  assign new_new_n27344__ = ~new_new_n27336__ & ~new_new_n27343__;
  assign new_new_n27345__ = new_new_n26774__ & ~new_new_n27344__;
  assign new_new_n27346__ = ~new_new_n27333__ & ~new_new_n27339__;
  assign new_new_n27347__ = ~new_new_n27342__ & ~new_new_n27345__;
  assign new_new_n27348__ = new_new_n27346__ & new_new_n27347__;
  assign new_new_n27349__ = new_new_n26722__ & ~new_new_n27348__;
  assign new_new_n27350__ = ~new_new_n26722__ & new_new_n27348__;
  assign new_new_n27351__ = ~new_new_n27349__ & ~new_new_n27350__;
  assign new_new_n27352__ = ~new_new_n27323__ & ~new_new_n27351__;
  assign new_new_n27353__ = ~new_new_n27242__ & ~new_new_n27352__;
  assign new_new_n27354__ = new_new_n11469__ & new_new_n27353__;
  assign new_new_n27355__ = new_new_n27320__ & ~new_new_n27354__;
  assign new_new_n27356__ = pi05 & ~new_new_n27355__;
  assign new_new_n27357__ = pi04 & new_new_n27242__;
  assign new_new_n27358__ = ~pi04 & ~new_new_n27242__;
  assign new_new_n27359__ = ~new_new_n11482__ & ~new_new_n27357__;
  assign new_new_n27360__ = ~new_new_n27358__ & new_new_n27359__;
  assign new_new_n27361__ = new_new_n27352__ & new_new_n27360__;
  assign new_new_n27362__ = new_new_n27242__ & ~new_new_n27352__;
  assign new_new_n27363__ = new_new_n11469__ & ~new_new_n27362__;
  assign new_new_n27364__ = ~pi05 & ~new_new_n27363__;
  assign new_new_n27365__ = ~new_new_n27361__ & ~new_new_n27364__;
  assign new_new_n27366__ = new_new_n27320__ & ~new_new_n27365__;
  assign new_new_n27367__ = ~new_new_n27356__ & ~new_new_n27366__;
  assign new_new_n27368__ = new_new_n26774__ & ~new_new_n26810__;
  assign new_new_n27369__ = ~new_new_n26774__ & new_new_n26810__;
  assign new_new_n27370__ = ~new_new_n27368__ & ~new_new_n27369__;
  assign new_new_n27371__ = ~new_new_n27330__ & new_new_n27370__;
  assign new_new_n27372__ = new_new_n27330__ & ~new_new_n27370__;
  assign new_new_n27373__ = ~new_new_n27371__ & ~new_new_n27372__;
  assign new_new_n27374__ = new_new_n11378__ & ~new_new_n27373__;
  assign new_new_n27375__ = ~new_new_n11409__ & ~new_new_n26802__;
  assign new_new_n27376__ = new_new_n10702__ & new_new_n26810__;
  assign new_new_n27377__ = ~new_new_n27375__ & ~new_new_n27376__;
  assign new_new_n27378__ = ~new_new_n27374__ & new_new_n27377__;
  assign new_new_n27379__ = new_new_n10694__ & new_new_n26774__;
  assign new_new_n27380__ = pi08 & ~new_new_n27379__;
  assign new_new_n27381__ = new_new_n12121__ & new_new_n26774__;
  assign new_new_n27382__ = ~new_new_n27380__ & ~new_new_n27381__;
  assign new_new_n27383__ = new_new_n27378__ & ~new_new_n27382__;
  assign new_new_n27384__ = ~pi08 & ~new_new_n27378__;
  assign new_new_n27385__ = ~new_new_n27383__ & ~new_new_n27384__;
  assign new_new_n27386__ = ~new_new_n27326__ & ~new_new_n27327__;
  assign new_new_n27387__ = new_new_n26802__ & ~new_new_n27386__;
  assign new_new_n27388__ = new_new_n26741__ & ~new_new_n27226__;
  assign new_new_n27389__ = new_new_n26810__ & ~new_new_n27388__;
  assign new_new_n27390__ = ~new_new_n27325__ & ~new_new_n27388__;
  assign new_new_n27391__ = new_new_n26802__ & ~new_new_n27390__;
  assign new_new_n27392__ = new_new_n27327__ & ~new_new_n27390__;
  assign new_new_n27393__ = ~new_new_n27389__ & ~new_new_n27391__;
  assign new_new_n27394__ = ~new_new_n27392__ & new_new_n27393__;
  assign new_new_n27395__ = ~new_new_n27387__ & ~new_new_n27394__;
  assign new_new_n27396__ = new_new_n11378__ & new_new_n27395__;
  assign new_new_n27397__ = ~new_new_n11409__ & ~new_new_n26741__;
  assign new_new_n27398__ = new_new_n10702__ & ~new_new_n26802__;
  assign new_new_n27399__ = new_new_n10698__ & new_new_n26810__;
  assign new_new_n27400__ = ~new_new_n27397__ & ~new_new_n27398__;
  assign new_new_n27401__ = ~new_new_n27399__ & new_new_n27400__;
  assign new_new_n27402__ = ~new_new_n27396__ & new_new_n27401__;
  assign new_new_n27403__ = ~pi08 & new_new_n27402__;
  assign new_new_n27404__ = pi08 & ~new_new_n27402__;
  assign new_new_n27405__ = ~new_new_n27403__ & ~new_new_n27404__;
  assign new_new_n27406__ = new_new_n8858__ & ~new_new_n27221__;
  assign new_new_n27407__ = ~new_new_n8479__ & new_new_n26847__;
  assign new_new_n27408__ = new_new_n8474__ & ~new_new_n26823__;
  assign new_new_n27409__ = ~new_new_n27191__ & ~new_new_n27221__;
  assign new_new_n27410__ = new_new_n27191__ & new_new_n27221__;
  assign new_new_n27411__ = ~new_new_n27409__ & ~new_new_n27410__;
  assign new_new_n27412__ = new_new_n8470__ & new_new_n27411__;
  assign new_new_n27413__ = ~new_new_n27407__ & ~new_new_n27408__;
  assign new_new_n27414__ = ~new_new_n27406__ & new_new_n27413__;
  assign new_new_n27415__ = ~new_new_n27412__ & new_new_n27414__;
  assign new_new_n27416__ = new_new_n6991__ & new_new_n26922__;
  assign new_new_n27417__ = new_new_n6985__ & ~new_new_n26888__;
  assign new_new_n27418__ = ~new_new_n27416__ & ~new_new_n27417__;
  assign new_new_n27419__ = ~new_new_n26888__ & ~new_new_n27176__;
  assign new_new_n27420__ = new_new_n26888__ & ~new_new_n27175__;
  assign new_new_n27421__ = ~new_new_n27419__ & ~new_new_n27420__;
  assign new_new_n27422__ = new_new_n26854__ & ~new_new_n27421__;
  assign new_new_n27423__ = new_new_n6994__ & ~new_new_n27422__;
  assign new_new_n27424__ = ~new_new_n26854__ & ~new_new_n27421__;
  assign new_new_n27425__ = new_new_n27423__ & new_new_n27424__;
  assign new_new_n27426__ = new_new_n27418__ & ~new_new_n27425__;
  assign new_new_n27427__ = ~pi14 & ~new_new_n27426__;
  assign new_new_n27428__ = pi13 & ~new_new_n26854__;
  assign new_new_n27429__ = new_new_n26854__ & new_new_n27421__;
  assign new_new_n27430__ = ~new_new_n27424__ & ~new_new_n27429__;
  assign new_new_n27431__ = ~pi13 & ~new_new_n27430__;
  assign new_new_n27432__ = new_new_n27423__ & ~new_new_n27428__;
  assign new_new_n27433__ = ~new_new_n27431__ & new_new_n27432__;
  assign new_new_n27434__ = pi14 & new_new_n27418__;
  assign new_new_n27435__ = ~new_new_n27423__ & new_new_n27434__;
  assign new_new_n27436__ = ~new_new_n27433__ & ~new_new_n27435__;
  assign new_new_n27437__ = ~new_new_n27427__ & new_new_n27436__;
  assign new_new_n27438__ = new_new_n7935__ & new_new_n26917__;
  assign new_new_n27439__ = new_new_n6968__ & new_new_n26928__;
  assign new_new_n27440__ = new_new_n6964__ & ~new_new_n26941__;
  assign new_new_n27441__ = new_new_n26928__ & ~new_new_n26941__;
  assign new_new_n27442__ = ~new_new_n27159__ & ~new_new_n27441__;
  assign new_new_n27443__ = new_new_n26917__ & ~new_new_n27442__;
  assign new_new_n27444__ = new_new_n26917__ & new_new_n27153__;
  assign new_new_n27445__ = new_new_n26928__ & ~new_new_n27128__;
  assign new_new_n27446__ = new_new_n26942__ & new_new_n27445__;
  assign new_new_n27447__ = ~new_new_n27444__ & ~new_new_n27446__;
  assign new_new_n27448__ = new_new_n26937__ & ~new_new_n27447__;
  assign new_new_n27449__ = new_new_n26929__ & ~new_new_n26941__;
  assign new_new_n27450__ = new_new_n27128__ & new_new_n27449__;
  assign new_new_n27451__ = new_new_n26917__ & new_new_n26928__;
  assign new_new_n27452__ = new_new_n27152__ & new_new_n27451__;
  assign new_new_n27453__ = ~new_new_n27450__ & ~new_new_n27452__;
  assign new_new_n27454__ = ~new_new_n26937__ & ~new_new_n27453__;
  assign new_new_n27455__ = new_new_n27128__ & new_new_n27451__;
  assign new_new_n27456__ = ~new_new_n27449__ & ~new_new_n27455__;
  assign new_new_n27457__ = new_new_n27152__ & ~new_new_n27456__;
  assign new_new_n27458__ = ~new_new_n26929__ & new_new_n27158__;
  assign new_new_n27459__ = ~new_new_n27448__ & ~new_new_n27457__;
  assign new_new_n27460__ = ~new_new_n27458__ & new_new_n27459__;
  assign new_new_n27461__ = ~new_new_n27454__ & new_new_n27460__;
  assign new_new_n27462__ = ~new_new_n27443__ & new_new_n27461__;
  assign new_new_n27463__ = new_new_n6959__ & ~new_new_n27462__;
  assign new_new_n27464__ = ~new_new_n27439__ & ~new_new_n27440__;
  assign new_new_n27465__ = ~new_new_n27438__ & new_new_n27464__;
  assign new_new_n27466__ = ~new_new_n27463__ & new_new_n27465__;
  assign new_new_n27467__ = pi17 & ~new_new_n27466__;
  assign new_new_n27468__ = ~pi17 & new_new_n27466__;
  assign new_new_n27469__ = ~new_new_n27467__ & ~new_new_n27468__;
  assign new_new_n27470__ = new_new_n6964__ & new_new_n27152__;
  assign new_new_n27471__ = new_new_n6968__ & ~new_new_n26941__;
  assign new_new_n27472__ = new_new_n7935__ & new_new_n26928__;
  assign new_new_n27473__ = ~new_new_n27470__ & ~new_new_n27471__;
  assign new_new_n27474__ = ~new_new_n27472__ & new_new_n27473__;
  assign new_new_n27475__ = new_new_n26937__ & ~new_new_n27128__;
  assign new_new_n27476__ = ~new_new_n26937__ & ~new_new_n27124__;
  assign new_new_n27477__ = ~new_new_n27475__ & ~new_new_n27476__;
  assign new_new_n27478__ = new_new_n27128__ & ~new_new_n27152__;
  assign new_new_n27479__ = ~new_new_n27128__ & new_new_n27152__;
  assign new_new_n27480__ = ~new_new_n27478__ & ~new_new_n27479__;
  assign new_new_n27481__ = ~new_new_n27477__ & ~new_new_n27480__;
  assign new_new_n27482__ = ~new_new_n26941__ & new_new_n27481__;
  assign new_new_n27483__ = ~new_new_n27152__ & ~new_new_n27482__;
  assign new_new_n27484__ = new_new_n26941__ & new_new_n27481__;
  assign new_new_n27485__ = ~new_new_n27483__ & ~new_new_n27484__;
  assign new_new_n27486__ = new_new_n27442__ & new_new_n27485__;
  assign new_new_n27487__ = ~new_new_n27442__ & ~new_new_n27485__;
  assign new_new_n27488__ = ~new_new_n27486__ & ~new_new_n27487__;
  assign new_new_n27489__ = new_new_n6958__ & new_new_n27488__;
  assign new_new_n27490__ = ~pi17 & ~new_new_n27489__;
  assign new_new_n27491__ = new_new_n8160__ & new_new_n27488__;
  assign new_new_n27492__ = ~new_new_n27490__ & ~new_new_n27491__;
  assign new_new_n27493__ = new_new_n27474__ & ~new_new_n27492__;
  assign new_new_n27494__ = pi17 & ~new_new_n27474__;
  assign new_new_n27495__ = ~new_new_n27493__ & ~new_new_n27494__;
  assign new_new_n27496__ = new_new_n6968__ & new_new_n27152__;
  assign new_new_n27497__ = new_new_n6964__ & ~new_new_n26937__;
  assign new_new_n27498__ = new_new_n7935__ & ~new_new_n26941__;
  assign new_new_n27499__ = ~new_new_n27497__ & ~new_new_n27498__;
  assign new_new_n27500__ = ~new_new_n27496__ & new_new_n27499__;
  assign new_new_n27501__ = ~new_new_n26941__ & ~new_new_n27481__;
  assign new_new_n27502__ = ~new_new_n27484__ & ~new_new_n27501__;
  assign new_new_n27503__ = new_new_n6958__ & ~new_new_n27502__;
  assign new_new_n27504__ = pi17 & ~new_new_n27503__;
  assign new_new_n27505__ = new_new_n7942__ & ~new_new_n27502__;
  assign new_new_n27506__ = ~new_new_n27504__ & ~new_new_n27505__;
  assign new_new_n27507__ = new_new_n27500__ & ~new_new_n27506__;
  assign new_new_n27508__ = ~pi17 & ~new_new_n27500__;
  assign new_new_n27509__ = ~new_new_n27507__ & ~new_new_n27508__;
  assign new_new_n27510__ = ~pi17 & new_new_n7942__;
  assign new_new_n27511__ = new_new_n27152__ & new_new_n27510__;
  assign new_new_n27512__ = new_new_n7935__ & new_new_n27152__;
  assign new_new_n27513__ = new_new_n6964__ & new_new_n26971__;
  assign new_new_n27514__ = new_new_n6968__ & ~new_new_n26937__;
  assign new_new_n27515__ = ~new_new_n27513__ & ~new_new_n27514__;
  assign new_new_n27516__ = ~new_new_n27512__ & new_new_n27515__;
  assign new_new_n27517__ = pi17 & ~new_new_n27152__;
  assign new_new_n27518__ = new_new_n27516__ & new_new_n27517__;
  assign new_new_n27519__ = ~new_new_n27511__ & ~new_new_n27518__;
  assign new_new_n27520__ = ~new_new_n27477__ & ~new_new_n27519__;
  assign new_new_n27521__ = ~new_new_n27152__ & new_new_n27510__;
  assign new_new_n27522__ = pi17 & new_new_n27152__;
  assign new_new_n27523__ = new_new_n27516__ & new_new_n27522__;
  assign new_new_n27524__ = ~new_new_n27521__ & ~new_new_n27523__;
  assign new_new_n27525__ = new_new_n27477__ & ~new_new_n27524__;
  assign new_new_n27526__ = ~pi17 & ~new_new_n27516__;
  assign new_new_n27527__ = pi17 & ~new_new_n8160__;
  assign new_new_n27528__ = new_new_n27516__ & new_new_n27527__;
  assign new_new_n27529__ = ~new_new_n27526__ & ~new_new_n27528__;
  assign new_new_n27530__ = ~new_new_n27520__ & new_new_n27529__;
  assign new_new_n27531__ = ~new_new_n27525__ & new_new_n27530__;
  assign new_new_n27532__ = new_new_n5191__ & new_new_n27041__;
  assign new_new_n27533__ = new_new_n5183__ & ~new_new_n27054__;
  assign new_new_n27534__ = ~new_new_n27532__ & ~new_new_n27533__;
  assign new_new_n27535__ = new_new_n27033__ & new_new_n27102__;
  assign new_new_n27536__ = new_new_n5195__ & ~new_new_n27535__;
  assign new_new_n27537__ = pi23 & ~new_new_n27536__;
  assign new_new_n27538__ = ~pi22 & new_new_n27033__;
  assign new_new_n27539__ = pi22 & ~new_new_n27033__;
  assign new_new_n27540__ = new_new_n5195__ & ~new_new_n27538__;
  assign new_new_n27541__ = ~new_new_n27539__ & new_new_n27540__;
  assign new_new_n27542__ = ~new_new_n27102__ & new_new_n27541__;
  assign new_new_n27543__ = ~new_new_n27537__ & ~new_new_n27542__;
  assign new_new_n27544__ = new_new_n27534__ & ~new_new_n27543__;
  assign new_new_n27545__ = ~new_new_n27033__ & new_new_n27102__;
  assign new_new_n27546__ = new_new_n5195__ & new_new_n27545__;
  assign new_new_n27547__ = new_new_n27534__ & ~new_new_n27546__;
  assign new_new_n27548__ = ~pi23 & ~new_new_n27547__;
  assign new_new_n27549__ = ~new_new_n27544__ & ~new_new_n27548__;
  assign new_new_n27550__ = new_new_n5213__ & new_new_n27041__;
  assign new_new_n27551__ = new_new_n5183__ & ~new_new_n27071__;
  assign new_new_n27552__ = new_new_n5191__ & new_new_n27059__;
  assign new_new_n27553__ = ~new_new_n27059__ & new_new_n27075__;
  assign new_new_n27554__ = new_new_n26118__ & ~new_new_n27553__;
  assign new_new_n27555__ = new_new_n27071__ & new_new_n27554__;
  assign new_new_n27556__ = ~new_new_n27071__ & ~new_new_n27554__;
  assign new_new_n27557__ = ~new_new_n27555__ & ~new_new_n27556__;
  assign new_new_n27558__ = ~new_new_n27041__ & new_new_n27557__;
  assign new_new_n27559__ = ~new_new_n27041__ & new_new_n27554__;
  assign new_new_n27560__ = new_new_n27041__ & new_new_n27556__;
  assign new_new_n27561__ = ~new_new_n27559__ & ~new_new_n27560__;
  assign new_new_n27562__ = ~new_new_n27059__ & ~new_new_n27561__;
  assign new_new_n27563__ = new_new_n27041__ & ~new_new_n27555__;
  assign new_new_n27564__ = new_new_n27059__ & ~new_new_n27559__;
  assign new_new_n27565__ = ~new_new_n27563__ & new_new_n27564__;
  assign new_new_n27566__ = ~new_new_n27562__ & ~new_new_n27565__;
  assign new_new_n27567__ = ~new_new_n27558__ & new_new_n27566__;
  assign new_new_n27568__ = new_new_n5215__ & new_new_n27567__;
  assign new_new_n27569__ = ~new_new_n27550__ & ~new_new_n27552__;
  assign new_new_n27570__ = ~new_new_n27551__ & new_new_n27569__;
  assign new_new_n27571__ = ~new_new_n27568__ & new_new_n27570__;
  assign new_new_n27572__ = pi23 & ~new_new_n27571__;
  assign new_new_n27573__ = ~pi23 & new_new_n27571__;
  assign new_new_n27574__ = ~new_new_n27572__ & ~new_new_n27573__;
  assign new_new_n27575__ = ~new_new_n110__ & ~new_new_n27075__;
  assign new_new_n27576__ = new_new_n5183__ & ~new_new_n27075__;
  assign new_new_n27577__ = ~new_new_n26118__ & new_new_n27075__;
  assign new_new_n27578__ = new_new_n5195__ & ~new_new_n27577__;
  assign new_new_n27579__ = ~new_new_n27576__ & ~new_new_n27578__;
  assign new_new_n27580__ = new_new_n5191__ & ~new_new_n27075__;
  assign new_new_n27581__ = new_new_n5183__ & new_new_n26118__;
  assign new_new_n27582__ = new_new_n26118__ & new_new_n27075__;
  assign new_new_n27583__ = new_new_n5212__ & new_new_n27582__;
  assign new_new_n27584__ = ~new_new_n27059__ & ~new_new_n27583__;
  assign new_new_n27585__ = new_new_n27059__ & new_new_n27583__;
  assign new_new_n27586__ = new_new_n5195__ & ~new_new_n27584__;
  assign new_new_n27587__ = ~new_new_n27585__ & new_new_n27586__;
  assign new_new_n27588__ = ~new_new_n27580__ & ~new_new_n27581__;
  assign new_new_n27589__ = ~new_new_n27587__ & new_new_n27588__;
  assign new_new_n27590__ = pi23 & new_new_n27579__;
  assign new_new_n27591__ = new_new_n27589__ & new_new_n27590__;
  assign new_new_n27592__ = ~new_new_n27575__ & ~new_new_n27591__;
  assign new_new_n27593__ = new_new_n5213__ & ~new_new_n27071__;
  assign new_new_n27594__ = new_new_n5191__ & new_new_n26118__;
  assign new_new_n27595__ = new_new_n5183__ & new_new_n27059__;
  assign new_new_n27596__ = ~new_new_n27594__ & ~new_new_n27595__;
  assign new_new_n27597__ = ~new_new_n27593__ & new_new_n27596__;
  assign new_new_n27598__ = new_new_n27059__ & ~new_new_n27557__;
  assign new_new_n27599__ = ~new_new_n27059__ & new_new_n27557__;
  assign new_new_n27600__ = ~new_new_n27598__ & ~new_new_n27599__;
  assign new_new_n27601__ = new_new_n5195__ & new_new_n27600__;
  assign new_new_n27602__ = ~pi23 & ~new_new_n27601__;
  assign new_new_n27603__ = new_new_n5974__ & new_new_n27600__;
  assign new_new_n27604__ = ~new_new_n27602__ & ~new_new_n27603__;
  assign new_new_n27605__ = new_new_n27597__ & ~new_new_n27604__;
  assign new_new_n27606__ = pi23 & ~new_new_n27597__;
  assign new_new_n27607__ = ~new_new_n27605__ & ~new_new_n27606__;
  assign new_new_n27608__ = ~new_new_n27592__ & new_new_n27607__;
  assign new_new_n27609__ = ~new_new_n27574__ & ~new_new_n27608__;
  assign new_new_n27610__ = new_new_n419__ & new_new_n27087__;
  assign new_new_n27611__ = ~new_new_n104__ & new_new_n26118__;
  assign new_new_n27612__ = new_new_n389__ & ~new_new_n27611__;
  assign new_new_n27613__ = new_new_n110__ & new_new_n27582__;
  assign new_new_n27614__ = ~new_new_n146__ & ~new_new_n27577__;
  assign new_new_n27615__ = ~new_new_n27610__ & new_new_n27614__;
  assign new_new_n27616__ = ~new_new_n27612__ & ~new_new_n27613__;
  assign new_new_n27617__ = new_new_n27615__ & new_new_n27616__;
  assign new_new_n27618__ = new_new_n27574__ & new_new_n27608__;
  assign new_new_n27619__ = ~new_new_n27609__ & ~new_new_n27618__;
  assign new_new_n27620__ = ~new_new_n27617__ & new_new_n27619__;
  assign new_new_n27621__ = ~new_new_n27609__ & ~new_new_n27620__;
  assign new_new_n27622__ = new_new_n5213__ & ~new_new_n27054__;
  assign new_new_n27623__ = new_new_n5191__ & ~new_new_n27071__;
  assign new_new_n27624__ = new_new_n5183__ & new_new_n27041__;
  assign new_new_n27625__ = ~new_new_n27623__ & ~new_new_n27624__;
  assign new_new_n27626__ = ~new_new_n27622__ & new_new_n27625__;
  assign new_new_n27627__ = new_new_n5195__ & ~new_new_n27094__;
  assign new_new_n27628__ = pi23 & ~new_new_n27627__;
  assign new_new_n27629__ = new_new_n7878__ & ~new_new_n27094__;
  assign new_new_n27630__ = ~new_new_n27628__ & ~new_new_n27629__;
  assign new_new_n27631__ = new_new_n27626__ & ~new_new_n27630__;
  assign new_new_n27632__ = ~pi23 & ~new_new_n27626__;
  assign new_new_n27633__ = ~new_new_n27631__ & ~new_new_n27632__;
  assign new_new_n27634__ = ~new_new_n27621__ & new_new_n27633__;
  assign new_new_n27635__ = new_new_n873__ & ~new_new_n27075__;
  assign new_new_n27636__ = new_new_n801__ & ~new_new_n27577__;
  assign new_new_n27637__ = ~new_new_n27635__ & ~new_new_n27636__;
  assign new_new_n27638__ = pi26 & ~new_new_n27637__;
  assign new_new_n27639__ = ~new_new_n333__ & ~new_new_n27075__;
  assign new_new_n27640__ = new_new_n873__ & new_new_n26118__;
  assign new_new_n27641__ = ~new_new_n447__ & new_new_n27582__;
  assign new_new_n27642__ = ~new_new_n27059__ & ~new_new_n27641__;
  assign new_new_n27643__ = new_new_n27059__ & new_new_n27641__;
  assign new_new_n27644__ = new_new_n801__ & ~new_new_n27642__;
  assign new_new_n27645__ = ~new_new_n27643__ & new_new_n27644__;
  assign new_new_n27646__ = ~new_new_n27639__ & ~new_new_n27640__;
  assign new_new_n27647__ = ~new_new_n27645__ & new_new_n27646__;
  assign new_new_n27648__ = ~new_new_n27638__ & new_new_n27647__;
  assign new_new_n27649__ = new_new_n27638__ & ~new_new_n27647__;
  assign new_new_n27650__ = ~new_new_n27648__ & ~new_new_n27649__;
  assign new_new_n27651__ = new_new_n27621__ & ~new_new_n27633__;
  assign new_new_n27652__ = ~new_new_n27650__ & ~new_new_n27651__;
  assign new_new_n27653__ = ~new_new_n27634__ & ~new_new_n27652__;
  assign new_new_n27654__ = new_new_n27549__ & ~new_new_n27653__;
  assign new_new_n27655__ = ~new_new_n27549__ & new_new_n27653__;
  assign new_new_n27656__ = new_new_n4214__ & ~new_new_n27075__;
  assign new_new_n27657__ = new_new_n3311__ & ~new_new_n27071__;
  assign new_new_n27658__ = new_new_n873__ & new_new_n27059__;
  assign new_new_n27659__ = ~new_new_n4900__ & new_new_n27600__;
  assign new_new_n27660__ = ~new_new_n27657__ & ~new_new_n27658__;
  assign new_new_n27661__ = ~new_new_n27659__ & new_new_n27660__;
  assign new_new_n27662__ = ~pi26 & ~new_new_n27661__;
  assign new_new_n27663__ = new_new_n349__ & new_new_n26118__;
  assign new_new_n27664__ = pi26 & ~new_new_n27663__;
  assign new_new_n27665__ = new_new_n146__ & new_new_n26118__;
  assign new_new_n27666__ = ~new_new_n27664__ & ~new_new_n27665__;
  assign new_new_n27667__ = new_new_n27661__ & ~new_new_n27666__;
  assign new_new_n27668__ = ~new_new_n27662__ & ~new_new_n27667__;
  assign new_new_n27669__ = pi26 & new_new_n27648__;
  assign new_new_n27670__ = ~new_new_n27668__ & ~new_new_n27669__;
  assign new_new_n27671__ = new_new_n27656__ & ~new_new_n27670__;
  assign new_new_n27672__ = new_new_n27656__ & ~new_new_n27668__;
  assign new_new_n27673__ = ~new_new_n27668__ & new_new_n27669__;
  assign new_new_n27674__ = ~new_new_n27672__ & ~new_new_n27673__;
  assign new_new_n27675__ = new_new_n27668__ & ~new_new_n27669__;
  assign new_new_n27676__ = new_new_n27674__ & ~new_new_n27675__;
  assign new_new_n27677__ = ~new_new_n27671__ & ~new_new_n27676__;
  assign new_new_n27678__ = ~new_new_n27655__ & new_new_n27677__;
  assign new_new_n27679__ = ~new_new_n27654__ & ~new_new_n27678__;
  assign new_new_n27680__ = new_new_n5183__ & ~new_new_n27033__;
  assign new_new_n27681__ = new_new_n5191__ & ~new_new_n27054__;
  assign new_new_n27682__ = ~new_new_n27680__ & ~new_new_n27681__;
  assign new_new_n27683__ = new_new_n27033__ & new_new_n27054__;
  assign new_new_n27684__ = ~new_new_n27033__ & ~new_new_n27054__;
  assign new_new_n27685__ = ~new_new_n27683__ & ~new_new_n27684__;
  assign new_new_n27686__ = new_new_n27102__ & new_new_n27685__;
  assign new_new_n27687__ = new_new_n27111__ & ~new_new_n27686__;
  assign new_new_n27688__ = new_new_n5195__ & new_new_n27687__;
  assign new_new_n27689__ = new_new_n27682__ & ~new_new_n27688__;
  assign new_new_n27690__ = pi23 & ~new_new_n27689__;
  assign new_new_n27691__ = ~new_new_n27111__ & ~new_new_n27686__;
  assign new_new_n27692__ = new_new_n5195__ & ~new_new_n27691__;
  assign new_new_n27693__ = ~pi23 & ~new_new_n27692__;
  assign new_new_n27694__ = ~pi22 & new_new_n27111__;
  assign new_new_n27695__ = pi22 & ~new_new_n27111__;
  assign new_new_n27696__ = new_new_n5195__ & ~new_new_n27694__;
  assign new_new_n27697__ = ~new_new_n27695__ & new_new_n27696__;
  assign new_new_n27698__ = new_new_n27686__ & new_new_n27697__;
  assign new_new_n27699__ = ~new_new_n27693__ & ~new_new_n27698__;
  assign new_new_n27700__ = new_new_n27682__ & ~new_new_n27699__;
  assign new_new_n27701__ = ~new_new_n27690__ & ~new_new_n27700__;
  assign new_new_n27702__ = new_new_n3311__ & new_new_n27041__;
  assign new_new_n27703__ = ~new_new_n333__ & new_new_n27059__;
  assign new_new_n27704__ = new_new_n873__ & ~new_new_n27071__;
  assign new_new_n27705__ = ~new_new_n27702__ & ~new_new_n27703__;
  assign new_new_n27706__ = ~new_new_n27704__ & new_new_n27705__;
  assign new_new_n27707__ = new_new_n512__ & new_new_n27567__;
  assign new_new_n27708__ = new_new_n801__ & new_new_n27567__;
  assign new_new_n27709__ = pi26 & ~new_new_n27708__;
  assign new_new_n27710__ = ~new_new_n27707__ & ~new_new_n27709__;
  assign new_new_n27711__ = new_new_n27706__ & ~new_new_n27710__;
  assign new_new_n27712__ = new_new_n27669__ & ~new_new_n27711__;
  assign new_new_n27713__ = ~pi26 & ~new_new_n27706__;
  assign new_new_n27714__ = ~new_new_n27711__ & ~new_new_n27713__;
  assign new_new_n27715__ = new_new_n4210__ & new_new_n27087__;
  assign new_new_n27716__ = ~new_new_n4214__ & new_new_n27582__;
  assign new_new_n27717__ = ~new_new_n4209__ & new_new_n26118__;
  assign new_new_n27718__ = new_new_n4211__ & ~new_new_n27717__;
  assign new_new_n27719__ = ~new_new_n66__ & ~new_new_n27577__;
  assign new_new_n27720__ = ~new_new_n27715__ & new_new_n27719__;
  assign new_new_n27721__ = ~new_new_n27716__ & ~new_new_n27718__;
  assign new_new_n27722__ = new_new_n27720__ & new_new_n27721__;
  assign new_new_n27723__ = new_new_n27714__ & ~new_new_n27722__;
  assign new_new_n27724__ = ~new_new_n27714__ & new_new_n27722__;
  assign new_new_n27725__ = ~new_new_n27723__ & ~new_new_n27724__;
  assign new_new_n27726__ = ~new_new_n27674__ & ~new_new_n27712__;
  assign new_new_n27727__ = new_new_n27725__ & new_new_n27726__;
  assign new_new_n27728__ = new_new_n27674__ & ~new_new_n27725__;
  assign new_new_n27729__ = ~new_new_n27727__ & ~new_new_n27728__;
  assign new_new_n27730__ = ~new_new_n27701__ & ~new_new_n27729__;
  assign new_new_n27731__ = new_new_n27701__ & new_new_n27729__;
  assign new_new_n27732__ = ~new_new_n27730__ & ~new_new_n27731__;
  assign new_new_n27733__ = new_new_n27679__ & ~new_new_n27732__;
  assign new_new_n27734__ = ~new_new_n27679__ & new_new_n27732__;
  assign new_new_n27735__ = ~new_new_n27733__ & ~new_new_n27734__;
  assign new_new_n27736__ = new_new_n6629__ & ~new_new_n27021__;
  assign new_new_n27737__ = ~new_new_n6625__ & new_new_n27111__;
  assign new_new_n27738__ = new_new_n6634__ & ~new_new_n27029__;
  assign new_new_n27739__ = ~new_new_n27736__ & ~new_new_n27737__;
  assign new_new_n27740__ = ~new_new_n27738__ & new_new_n27739__;
  assign new_new_n27741__ = new_new_n27033__ & new_new_n27111__;
  assign new_new_n27742__ = ~new_new_n27033__ & ~new_new_n27111__;
  assign new_new_n27743__ = ~new_new_n27741__ & ~new_new_n27742__;
  assign new_new_n27744__ = new_new_n27021__ & new_new_n27033__;
  assign new_new_n27745__ = ~new_new_n27021__ & ~new_new_n27033__;
  assign new_new_n27746__ = ~new_new_n27744__ & ~new_new_n27745__;
  assign new_new_n27747__ = new_new_n27743__ & new_new_n27746__;
  assign new_new_n27748__ = new_new_n27021__ & new_new_n27111__;
  assign new_new_n27749__ = ~new_new_n27054__ & new_new_n27748__;
  assign new_new_n27750__ = ~new_new_n27021__ & ~new_new_n27111__;
  assign new_new_n27751__ = new_new_n27054__ & new_new_n27750__;
  assign new_new_n27752__ = ~new_new_n27749__ & ~new_new_n27751__;
  assign new_new_n27753__ = new_new_n27102__ & ~new_new_n27752__;
  assign new_new_n27754__ = ~new_new_n27747__ & ~new_new_n27753__;
  assign new_new_n27755__ = ~new_new_n27029__ & ~new_new_n27754__;
  assign new_new_n27756__ = ~new_new_n27111__ & ~new_new_n27684__;
  assign new_new_n27757__ = new_new_n27021__ & ~new_new_n27683__;
  assign new_new_n27758__ = ~new_new_n27756__ & ~new_new_n27757__;
  assign new_new_n27759__ = new_new_n27021__ & ~new_new_n27111__;
  assign new_new_n27760__ = ~new_new_n27102__ & ~new_new_n27746__;
  assign new_new_n27761__ = ~new_new_n27758__ & ~new_new_n27759__;
  assign new_new_n27762__ = ~new_new_n27760__ & new_new_n27761__;
  assign new_new_n27763__ = new_new_n27029__ & ~new_new_n27762__;
  assign new_new_n27764__ = ~new_new_n27755__ & ~new_new_n27763__;
  assign new_new_n27765__ = new_new_n6631__ & new_new_n27764__;
  assign new_new_n27766__ = pi20 & ~new_new_n27765__;
  assign new_new_n27767__ = new_new_n6640__ & new_new_n27764__;
  assign new_new_n27768__ = ~new_new_n27766__ & ~new_new_n27767__;
  assign new_new_n27769__ = new_new_n27740__ & ~new_new_n27768__;
  assign new_new_n27770__ = ~pi20 & ~new_new_n27740__;
  assign new_new_n27771__ = ~new_new_n27769__ & ~new_new_n27770__;
  assign new_new_n27772__ = new_new_n6629__ & new_new_n27111__;
  assign new_new_n27773__ = ~new_new_n6625__ & ~new_new_n27033__;
  assign new_new_n27774__ = new_new_n6634__ & ~new_new_n27021__;
  assign new_new_n27775__ = ~new_new_n27772__ & ~new_new_n27773__;
  assign new_new_n27776__ = ~new_new_n27774__ & new_new_n27775__;
  assign new_new_n27777__ = new_new_n27021__ & new_new_n27743__;
  assign new_new_n27778__ = ~new_new_n27033__ & new_new_n27750__;
  assign new_new_n27779__ = new_new_n27097__ & new_new_n27778__;
  assign new_new_n27780__ = ~new_new_n27749__ & ~new_new_n27779__;
  assign new_new_n27781__ = new_new_n27041__ & ~new_new_n27780__;
  assign new_new_n27782__ = ~new_new_n27021__ & new_new_n27741__;
  assign new_new_n27783__ = ~new_new_n27097__ & new_new_n27759__;
  assign new_new_n27784__ = ~new_new_n27782__ & ~new_new_n27783__;
  assign new_new_n27785__ = new_new_n27054__ & ~new_new_n27784__;
  assign new_new_n27786__ = new_new_n27054__ & new_new_n27759__;
  assign new_new_n27787__ = ~new_new_n27097__ & new_new_n27782__;
  assign new_new_n27788__ = ~new_new_n27786__ & ~new_new_n27787__;
  assign new_new_n27789__ = ~new_new_n27041__ & ~new_new_n27788__;
  assign new_new_n27790__ = new_new_n27097__ & new_new_n27748__;
  assign new_new_n27791__ = ~new_new_n27778__ & ~new_new_n27790__;
  assign new_new_n27792__ = ~new_new_n27054__ & ~new_new_n27791__;
  assign new_new_n27793__ = ~new_new_n27785__ & ~new_new_n27789__;
  assign new_new_n27794__ = ~new_new_n27792__ & new_new_n27793__;
  assign new_new_n27795__ = ~new_new_n27781__ & new_new_n27794__;
  assign new_new_n27796__ = ~new_new_n27777__ & new_new_n27795__;
  assign new_new_n27797__ = new_new_n6631__ & new_new_n27796__;
  assign new_new_n27798__ = ~pi20 & ~new_new_n27797__;
  assign new_new_n27799__ = new_new_n7015__ & new_new_n27796__;
  assign new_new_n27800__ = ~new_new_n27798__ & ~new_new_n27799__;
  assign new_new_n27801__ = new_new_n27776__ & ~new_new_n27800__;
  assign new_new_n27802__ = pi20 & ~new_new_n27776__;
  assign new_new_n27803__ = ~new_new_n27801__ & ~new_new_n27802__;
  assign new_new_n27804__ = new_new_n6629__ & ~new_new_n27054__;
  assign new_new_n27805__ = ~new_new_n6625__ & new_new_n27041__;
  assign new_new_n27806__ = ~new_new_n6633__ & ~new_new_n27102__;
  assign new_new_n27807__ = new_new_n27033__ & ~new_new_n27806__;
  assign new_new_n27808__ = ~new_new_n27033__ & new_new_n27806__;
  assign new_new_n27809__ = new_new_n6631__ & ~new_new_n27807__;
  assign new_new_n27810__ = ~new_new_n27808__ & new_new_n27809__;
  assign new_new_n27811__ = ~new_new_n27804__ & ~new_new_n27805__;
  assign new_new_n27812__ = ~new_new_n27810__ & new_new_n27811__;
  assign new_new_n27813__ = ~pi20 & ~new_new_n27812__;
  assign new_new_n27814__ = pi20 & new_new_n27812__;
  assign new_new_n27815__ = ~new_new_n27813__ & ~new_new_n27814__;
  assign new_new_n27816__ = new_new_n27575__ & ~new_new_n27607__;
  assign new_new_n27817__ = ~new_new_n27575__ & new_new_n27607__;
  assign new_new_n27818__ = new_new_n27591__ & ~new_new_n27817__;
  assign new_new_n27819__ = new_new_n26508__ & ~new_new_n27577__;
  assign new_new_n27820__ = new_new_n27589__ & ~new_new_n27819__;
  assign new_new_n27821__ = pi23 & ~new_new_n27579__;
  assign new_new_n27822__ = ~new_new_n27589__ & new_new_n27821__;
  assign new_new_n27823__ = ~new_new_n27820__ & ~new_new_n27822__;
  assign new_new_n27824__ = new_new_n6634__ & ~new_new_n27054__;
  assign new_new_n27825__ = ~new_new_n6625__ & ~new_new_n27071__;
  assign new_new_n27826__ = new_new_n6629__ & new_new_n27041__;
  assign new_new_n27827__ = new_new_n6936__ & ~new_new_n27094__;
  assign new_new_n27828__ = ~new_new_n27825__ & ~new_new_n27826__;
  assign new_new_n27829__ = ~new_new_n27824__ & new_new_n27828__;
  assign new_new_n27830__ = ~new_new_n27827__ & new_new_n27829__;
  assign new_new_n27831__ = new_new_n6629__ & ~new_new_n27071__;
  assign new_new_n27832__ = ~new_new_n6625__ & new_new_n27059__;
  assign new_new_n27833__ = new_new_n6634__ & new_new_n27041__;
  assign new_new_n27834__ = ~new_new_n27831__ & ~new_new_n27832__;
  assign new_new_n27835__ = ~new_new_n27833__ & new_new_n27834__;
  assign new_new_n27836__ = new_new_n6631__ & new_new_n27567__;
  assign new_new_n27837__ = ~pi20 & ~new_new_n27836__;
  assign new_new_n27838__ = new_new_n7015__ & new_new_n27567__;
  assign new_new_n27839__ = ~new_new_n27837__ & ~new_new_n27838__;
  assign new_new_n27840__ = new_new_n27835__ & ~new_new_n27839__;
  assign new_new_n27841__ = pi20 & ~new_new_n27835__;
  assign new_new_n27842__ = ~new_new_n27840__ & ~new_new_n27841__;
  assign new_new_n27843__ = new_new_n9921__ & ~new_new_n27577__;
  assign new_new_n27844__ = ~new_new_n6633__ & new_new_n26118__;
  assign new_new_n27845__ = new_new_n27059__ & ~new_new_n27844__;
  assign new_new_n27846__ = ~new_new_n27059__ & new_new_n27582__;
  assign new_new_n27847__ = ~new_new_n6633__ & new_new_n27846__;
  assign new_new_n27848__ = ~new_new_n27845__ & ~new_new_n27847__;
  assign new_new_n27849__ = new_new_n6631__ & ~new_new_n27848__;
  assign new_new_n27850__ = new_new_n6631__ & new_new_n27059__;
  assign new_new_n27851__ = new_new_n6625__ & ~new_new_n27850__;
  assign new_new_n27852__ = ~new_new_n27075__ & ~new_new_n27851__;
  assign new_new_n27853__ = ~new_new_n27849__ & ~new_new_n27852__;
  assign new_new_n27854__ = ~new_new_n27843__ & new_new_n27853__;
  assign new_new_n27855__ = ~pi21 & ~new_new_n27075__;
  assign new_new_n27856__ = ~new_new_n27854__ & ~new_new_n27855__;
  assign new_new_n27857__ = ~new_new_n6625__ & new_new_n26118__;
  assign new_new_n27858__ = new_new_n6629__ & new_new_n27059__;
  assign new_new_n27859__ = ~new_new_n6633__ & ~new_new_n27600__;
  assign new_new_n27860__ = new_new_n6633__ & new_new_n27071__;
  assign new_new_n27861__ = new_new_n6631__ & ~new_new_n27860__;
  assign new_new_n27862__ = ~new_new_n27859__ & new_new_n27861__;
  assign new_new_n27863__ = ~new_new_n27857__ & ~new_new_n27858__;
  assign new_new_n27864__ = ~new_new_n27862__ & new_new_n27863__;
  assign new_new_n27865__ = pi20 & ~new_new_n27856__;
  assign new_new_n27866__ = new_new_n27864__ & new_new_n27865__;
  assign new_new_n27867__ = ~pi20 & pi21;
  assign new_new_n27868__ = ~new_new_n27075__ & new_new_n27867__;
  assign new_new_n27869__ = ~new_new_n27864__ & new_new_n27868__;
  assign new_new_n27870__ = ~new_new_n27866__ & ~new_new_n27869__;
  assign new_new_n27871__ = ~new_new_n27842__ & new_new_n27870__;
  assign new_new_n27872__ = new_new_n27842__ & ~new_new_n27870__;
  assign new_new_n27873__ = new_new_n5180__ & new_new_n27087__;
  assign new_new_n27874__ = ~new_new_n5195__ & new_new_n27582__;
  assign new_new_n27875__ = ~new_new_n5179__ & new_new_n26118__;
  assign new_new_n27876__ = new_new_n5182__ & ~new_new_n27875__;
  assign new_new_n27877__ = ~new_new_n5189__ & ~new_new_n27577__;
  assign new_new_n27878__ = ~new_new_n27873__ & new_new_n27877__;
  assign new_new_n27879__ = ~new_new_n27874__ & ~new_new_n27876__;
  assign new_new_n27880__ = new_new_n27878__ & new_new_n27879__;
  assign new_new_n27881__ = ~new_new_n27872__ & ~new_new_n27880__;
  assign new_new_n27882__ = ~new_new_n27871__ & ~new_new_n27881__;
  assign new_new_n27883__ = pi20 & ~new_new_n27823__;
  assign new_new_n27884__ = ~pi20 & new_new_n27823__;
  assign new_new_n27885__ = ~new_new_n27883__ & ~new_new_n27884__;
  assign new_new_n27886__ = new_new_n27882__ & ~new_new_n27885__;
  assign new_new_n27887__ = ~new_new_n27882__ & new_new_n27885__;
  assign new_new_n27888__ = ~new_new_n27886__ & ~new_new_n27887__;
  assign new_new_n27889__ = new_new_n27830__ & new_new_n27888__;
  assign new_new_n27890__ = ~new_new_n27830__ & ~new_new_n27888__;
  assign new_new_n27891__ = ~new_new_n27889__ & ~new_new_n27890__;
  assign new_new_n27892__ = ~new_new_n27823__ & ~new_new_n27891__;
  assign new_new_n27893__ = new_new_n27823__ & new_new_n27891__;
  assign new_new_n27894__ = ~new_new_n27882__ & ~new_new_n27893__;
  assign new_new_n27895__ = ~new_new_n27892__ & ~new_new_n27894__;
  assign new_new_n27896__ = ~new_new_n27816__ & ~new_new_n27818__;
  assign new_new_n27897__ = ~new_new_n27895__ & new_new_n27896__;
  assign new_new_n27898__ = ~new_new_n27815__ & ~new_new_n27897__;
  assign new_new_n27899__ = new_new_n27815__ & ~new_new_n27895__;
  assign new_new_n27900__ = new_new_n27817__ & ~new_new_n27899__;
  assign new_new_n27901__ = new_new_n27816__ & new_new_n27895__;
  assign new_new_n27902__ = ~new_new_n27900__ & ~new_new_n27901__;
  assign new_new_n27903__ = ~new_new_n27591__ & ~new_new_n27902__;
  assign new_new_n27904__ = ~new_new_n27898__ & ~new_new_n27903__;
  assign new_new_n27905__ = new_new_n27617__ & ~new_new_n27619__;
  assign new_new_n27906__ = ~new_new_n27620__ & ~new_new_n27905__;
  assign new_new_n27907__ = ~new_new_n27904__ & ~new_new_n27906__;
  assign new_new_n27908__ = new_new_n27904__ & new_new_n27906__;
  assign new_new_n27909__ = ~new_new_n6625__ & ~new_new_n27054__;
  assign new_new_n27910__ = new_new_n6629__ & ~new_new_n27033__;
  assign new_new_n27911__ = ~new_new_n6633__ & new_new_n27686__;
  assign new_new_n27912__ = new_new_n27111__ & new_new_n27911__;
  assign new_new_n27913__ = ~new_new_n27111__ & ~new_new_n27911__;
  assign new_new_n27914__ = new_new_n6631__ & ~new_new_n27912__;
  assign new_new_n27915__ = ~new_new_n27913__ & new_new_n27914__;
  assign new_new_n27916__ = ~new_new_n27909__ & ~new_new_n27910__;
  assign new_new_n27917__ = ~new_new_n27915__ & new_new_n27916__;
  assign new_new_n27918__ = pi20 & ~new_new_n27917__;
  assign new_new_n27919__ = ~pi20 & new_new_n27917__;
  assign new_new_n27920__ = ~new_new_n27918__ & ~new_new_n27919__;
  assign new_new_n27921__ = ~new_new_n27908__ & new_new_n27920__;
  assign new_new_n27922__ = ~new_new_n27907__ & ~new_new_n27921__;
  assign new_new_n27923__ = new_new_n27803__ & ~new_new_n27922__;
  assign new_new_n27924__ = ~new_new_n27803__ & new_new_n27922__;
  assign new_new_n27925__ = ~new_new_n27634__ & ~new_new_n27651__;
  assign new_new_n27926__ = new_new_n27650__ & new_new_n27925__;
  assign new_new_n27927__ = ~new_new_n27650__ & ~new_new_n27925__;
  assign new_new_n27928__ = ~new_new_n27926__ & ~new_new_n27927__;
  assign new_new_n27929__ = ~new_new_n27924__ & new_new_n27928__;
  assign new_new_n27930__ = ~new_new_n27923__ & ~new_new_n27929__;
  assign new_new_n27931__ = ~new_new_n27771__ & ~new_new_n27930__;
  assign new_new_n27932__ = new_new_n27771__ & new_new_n27930__;
  assign new_new_n27933__ = ~new_new_n27654__ & ~new_new_n27655__;
  assign new_new_n27934__ = ~new_new_n27677__ & ~new_new_n27933__;
  assign new_new_n27935__ = new_new_n27677__ & new_new_n27933__;
  assign new_new_n27936__ = ~new_new_n27934__ & ~new_new_n27935__;
  assign new_new_n27937__ = ~new_new_n27932__ & ~new_new_n27936__;
  assign new_new_n27938__ = ~new_new_n27931__ & ~new_new_n27937__;
  assign new_new_n27939__ = new_new_n6634__ & ~new_new_n27003__;
  assign new_new_n27940__ = ~new_new_n6625__ & ~new_new_n27021__;
  assign new_new_n27941__ = new_new_n6629__ & ~new_new_n27029__;
  assign new_new_n27942__ = new_new_n27021__ & new_new_n27029__;
  assign new_new_n27943__ = ~new_new_n27118__ & ~new_new_n27942__;
  assign new_new_n27944__ = new_new_n27003__ & ~new_new_n27943__;
  assign new_new_n27945__ = new_new_n27112__ & ~new_new_n27113__;
  assign new_new_n27946__ = new_new_n27021__ & new_new_n27113__;
  assign new_new_n27947__ = new_new_n27003__ & new_new_n27029__;
  assign new_new_n27948__ = ~new_new_n27105__ & new_new_n27947__;
  assign new_new_n27949__ = ~new_new_n27946__ & ~new_new_n27948__;
  assign new_new_n27950__ = ~new_new_n27111__ & ~new_new_n27949__;
  assign new_new_n27951__ = ~new_new_n27111__ & new_new_n27947__;
  assign new_new_n27952__ = ~new_new_n27105__ & new_new_n27946__;
  assign new_new_n27953__ = new_new_n27033__ & ~new_new_n27951__;
  assign new_new_n27954__ = ~new_new_n27952__ & new_new_n27953__;
  assign new_new_n27955__ = new_new_n27029__ & new_new_n27115__;
  assign new_new_n27956__ = new_new_n27003__ & new_new_n27114__;
  assign new_new_n27957__ = ~new_new_n27033__ & ~new_new_n27956__;
  assign new_new_n27958__ = ~new_new_n27955__ & new_new_n27957__;
  assign new_new_n27959__ = ~new_new_n27954__ & ~new_new_n27958__;
  assign new_new_n27960__ = ~new_new_n27944__ & ~new_new_n27945__;
  assign new_new_n27961__ = ~new_new_n27950__ & new_new_n27960__;
  assign new_new_n27962__ = ~new_new_n27959__ & new_new_n27961__;
  assign new_new_n27963__ = new_new_n6936__ & new_new_n27962__;
  assign new_new_n27964__ = ~new_new_n27940__ & ~new_new_n27941__;
  assign new_new_n27965__ = ~new_new_n27939__ & new_new_n27964__;
  assign new_new_n27966__ = ~new_new_n27963__ & new_new_n27965__;
  assign new_new_n27967__ = pi20 & ~new_new_n27966__;
  assign new_new_n27968__ = ~pi20 & new_new_n27966__;
  assign new_new_n27969__ = ~new_new_n27967__ & ~new_new_n27968__;
  assign new_new_n27970__ = new_new_n27938__ & new_new_n27969__;
  assign new_new_n27971__ = ~new_new_n27938__ & ~new_new_n27969__;
  assign new_new_n27972__ = ~new_new_n27970__ & ~new_new_n27971__;
  assign new_new_n27973__ = ~new_new_n27735__ & ~new_new_n27972__;
  assign new_new_n27974__ = new_new_n27735__ & new_new_n27972__;
  assign new_new_n27975__ = ~new_new_n27973__ & ~new_new_n27974__;
  assign new_new_n27976__ = new_new_n6968__ & new_new_n26971__;
  assign new_new_n27977__ = new_new_n6964__ & ~new_new_n26978__;
  assign new_new_n27978__ = new_new_n7935__ & ~new_new_n26937__;
  assign new_new_n27979__ = ~new_new_n27976__ & ~new_new_n27977__;
  assign new_new_n27980__ = ~new_new_n27978__ & new_new_n27979__;
  assign new_new_n27981__ = new_new_n26978__ & new_new_n27003__;
  assign new_new_n27982__ = ~new_new_n26978__ & ~new_new_n27003__;
  assign new_new_n27983__ = ~new_new_n27981__ & ~new_new_n27982__;
  assign new_new_n27984__ = ~new_new_n27121__ & new_new_n27983__;
  assign new_new_n27985__ = new_new_n27121__ & ~new_new_n27983__;
  assign new_new_n27986__ = ~new_new_n27984__ & ~new_new_n27985__;
  assign new_new_n27987__ = ~new_new_n27003__ & new_new_n27125__;
  assign new_new_n27988__ = ~new_new_n26971__ & ~new_new_n26978__;
  assign new_new_n27989__ = ~new_new_n26937__ & new_new_n27988__;
  assign new_new_n27990__ = ~new_new_n27987__ & ~new_new_n27989__;
  assign new_new_n27991__ = ~new_new_n27986__ & ~new_new_n27990__;
  assign new_new_n27992__ = ~new_new_n26978__ & new_new_n27986__;
  assign new_new_n27993__ = ~new_new_n26971__ & ~new_new_n27992__;
  assign new_new_n27994__ = new_new_n27121__ & ~new_new_n27993__;
  assign new_new_n27995__ = ~new_new_n26979__ & ~new_new_n27125__;
  assign new_new_n27996__ = new_new_n26978__ & ~new_new_n27986__;
  assign new_new_n27997__ = new_new_n26971__ & ~new_new_n27996__;
  assign new_new_n27998__ = ~new_new_n27994__ & ~new_new_n27997__;
  assign new_new_n27999__ = new_new_n27995__ & new_new_n27998__;
  assign new_new_n28000__ = ~new_new_n26971__ & new_new_n26978__;
  assign new_new_n28001__ = ~new_new_n26971__ & ~new_new_n27003__;
  assign new_new_n28002__ = ~new_new_n28000__ & ~new_new_n28001__;
  assign new_new_n28003__ = ~new_new_n27995__ & new_new_n28002__;
  assign new_new_n28004__ = ~new_new_n27999__ & ~new_new_n28003__;
  assign new_new_n28005__ = ~new_new_n27991__ & ~new_new_n28004__;
  assign new_new_n28006__ = new_new_n6958__ & new_new_n28005__;
  assign new_new_n28007__ = ~pi17 & ~new_new_n28006__;
  assign new_new_n28008__ = new_new_n8160__ & new_new_n28005__;
  assign new_new_n28009__ = ~new_new_n28007__ & ~new_new_n28008__;
  assign new_new_n28010__ = new_new_n27980__ & ~new_new_n28009__;
  assign new_new_n28011__ = pi17 & ~new_new_n27980__;
  assign new_new_n28012__ = ~new_new_n28010__ & ~new_new_n28011__;
  assign new_new_n28013__ = ~new_new_n27975__ & ~new_new_n28012__;
  assign new_new_n28014__ = new_new_n27975__ & new_new_n28012__;
  assign new_new_n28015__ = ~new_new_n27923__ & ~new_new_n27924__;
  assign new_new_n28016__ = ~new_new_n27928__ & new_new_n28015__;
  assign new_new_n28017__ = new_new_n27928__ & ~new_new_n28015__;
  assign new_new_n28018__ = ~new_new_n28016__ & ~new_new_n28017__;
  assign new_new_n28019__ = new_new_n7935__ & ~new_new_n27003__;
  assign new_new_n28020__ = new_new_n6968__ & ~new_new_n27029__;
  assign new_new_n28021__ = new_new_n6964__ & ~new_new_n27021__;
  assign new_new_n28022__ = new_new_n6959__ & new_new_n27962__;
  assign new_new_n28023__ = ~new_new_n28020__ & ~new_new_n28021__;
  assign new_new_n28024__ = ~new_new_n28019__ & new_new_n28023__;
  assign new_new_n28025__ = ~new_new_n28022__ & new_new_n28024__;
  assign new_new_n28026__ = pi17 & ~new_new_n28025__;
  assign new_new_n28027__ = ~pi17 & new_new_n28025__;
  assign new_new_n28028__ = ~new_new_n28026__ & ~new_new_n28027__;
  assign new_new_n28029__ = ~new_new_n27815__ & new_new_n27895__;
  assign new_new_n28030__ = ~new_new_n27899__ & ~new_new_n28029__;
  assign new_new_n28031__ = ~new_new_n27575__ & ~new_new_n27607__;
  assign new_new_n28032__ = ~new_new_n27608__ & ~new_new_n28031__;
  assign new_new_n28033__ = ~new_new_n27815__ & new_new_n27818__;
  assign new_new_n28034__ = ~new_new_n28032__ & ~new_new_n28033__;
  assign new_new_n28035__ = new_new_n28030__ & ~new_new_n28034__;
  assign new_new_n28036__ = ~new_new_n27818__ & ~new_new_n28032__;
  assign new_new_n28037__ = ~new_new_n28030__ & new_new_n28036__;
  assign new_new_n28038__ = ~new_new_n28035__ & ~new_new_n28037__;
  assign new_new_n28039__ = new_new_n6964__ & new_new_n27041__;
  assign new_new_n28040__ = new_new_n6968__ & ~new_new_n27054__;
  assign new_new_n28041__ = ~new_new_n28039__ & ~new_new_n28040__;
  assign new_new_n28042__ = new_new_n6958__ & ~new_new_n27535__;
  assign new_new_n28043__ = pi17 & ~new_new_n28042__;
  assign new_new_n28044__ = ~pi16 & new_new_n27033__;
  assign new_new_n28045__ = pi16 & ~new_new_n27033__;
  assign new_new_n28046__ = new_new_n6958__ & ~new_new_n28044__;
  assign new_new_n28047__ = ~new_new_n28045__ & new_new_n28046__;
  assign new_new_n28048__ = ~new_new_n27102__ & new_new_n28047__;
  assign new_new_n28049__ = ~new_new_n28043__ & ~new_new_n28048__;
  assign new_new_n28050__ = new_new_n28041__ & ~new_new_n28049__;
  assign new_new_n28051__ = new_new_n6958__ & new_new_n27545__;
  assign new_new_n28052__ = new_new_n28041__ & ~new_new_n28051__;
  assign new_new_n28053__ = ~pi17 & ~new_new_n28052__;
  assign new_new_n28054__ = ~new_new_n28050__ & ~new_new_n28053__;
  assign new_new_n28055__ = new_new_n6631__ & ~new_new_n27577__;
  assign new_new_n28056__ = new_new_n27853__ & new_new_n28055__;
  assign new_new_n28057__ = new_new_n6629__ & ~new_new_n27075__;
  assign new_new_n28058__ = ~new_new_n26118__ & new_new_n28057__;
  assign new_new_n28059__ = ~new_new_n28056__ & ~new_new_n28058__;
  assign new_new_n28060__ = pi20 & ~new_new_n28059__;
  assign new_new_n28061__ = pi20 & new_new_n28055__;
  assign new_new_n28062__ = ~new_new_n27853__ & ~new_new_n28061__;
  assign new_new_n28063__ = pi20 & ~new_new_n27075__;
  assign new_new_n28064__ = new_new_n6629__ & ~new_new_n28063__;
  assign new_new_n28065__ = new_new_n26118__ & new_new_n28064__;
  assign new_new_n28066__ = ~new_new_n28062__ & ~new_new_n28065__;
  assign new_new_n28067__ = ~new_new_n28060__ & new_new_n28066__;
  assign new_new_n28068__ = new_new_n7935__ & ~new_new_n27054__;
  assign new_new_n28069__ = new_new_n6964__ & ~new_new_n27071__;
  assign new_new_n28070__ = new_new_n6968__ & new_new_n27041__;
  assign new_new_n28071__ = ~new_new_n28069__ & ~new_new_n28070__;
  assign new_new_n28072__ = ~new_new_n28068__ & new_new_n28071__;
  assign new_new_n28073__ = new_new_n6958__ & ~new_new_n27094__;
  assign new_new_n28074__ = ~pi17 & ~new_new_n28073__;
  assign new_new_n28075__ = new_new_n8160__ & ~new_new_n27094__;
  assign new_new_n28076__ = ~new_new_n28074__ & ~new_new_n28075__;
  assign new_new_n28077__ = new_new_n28072__ & ~new_new_n28076__;
  assign new_new_n28078__ = pi17 & ~new_new_n28072__;
  assign new_new_n28079__ = ~new_new_n28077__ & ~new_new_n28078__;
  assign new_new_n28080__ = new_new_n28067__ & ~new_new_n28079__;
  assign new_new_n28081__ = new_new_n6968__ & ~new_new_n27071__;
  assign new_new_n28082__ = new_new_n6964__ & new_new_n27059__;
  assign new_new_n28083__ = ~new_new_n28081__ & ~new_new_n28082__;
  assign new_new_n28084__ = new_new_n6958__ & new_new_n27041__;
  assign new_new_n28085__ = new_new_n27567__ & new_new_n28084__;
  assign new_new_n28086__ = new_new_n28083__ & ~new_new_n28085__;
  assign new_new_n28087__ = pi17 & ~new_new_n28086__;
  assign new_new_n28088__ = ~new_new_n27041__ & ~new_new_n27567__;
  assign new_new_n28089__ = new_new_n6958__ & ~new_new_n28088__;
  assign new_new_n28090__ = ~pi17 & ~new_new_n28089__;
  assign new_new_n28091__ = ~new_new_n27041__ & new_new_n27567__;
  assign new_new_n28092__ = ~pi16 & ~new_new_n28091__;
  assign new_new_n28093__ = new_new_n27041__ & ~new_new_n27566__;
  assign new_new_n28094__ = pi16 & ~new_new_n28093__;
  assign new_new_n28095__ = new_new_n6958__ & ~new_new_n28094__;
  assign new_new_n28096__ = ~new_new_n28092__ & new_new_n28095__;
  assign new_new_n28097__ = ~new_new_n28090__ & ~new_new_n28096__;
  assign new_new_n28098__ = new_new_n28083__ & ~new_new_n28097__;
  assign new_new_n28099__ = ~new_new_n28087__ & ~new_new_n28098__;
  assign new_new_n28100__ = new_new_n6631__ & new_new_n26118__;
  assign new_new_n28101__ = ~new_new_n28099__ & new_new_n28100__;
  assign new_new_n28102__ = new_new_n28099__ & ~new_new_n28100__;
  assign new_new_n28103__ = ~new_new_n28101__ & ~new_new_n28102__;
  assign new_new_n28104__ = new_new_n27075__ & ~new_new_n28103__;
  assign new_new_n28105__ = ~new_new_n6622__ & new_new_n26118__;
  assign new_new_n28106__ = ~new_new_n6619__ & ~new_new_n28105__;
  assign new_new_n28107__ = pi19 & new_new_n28099__;
  assign new_new_n28108__ = ~pi19 & ~new_new_n28099__;
  assign new_new_n28109__ = new_new_n28106__ & ~new_new_n28107__;
  assign new_new_n28110__ = ~new_new_n28108__ & new_new_n28109__;
  assign new_new_n28111__ = ~new_new_n9920__ & ~new_new_n28110__;
  assign new_new_n28112__ = new_new_n28099__ & ~new_new_n28111__;
  assign new_new_n28113__ = new_new_n28105__ & new_new_n28107__;
  assign new_new_n28114__ = ~new_new_n28106__ & new_new_n28108__;
  assign new_new_n28115__ = ~new_new_n28113__ & ~new_new_n28114__;
  assign new_new_n28116__ = ~new_new_n28110__ & new_new_n28115__;
  assign new_new_n28117__ = ~new_new_n27075__ & ~new_new_n28116__;
  assign new_new_n28118__ = ~new_new_n28104__ & ~new_new_n28112__;
  assign new_new_n28119__ = ~new_new_n28117__ & new_new_n28118__;
  assign new_new_n28120__ = new_new_n28099__ & new_new_n28119__;
  assign new_new_n28121__ = new_new_n6631__ & ~new_new_n27075__;
  assign new_new_n28122__ = new_new_n6958__ & new_new_n26118__;
  assign new_new_n28123__ = new_new_n27075__ & ~new_new_n28122__;
  assign new_new_n28124__ = new_new_n6963__ & ~new_new_n28123__;
  assign new_new_n28125__ = new_new_n6964__ & ~new_new_n27075__;
  assign new_new_n28126__ = new_new_n6968__ & new_new_n26118__;
  assign new_new_n28127__ = new_new_n6955__ & new_new_n27582__;
  assign new_new_n28128__ = ~new_new_n27059__ & ~new_new_n28127__;
  assign new_new_n28129__ = new_new_n27059__ & new_new_n28127__;
  assign new_new_n28130__ = new_new_n6958__ & ~new_new_n28128__;
  assign new_new_n28131__ = ~new_new_n28129__ & new_new_n28130__;
  assign new_new_n28132__ = ~new_new_n28125__ & ~new_new_n28126__;
  assign new_new_n28133__ = ~new_new_n28131__ & new_new_n28132__;
  assign new_new_n28134__ = pi17 & ~new_new_n28124__;
  assign new_new_n28135__ = new_new_n28133__ & new_new_n28134__;
  assign new_new_n28136__ = ~new_new_n28121__ & ~new_new_n28135__;
  assign new_new_n28137__ = new_new_n7935__ & ~new_new_n27071__;
  assign new_new_n28138__ = new_new_n6968__ & new_new_n27059__;
  assign new_new_n28139__ = new_new_n6959__ & new_new_n27600__;
  assign new_new_n28140__ = ~new_new_n28137__ & ~new_new_n28138__;
  assign new_new_n28141__ = ~new_new_n28139__ & new_new_n28140__;
  assign new_new_n28142__ = new_new_n10337__ & new_new_n26118__;
  assign new_new_n28143__ = pi17 & ~new_new_n28142__;
  assign new_new_n28144__ = new_new_n10340__ & new_new_n26118__;
  assign new_new_n28145__ = ~pi17 & ~new_new_n28144__;
  assign new_new_n28146__ = pi14 & ~new_new_n28145__;
  assign new_new_n28147__ = ~new_new_n28143__ & ~new_new_n28146__;
  assign new_new_n28148__ = new_new_n28141__ & ~new_new_n28147__;
  assign new_new_n28149__ = ~pi17 & ~new_new_n28141__;
  assign new_new_n28150__ = ~new_new_n28148__ & ~new_new_n28149__;
  assign new_new_n28151__ = ~new_new_n28136__ & ~new_new_n28150__;
  assign new_new_n28152__ = ~new_new_n28119__ & new_new_n28151__;
  assign new_new_n28153__ = ~new_new_n28120__ & ~new_new_n28152__;
  assign new_new_n28154__ = ~new_new_n28067__ & new_new_n28079__;
  assign new_new_n28155__ = ~new_new_n28080__ & ~new_new_n28154__;
  assign new_new_n28156__ = new_new_n28153__ & new_new_n28155__;
  assign new_new_n28157__ = ~new_new_n28080__ & ~new_new_n28156__;
  assign new_new_n28158__ = new_new_n28054__ & ~new_new_n28157__;
  assign new_new_n28159__ = ~new_new_n28054__ & new_new_n28157__;
  assign new_new_n28160__ = pi20 & new_new_n27856__;
  assign new_new_n28161__ = pi20 & ~new_new_n27854__;
  assign new_new_n28162__ = new_new_n5195__ & ~new_new_n27075__;
  assign new_new_n28163__ = ~new_new_n28161__ & new_new_n28162__;
  assign new_new_n28164__ = ~new_new_n28160__ & ~new_new_n28163__;
  assign new_new_n28165__ = new_new_n27864__ & new_new_n28164__;
  assign new_new_n28166__ = ~pi20 & new_new_n27075__;
  assign new_new_n28167__ = new_new_n27856__ & ~new_new_n28166__;
  assign new_new_n28168__ = ~new_new_n27864__ & new_new_n28167__;
  assign new_new_n28169__ = ~new_new_n28165__ & ~new_new_n28168__;
  assign new_new_n28170__ = ~new_new_n28159__ & ~new_new_n28169__;
  assign new_new_n28171__ = ~new_new_n28158__ & ~new_new_n28170__;
  assign new_new_n28172__ = new_new_n6968__ & ~new_new_n27033__;
  assign new_new_n28173__ = new_new_n6964__ & ~new_new_n27054__;
  assign new_new_n28174__ = new_new_n6955__ & new_new_n27686__;
  assign new_new_n28175__ = ~new_new_n27111__ & ~new_new_n28174__;
  assign new_new_n28176__ = new_new_n27111__ & new_new_n28174__;
  assign new_new_n28177__ = new_new_n6958__ & ~new_new_n28175__;
  assign new_new_n28178__ = ~new_new_n28176__ & new_new_n28177__;
  assign new_new_n28179__ = ~new_new_n28172__ & ~new_new_n28173__;
  assign new_new_n28180__ = ~new_new_n28178__ & new_new_n28179__;
  assign new_new_n28181__ = pi17 & ~new_new_n28180__;
  assign new_new_n28182__ = ~pi17 & new_new_n28180__;
  assign new_new_n28183__ = ~new_new_n28181__ & ~new_new_n28182__;
  assign new_new_n28184__ = ~new_new_n28171__ & ~new_new_n28183__;
  assign new_new_n28185__ = new_new_n28171__ & new_new_n28183__;
  assign new_new_n28186__ = ~new_new_n27871__ & ~new_new_n27872__;
  assign new_new_n28187__ = new_new_n27880__ & ~new_new_n28186__;
  assign new_new_n28188__ = ~new_new_n27880__ & new_new_n28186__;
  assign new_new_n28189__ = ~new_new_n28187__ & ~new_new_n28188__;
  assign new_new_n28190__ = ~new_new_n28185__ & new_new_n28189__;
  assign new_new_n28191__ = ~new_new_n28184__ & ~new_new_n28190__;
  assign new_new_n28192__ = new_new_n27891__ & ~new_new_n28191__;
  assign new_new_n28193__ = ~new_new_n27891__ & new_new_n28191__;
  assign new_new_n28194__ = new_new_n7935__ & ~new_new_n27021__;
  assign new_new_n28195__ = new_new_n6968__ & new_new_n27111__;
  assign new_new_n28196__ = new_new_n6964__ & ~new_new_n27033__;
  assign new_new_n28197__ = new_new_n6959__ & new_new_n27796__;
  assign new_new_n28198__ = ~new_new_n28195__ & ~new_new_n28196__;
  assign new_new_n28199__ = ~new_new_n28194__ & new_new_n28198__;
  assign new_new_n28200__ = ~new_new_n28197__ & new_new_n28199__;
  assign new_new_n28201__ = ~new_new_n28192__ & ~new_new_n28193__;
  assign new_new_n28202__ = pi17 & ~new_new_n28201__;
  assign new_new_n28203__ = ~pi17 & new_new_n28201__;
  assign new_new_n28204__ = ~new_new_n28202__ & ~new_new_n28203__;
  assign new_new_n28205__ = new_new_n28200__ & new_new_n28204__;
  assign new_new_n28206__ = ~new_new_n28200__ & ~new_new_n28204__;
  assign new_new_n28207__ = ~new_new_n28205__ & ~new_new_n28206__;
  assign new_new_n28208__ = ~new_new_n28193__ & new_new_n28207__;
  assign new_new_n28209__ = ~new_new_n28192__ & ~new_new_n28208__;
  assign new_new_n28210__ = new_new_n28038__ & new_new_n28209__;
  assign new_new_n28211__ = ~new_new_n28038__ & ~new_new_n28209__;
  assign new_new_n28212__ = new_new_n7935__ & ~new_new_n27029__;
  assign new_new_n28213__ = new_new_n6968__ & ~new_new_n27021__;
  assign new_new_n28214__ = new_new_n6964__ & new_new_n27111__;
  assign new_new_n28215__ = new_new_n6959__ & new_new_n27764__;
  assign new_new_n28216__ = ~new_new_n28213__ & ~new_new_n28214__;
  assign new_new_n28217__ = ~new_new_n28212__ & new_new_n28216__;
  assign new_new_n28218__ = ~new_new_n28215__ & new_new_n28217__;
  assign new_new_n28219__ = pi17 & ~new_new_n28218__;
  assign new_new_n28220__ = ~pi17 & new_new_n28218__;
  assign new_new_n28221__ = ~new_new_n28219__ & ~new_new_n28220__;
  assign new_new_n28222__ = ~new_new_n28211__ & new_new_n28221__;
  assign new_new_n28223__ = ~new_new_n28210__ & ~new_new_n28222__;
  assign new_new_n28224__ = new_new_n28028__ & ~new_new_n28223__;
  assign new_new_n28225__ = ~new_new_n28028__ & new_new_n28223__;
  assign new_new_n28226__ = ~new_new_n27907__ & ~new_new_n27908__;
  assign new_new_n28227__ = ~new_new_n27920__ & new_new_n28226__;
  assign new_new_n28228__ = new_new_n27920__ & ~new_new_n28226__;
  assign new_new_n28229__ = ~new_new_n28227__ & ~new_new_n28228__;
  assign new_new_n28230__ = ~new_new_n28225__ & ~new_new_n28229__;
  assign new_new_n28231__ = ~new_new_n28224__ & ~new_new_n28230__;
  assign new_new_n28232__ = new_new_n28018__ & new_new_n28231__;
  assign new_new_n28233__ = ~new_new_n28018__ & ~new_new_n28231__;
  assign new_new_n28234__ = new_new_n6968__ & ~new_new_n27003__;
  assign new_new_n28235__ = new_new_n6964__ & ~new_new_n27029__;
  assign new_new_n28236__ = new_new_n7935__ & ~new_new_n26978__;
  assign new_new_n28237__ = ~new_new_n28234__ & ~new_new_n28235__;
  assign new_new_n28238__ = ~new_new_n28236__ & new_new_n28237__;
  assign new_new_n28239__ = new_new_n6958__ & new_new_n27986__;
  assign new_new_n28240__ = ~pi17 & ~new_new_n28239__;
  assign new_new_n28241__ = new_new_n8160__ & new_new_n27986__;
  assign new_new_n28242__ = ~new_new_n28240__ & ~new_new_n28241__;
  assign new_new_n28243__ = new_new_n28238__ & ~new_new_n28242__;
  assign new_new_n28244__ = pi17 & ~new_new_n28238__;
  assign new_new_n28245__ = ~new_new_n28243__ & ~new_new_n28244__;
  assign new_new_n28246__ = ~new_new_n28233__ & ~new_new_n28245__;
  assign new_new_n28247__ = ~new_new_n28232__ & ~new_new_n28246__;
  assign new_new_n28248__ = ~new_new_n27931__ & ~new_new_n27932__;
  assign new_new_n28249__ = ~new_new_n27936__ & new_new_n28248__;
  assign new_new_n28250__ = new_new_n27936__ & ~new_new_n28248__;
  assign new_new_n28251__ = ~new_new_n28249__ & ~new_new_n28250__;
  assign new_new_n28252__ = ~new_new_n28247__ & ~new_new_n28251__;
  assign new_new_n28253__ = new_new_n28247__ & new_new_n28251__;
  assign new_new_n28254__ = ~new_new_n27029__ & new_new_n27988__;
  assign new_new_n28255__ = new_new_n26971__ & ~new_new_n27003__;
  assign new_new_n28256__ = new_new_n26978__ & new_new_n28255__;
  assign new_new_n28257__ = ~new_new_n27764__ & new_new_n28256__;
  assign new_new_n28258__ = ~new_new_n28254__ & ~new_new_n28257__;
  assign new_new_n28259__ = ~new_new_n27021__ & ~new_new_n28258__;
  assign new_new_n28260__ = ~new_new_n26971__ & ~new_new_n27983__;
  assign new_new_n28261__ = ~new_new_n27764__ & new_new_n27988__;
  assign new_new_n28262__ = ~new_new_n28256__ & ~new_new_n28261__;
  assign new_new_n28263__ = ~new_new_n27029__ & ~new_new_n28262__;
  assign new_new_n28264__ = new_new_n27764__ & new_new_n28000__;
  assign new_new_n28265__ = new_new_n26971__ & ~new_new_n26978__;
  assign new_new_n28266__ = new_new_n27003__ & new_new_n28265__;
  assign new_new_n28267__ = ~new_new_n28264__ & ~new_new_n28266__;
  assign new_new_n28268__ = new_new_n27029__ & ~new_new_n28267__;
  assign new_new_n28269__ = new_new_n27029__ & new_new_n28000__;
  assign new_new_n28270__ = new_new_n27003__ & new_new_n27764__;
  assign new_new_n28271__ = new_new_n28265__ & new_new_n28270__;
  assign new_new_n28272__ = ~new_new_n28269__ & ~new_new_n28271__;
  assign new_new_n28273__ = new_new_n27021__ & ~new_new_n28272__;
  assign new_new_n28274__ = ~new_new_n28260__ & ~new_new_n28263__;
  assign new_new_n28275__ = ~new_new_n28268__ & ~new_new_n28273__;
  assign new_new_n28276__ = new_new_n28274__ & new_new_n28275__;
  assign new_new_n28277__ = ~new_new_n28259__ & new_new_n28276__;
  assign new_new_n28278__ = new_new_n6959__ & new_new_n28277__;
  assign new_new_n28279__ = new_new_n6964__ & ~new_new_n27003__;
  assign new_new_n28280__ = new_new_n6968__ & ~new_new_n26978__;
  assign new_new_n28281__ = ~new_new_n28279__ & ~new_new_n28280__;
  assign new_new_n28282__ = ~new_new_n28278__ & new_new_n28281__;
  assign new_new_n28283__ = new_new_n6958__ & new_new_n26971__;
  assign new_new_n28284__ = ~pi17 & ~new_new_n28283__;
  assign new_new_n28285__ = new_new_n7942__ & new_new_n26971__;
  assign new_new_n28286__ = ~new_new_n28284__ & ~new_new_n28285__;
  assign new_new_n28287__ = new_new_n28282__ & ~new_new_n28286__;
  assign new_new_n28288__ = pi17 & ~new_new_n28282__;
  assign new_new_n28289__ = ~new_new_n28287__ & ~new_new_n28288__;
  assign new_new_n28290__ = ~new_new_n28253__ & ~new_new_n28289__;
  assign new_new_n28291__ = ~new_new_n28252__ & ~new_new_n28290__;
  assign new_new_n28292__ = ~new_new_n28014__ & ~new_new_n28291__;
  assign new_new_n28293__ = ~new_new_n28013__ & ~new_new_n28292__;
  assign new_new_n28294__ = ~new_new_n27531__ & new_new_n28293__;
  assign new_new_n28295__ = new_new_n27531__ & ~new_new_n28293__;
  assign new_new_n28296__ = new_new_n27075__ & ~new_new_n27717__;
  assign new_new_n28297__ = ~pi28 & ~new_new_n27075__;
  assign new_new_n28298__ = new_new_n3889__ & ~new_new_n28297__;
  assign new_new_n28299__ = ~new_new_n68__ & ~new_new_n28298__;
  assign new_new_n28300__ = ~new_new_n28296__ & new_new_n28299__;
  assign new_new_n28301__ = pi29 & ~new_new_n28300__;
  assign new_new_n28302__ = new_new_n66__ & ~new_new_n27075__;
  assign new_new_n28303__ = new_new_n4221__ & ~new_new_n27075__;
  assign new_new_n28304__ = pi29 & ~new_new_n28303__;
  assign new_new_n28305__ = ~new_new_n28302__ & ~new_new_n28304__;
  assign new_new_n28306__ = ~pi28 & new_new_n3889__;
  assign new_new_n28307__ = ~pi26 & new_new_n77__;
  assign new_new_n28308__ = new_new_n4813__ & new_new_n27553__;
  assign new_new_n28309__ = ~new_new_n28306__ & ~new_new_n28307__;
  assign new_new_n28310__ = ~new_new_n28308__ & new_new_n28309__;
  assign new_new_n28311__ = new_new_n26118__ & ~new_new_n28310__;
  assign new_new_n28312__ = ~new_new_n4215__ & new_new_n27582__;
  assign new_new_n28313__ = new_new_n4214__ & ~new_new_n28312__;
  assign new_new_n28314__ = new_new_n27059__ & new_new_n28313__;
  assign new_new_n28315__ = ~new_new_n28311__ & ~new_new_n28314__;
  assign new_new_n28316__ = ~new_new_n28305__ & new_new_n28315__;
  assign new_new_n28317__ = ~pi29 & ~new_new_n28315__;
  assign new_new_n28318__ = ~new_new_n28316__ & ~new_new_n28317__;
  assign new_new_n28319__ = ~new_new_n28301__ & ~new_new_n28318__;
  assign new_new_n28320__ = new_new_n28301__ & ~new_new_n28316__;
  assign new_new_n28321__ = ~new_new_n28319__ & ~new_new_n28320__;
  assign new_new_n28322__ = new_new_n3311__ & ~new_new_n27054__;
  assign new_new_n28323__ = ~new_new_n333__ & ~new_new_n27071__;
  assign new_new_n28324__ = new_new_n873__ & new_new_n27041__;
  assign new_new_n28325__ = ~new_new_n28323__ & ~new_new_n28324__;
  assign new_new_n28326__ = ~new_new_n28322__ & new_new_n28325__;
  assign new_new_n28327__ = ~pi26 & ~new_new_n28326__;
  assign new_new_n28328__ = new_new_n512__ & ~new_new_n27094__;
  assign new_new_n28329__ = new_new_n801__ & ~new_new_n27094__;
  assign new_new_n28330__ = pi26 & ~new_new_n28329__;
  assign new_new_n28331__ = ~new_new_n28328__ & ~new_new_n28330__;
  assign new_new_n28332__ = new_new_n28326__ & ~new_new_n28331__;
  assign new_new_n28333__ = ~new_new_n28327__ & ~new_new_n28332__;
  assign new_new_n28334__ = ~new_new_n28319__ & new_new_n28333__;
  assign new_new_n28335__ = ~new_new_n28321__ & ~new_new_n28334__;
  assign new_new_n28336__ = new_new_n27674__ & ~new_new_n27722__;
  assign new_new_n28337__ = ~new_new_n27714__ & ~new_new_n28336__;
  assign new_new_n28338__ = new_new_n27672__ & new_new_n27722__;
  assign new_new_n28339__ = ~new_new_n28337__ & ~new_new_n28338__;
  assign new_new_n28340__ = new_new_n28333__ & new_new_n28339__;
  assign new_new_n28341__ = ~new_new_n28333__ & ~new_new_n28339__;
  assign new_new_n28342__ = ~new_new_n28340__ & ~new_new_n28341__;
  assign new_new_n28343__ = new_new_n28335__ & new_new_n28342__;
  assign new_new_n28344__ = new_new_n5213__ & ~new_new_n27021__;
  assign new_new_n28345__ = new_new_n5191__ & ~new_new_n27033__;
  assign new_new_n28346__ = new_new_n5183__ & new_new_n27111__;
  assign new_new_n28347__ = ~new_new_n28345__ & ~new_new_n28346__;
  assign new_new_n28348__ = ~new_new_n28344__ & new_new_n28347__;
  assign new_new_n28349__ = new_new_n5195__ & new_new_n27796__;
  assign new_new_n28350__ = pi23 & ~new_new_n28349__;
  assign new_new_n28351__ = new_new_n7878__ & new_new_n27796__;
  assign new_new_n28352__ = ~new_new_n28350__ & ~new_new_n28351__;
  assign new_new_n28353__ = new_new_n28348__ & ~new_new_n28352__;
  assign new_new_n28354__ = ~pi23 & ~new_new_n28348__;
  assign new_new_n28355__ = ~new_new_n28353__ & ~new_new_n28354__;
  assign new_new_n28356__ = ~new_new_n27679__ & ~new_new_n27731__;
  assign new_new_n28357__ = ~new_new_n27730__ & ~new_new_n28356__;
  assign new_new_n28358__ = ~new_new_n28355__ & new_new_n28357__;
  assign new_new_n28359__ = new_new_n28355__ & ~new_new_n28357__;
  assign new_new_n28360__ = ~new_new_n28358__ & ~new_new_n28359__;
  assign new_new_n28361__ = new_new_n28321__ & ~new_new_n28342__;
  assign new_new_n28362__ = ~new_new_n28343__ & ~new_new_n28361__;
  assign new_new_n28363__ = ~new_new_n28360__ & new_new_n28362__;
  assign new_new_n28364__ = ~new_new_n28318__ & new_new_n28339__;
  assign new_new_n28365__ = new_new_n28301__ & ~new_new_n28364__;
  assign new_new_n28366__ = new_new_n28318__ & ~new_new_n28339__;
  assign new_new_n28367__ = ~new_new_n28364__ & ~new_new_n28366__;
  assign new_new_n28368__ = ~new_new_n28301__ & ~new_new_n28367__;
  assign new_new_n28369__ = ~new_new_n28365__ & ~new_new_n28368__;
  assign new_new_n28370__ = ~new_new_n28333__ & new_new_n28369__;
  assign new_new_n28371__ = new_new_n28320__ & ~new_new_n28339__;
  assign new_new_n28372__ = ~new_new_n28357__ & new_new_n28371__;
  assign new_new_n28373__ = new_new_n28301__ & new_new_n28316__;
  assign new_new_n28374__ = ~new_new_n28367__ & ~new_new_n28373__;
  assign new_new_n28375__ = ~new_new_n28365__ & ~new_new_n28374__;
  assign new_new_n28376__ = new_new_n28333__ & ~new_new_n28375__;
  assign new_new_n28377__ = ~new_new_n28370__ & ~new_new_n28376__;
  assign new_new_n28378__ = ~new_new_n28372__ & new_new_n28377__;
  assign new_new_n28379__ = new_new_n28360__ & new_new_n28378__;
  assign new_new_n28380__ = ~new_new_n28363__ & ~new_new_n28379__;
  assign new_new_n28381__ = ~new_new_n27938__ & new_new_n27969__;
  assign new_new_n28382__ = ~new_new_n27973__ & ~new_new_n28381__;
  assign new_new_n28383__ = new_new_n6629__ & ~new_new_n27003__;
  assign new_new_n28384__ = ~new_new_n6625__ & ~new_new_n27029__;
  assign new_new_n28385__ = new_new_n6634__ & ~new_new_n26978__;
  assign new_new_n28386__ = ~new_new_n28383__ & ~new_new_n28384__;
  assign new_new_n28387__ = ~new_new_n28385__ & new_new_n28386__;
  assign new_new_n28388__ = new_new_n6631__ & new_new_n27986__;
  assign new_new_n28389__ = pi20 & ~new_new_n28388__;
  assign new_new_n28390__ = new_new_n6640__ & new_new_n27986__;
  assign new_new_n28391__ = ~new_new_n28389__ & ~new_new_n28390__;
  assign new_new_n28392__ = new_new_n28387__ & ~new_new_n28391__;
  assign new_new_n28393__ = ~pi20 & ~new_new_n28387__;
  assign new_new_n28394__ = ~new_new_n28392__ & ~new_new_n28393__;
  assign new_new_n28395__ = new_new_n28382__ & new_new_n28394__;
  assign new_new_n28396__ = ~new_new_n28382__ & ~new_new_n28394__;
  assign new_new_n28397__ = ~new_new_n28395__ & ~new_new_n28396__;
  assign new_new_n28398__ = ~new_new_n28380__ & new_new_n28397__;
  assign new_new_n28399__ = new_new_n28380__ & ~new_new_n28397__;
  assign new_new_n28400__ = ~new_new_n28398__ & ~new_new_n28399__;
  assign new_new_n28401__ = ~new_new_n28295__ & new_new_n28400__;
  assign new_new_n28402__ = ~new_new_n28294__ & ~new_new_n28401__;
  assign new_new_n28403__ = ~new_new_n27509__ & ~new_new_n28402__;
  assign new_new_n28404__ = new_new_n27509__ & new_new_n28402__;
  assign new_new_n28405__ = new_new_n6634__ & new_new_n26971__;
  assign new_new_n28406__ = new_new_n6629__ & ~new_new_n26978__;
  assign new_new_n28407__ = ~new_new_n6625__ & ~new_new_n27003__;
  assign new_new_n28408__ = new_new_n6936__ & new_new_n28277__;
  assign new_new_n28409__ = ~new_new_n28406__ & ~new_new_n28407__;
  assign new_new_n28410__ = ~new_new_n28405__ & new_new_n28409__;
  assign new_new_n28411__ = ~new_new_n28408__ & new_new_n28410__;
  assign new_new_n28412__ = pi20 & ~new_new_n28411__;
  assign new_new_n28413__ = ~pi20 & new_new_n28411__;
  assign new_new_n28414__ = ~new_new_n28412__ & ~new_new_n28413__;
  assign new_new_n28415__ = new_new_n5213__ & ~new_new_n27029__;
  assign new_new_n28416__ = new_new_n5183__ & ~new_new_n27021__;
  assign new_new_n28417__ = new_new_n5191__ & new_new_n27111__;
  assign new_new_n28418__ = new_new_n5215__ & new_new_n27764__;
  assign new_new_n28419__ = ~new_new_n28416__ & ~new_new_n28417__;
  assign new_new_n28420__ = ~new_new_n28415__ & new_new_n28419__;
  assign new_new_n28421__ = ~new_new_n28418__ & new_new_n28420__;
  assign new_new_n28422__ = ~new_new_n333__ & new_new_n27041__;
  assign new_new_n28423__ = new_new_n873__ & ~new_new_n27054__;
  assign new_new_n28424__ = ~new_new_n28422__ & ~new_new_n28423__;
  assign new_new_n28425__ = new_new_n801__ & new_new_n27545__;
  assign new_new_n28426__ = new_new_n28424__ & ~new_new_n28425__;
  assign new_new_n28427__ = pi26 & ~new_new_n28426__;
  assign new_new_n28428__ = new_new_n801__ & ~new_new_n27535__;
  assign new_new_n28429__ = ~pi26 & ~new_new_n28428__;
  assign new_new_n28430__ = ~pi25 & ~new_new_n27033__;
  assign new_new_n28431__ = pi25 & new_new_n27033__;
  assign new_new_n28432__ = ~new_new_n110__ & ~new_new_n28430__;
  assign new_new_n28433__ = ~new_new_n28431__ & new_new_n28432__;
  assign new_new_n28434__ = ~new_new_n27102__ & new_new_n28433__;
  assign new_new_n28435__ = ~new_new_n28429__ & ~new_new_n28434__;
  assign new_new_n28436__ = new_new_n28424__ & ~new_new_n28435__;
  assign new_new_n28437__ = ~new_new_n28427__ & ~new_new_n28436__;
  assign new_new_n28438__ = ~pi30 & ~new_new_n27075__;
  assign new_new_n28439__ = new_new_n28373__ & new_new_n28438__;
  assign new_new_n28440__ = new_new_n4815__ & ~new_new_n27071__;
  assign new_new_n28441__ = ~new_new_n27084__ & ~new_new_n27088__;
  assign new_new_n28442__ = ~new_new_n27071__ & ~new_new_n28441__;
  assign new_new_n28443__ = new_new_n27071__ & new_new_n28441__;
  assign new_new_n28444__ = ~new_new_n4215__ & new_new_n28443__;
  assign new_new_n28445__ = ~new_new_n28442__ & ~new_new_n28444__;
  assign new_new_n28446__ = new_new_n4214__ & ~new_new_n28445__;
  assign new_new_n28447__ = new_new_n4212__ & new_new_n27059__;
  assign new_new_n28448__ = ~new_new_n28440__ & ~new_new_n28447__;
  assign new_new_n28449__ = ~new_new_n28446__ & new_new_n28448__;
  assign new_new_n28450__ = ~pi29 & ~new_new_n28449__;
  assign new_new_n28451__ = new_new_n4221__ & new_new_n26118__;
  assign new_new_n28452__ = pi29 & ~new_new_n28451__;
  assign new_new_n28453__ = new_new_n66__ & new_new_n26118__;
  assign new_new_n28454__ = ~new_new_n28452__ & ~new_new_n28453__;
  assign new_new_n28455__ = new_new_n28449__ & ~new_new_n28454__;
  assign new_new_n28456__ = ~new_new_n28450__ & ~new_new_n28455__;
  assign new_new_n28457__ = new_new_n765__ & ~new_new_n27075__;
  assign new_new_n28458__ = ~new_new_n28373__ & ~new_new_n28457__;
  assign new_new_n28459__ = ~new_new_n28456__ & ~new_new_n28458__;
  assign new_new_n28460__ = new_new_n28456__ & new_new_n28458__;
  assign new_new_n28461__ = ~new_new_n28459__ & ~new_new_n28460__;
  assign new_new_n28462__ = ~new_new_n28439__ & ~new_new_n28461__;
  assign new_new_n28463__ = new_new_n28437__ & ~new_new_n28462__;
  assign new_new_n28464__ = ~new_new_n28437__ & new_new_n28462__;
  assign new_new_n28465__ = ~new_new_n28463__ & ~new_new_n28464__;
  assign new_new_n28466__ = new_new_n28335__ & ~new_new_n28340__;
  assign new_new_n28467__ = ~new_new_n28341__ & ~new_new_n28466__;
  assign new_new_n28468__ = ~new_new_n28465__ & new_new_n28467__;
  assign new_new_n28469__ = new_new_n28301__ & ~new_new_n28333__;
  assign new_new_n28470__ = new_new_n28318__ & ~new_new_n28469__;
  assign new_new_n28471__ = ~new_new_n28341__ & new_new_n28470__;
  assign new_new_n28472__ = ~new_new_n28340__ & ~new_new_n28471__;
  assign new_new_n28473__ = new_new_n28465__ & new_new_n28472__;
  assign new_new_n28474__ = ~new_new_n28468__ & ~new_new_n28473__;
  assign new_new_n28475__ = new_new_n28333__ & new_new_n28437__;
  assign new_new_n28476__ = ~new_new_n28318__ & ~new_new_n28437__;
  assign new_new_n28477__ = ~new_new_n28364__ & ~new_new_n28475__;
  assign new_new_n28478__ = ~new_new_n28476__ & new_new_n28477__;
  assign new_new_n28479__ = new_new_n28301__ & new_new_n28465__;
  assign new_new_n28480__ = ~new_new_n28478__ & new_new_n28479__;
  assign new_new_n28481__ = ~new_new_n28474__ & ~new_new_n28480__;
  assign new_new_n28482__ = new_new_n28333__ & new_new_n28369__;
  assign new_new_n28483__ = ~new_new_n28358__ & new_new_n28482__;
  assign new_new_n28484__ = new_new_n28355__ & ~new_new_n28375__;
  assign new_new_n28485__ = ~new_new_n28317__ & new_new_n28371__;
  assign new_new_n28486__ = ~new_new_n28369__ & ~new_new_n28485__;
  assign new_new_n28487__ = ~new_new_n28357__ & new_new_n28486__;
  assign new_new_n28488__ = ~new_new_n28484__ & ~new_new_n28487__;
  assign new_new_n28489__ = ~new_new_n28333__ & ~new_new_n28488__;
  assign new_new_n28490__ = ~new_new_n28359__ & ~new_new_n28483__;
  assign new_new_n28491__ = ~new_new_n28489__ & new_new_n28490__;
  assign new_new_n28492__ = ~new_new_n28481__ & new_new_n28491__;
  assign new_new_n28493__ = new_new_n28481__ & ~new_new_n28491__;
  assign new_new_n28494__ = ~new_new_n28492__ & ~new_new_n28493__;
  assign new_new_n28495__ = pi23 & ~new_new_n28494__;
  assign new_new_n28496__ = ~pi23 & new_new_n28494__;
  assign new_new_n28497__ = ~new_new_n28495__ & ~new_new_n28496__;
  assign new_new_n28498__ = new_new_n28421__ & new_new_n28497__;
  assign new_new_n28499__ = ~new_new_n28421__ & ~new_new_n28497__;
  assign new_new_n28500__ = ~new_new_n28498__ & ~new_new_n28499__;
  assign new_new_n28501__ = new_new_n28380__ & ~new_new_n28396__;
  assign new_new_n28502__ = ~new_new_n28395__ & ~new_new_n28501__;
  assign new_new_n28503__ = new_new_n28500__ & new_new_n28502__;
  assign new_new_n28504__ = ~new_new_n28500__ & ~new_new_n28502__;
  assign new_new_n28505__ = ~new_new_n28503__ & ~new_new_n28504__;
  assign new_new_n28506__ = ~new_new_n28414__ & new_new_n28505__;
  assign new_new_n28507__ = new_new_n28414__ & ~new_new_n28505__;
  assign new_new_n28508__ = ~new_new_n28506__ & ~new_new_n28507__;
  assign new_new_n28509__ = ~new_new_n28404__ & ~new_new_n28508__;
  assign new_new_n28510__ = ~new_new_n28403__ & ~new_new_n28509__;
  assign new_new_n28511__ = ~new_new_n27495__ & new_new_n28510__;
  assign new_new_n28512__ = new_new_n27495__ & ~new_new_n28510__;
  assign new_new_n28513__ = new_new_n6629__ & new_new_n26971__;
  assign new_new_n28514__ = ~new_new_n6625__ & ~new_new_n26978__;
  assign new_new_n28515__ = new_new_n6936__ & new_new_n28005__;
  assign new_new_n28516__ = ~new_new_n28513__ & ~new_new_n28514__;
  assign new_new_n28517__ = ~new_new_n28515__ & new_new_n28516__;
  assign new_new_n28518__ = new_new_n6631__ & ~new_new_n26937__;
  assign new_new_n28519__ = pi20 & ~new_new_n28518__;
  assign new_new_n28520__ = new_new_n7015__ & ~new_new_n26937__;
  assign new_new_n28521__ = ~new_new_n28519__ & ~new_new_n28520__;
  assign new_new_n28522__ = new_new_n28517__ & ~new_new_n28521__;
  assign new_new_n28523__ = ~pi20 & ~new_new_n28517__;
  assign new_new_n28524__ = ~new_new_n28522__ & ~new_new_n28523__;
  assign new_new_n28525__ = new_new_n28414__ & ~new_new_n28504__;
  assign new_new_n28526__ = ~new_new_n28503__ & ~new_new_n28525__;
  assign new_new_n28527__ = ~new_new_n333__ & ~new_new_n27054__;
  assign new_new_n28528__ = new_new_n873__ & ~new_new_n27033__;
  assign new_new_n28529__ = ~new_new_n447__ & new_new_n27686__;
  assign new_new_n28530__ = ~new_new_n27111__ & ~new_new_n28529__;
  assign new_new_n28531__ = new_new_n27111__ & new_new_n28529__;
  assign new_new_n28532__ = new_new_n801__ & ~new_new_n28530__;
  assign new_new_n28533__ = ~new_new_n28531__ & new_new_n28532__;
  assign new_new_n28534__ = ~new_new_n28527__ & ~new_new_n28528__;
  assign new_new_n28535__ = ~new_new_n28533__ & new_new_n28534__;
  assign new_new_n28536__ = pi26 & ~new_new_n28535__;
  assign new_new_n28537__ = ~pi26 & new_new_n28535__;
  assign new_new_n28538__ = ~new_new_n28536__ & ~new_new_n28537__;
  assign new_new_n28539__ = new_new_n28341__ & ~new_new_n28476__;
  assign new_new_n28540__ = ~new_new_n28463__ & ~new_new_n28466__;
  assign new_new_n28541__ = ~new_new_n28539__ & new_new_n28540__;
  assign new_new_n28542__ = ~new_new_n28464__ & ~new_new_n28541__;
  assign new_new_n28543__ = new_new_n4813__ & new_new_n27567__;
  assign new_new_n28544__ = ~new_new_n4818__ & new_new_n27059__;
  assign new_new_n28545__ = new_new_n4212__ & ~new_new_n27071__;
  assign new_new_n28546__ = ~new_new_n28544__ & ~new_new_n28545__;
  assign new_new_n28547__ = ~new_new_n28543__ & new_new_n28546__;
  assign new_new_n28548__ = new_new_n4214__ & new_new_n27041__;
  assign new_new_n28549__ = pi29 & ~new_new_n28548__;
  assign new_new_n28550__ = new_new_n5732__ & new_new_n27041__;
  assign new_new_n28551__ = ~new_new_n28549__ & ~new_new_n28550__;
  assign new_new_n28552__ = new_new_n28547__ & ~new_new_n28551__;
  assign new_new_n28553__ = ~pi29 & ~new_new_n28547__;
  assign new_new_n28554__ = ~new_new_n28552__ & ~new_new_n28553__;
  assign new_new_n28555__ = new_new_n28459__ & ~new_new_n28554__;
  assign new_new_n28556__ = ~new_new_n28459__ & new_new_n28554__;
  assign new_new_n28557__ = ~new_new_n28555__ & ~new_new_n28556__;
  assign new_new_n28558__ = ~new_new_n282__ & ~new_new_n312__;
  assign new_new_n28559__ = new_new_n83__ & ~new_new_n160__;
  assign new_new_n28560__ = ~new_new_n390__ & new_new_n1332__;
  assign new_new_n28561__ = ~new_new_n1506__ & new_new_n4314__;
  assign new_new_n28562__ = new_new_n19270__ & new_new_n28558__;
  assign new_new_n28563__ = new_new_n28561__ & new_new_n28562__;
  assign new_new_n28564__ = new_new_n28559__ & new_new_n28560__;
  assign new_new_n28565__ = new_new_n1037__ & ~new_new_n1105__;
  assign new_new_n28566__ = new_new_n2341__ & new_new_n5623__;
  assign new_new_n28567__ = new_new_n7400__ & new_new_n28566__;
  assign new_new_n28568__ = new_new_n28564__ & new_new_n28565__;
  assign new_new_n28569__ = new_new_n17260__ & new_new_n28563__;
  assign new_new_n28570__ = new_new_n28568__ & new_new_n28569__;
  assign new_new_n28571__ = new_new_n5697__ & new_new_n28567__;
  assign new_new_n28572__ = new_new_n28570__ & new_new_n28571__;
  assign new_new_n28573__ = ~new_new_n1064__ & new_new_n1627__;
  assign new_new_n28574__ = ~new_new_n441__ & ~new_new_n656__;
  assign new_new_n28575__ = ~new_new_n937__ & ~new_new_n1176__;
  assign new_new_n28576__ = ~new_new_n1210__ & new_new_n28575__;
  assign new_new_n28577__ = new_new_n2754__ & new_new_n28574__;
  assign new_new_n28578__ = new_new_n28576__ & new_new_n28577__;
  assign new_new_n28579__ = new_new_n1164__ & new_new_n3583__;
  assign new_new_n28580__ = new_new_n19013__ & new_new_n28579__;
  assign new_new_n28581__ = ~new_new_n895__ & new_new_n28578__;
  assign new_new_n28582__ = new_new_n28580__ & new_new_n28581__;
  assign new_new_n28583__ = new_new_n28573__ & new_new_n28582__;
  assign new_new_n28584__ = ~new_new_n130__ & ~new_new_n315__;
  assign new_new_n28585__ = ~new_new_n445__ & ~new_new_n584__;
  assign new_new_n28586__ = new_new_n28584__ & new_new_n28585__;
  assign new_new_n28587__ = ~new_new_n835__ & new_new_n1742__;
  assign new_new_n28588__ = new_new_n3805__ & new_new_n28587__;
  assign new_new_n28589__ = new_new_n1341__ & new_new_n28586__;
  assign new_new_n28590__ = new_new_n1516__ & new_new_n2378__;
  assign new_new_n28591__ = new_new_n2850__ & new_new_n7523__;
  assign new_new_n28592__ = new_new_n18481__ & new_new_n28591__;
  assign new_new_n28593__ = new_new_n28589__ & new_new_n28590__;
  assign new_new_n28594__ = new_new_n2641__ & new_new_n28588__;
  assign new_new_n28595__ = new_new_n19326__ & new_new_n28594__;
  assign new_new_n28596__ = new_new_n28592__ & new_new_n28593__;
  assign new_new_n28597__ = new_new_n1635__ & new_new_n28596__;
  assign new_new_n28598__ = new_new_n28595__ & new_new_n28597__;
  assign new_new_n28599__ = new_new_n28572__ & new_new_n28583__;
  assign new_new_n28600__ = new_new_n28598__ & new_new_n28599__;
  assign new_new_n28601__ = new_new_n19157__ & new_new_n28600__;
  assign new_new_n28602__ = new_new_n5059__ & new_new_n28601__;
  assign new_new_n28603__ = pi31 & new_new_n28601__;
  assign new_new_n28604__ = ~pi31 & ~new_new_n28601__;
  assign new_new_n28605__ = ~new_new_n28603__ & ~new_new_n28604__;
  assign new_new_n28606__ = ~new_new_n71__ & new_new_n26118__;
  assign new_new_n28607__ = ~new_new_n28605__ & new_new_n28606__;
  assign new_new_n28608__ = new_new_n161__ & new_new_n28604__;
  assign new_new_n28609__ = ~new_new_n28607__ & ~new_new_n28608__;
  assign new_new_n28610__ = ~new_new_n27075__ & ~new_new_n28609__;
  assign new_new_n28611__ = new_new_n27075__ & ~new_new_n28601__;
  assign new_new_n28612__ = ~new_new_n161__ & new_new_n28605__;
  assign new_new_n28613__ = ~new_new_n28611__ & new_new_n28612__;
  assign new_new_n28614__ = ~new_new_n28606__ & new_new_n28613__;
  assign new_new_n28615__ = new_new_n765__ & new_new_n26118__;
  assign new_new_n28616__ = ~new_new_n28601__ & ~new_new_n28615__;
  assign new_new_n28617__ = new_new_n28601__ & new_new_n28615__;
  assign new_new_n28618__ = new_new_n27075__ & ~new_new_n28616__;
  assign new_new_n28619__ = ~new_new_n28617__ & new_new_n28618__;
  assign new_new_n28620__ = ~new_new_n28602__ & ~new_new_n28614__;
  assign new_new_n28621__ = ~new_new_n28610__ & new_new_n28620__;
  assign new_new_n28622__ = ~new_new_n28619__ & new_new_n28621__;
  assign new_new_n28623__ = ~new_new_n28557__ & new_new_n28622__;
  assign new_new_n28624__ = new_new_n28557__ & ~new_new_n28622__;
  assign new_new_n28625__ = ~new_new_n28623__ & ~new_new_n28624__;
  assign new_new_n28626__ = new_new_n28542__ & ~new_new_n28625__;
  assign new_new_n28627__ = ~new_new_n28542__ & new_new_n28625__;
  assign new_new_n28628__ = ~new_new_n28626__ & ~new_new_n28627__;
  assign new_new_n28629__ = new_new_n28538__ & ~new_new_n28628__;
  assign new_new_n28630__ = ~new_new_n28538__ & new_new_n28628__;
  assign new_new_n28631__ = ~new_new_n28629__ & ~new_new_n28630__;
  assign new_new_n28632__ = new_new_n5213__ & ~new_new_n27003__;
  assign new_new_n28633__ = new_new_n5191__ & ~new_new_n27021__;
  assign new_new_n28634__ = new_new_n5183__ & ~new_new_n27029__;
  assign new_new_n28635__ = ~new_new_n28633__ & ~new_new_n28634__;
  assign new_new_n28636__ = ~new_new_n28632__ & new_new_n28635__;
  assign new_new_n28637__ = new_new_n5195__ & new_new_n27962__;
  assign new_new_n28638__ = pi23 & ~new_new_n28637__;
  assign new_new_n28639__ = new_new_n7878__ & new_new_n27962__;
  assign new_new_n28640__ = ~new_new_n28638__ & ~new_new_n28639__;
  assign new_new_n28641__ = new_new_n28636__ & ~new_new_n28640__;
  assign new_new_n28642__ = ~pi23 & ~new_new_n28636__;
  assign new_new_n28643__ = ~new_new_n28641__ & ~new_new_n28642__;
  assign new_new_n28644__ = ~new_new_n28493__ & ~new_new_n28500__;
  assign new_new_n28645__ = ~new_new_n28492__ & ~new_new_n28644__;
  assign new_new_n28646__ = ~new_new_n28643__ & ~new_new_n28645__;
  assign new_new_n28647__ = new_new_n28643__ & new_new_n28645__;
  assign new_new_n28648__ = ~new_new_n28646__ & ~new_new_n28647__;
  assign new_new_n28649__ = ~new_new_n28631__ & new_new_n28648__;
  assign new_new_n28650__ = new_new_n28631__ & ~new_new_n28648__;
  assign new_new_n28651__ = ~new_new_n28649__ & ~new_new_n28650__;
  assign new_new_n28652__ = new_new_n28526__ & ~new_new_n28651__;
  assign new_new_n28653__ = ~new_new_n28526__ & new_new_n28651__;
  assign new_new_n28654__ = ~new_new_n28652__ & ~new_new_n28653__;
  assign new_new_n28655__ = ~new_new_n28524__ & new_new_n28654__;
  assign new_new_n28656__ = new_new_n28524__ & ~new_new_n28654__;
  assign new_new_n28657__ = ~new_new_n28655__ & ~new_new_n28656__;
  assign new_new_n28658__ = ~new_new_n28512__ & ~new_new_n28657__;
  assign new_new_n28659__ = ~new_new_n28511__ & ~new_new_n28658__;
  assign new_new_n28660__ = new_new_n27469__ & new_new_n28659__;
  assign new_new_n28661__ = new_new_n6634__ & new_new_n27152__;
  assign new_new_n28662__ = ~new_new_n6625__ & new_new_n26971__;
  assign new_new_n28663__ = new_new_n6629__ & ~new_new_n26937__;
  assign new_new_n28664__ = new_new_n27152__ & ~new_new_n27477__;
  assign new_new_n28665__ = ~new_new_n27152__ & new_new_n27477__;
  assign new_new_n28666__ = ~new_new_n28664__ & ~new_new_n28665__;
  assign new_new_n28667__ = new_new_n6936__ & ~new_new_n28666__;
  assign new_new_n28668__ = ~new_new_n28662__ & ~new_new_n28663__;
  assign new_new_n28669__ = ~new_new_n28661__ & new_new_n28668__;
  assign new_new_n28670__ = ~new_new_n28667__ & new_new_n28669__;
  assign new_new_n28671__ = ~pi20 & new_new_n28670__;
  assign new_new_n28672__ = pi20 & ~new_new_n28670__;
  assign new_new_n28673__ = ~new_new_n28671__ & ~new_new_n28672__;
  assign new_new_n28674__ = new_new_n5191__ & ~new_new_n27029__;
  assign new_new_n28675__ = new_new_n5183__ & ~new_new_n27003__;
  assign new_new_n28676__ = ~new_new_n5212__ & new_new_n26978__;
  assign new_new_n28677__ = new_new_n5212__ & ~new_new_n27986__;
  assign new_new_n28678__ = new_new_n5195__ & ~new_new_n28676__;
  assign new_new_n28679__ = ~new_new_n28677__ & new_new_n28678__;
  assign new_new_n28680__ = ~new_new_n28674__ & ~new_new_n28675__;
  assign new_new_n28681__ = ~new_new_n28679__ & new_new_n28680__;
  assign new_new_n28682__ = pi23 & ~new_new_n28681__;
  assign new_new_n28683__ = ~pi23 & new_new_n28681__;
  assign new_new_n28684__ = ~new_new_n28682__ & ~new_new_n28683__;
  assign new_new_n28685__ = ~new_new_n28631__ & ~new_new_n28647__;
  assign new_new_n28686__ = ~new_new_n28646__ & ~new_new_n28685__;
  assign new_new_n28687__ = ~new_new_n28538__ & ~new_new_n28626__;
  assign new_new_n28688__ = ~new_new_n28627__ & ~new_new_n28687__;
  assign new_new_n28689__ = new_new_n8646__ & ~new_new_n27075__;
  assign new_new_n28690__ = ~new_new_n28615__ & new_new_n28689__;
  assign new_new_n28691__ = new_new_n28615__ & ~new_new_n28689__;
  assign new_new_n28692__ = ~new_new_n28690__ & ~new_new_n28691__;
  assign new_new_n28693__ = ~new_new_n28601__ & ~new_new_n28692__;
  assign new_new_n28694__ = ~new_new_n259__ & ~new_new_n772__;
  assign new_new_n28695__ = ~new_new_n1176__ & new_new_n28694__;
  assign new_new_n28696__ = ~new_new_n427__ & new_new_n3440__;
  assign new_new_n28697__ = ~new_new_n747__ & new_new_n1563__;
  assign new_new_n28698__ = new_new_n1741__ & new_new_n3258__;
  assign new_new_n28699__ = new_new_n3625__ & new_new_n16470__;
  assign new_new_n28700__ = new_new_n28698__ & new_new_n28699__;
  assign new_new_n28701__ = new_new_n28696__ & new_new_n28697__;
  assign new_new_n28702__ = new_new_n323__ & new_new_n28695__;
  assign new_new_n28703__ = new_new_n633__ & new_new_n941__;
  assign new_new_n28704__ = new_new_n3368__ & new_new_n28703__;
  assign new_new_n28705__ = new_new_n28701__ & new_new_n28702__;
  assign new_new_n28706__ = new_new_n1562__ & new_new_n28700__;
  assign new_new_n28707__ = new_new_n3959__ & new_new_n28706__;
  assign new_new_n28708__ = new_new_n28704__ & new_new_n28705__;
  assign new_new_n28709__ = new_new_n4959__ & new_new_n28708__;
  assign new_new_n28710__ = new_new_n6255__ & new_new_n28707__;
  assign new_new_n28711__ = new_new_n28709__ & new_new_n28710__;
  assign new_new_n28712__ = new_new_n7490__ & new_new_n28711__;
  assign new_new_n28713__ = new_new_n19157__ & new_new_n28712__;
  assign new_new_n28714__ = new_new_n28693__ & ~new_new_n28713__;
  assign new_new_n28715__ = new_new_n1424__ & new_new_n28713__;
  assign new_new_n28716__ = ~new_new_n28693__ & new_new_n28715__;
  assign new_new_n28717__ = ~new_new_n28714__ & ~new_new_n28716__;
  assign new_new_n28718__ = ~new_new_n26118__ & new_new_n27059__;
  assign new_new_n28719__ = new_new_n765__ & new_new_n28718__;
  assign new_new_n28720__ = ~new_new_n161__ & ~new_new_n27059__;
  assign new_new_n28721__ = new_new_n4876__ & ~new_new_n28720__;
  assign new_new_n28722__ = new_new_n27059__ & ~new_new_n27075__;
  assign new_new_n28723__ = ~new_new_n161__ & new_new_n27553__;
  assign new_new_n28724__ = ~new_new_n71__ & ~new_new_n28722__;
  assign new_new_n28725__ = ~new_new_n28723__ & new_new_n28724__;
  assign new_new_n28726__ = pi31 & ~new_new_n28725__;
  assign new_new_n28727__ = ~new_new_n28721__ & ~new_new_n28726__;
  assign new_new_n28728__ = new_new_n26118__ & ~new_new_n28727__;
  assign new_new_n28729__ = new_new_n5059__ & ~new_new_n27075__;
  assign new_new_n28730__ = ~new_new_n28719__ & ~new_new_n28729__;
  assign new_new_n28731__ = ~new_new_n28728__ & new_new_n28730__;
  assign new_new_n28732__ = ~new_new_n28717__ & new_new_n28731__;
  assign new_new_n28733__ = new_new_n28717__ & ~new_new_n28731__;
  assign new_new_n28734__ = ~new_new_n28732__ & ~new_new_n28733__;
  assign new_new_n28735__ = new_new_n4815__ & ~new_new_n27054__;
  assign new_new_n28736__ = ~new_new_n4818__ & ~new_new_n27071__;
  assign new_new_n28737__ = new_new_n4212__ & new_new_n27041__;
  assign new_new_n28738__ = ~new_new_n28736__ & ~new_new_n28737__;
  assign new_new_n28739__ = ~new_new_n28735__ & new_new_n28738__;
  assign new_new_n28740__ = new_new_n4214__ & ~new_new_n27094__;
  assign new_new_n28741__ = ~pi29 & ~new_new_n28740__;
  assign new_new_n28742__ = new_new_n5732__ & ~new_new_n27094__;
  assign new_new_n28743__ = ~new_new_n28741__ & ~new_new_n28742__;
  assign new_new_n28744__ = new_new_n28739__ & ~new_new_n28743__;
  assign new_new_n28745__ = pi29 & ~new_new_n28739__;
  assign new_new_n28746__ = ~new_new_n28744__ & ~new_new_n28745__;
  assign new_new_n28747__ = new_new_n28734__ & new_new_n28746__;
  assign new_new_n28748__ = ~new_new_n28734__ & ~new_new_n28746__;
  assign new_new_n28749__ = ~new_new_n28747__ & ~new_new_n28748__;
  assign new_new_n28750__ = ~new_new_n28556__ & new_new_n28622__;
  assign new_new_n28751__ = ~new_new_n28555__ & ~new_new_n28750__;
  assign new_new_n28752__ = new_new_n28749__ & ~new_new_n28751__;
  assign new_new_n28753__ = ~new_new_n28749__ & new_new_n28751__;
  assign new_new_n28754__ = ~new_new_n28752__ & ~new_new_n28753__;
  assign new_new_n28755__ = new_new_n3311__ & ~new_new_n27021__;
  assign new_new_n28756__ = new_new_n873__ & new_new_n27111__;
  assign new_new_n28757__ = ~new_new_n333__ & ~new_new_n27033__;
  assign new_new_n28758__ = ~new_new_n4900__ & new_new_n27796__;
  assign new_new_n28759__ = ~new_new_n28756__ & ~new_new_n28757__;
  assign new_new_n28760__ = ~new_new_n28755__ & new_new_n28759__;
  assign new_new_n28761__ = ~new_new_n28758__ & new_new_n28760__;
  assign new_new_n28762__ = pi26 & ~new_new_n28761__;
  assign new_new_n28763__ = ~pi26 & new_new_n28761__;
  assign new_new_n28764__ = ~new_new_n28762__ & ~new_new_n28763__;
  assign new_new_n28765__ = new_new_n28754__ & new_new_n28764__;
  assign new_new_n28766__ = ~new_new_n28754__ & ~new_new_n28764__;
  assign new_new_n28767__ = ~new_new_n28765__ & ~new_new_n28766__;
  assign new_new_n28768__ = new_new_n28688__ & new_new_n28767__;
  assign new_new_n28769__ = ~new_new_n28688__ & ~new_new_n28767__;
  assign new_new_n28770__ = ~new_new_n28768__ & ~new_new_n28769__;
  assign new_new_n28771__ = new_new_n28686__ & ~new_new_n28770__;
  assign new_new_n28772__ = ~new_new_n28686__ & new_new_n28770__;
  assign new_new_n28773__ = ~new_new_n28771__ & ~new_new_n28772__;
  assign new_new_n28774__ = new_new_n28684__ & new_new_n28773__;
  assign new_new_n28775__ = ~new_new_n28684__ & ~new_new_n28773__;
  assign new_new_n28776__ = ~new_new_n28774__ & ~new_new_n28775__;
  assign new_new_n28777__ = new_new_n28673__ & new_new_n28776__;
  assign new_new_n28778__ = ~new_new_n28673__ & ~new_new_n28776__;
  assign new_new_n28779__ = ~new_new_n28777__ & ~new_new_n28778__;
  assign new_new_n28780__ = new_new_n28524__ & ~new_new_n28653__;
  assign new_new_n28781__ = ~new_new_n28652__ & ~new_new_n28780__;
  assign new_new_n28782__ = ~new_new_n28779__ & new_new_n28781__;
  assign new_new_n28783__ = new_new_n28779__ & ~new_new_n28781__;
  assign new_new_n28784__ = ~new_new_n28782__ & ~new_new_n28783__;
  assign new_new_n28785__ = ~new_new_n27469__ & ~new_new_n28659__;
  assign new_new_n28786__ = ~new_new_n28660__ & ~new_new_n28785__;
  assign new_new_n28787__ = ~new_new_n28784__ & new_new_n28786__;
  assign new_new_n28788__ = ~new_new_n28660__ & ~new_new_n28787__;
  assign new_new_n28789__ = new_new_n6968__ & new_new_n26917__;
  assign new_new_n28790__ = new_new_n6964__ & new_new_n26928__;
  assign new_new_n28791__ = new_new_n7935__ & ~new_new_n27168__;
  assign new_new_n28792__ = ~new_new_n28790__ & ~new_new_n28791__;
  assign new_new_n28793__ = ~new_new_n28789__ & new_new_n28792__;
  assign new_new_n28794__ = ~new_new_n27162__ & new_new_n27168__;
  assign new_new_n28795__ = new_new_n27162__ & ~new_new_n27168__;
  assign new_new_n28796__ = ~new_new_n28794__ & ~new_new_n28795__;
  assign new_new_n28797__ = new_new_n26917__ & ~new_new_n28796__;
  assign new_new_n28798__ = ~new_new_n26917__ & new_new_n28796__;
  assign new_new_n28799__ = ~new_new_n28797__ & ~new_new_n28798__;
  assign new_new_n28800__ = new_new_n6958__ & ~new_new_n28799__;
  assign new_new_n28801__ = pi17 & ~new_new_n28800__;
  assign new_new_n28802__ = new_new_n7942__ & ~new_new_n28799__;
  assign new_new_n28803__ = ~new_new_n28801__ & ~new_new_n28802__;
  assign new_new_n28804__ = new_new_n28793__ & ~new_new_n28803__;
  assign new_new_n28805__ = ~pi17 & ~new_new_n28793__;
  assign new_new_n28806__ = ~new_new_n28804__ & ~new_new_n28805__;
  assign new_new_n28807__ = ~new_new_n28788__ & ~new_new_n28806__;
  assign new_new_n28808__ = new_new_n28788__ & new_new_n28806__;
  assign new_new_n28809__ = ~new_new_n28807__ & ~new_new_n28808__;
  assign new_new_n28810__ = new_new_n5215__ & new_new_n28277__;
  assign new_new_n28811__ = new_new_n5191__ & ~new_new_n27003__;
  assign new_new_n28812__ = new_new_n5183__ & ~new_new_n26978__;
  assign new_new_n28813__ = ~new_new_n28811__ & ~new_new_n28812__;
  assign new_new_n28814__ = ~new_new_n28810__ & new_new_n28813__;
  assign new_new_n28815__ = new_new_n5195__ & new_new_n26971__;
  assign new_new_n28816__ = pi23 & ~new_new_n28815__;
  assign new_new_n28817__ = new_new_n5974__ & new_new_n26971__;
  assign new_new_n28818__ = ~new_new_n28816__ & ~new_new_n28817__;
  assign new_new_n28819__ = new_new_n28814__ & ~new_new_n28818__;
  assign new_new_n28820__ = ~pi23 & ~new_new_n28814__;
  assign new_new_n28821__ = ~new_new_n28819__ & ~new_new_n28820__;
  assign new_new_n28822__ = new_new_n3311__ & ~new_new_n27029__;
  assign new_new_n28823__ = new_new_n873__ & ~new_new_n27021__;
  assign new_new_n28824__ = ~new_new_n333__ & new_new_n27111__;
  assign new_new_n28825__ = ~new_new_n4900__ & new_new_n27764__;
  assign new_new_n28826__ = ~new_new_n28823__ & ~new_new_n28824__;
  assign new_new_n28827__ = ~new_new_n28822__ & new_new_n28826__;
  assign new_new_n28828__ = ~new_new_n28825__ & new_new_n28827__;
  assign new_new_n28829__ = pi26 & ~new_new_n28828__;
  assign new_new_n28830__ = ~pi26 & new_new_n28828__;
  assign new_new_n28831__ = ~new_new_n28829__ & ~new_new_n28830__;
  assign new_new_n28832__ = ~new_new_n28765__ & ~new_new_n28768__;
  assign new_new_n28833__ = new_new_n28831__ & ~new_new_n28832__;
  assign new_new_n28834__ = ~new_new_n28831__ & new_new_n28832__;
  assign new_new_n28835__ = ~new_new_n28833__ & ~new_new_n28834__;
  assign new_new_n28836__ = ~new_new_n4818__ & new_new_n27041__;
  assign new_new_n28837__ = new_new_n4212__ & ~new_new_n27054__;
  assign new_new_n28838__ = ~new_new_n28836__ & ~new_new_n28837__;
  assign new_new_n28839__ = new_new_n4214__ & ~new_new_n27535__;
  assign new_new_n28840__ = pi29 & ~new_new_n28839__;
  assign new_new_n28841__ = ~pi28 & new_new_n27033__;
  assign new_new_n28842__ = pi28 & ~new_new_n27033__;
  assign new_new_n28843__ = new_new_n4214__ & ~new_new_n28841__;
  assign new_new_n28844__ = ~new_new_n28842__ & new_new_n28843__;
  assign new_new_n28845__ = ~new_new_n27102__ & new_new_n28844__;
  assign new_new_n28846__ = ~new_new_n28840__ & ~new_new_n28845__;
  assign new_new_n28847__ = new_new_n28838__ & ~new_new_n28846__;
  assign new_new_n28848__ = new_new_n4214__ & new_new_n27545__;
  assign new_new_n28849__ = new_new_n28838__ & ~new_new_n28848__;
  assign new_new_n28850__ = ~pi29 & ~new_new_n28849__;
  assign new_new_n28851__ = ~new_new_n28847__ & ~new_new_n28850__;
  assign new_new_n28852__ = ~new_new_n71__ & ~new_new_n27071__;
  assign new_new_n28853__ = ~new_new_n28606__ & ~new_new_n28852__;
  assign new_new_n28854__ = new_new_n27071__ & ~new_new_n27075__;
  assign new_new_n28855__ = ~new_new_n27071__ & ~new_new_n27087__;
  assign new_new_n28856__ = ~new_new_n161__ & ~new_new_n28854__;
  assign new_new_n28857__ = ~new_new_n28855__ & new_new_n28856__;
  assign new_new_n28858__ = ~new_new_n28853__ & ~new_new_n28857__;
  assign new_new_n28859__ = ~new_new_n27059__ & ~new_new_n28858__;
  assign new_new_n28860__ = new_new_n161__ & ~new_new_n26118__;
  assign new_new_n28861__ = ~new_new_n161__ & new_new_n27071__;
  assign new_new_n28862__ = new_new_n26118__ & ~new_new_n28861__;
  assign new_new_n28863__ = new_new_n27059__ & ~new_new_n28853__;
  assign new_new_n28864__ = ~new_new_n28862__ & new_new_n28863__;
  assign new_new_n28865__ = pi31 & ~new_new_n28860__;
  assign new_new_n28866__ = ~new_new_n28864__ & new_new_n28865__;
  assign new_new_n28867__ = ~new_new_n28859__ & new_new_n28866__;
  assign new_new_n28868__ = new_new_n161__ & new_new_n27059__;
  assign new_new_n28869__ = new_new_n765__ & ~new_new_n27071__;
  assign new_new_n28870__ = ~new_new_n28868__ & ~new_new_n28869__;
  assign new_new_n28871__ = ~pi31 & ~new_new_n28870__;
  assign new_new_n28872__ = ~new_new_n28867__ & ~new_new_n28871__;
  assign new_new_n28873__ = ~new_new_n28714__ & ~new_new_n28733__;
  assign new_new_n28874__ = ~new_new_n28872__ & ~new_new_n28873__;
  assign new_new_n28875__ = new_new_n28872__ & new_new_n28873__;
  assign new_new_n28876__ = ~new_new_n28874__ & ~new_new_n28875__;
  assign new_new_n28877__ = ~new_new_n476__ & ~new_new_n853__;
  assign new_new_n28878__ = ~new_new_n1081__ & new_new_n28877__;
  assign new_new_n28879__ = new_new_n672__ & ~new_new_n919__;
  assign new_new_n28880__ = new_new_n1106__ & new_new_n2895__;
  assign new_new_n28881__ = new_new_n19384__ & new_new_n28880__;
  assign new_new_n28882__ = new_new_n28878__ & new_new_n28879__;
  assign new_new_n28883__ = new_new_n1097__ & new_new_n3793__;
  assign new_new_n28884__ = new_new_n28882__ & new_new_n28883__;
  assign new_new_n28885__ = new_new_n440__ & new_new_n28881__;
  assign new_new_n28886__ = new_new_n2165__ & new_new_n3634__;
  assign new_new_n28887__ = new_new_n28885__ & new_new_n28886__;
  assign new_new_n28888__ = new_new_n4986__ & new_new_n28884__;
  assign new_new_n28889__ = new_new_n28887__ & new_new_n28888__;
  assign new_new_n28890__ = new_new_n6195__ & new_new_n28889__;
  assign new_new_n28891__ = new_new_n1699__ & new_new_n28890__;
  assign new_new_n28892__ = new_new_n2466__ & new_new_n28891__;
  assign new_new_n28893__ = ~new_new_n28876__ & new_new_n28892__;
  assign new_new_n28894__ = new_new_n28876__ & ~new_new_n28892__;
  assign new_new_n28895__ = ~new_new_n28893__ & ~new_new_n28894__;
  assign new_new_n28896__ = ~new_new_n28748__ & ~new_new_n28751__;
  assign new_new_n28897__ = ~new_new_n28747__ & ~new_new_n28896__;
  assign new_new_n28898__ = new_new_n28895__ & ~new_new_n28897__;
  assign new_new_n28899__ = ~new_new_n28895__ & new_new_n28897__;
  assign new_new_n28900__ = ~new_new_n28898__ & ~new_new_n28899__;
  assign new_new_n28901__ = ~new_new_n28851__ & ~new_new_n28900__;
  assign new_new_n28902__ = new_new_n28851__ & new_new_n28900__;
  assign new_new_n28903__ = ~new_new_n28901__ & ~new_new_n28902__;
  assign new_new_n28904__ = ~new_new_n28835__ & new_new_n28903__;
  assign new_new_n28905__ = new_new_n28835__ & ~new_new_n28903__;
  assign new_new_n28906__ = ~new_new_n28904__ & ~new_new_n28905__;
  assign new_new_n28907__ = new_new_n28821__ & ~new_new_n28906__;
  assign new_new_n28908__ = ~new_new_n28821__ & new_new_n28906__;
  assign new_new_n28909__ = ~new_new_n28907__ & ~new_new_n28908__;
  assign new_new_n28910__ = new_new_n28684__ & ~new_new_n28771__;
  assign new_new_n28911__ = ~new_new_n28772__ & ~new_new_n28910__;
  assign new_new_n28912__ = ~new_new_n28909__ & new_new_n28911__;
  assign new_new_n28913__ = new_new_n28909__ & ~new_new_n28911__;
  assign new_new_n28914__ = ~new_new_n28912__ & ~new_new_n28913__;
  assign new_new_n28915__ = ~new_new_n28777__ & ~new_new_n28781__;
  assign new_new_n28916__ = ~new_new_n28778__ & ~new_new_n28915__;
  assign new_new_n28917__ = new_new_n28914__ & new_new_n28916__;
  assign new_new_n28918__ = ~new_new_n28914__ & ~new_new_n28916__;
  assign new_new_n28919__ = ~new_new_n28917__ & ~new_new_n28918__;
  assign new_new_n28920__ = new_new_n6629__ & new_new_n27152__;
  assign new_new_n28921__ = ~new_new_n6625__ & ~new_new_n26937__;
  assign new_new_n28922__ = new_new_n6634__ & ~new_new_n26941__;
  assign new_new_n28923__ = ~new_new_n28921__ & ~new_new_n28922__;
  assign new_new_n28924__ = ~new_new_n28920__ & new_new_n28923__;
  assign new_new_n28925__ = new_new_n6631__ & ~new_new_n27502__;
  assign new_new_n28926__ = ~pi20 & ~new_new_n28925__;
  assign new_new_n28927__ = new_new_n7015__ & ~new_new_n27502__;
  assign new_new_n28928__ = ~new_new_n28926__ & ~new_new_n28927__;
  assign new_new_n28929__ = new_new_n28924__ & ~new_new_n28928__;
  assign new_new_n28930__ = pi20 & ~new_new_n28924__;
  assign new_new_n28931__ = ~new_new_n28929__ & ~new_new_n28930__;
  assign new_new_n28932__ = ~new_new_n28919__ & new_new_n28931__;
  assign new_new_n28933__ = new_new_n28919__ & ~new_new_n28931__;
  assign new_new_n28934__ = ~new_new_n28932__ & ~new_new_n28933__;
  assign new_new_n28935__ = new_new_n28809__ & new_new_n28934__;
  assign new_new_n28936__ = ~new_new_n28809__ & ~new_new_n28934__;
  assign new_new_n28937__ = ~new_new_n28935__ & ~new_new_n28936__;
  assign new_new_n28938__ = ~new_new_n27437__ & ~new_new_n28937__;
  assign new_new_n28939__ = new_new_n27437__ & new_new_n28937__;
  assign new_new_n28940__ = ~new_new_n28938__ & ~new_new_n28939__;
  assign new_new_n28941__ = new_new_n28784__ & ~new_new_n28786__;
  assign new_new_n28942__ = ~new_new_n28787__ & ~new_new_n28941__;
  assign new_new_n28943__ = ~new_new_n28403__ & ~new_new_n28404__;
  assign new_new_n28944__ = new_new_n28508__ & ~new_new_n28943__;
  assign new_new_n28945__ = ~new_new_n28508__ & new_new_n28943__;
  assign new_new_n28946__ = ~new_new_n28944__ & ~new_new_n28945__;
  assign new_new_n28947__ = new_new_n6991__ & ~new_new_n26941__;
  assign new_new_n28948__ = new_new_n6985__ & new_new_n26928__;
  assign new_new_n28949__ = ~new_new_n28947__ & ~new_new_n28948__;
  assign new_new_n28950__ = new_new_n6994__ & new_new_n26917__;
  assign new_new_n28951__ = ~new_new_n27462__ & new_new_n28950__;
  assign new_new_n28952__ = new_new_n28949__ & ~new_new_n28951__;
  assign new_new_n28953__ = pi14 & ~new_new_n28952__;
  assign new_new_n28954__ = ~pi13 & new_new_n26917__;
  assign new_new_n28955__ = ~new_new_n26917__ & new_new_n27461__;
  assign new_new_n28956__ = new_new_n6994__ & ~new_new_n28955__;
  assign new_new_n28957__ = pi13 & ~new_new_n27462__;
  assign new_new_n28958__ = ~new_new_n28954__ & new_new_n28956__;
  assign new_new_n28959__ = ~new_new_n28957__ & new_new_n28958__;
  assign new_new_n28960__ = ~pi14 & new_new_n28949__;
  assign new_new_n28961__ = ~new_new_n28956__ & new_new_n28960__;
  assign new_new_n28962__ = ~new_new_n28953__ & ~new_new_n28961__;
  assign new_new_n28963__ = ~new_new_n28959__ & new_new_n28962__;
  assign new_new_n28964__ = ~new_new_n28294__ & ~new_new_n28295__;
  assign new_new_n28965__ = new_new_n28400__ & new_new_n28964__;
  assign new_new_n28966__ = ~new_new_n28400__ & ~new_new_n28964__;
  assign new_new_n28967__ = ~new_new_n28965__ & ~new_new_n28966__;
  assign new_new_n28968__ = new_new_n28963__ & new_new_n28967__;
  assign new_new_n28969__ = ~new_new_n28963__ & ~new_new_n28967__;
  assign new_new_n28970__ = new_new_n6985__ & new_new_n27152__;
  assign new_new_n28971__ = new_new_n6991__ & ~new_new_n26937__;
  assign new_new_n28972__ = ~new_new_n28970__ & ~new_new_n28971__;
  assign new_new_n28973__ = new_new_n6994__ & new_new_n27501__;
  assign new_new_n28974__ = new_new_n28972__ & ~new_new_n28973__;
  assign new_new_n28975__ = pi14 & ~new_new_n28974__;
  assign new_new_n28976__ = ~pi13 & ~new_new_n27484__;
  assign new_new_n28977__ = pi13 & ~new_new_n27482__;
  assign new_new_n28978__ = new_new_n6994__ & ~new_new_n28976__;
  assign new_new_n28979__ = ~new_new_n28977__ & new_new_n28978__;
  assign new_new_n28980__ = new_new_n26941__ & ~new_new_n27481__;
  assign new_new_n28981__ = new_new_n6994__ & ~new_new_n28980__;
  assign new_new_n28982__ = ~pi14 & new_new_n28972__;
  assign new_new_n28983__ = ~new_new_n28981__ & new_new_n28982__;
  assign new_new_n28984__ = ~new_new_n28975__ & ~new_new_n28983__;
  assign new_new_n28985__ = ~new_new_n28979__ & new_new_n28984__;
  assign new_new_n28986__ = new_new_n6985__ & new_new_n26971__;
  assign new_new_n28987__ = new_new_n6991__ & ~new_new_n26978__;
  assign new_new_n28988__ = ~new_new_n28986__ & ~new_new_n28987__;
  assign new_new_n28989__ = new_new_n6994__ & ~new_new_n26937__;
  assign new_new_n28990__ = new_new_n28005__ & new_new_n28989__;
  assign new_new_n28991__ = new_new_n28988__ & ~new_new_n28990__;
  assign new_new_n28992__ = ~pi14 & ~new_new_n28991__;
  assign new_new_n28993__ = ~pi13 & new_new_n28005__;
  assign new_new_n28994__ = new_new_n26937__ & ~new_new_n28005__;
  assign new_new_n28995__ = new_new_n6994__ & ~new_new_n28994__;
  assign new_new_n28996__ = pi13 & ~new_new_n26937__;
  assign new_new_n28997__ = ~new_new_n28993__ & ~new_new_n28996__;
  assign new_new_n28998__ = new_new_n28995__ & new_new_n28997__;
  assign new_new_n28999__ = pi14 & new_new_n28988__;
  assign new_new_n29000__ = ~new_new_n28995__ & new_new_n28999__;
  assign new_new_n29001__ = ~new_new_n28992__ & ~new_new_n28998__;
  assign new_new_n29002__ = ~new_new_n29000__ & new_new_n29001__;
  assign new_new_n29003__ = ~new_new_n28210__ & ~new_new_n28211__;
  assign new_new_n29004__ = ~new_new_n28221__ & new_new_n29003__;
  assign new_new_n29005__ = new_new_n28221__ & ~new_new_n29003__;
  assign new_new_n29006__ = ~new_new_n29004__ & ~new_new_n29005__;
  assign new_new_n29007__ = new_new_n6991__ & ~new_new_n27003__;
  assign new_new_n29008__ = new_new_n6985__ & ~new_new_n26978__;
  assign new_new_n29009__ = ~new_new_n29007__ & ~new_new_n29008__;
  assign new_new_n29010__ = new_new_n6994__ & new_new_n26971__;
  assign new_new_n29011__ = new_new_n28277__ & new_new_n29010__;
  assign new_new_n29012__ = new_new_n29009__ & ~new_new_n29011__;
  assign new_new_n29013__ = pi14 & ~new_new_n29012__;
  assign new_new_n29014__ = ~new_new_n26971__ & ~new_new_n28277__;
  assign new_new_n29015__ = new_new_n6994__ & ~new_new_n29014__;
  assign new_new_n29016__ = ~pi14 & new_new_n29009__;
  assign new_new_n29017__ = ~new_new_n29015__ & new_new_n29016__;
  assign new_new_n29018__ = ~pi13 & new_new_n26971__;
  assign new_new_n29019__ = pi13 & new_new_n28277__;
  assign new_new_n29020__ = ~new_new_n29018__ & ~new_new_n29019__;
  assign new_new_n29021__ = new_new_n29015__ & new_new_n29020__;
  assign new_new_n29022__ = ~new_new_n29013__ & ~new_new_n29017__;
  assign new_new_n29023__ = ~new_new_n29021__ & new_new_n29022__;
  assign new_new_n29024__ = ~new_new_n29006__ & new_new_n29023__;
  assign new_new_n29025__ = new_new_n29006__ & ~new_new_n29023__;
  assign new_new_n29026__ = new_new_n6991__ & ~new_new_n27029__;
  assign new_new_n29027__ = new_new_n6985__ & ~new_new_n27003__;
  assign new_new_n29028__ = ~new_new_n29026__ & ~new_new_n29027__;
  assign new_new_n29029__ = new_new_n6994__ & new_new_n27992__;
  assign new_new_n29030__ = new_new_n29028__ & ~new_new_n29029__;
  assign new_new_n29031__ = ~pi14 & ~new_new_n29030__;
  assign new_new_n29032__ = ~new_new_n26978__ & ~new_new_n27986__;
  assign new_new_n29033__ = ~pi13 & ~new_new_n29032__;
  assign new_new_n29034__ = new_new_n26978__ & new_new_n27986__;
  assign new_new_n29035__ = pi13 & ~new_new_n29034__;
  assign new_new_n29036__ = new_new_n6994__ & ~new_new_n29033__;
  assign new_new_n29037__ = ~new_new_n29035__ & new_new_n29036__;
  assign new_new_n29038__ = new_new_n6994__ & ~new_new_n27996__;
  assign new_new_n29039__ = pi14 & new_new_n29028__;
  assign new_new_n29040__ = ~new_new_n29038__ & new_new_n29039__;
  assign new_new_n29041__ = ~new_new_n29031__ & ~new_new_n29040__;
  assign new_new_n29042__ = ~new_new_n29037__ & new_new_n29041__;
  assign new_new_n29043__ = new_new_n6991__ & ~new_new_n27021__;
  assign new_new_n29044__ = new_new_n6985__ & ~new_new_n27029__;
  assign new_new_n29045__ = ~new_new_n29043__ & ~new_new_n29044__;
  assign new_new_n29046__ = new_new_n6994__ & ~new_new_n27003__;
  assign new_new_n29047__ = new_new_n27962__ & new_new_n29046__;
  assign new_new_n29048__ = new_new_n29045__ & ~new_new_n29047__;
  assign new_new_n29049__ = ~pi14 & ~new_new_n29048__;
  assign new_new_n29050__ = ~pi13 & new_new_n27962__;
  assign new_new_n29051__ = new_new_n27003__ & ~new_new_n27962__;
  assign new_new_n29052__ = new_new_n6994__ & ~new_new_n29051__;
  assign new_new_n29053__ = pi13 & ~new_new_n27003__;
  assign new_new_n29054__ = ~new_new_n29050__ & ~new_new_n29053__;
  assign new_new_n29055__ = new_new_n29052__ & new_new_n29054__;
  assign new_new_n29056__ = pi14 & new_new_n29045__;
  assign new_new_n29057__ = ~new_new_n29052__ & new_new_n29056__;
  assign new_new_n29058__ = ~new_new_n29049__ & ~new_new_n29055__;
  assign new_new_n29059__ = ~new_new_n29057__ & new_new_n29058__;
  assign new_new_n29060__ = ~new_new_n28184__ & ~new_new_n28185__;
  assign new_new_n29061__ = new_new_n28189__ & new_new_n29060__;
  assign new_new_n29062__ = ~new_new_n28189__ & ~new_new_n29060__;
  assign new_new_n29063__ = ~new_new_n29061__ & ~new_new_n29062__;
  assign new_new_n29064__ = new_new_n29059__ & new_new_n29063__;
  assign new_new_n29065__ = ~new_new_n29059__ & ~new_new_n29063__;
  assign new_new_n29066__ = ~new_new_n28158__ & ~new_new_n28159__;
  assign new_new_n29067__ = new_new_n28169__ & ~new_new_n29066__;
  assign new_new_n29068__ = ~new_new_n28169__ & new_new_n29066__;
  assign new_new_n29069__ = ~new_new_n29067__ & ~new_new_n29068__;
  assign new_new_n29070__ = ~new_new_n28153__ & ~new_new_n28155__;
  assign new_new_n29071__ = ~new_new_n28156__ & ~new_new_n29070__;
  assign new_new_n29072__ = new_new_n6985__ & ~new_new_n27033__;
  assign new_new_n29073__ = new_new_n6991__ & ~new_new_n27054__;
  assign new_new_n29074__ = ~new_new_n29072__ & ~new_new_n29073__;
  assign new_new_n29075__ = new_new_n6994__ & ~new_new_n27691__;
  assign new_new_n29076__ = pi14 & ~new_new_n29075__;
  assign new_new_n29077__ = new_new_n6994__ & new_new_n27111__;
  assign new_new_n29078__ = ~pi13 & new_new_n29077__;
  assign new_new_n29079__ = new_new_n27686__ & new_new_n29078__;
  assign new_new_n29080__ = ~new_new_n29076__ & ~new_new_n29079__;
  assign new_new_n29081__ = new_new_n29074__ & ~new_new_n29080__;
  assign new_new_n29082__ = ~new_new_n27686__ & new_new_n29077__;
  assign new_new_n29083__ = new_new_n29074__ & ~new_new_n29082__;
  assign new_new_n29084__ = ~pi14 & ~new_new_n29083__;
  assign new_new_n29085__ = new_new_n8820__ & ~new_new_n27111__;
  assign new_new_n29086__ = new_new_n27686__ & new_new_n29085__;
  assign new_new_n29087__ = ~new_new_n29084__ & ~new_new_n29086__;
  assign new_new_n29088__ = ~new_new_n29081__ & new_new_n29087__;
  assign new_new_n29089__ = new_new_n8388__ & new_new_n27103__;
  assign new_new_n29090__ = new_new_n6991__ & new_new_n27041__;
  assign new_new_n29091__ = new_new_n6985__ & ~new_new_n27054__;
  assign new_new_n29092__ = ~new_new_n29090__ & ~new_new_n29091__;
  assign new_new_n29093__ = new_new_n6994__ & ~new_new_n27535__;
  assign new_new_n29094__ = ~pi14 & ~new_new_n29093__;
  assign new_new_n29095__ = ~new_new_n27033__ & ~new_new_n27102__;
  assign new_new_n29096__ = new_new_n8820__ & new_new_n29095__;
  assign new_new_n29097__ = ~new_new_n29094__ & ~new_new_n29096__;
  assign new_new_n29098__ = new_new_n29092__ & ~new_new_n29097__;
  assign new_new_n29099__ = new_new_n6994__ & new_new_n27545__;
  assign new_new_n29100__ = new_new_n29092__ & ~new_new_n29099__;
  assign new_new_n29101__ = pi14 & ~new_new_n29100__;
  assign new_new_n29102__ = ~new_new_n29089__ & ~new_new_n29101__;
  assign new_new_n29103__ = ~new_new_n29098__ & new_new_n29102__;
  assign new_new_n29104__ = new_new_n6991__ & ~new_new_n27071__;
  assign new_new_n29105__ = new_new_n6985__ & new_new_n27041__;
  assign new_new_n29106__ = ~new_new_n29104__ & ~new_new_n29105__;
  assign new_new_n29107__ = new_new_n6994__ & ~new_new_n27054__;
  assign new_new_n29108__ = ~new_new_n27094__ & new_new_n29107__;
  assign new_new_n29109__ = new_new_n29106__ & ~new_new_n29108__;
  assign new_new_n29110__ = pi14 & ~new_new_n29109__;
  assign new_new_n29111__ = ~pi13 & ~new_new_n27054__;
  assign new_new_n29112__ = new_new_n27054__ & new_new_n27094__;
  assign new_new_n29113__ = new_new_n6994__ & ~new_new_n29112__;
  assign new_new_n29114__ = pi13 & ~new_new_n27094__;
  assign new_new_n29115__ = ~new_new_n29111__ & ~new_new_n29114__;
  assign new_new_n29116__ = new_new_n29113__ & new_new_n29115__;
  assign new_new_n29117__ = ~pi14 & new_new_n29106__;
  assign new_new_n29118__ = ~new_new_n29113__ & new_new_n29117__;
  assign new_new_n29119__ = ~new_new_n29110__ & ~new_new_n29116__;
  assign new_new_n29120__ = ~new_new_n29118__ & new_new_n29119__;
  assign new_new_n29121__ = new_new_n6985__ & ~new_new_n27071__;
  assign new_new_n29122__ = new_new_n6991__ & new_new_n27059__;
  assign new_new_n29123__ = ~new_new_n29121__ & ~new_new_n29122__;
  assign new_new_n29124__ = new_new_n6994__ & new_new_n27041__;
  assign new_new_n29125__ = new_new_n27567__ & new_new_n29124__;
  assign new_new_n29126__ = new_new_n29123__ & ~new_new_n29125__;
  assign new_new_n29127__ = ~pi14 & ~new_new_n29126__;
  assign new_new_n29128__ = new_new_n6994__ & ~new_new_n28088__;
  assign new_new_n29129__ = pi14 & new_new_n29123__;
  assign new_new_n29130__ = ~new_new_n29128__ & new_new_n29129__;
  assign new_new_n29131__ = pi13 & ~new_new_n28091__;
  assign new_new_n29132__ = ~pi13 & ~new_new_n28093__;
  assign new_new_n29133__ = new_new_n6994__ & ~new_new_n29132__;
  assign new_new_n29134__ = ~new_new_n29131__ & new_new_n29133__;
  assign new_new_n29135__ = ~new_new_n29127__ & ~new_new_n29130__;
  assign new_new_n29136__ = ~new_new_n29134__ & new_new_n29135__;
  assign new_new_n29137__ = new_new_n8388__ & new_new_n27846__;
  assign new_new_n29138__ = new_new_n6991__ & ~new_new_n27075__;
  assign new_new_n29139__ = new_new_n6985__ & new_new_n26118__;
  assign new_new_n29140__ = ~new_new_n29138__ & ~new_new_n29139__;
  assign new_new_n29141__ = ~new_new_n27059__ & ~new_new_n27582__;
  assign new_new_n29142__ = new_new_n6994__ & ~new_new_n29141__;
  assign new_new_n29143__ = ~pi14 & ~new_new_n29142__;
  assign new_new_n29144__ = new_new_n8820__ & new_new_n27582__;
  assign new_new_n29145__ = new_new_n27059__ & new_new_n29144__;
  assign new_new_n29146__ = ~new_new_n29143__ & ~new_new_n29145__;
  assign new_new_n29147__ = new_new_n29140__ & ~new_new_n29146__;
  assign new_new_n29148__ = new_new_n6994__ & ~new_new_n27582__;
  assign new_new_n29149__ = new_new_n27059__ & new_new_n29148__;
  assign new_new_n29150__ = new_new_n29140__ & ~new_new_n29149__;
  assign new_new_n29151__ = pi14 & ~new_new_n29150__;
  assign new_new_n29152__ = ~new_new_n29137__ & ~new_new_n29151__;
  assign new_new_n29153__ = ~new_new_n29147__ & new_new_n29152__;
  assign new_new_n29154__ = new_new_n6994__ & ~new_new_n27577__;
  assign new_new_n29155__ = new_new_n19825__ & ~new_new_n27075__;
  assign new_new_n29156__ = pi14 & ~new_new_n29155__;
  assign new_new_n29157__ = ~new_new_n29154__ & new_new_n29156__;
  assign new_new_n29158__ = new_new_n29153__ & new_new_n29157__;
  assign new_new_n29159__ = new_new_n6958__ & ~new_new_n27075__;
  assign new_new_n29160__ = ~new_new_n29158__ & ~new_new_n29159__;
  assign new_new_n29161__ = new_new_n6991__ & new_new_n26118__;
  assign new_new_n29162__ = new_new_n6985__ & new_new_n27059__;
  assign new_new_n29163__ = ~new_new_n29161__ & ~new_new_n29162__;
  assign new_new_n29164__ = new_new_n6994__ & new_new_n28442__;
  assign new_new_n29165__ = new_new_n29163__ & ~new_new_n29164__;
  assign new_new_n29166__ = ~pi14 & ~new_new_n29165__;
  assign new_new_n29167__ = ~pi13 & new_new_n27600__;
  assign new_new_n29168__ = new_new_n27071__ & ~new_new_n28441__;
  assign new_new_n29169__ = new_new_n6994__ & ~new_new_n29168__;
  assign new_new_n29170__ = pi13 & ~new_new_n27071__;
  assign new_new_n29171__ = new_new_n29169__ & ~new_new_n29170__;
  assign new_new_n29172__ = ~new_new_n29167__ & new_new_n29171__;
  assign new_new_n29173__ = pi14 & new_new_n29163__;
  assign new_new_n29174__ = ~new_new_n29169__ & new_new_n29173__;
  assign new_new_n29175__ = ~new_new_n29166__ & ~new_new_n29174__;
  assign new_new_n29176__ = ~new_new_n29172__ & new_new_n29175__;
  assign new_new_n29177__ = ~new_new_n29160__ & ~new_new_n29176__;
  assign new_new_n29178__ = new_new_n29136__ & ~new_new_n29177__;
  assign new_new_n29179__ = ~new_new_n29136__ & new_new_n29177__;
  assign new_new_n29180__ = new_new_n6966__ & new_new_n27087__;
  assign new_new_n29181__ = ~new_new_n6958__ & new_new_n27582__;
  assign new_new_n29182__ = ~new_new_n6956__ & new_new_n26118__;
  assign new_new_n29183__ = new_new_n6967__ & ~new_new_n29182__;
  assign new_new_n29184__ = ~new_new_n6962__ & ~new_new_n27577__;
  assign new_new_n29185__ = ~new_new_n29180__ & new_new_n29184__;
  assign new_new_n29186__ = ~new_new_n29181__ & ~new_new_n29183__;
  assign new_new_n29187__ = new_new_n29185__ & new_new_n29186__;
  assign new_new_n29188__ = ~new_new_n29179__ & ~new_new_n29187__;
  assign new_new_n29189__ = ~new_new_n29178__ & ~new_new_n29188__;
  assign new_new_n29190__ = ~new_new_n29120__ & ~new_new_n29189__;
  assign new_new_n29191__ = new_new_n29120__ & new_new_n29189__;
  assign new_new_n29192__ = ~new_new_n6963__ & ~new_new_n28122__;
  assign new_new_n29193__ = pi17 & ~new_new_n28123__;
  assign new_new_n29194__ = ~new_new_n29192__ & new_new_n29193__;
  assign new_new_n29195__ = ~new_new_n28133__ & ~new_new_n29194__;
  assign new_new_n29196__ = new_new_n28133__ & new_new_n29194__;
  assign new_new_n29197__ = ~new_new_n29195__ & ~new_new_n29196__;
  assign new_new_n29198__ = ~new_new_n29191__ & new_new_n29197__;
  assign new_new_n29199__ = ~new_new_n29190__ & ~new_new_n29198__;
  assign new_new_n29200__ = ~new_new_n29103__ & ~new_new_n29199__;
  assign new_new_n29201__ = ~new_new_n28121__ & new_new_n28150__;
  assign new_new_n29202__ = ~new_new_n28151__ & ~new_new_n29201__;
  assign new_new_n29203__ = ~new_new_n29200__ & new_new_n29202__;
  assign new_new_n29204__ = ~new_new_n28121__ & ~new_new_n28150__;
  assign new_new_n29205__ = new_new_n28135__ & ~new_new_n29204__;
  assign new_new_n29206__ = ~new_new_n29199__ & ~new_new_n29205__;
  assign new_new_n29207__ = new_new_n29103__ & ~new_new_n29206__;
  assign new_new_n29208__ = ~new_new_n29203__ & ~new_new_n29207__;
  assign new_new_n29209__ = new_new_n29088__ & new_new_n29208__;
  assign new_new_n29210__ = ~new_new_n29088__ & ~new_new_n29208__;
  assign new_new_n29211__ = new_new_n28119__ & ~new_new_n28151__;
  assign new_new_n29212__ = ~new_new_n28152__ & ~new_new_n29211__;
  assign new_new_n29213__ = ~new_new_n29210__ & ~new_new_n29212__;
  assign new_new_n29214__ = ~new_new_n29209__ & ~new_new_n29213__;
  assign new_new_n29215__ = new_new_n6991__ & ~new_new_n27033__;
  assign new_new_n29216__ = new_new_n6985__ & new_new_n27111__;
  assign new_new_n29217__ = ~new_new_n29215__ & ~new_new_n29216__;
  assign new_new_n29218__ = new_new_n6994__ & ~new_new_n27021__;
  assign new_new_n29219__ = new_new_n27796__ & new_new_n29218__;
  assign new_new_n29220__ = new_new_n29217__ & ~new_new_n29219__;
  assign new_new_n29221__ = pi14 & ~new_new_n29220__;
  assign new_new_n29222__ = ~new_new_n27021__ & ~new_new_n27795__;
  assign new_new_n29223__ = pi13 & ~new_new_n29222__;
  assign new_new_n29224__ = new_new_n27021__ & new_new_n27796__;
  assign new_new_n29225__ = ~pi13 & ~new_new_n29224__;
  assign new_new_n29226__ = new_new_n6994__ & ~new_new_n29223__;
  assign new_new_n29227__ = ~new_new_n29225__ & new_new_n29226__;
  assign new_new_n29228__ = new_new_n27021__ & ~new_new_n27796__;
  assign new_new_n29229__ = new_new_n6994__ & ~new_new_n29228__;
  assign new_new_n29230__ = ~pi14 & new_new_n29217__;
  assign new_new_n29231__ = ~new_new_n29229__ & new_new_n29230__;
  assign new_new_n29232__ = ~new_new_n29221__ & ~new_new_n29227__;
  assign new_new_n29233__ = ~new_new_n29231__ & new_new_n29232__;
  assign new_new_n29234__ = new_new_n29214__ & new_new_n29233__;
  assign new_new_n29235__ = new_new_n29071__ & ~new_new_n29234__;
  assign new_new_n29236__ = ~new_new_n29214__ & ~new_new_n29233__;
  assign new_new_n29237__ = ~new_new_n29235__ & ~new_new_n29236__;
  assign new_new_n29238__ = new_new_n29069__ & ~new_new_n29237__;
  assign new_new_n29239__ = ~new_new_n29069__ & new_new_n29237__;
  assign new_new_n29240__ = new_new_n6991__ & new_new_n27111__;
  assign new_new_n29241__ = new_new_n6985__ & ~new_new_n27021__;
  assign new_new_n29242__ = ~new_new_n10772__ & new_new_n27029__;
  assign new_new_n29243__ = new_new_n10772__ & ~new_new_n27764__;
  assign new_new_n29244__ = new_new_n6994__ & ~new_new_n29242__;
  assign new_new_n29245__ = ~new_new_n29243__ & new_new_n29244__;
  assign new_new_n29246__ = ~new_new_n29240__ & ~new_new_n29241__;
  assign new_new_n29247__ = ~new_new_n29245__ & new_new_n29246__;
  assign new_new_n29248__ = ~pi14 & ~new_new_n29247__;
  assign new_new_n29249__ = pi14 & new_new_n29247__;
  assign new_new_n29250__ = ~new_new_n29248__ & ~new_new_n29249__;
  assign new_new_n29251__ = ~new_new_n29239__ & new_new_n29250__;
  assign new_new_n29252__ = ~new_new_n29238__ & ~new_new_n29251__;
  assign new_new_n29253__ = ~new_new_n29065__ & ~new_new_n29252__;
  assign new_new_n29254__ = ~new_new_n29064__ & ~new_new_n29253__;
  assign new_new_n29255__ = ~new_new_n29042__ & new_new_n29254__;
  assign new_new_n29256__ = new_new_n29042__ & ~new_new_n29254__;
  assign new_new_n29257__ = new_new_n28207__ & ~new_new_n29256__;
  assign new_new_n29258__ = ~new_new_n29255__ & ~new_new_n29257__;
  assign new_new_n29259__ = ~new_new_n29025__ & ~new_new_n29258__;
  assign new_new_n29260__ = ~new_new_n29024__ & ~new_new_n29259__;
  assign new_new_n29261__ = ~new_new_n28224__ & ~new_new_n28225__;
  assign new_new_n29262__ = ~new_new_n28229__ & new_new_n29261__;
  assign new_new_n29263__ = new_new_n28229__ & ~new_new_n29261__;
  assign new_new_n29264__ = ~new_new_n29262__ & ~new_new_n29263__;
  assign new_new_n29265__ = new_new_n29260__ & new_new_n29264__;
  assign new_new_n29266__ = ~new_new_n29260__ & ~new_new_n29264__;
  assign new_new_n29267__ = ~new_new_n29265__ & ~new_new_n29266__;
  assign new_new_n29268__ = ~new_new_n29002__ & ~new_new_n29267__;
  assign new_new_n29269__ = ~new_new_n29260__ & new_new_n29264__;
  assign new_new_n29270__ = ~new_new_n29268__ & ~new_new_n29269__;
  assign new_new_n29271__ = ~pi13 & new_new_n27477__;
  assign new_new_n29272__ = ~pi14 & ~new_new_n27477__;
  assign new_new_n29273__ = ~new_new_n29271__ & ~new_new_n29272__;
  assign new_new_n29274__ = ~new_new_n27152__ & new_new_n29273__;
  assign new_new_n29275__ = new_new_n27152__ & ~new_new_n29273__;
  assign new_new_n29276__ = new_new_n6994__ & ~new_new_n29274__;
  assign new_new_n29277__ = ~new_new_n29275__ & new_new_n29276__;
  assign new_new_n29278__ = new_new_n20894__ & ~new_new_n26937__;
  assign new_new_n29279__ = new_new_n19823__ & new_new_n26971__;
  assign new_new_n29280__ = new_new_n19825__ & ~new_new_n26937__;
  assign new_new_n29281__ = ~pi12 & new_new_n29018__;
  assign new_new_n29282__ = pi14 & ~new_new_n29281__;
  assign new_new_n29283__ = ~new_new_n29280__ & new_new_n29282__;
  assign new_new_n29284__ = ~new_new_n6994__ & ~new_new_n29279__;
  assign new_new_n29285__ = ~new_new_n29278__ & new_new_n29284__;
  assign new_new_n29286__ = ~new_new_n29283__ & new_new_n29285__;
  assign new_new_n29287__ = ~new_new_n29277__ & ~new_new_n29286__;
  assign new_new_n29288__ = new_new_n29270__ & ~new_new_n29287__;
  assign new_new_n29289__ = ~new_new_n29270__ & new_new_n29287__;
  assign new_new_n29290__ = ~new_new_n28232__ & ~new_new_n28233__;
  assign new_new_n29291__ = new_new_n28245__ & new_new_n29290__;
  assign new_new_n29292__ = ~new_new_n28245__ & ~new_new_n29290__;
  assign new_new_n29293__ = ~new_new_n29291__ & ~new_new_n29292__;
  assign new_new_n29294__ = ~new_new_n29289__ & ~new_new_n29293__;
  assign new_new_n29295__ = ~new_new_n29288__ & ~new_new_n29294__;
  assign new_new_n29296__ = new_new_n28985__ & new_new_n29295__;
  assign new_new_n29297__ = ~new_new_n28985__ & ~new_new_n29295__;
  assign new_new_n29298__ = ~new_new_n28252__ & ~new_new_n28253__;
  assign new_new_n29299__ = ~new_new_n28289__ & new_new_n29298__;
  assign new_new_n29300__ = new_new_n28289__ & ~new_new_n29298__;
  assign new_new_n29301__ = ~new_new_n29299__ & ~new_new_n29300__;
  assign new_new_n29302__ = ~new_new_n29297__ & ~new_new_n29301__;
  assign new_new_n29303__ = ~new_new_n29296__ & ~new_new_n29302__;
  assign new_new_n29304__ = ~new_new_n28013__ & ~new_new_n28014__;
  assign new_new_n29305__ = new_new_n28291__ & ~new_new_n29304__;
  assign new_new_n29306__ = ~new_new_n28291__ & new_new_n29304__;
  assign new_new_n29307__ = ~new_new_n29305__ & ~new_new_n29306__;
  assign new_new_n29308__ = ~new_new_n29303__ & ~new_new_n29307__;
  assign new_new_n29309__ = new_new_n29303__ & new_new_n29307__;
  assign new_new_n29310__ = new_new_n6991__ & new_new_n27152__;
  assign new_new_n29311__ = new_new_n6985__ & ~new_new_n26941__;
  assign new_new_n29312__ = ~new_new_n29310__ & ~new_new_n29311__;
  assign new_new_n29313__ = new_new_n6994__ & new_new_n26928__;
  assign new_new_n29314__ = new_new_n27488__ & new_new_n29313__;
  assign new_new_n29315__ = new_new_n29312__ & ~new_new_n29314__;
  assign new_new_n29316__ = ~pi14 & ~new_new_n29315__;
  assign new_new_n29317__ = pi13 & new_new_n26928__;
  assign new_new_n29318__ = ~new_new_n26928__ & ~new_new_n27488__;
  assign new_new_n29319__ = new_new_n6994__ & ~new_new_n29318__;
  assign new_new_n29320__ = ~pi13 & new_new_n27488__;
  assign new_new_n29321__ = ~new_new_n29317__ & ~new_new_n29320__;
  assign new_new_n29322__ = new_new_n29319__ & new_new_n29321__;
  assign new_new_n29323__ = pi14 & new_new_n29312__;
  assign new_new_n29324__ = ~new_new_n29319__ & new_new_n29323__;
  assign new_new_n29325__ = ~new_new_n29316__ & ~new_new_n29322__;
  assign new_new_n29326__ = ~new_new_n29324__ & new_new_n29325__;
  assign new_new_n29327__ = ~new_new_n29309__ & ~new_new_n29326__;
  assign new_new_n29328__ = ~new_new_n29308__ & ~new_new_n29327__;
  assign new_new_n29329__ = ~new_new_n28969__ & ~new_new_n29328__;
  assign new_new_n29330__ = ~new_new_n28968__ & ~new_new_n29329__;
  assign new_new_n29331__ = new_new_n28946__ & ~new_new_n29330__;
  assign new_new_n29332__ = ~new_new_n28946__ & new_new_n29330__;
  assign new_new_n29333__ = new_new_n6991__ & new_new_n26928__;
  assign new_new_n29334__ = new_new_n6985__ & new_new_n26917__;
  assign new_new_n29335__ = ~new_new_n29333__ & ~new_new_n29334__;
  assign new_new_n29336__ = new_new_n6994__ & ~new_new_n27168__;
  assign new_new_n29337__ = ~new_new_n28799__ & new_new_n29336__;
  assign new_new_n29338__ = new_new_n29335__ & ~new_new_n29337__;
  assign new_new_n29339__ = ~pi14 & ~new_new_n29338__;
  assign new_new_n29340__ = pi13 & ~new_new_n27168__;
  assign new_new_n29341__ = new_new_n27168__ & new_new_n28799__;
  assign new_new_n29342__ = new_new_n6994__ & ~new_new_n29341__;
  assign new_new_n29343__ = ~pi13 & ~new_new_n28799__;
  assign new_new_n29344__ = ~new_new_n29340__ & ~new_new_n29343__;
  assign new_new_n29345__ = new_new_n29342__ & new_new_n29344__;
  assign new_new_n29346__ = pi14 & new_new_n29335__;
  assign new_new_n29347__ = ~new_new_n29342__ & new_new_n29346__;
  assign new_new_n29348__ = ~new_new_n29339__ & ~new_new_n29345__;
  assign new_new_n29349__ = ~new_new_n29347__ & new_new_n29348__;
  assign new_new_n29350__ = ~new_new_n29332__ & ~new_new_n29349__;
  assign new_new_n29351__ = ~new_new_n29331__ & ~new_new_n29350__;
  assign new_new_n29352__ = ~new_new_n28511__ & ~new_new_n28512__;
  assign new_new_n29353__ = ~new_new_n28657__ & new_new_n29352__;
  assign new_new_n29354__ = new_new_n28657__ & ~new_new_n29352__;
  assign new_new_n29355__ = ~new_new_n29353__ & ~new_new_n29354__;
  assign new_new_n29356__ = ~new_new_n29351__ & ~new_new_n29355__;
  assign new_new_n29357__ = new_new_n29351__ & new_new_n29355__;
  assign new_new_n29358__ = new_new_n6991__ & new_new_n26917__;
  assign new_new_n29359__ = new_new_n6985__ & ~new_new_n27168__;
  assign new_new_n29360__ = ~new_new_n10772__ & ~new_new_n26922__;
  assign new_new_n29361__ = ~new_new_n27163__ & ~new_new_n27170__;
  assign new_new_n29362__ = new_new_n26917__ & ~new_new_n28795__;
  assign new_new_n29363__ = ~new_new_n28794__ & ~new_new_n29362__;
  assign new_new_n29364__ = new_new_n29361__ & ~new_new_n29363__;
  assign new_new_n29365__ = ~new_new_n29361__ & new_new_n29363__;
  assign new_new_n29366__ = ~new_new_n29364__ & ~new_new_n29365__;
  assign new_new_n29367__ = new_new_n10772__ & new_new_n29366__;
  assign new_new_n29368__ = new_new_n6994__ & ~new_new_n29360__;
  assign new_new_n29369__ = ~new_new_n29367__ & new_new_n29368__;
  assign new_new_n29370__ = ~new_new_n29358__ & ~new_new_n29359__;
  assign new_new_n29371__ = ~new_new_n29369__ & new_new_n29370__;
  assign new_new_n29372__ = ~pi14 & ~new_new_n29371__;
  assign new_new_n29373__ = pi14 & new_new_n29371__;
  assign new_new_n29374__ = ~new_new_n29372__ & ~new_new_n29373__;
  assign new_new_n29375__ = ~new_new_n29357__ & ~new_new_n29374__;
  assign new_new_n29376__ = ~new_new_n29356__ & ~new_new_n29375__;
  assign new_new_n29377__ = new_new_n28942__ & ~new_new_n29376__;
  assign new_new_n29378__ = ~new_new_n28942__ & new_new_n29376__;
  assign new_new_n29379__ = new_new_n6991__ & ~new_new_n27168__;
  assign new_new_n29380__ = new_new_n6985__ & new_new_n26922__;
  assign new_new_n29381__ = ~new_new_n10772__ & new_new_n26888__;
  assign new_new_n29382__ = new_new_n10772__ & ~new_new_n27180__;
  assign new_new_n29383__ = new_new_n6994__ & ~new_new_n29381__;
  assign new_new_n29384__ = ~new_new_n29382__ & new_new_n29383__;
  assign new_new_n29385__ = ~new_new_n29379__ & ~new_new_n29380__;
  assign new_new_n29386__ = ~new_new_n29384__ & new_new_n29385__;
  assign new_new_n29387__ = ~pi14 & ~new_new_n29386__;
  assign new_new_n29388__ = pi14 & new_new_n29386__;
  assign new_new_n29389__ = ~new_new_n29387__ & ~new_new_n29388__;
  assign new_new_n29390__ = ~new_new_n29378__ & ~new_new_n29389__;
  assign new_new_n29391__ = ~new_new_n29377__ & ~new_new_n29390__;
  assign new_new_n29392__ = new_new_n28940__ & ~new_new_n29391__;
  assign new_new_n29393__ = ~new_new_n28940__ & new_new_n29391__;
  assign new_new_n29394__ = ~new_new_n29392__ & ~new_new_n29393__;
  assign new_new_n29395__ = new_new_n8474__ & new_new_n26847__;
  assign new_new_n29396__ = ~new_new_n8479__ & ~new_new_n26854__;
  assign new_new_n29397__ = ~new_new_n27187__ & ~new_new_n27189__;
  assign new_new_n29398__ = new_new_n26847__ & new_new_n29397__;
  assign new_new_n29399__ = ~new_new_n26847__ & ~new_new_n29397__;
  assign new_new_n29400__ = ~new_new_n29398__ & ~new_new_n29399__;
  assign new_new_n29401__ = new_new_n8470__ & ~new_new_n29400__;
  assign new_new_n29402__ = ~new_new_n29395__ & ~new_new_n29396__;
  assign new_new_n29403__ = ~new_new_n29401__ & new_new_n29402__;
  assign new_new_n29404__ = new_new_n8469__ & ~new_new_n26823__;
  assign new_new_n29405__ = pi11 & ~new_new_n29404__;
  assign new_new_n29406__ = new_new_n11368__ & ~new_new_n26823__;
  assign new_new_n29407__ = ~new_new_n29405__ & ~new_new_n29406__;
  assign new_new_n29408__ = new_new_n29403__ & ~new_new_n29407__;
  assign new_new_n29409__ = ~pi11 & ~new_new_n29403__;
  assign new_new_n29410__ = ~new_new_n29408__ & ~new_new_n29409__;
  assign new_new_n29411__ = new_new_n8474__ & ~new_new_n26854__;
  assign new_new_n29412__ = ~new_new_n8479__ & ~new_new_n26888__;
  assign new_new_n29413__ = new_new_n26855__ & new_new_n27420__;
  assign new_new_n29414__ = ~new_new_n26855__ & new_new_n27184__;
  assign new_new_n29415__ = ~new_new_n26854__ & new_new_n27175__;
  assign new_new_n29416__ = ~new_new_n26889__ & ~new_new_n29415__;
  assign new_new_n29417__ = ~new_new_n26855__ & ~new_new_n27180__;
  assign new_new_n29418__ = ~new_new_n29416__ & new_new_n29417__;
  assign new_new_n29419__ = ~new_new_n26854__ & new_new_n26888__;
  assign new_new_n29420__ = ~new_new_n27419__ & ~new_new_n29419__;
  assign new_new_n29421__ = ~new_new_n26847__ & new_new_n29420__;
  assign new_new_n29422__ = ~new_new_n29414__ & ~new_new_n29421__;
  assign new_new_n29423__ = ~new_new_n29418__ & new_new_n29422__;
  assign new_new_n29424__ = ~new_new_n29413__ & new_new_n29423__;
  assign new_new_n29425__ = new_new_n8470__ & new_new_n29424__;
  assign new_new_n29426__ = ~new_new_n29411__ & ~new_new_n29412__;
  assign new_new_n29427__ = ~new_new_n29425__ & new_new_n29426__;
  assign new_new_n29428__ = new_new_n8469__ & new_new_n26847__;
  assign new_new_n29429__ = ~pi11 & ~new_new_n29428__;
  assign new_new_n29430__ = new_new_n11530__ & new_new_n26847__;
  assign new_new_n29431__ = ~new_new_n29429__ & ~new_new_n29430__;
  assign new_new_n29432__ = new_new_n29427__ & ~new_new_n29431__;
  assign new_new_n29433__ = pi11 & ~new_new_n29427__;
  assign new_new_n29434__ = ~new_new_n29432__ & ~new_new_n29433__;
  assign new_new_n29435__ = new_new_n8858__ & ~new_new_n26854__;
  assign new_new_n29436__ = ~new_new_n8479__ & new_new_n26922__;
  assign new_new_n29437__ = new_new_n8474__ & ~new_new_n26888__;
  assign new_new_n29438__ = ~new_new_n29436__ & ~new_new_n29437__;
  assign new_new_n29439__ = ~new_new_n29435__ & new_new_n29438__;
  assign new_new_n29440__ = new_new_n8469__ & ~new_new_n27430__;
  assign new_new_n29441__ = pi11 & ~new_new_n29440__;
  assign new_new_n29442__ = new_new_n11530__ & ~new_new_n27430__;
  assign new_new_n29443__ = ~new_new_n29441__ & ~new_new_n29442__;
  assign new_new_n29444__ = new_new_n29439__ & ~new_new_n29443__;
  assign new_new_n29445__ = ~pi11 & ~new_new_n29439__;
  assign new_new_n29446__ = ~new_new_n29444__ & ~new_new_n29445__;
  assign new_new_n29447__ = new_new_n8470__ & ~new_new_n29366__;
  assign new_new_n29448__ = new_new_n8474__ & ~new_new_n27168__;
  assign new_new_n29449__ = ~new_new_n8479__ & new_new_n26917__;
  assign new_new_n29450__ = ~new_new_n29448__ & ~new_new_n29449__;
  assign new_new_n29451__ = ~new_new_n29447__ & new_new_n29450__;
  assign new_new_n29452__ = new_new_n8469__ & new_new_n26922__;
  assign new_new_n29453__ = pi11 & ~new_new_n29452__;
  assign new_new_n29454__ = new_new_n11368__ & new_new_n26922__;
  assign new_new_n29455__ = ~new_new_n29453__ & ~new_new_n29454__;
  assign new_new_n29456__ = new_new_n29451__ & ~new_new_n29455__;
  assign new_new_n29457__ = ~pi11 & ~new_new_n29451__;
  assign new_new_n29458__ = ~new_new_n29456__ & ~new_new_n29457__;
  assign new_new_n29459__ = ~new_new_n29296__ & ~new_new_n29297__;
  assign new_new_n29460__ = ~new_new_n29301__ & new_new_n29459__;
  assign new_new_n29461__ = new_new_n29301__ & ~new_new_n29459__;
  assign new_new_n29462__ = ~new_new_n29460__ & ~new_new_n29461__;
  assign new_new_n29463__ = ~new_new_n29288__ & ~new_new_n29289__;
  assign new_new_n29464__ = ~new_new_n29293__ & new_new_n29463__;
  assign new_new_n29465__ = new_new_n29293__ & ~new_new_n29463__;
  assign new_new_n29466__ = ~new_new_n29464__ & ~new_new_n29465__;
  assign new_new_n29467__ = new_new_n8858__ & new_new_n26928__;
  assign new_new_n29468__ = new_new_n8474__ & ~new_new_n26941__;
  assign new_new_n29469__ = ~new_new_n8479__ & new_new_n27152__;
  assign new_new_n29470__ = new_new_n8470__ & new_new_n27488__;
  assign new_new_n29471__ = ~new_new_n29468__ & ~new_new_n29469__;
  assign new_new_n29472__ = ~new_new_n29467__ & new_new_n29471__;
  assign new_new_n29473__ = ~new_new_n29470__ & new_new_n29472__;
  assign new_new_n29474__ = pi11 & ~new_new_n29473__;
  assign new_new_n29475__ = ~pi11 & new_new_n29473__;
  assign new_new_n29476__ = ~new_new_n29474__ & ~new_new_n29475__;
  assign new_new_n29477__ = new_new_n8858__ & ~new_new_n26941__;
  assign new_new_n29478__ = ~new_new_n8479__ & ~new_new_n26937__;
  assign new_new_n29479__ = new_new_n8474__ & new_new_n27152__;
  assign new_new_n29480__ = ~new_new_n29477__ & ~new_new_n29478__;
  assign new_new_n29481__ = ~new_new_n29479__ & new_new_n29480__;
  assign new_new_n29482__ = new_new_n8469__ & ~new_new_n27502__;
  assign new_new_n29483__ = ~pi11 & ~new_new_n29482__;
  assign new_new_n29484__ = new_new_n11368__ & ~new_new_n27502__;
  assign new_new_n29485__ = ~new_new_n29483__ & ~new_new_n29484__;
  assign new_new_n29486__ = new_new_n29481__ & ~new_new_n29485__;
  assign new_new_n29487__ = pi11 & ~new_new_n29481__;
  assign new_new_n29488__ = ~new_new_n29486__ & ~new_new_n29487__;
  assign new_new_n29489__ = new_new_n8858__ & new_new_n27152__;
  assign new_new_n29490__ = ~new_new_n8479__ & new_new_n26971__;
  assign new_new_n29491__ = new_new_n8474__ & ~new_new_n26937__;
  assign new_new_n29492__ = new_new_n8470__ & ~new_new_n28666__;
  assign new_new_n29493__ = ~new_new_n29490__ & ~new_new_n29491__;
  assign new_new_n29494__ = ~new_new_n29489__ & new_new_n29493__;
  assign new_new_n29495__ = ~new_new_n29492__ & new_new_n29494__;
  assign new_new_n29496__ = pi11 & ~new_new_n29495__;
  assign new_new_n29497__ = ~pi11 & new_new_n29495__;
  assign new_new_n29498__ = ~new_new_n29496__ & ~new_new_n29497__;
  assign new_new_n29499__ = ~new_new_n29255__ & ~new_new_n29256__;
  assign new_new_n29500__ = new_new_n28207__ & new_new_n29499__;
  assign new_new_n29501__ = ~new_new_n28207__ & ~new_new_n29499__;
  assign new_new_n29502__ = ~new_new_n29500__ & ~new_new_n29501__;
  assign new_new_n29503__ = ~new_new_n29498__ & ~new_new_n29502__;
  assign new_new_n29504__ = new_new_n29498__ & new_new_n29502__;
  assign new_new_n29505__ = ~new_new_n29064__ & ~new_new_n29065__;
  assign new_new_n29506__ = new_new_n29252__ & ~new_new_n29505__;
  assign new_new_n29507__ = ~new_new_n29252__ & new_new_n29505__;
  assign new_new_n29508__ = ~new_new_n29506__ & ~new_new_n29507__;
  assign new_new_n29509__ = new_new_n8474__ & ~new_new_n26978__;
  assign new_new_n29510__ = ~new_new_n8479__ & ~new_new_n27003__;
  assign new_new_n29511__ = new_new_n8470__ & new_new_n28277__;
  assign new_new_n29512__ = ~new_new_n29509__ & ~new_new_n29510__;
  assign new_new_n29513__ = ~new_new_n29511__ & new_new_n29512__;
  assign new_new_n29514__ = new_new_n8469__ & new_new_n26971__;
  assign new_new_n29515__ = ~pi11 & ~new_new_n29514__;
  assign new_new_n29516__ = new_new_n11530__ & new_new_n26971__;
  assign new_new_n29517__ = ~new_new_n29515__ & ~new_new_n29516__;
  assign new_new_n29518__ = new_new_n29513__ & ~new_new_n29517__;
  assign new_new_n29519__ = pi11 & ~new_new_n29513__;
  assign new_new_n29520__ = ~new_new_n29518__ & ~new_new_n29519__;
  assign new_new_n29521__ = new_new_n8858__ & ~new_new_n26978__;
  assign new_new_n29522__ = new_new_n8474__ & ~new_new_n27003__;
  assign new_new_n29523__ = new_new_n8470__ & new_new_n27986__;
  assign new_new_n29524__ = ~new_new_n29521__ & ~new_new_n29522__;
  assign new_new_n29525__ = ~new_new_n29523__ & new_new_n29524__;
  assign new_new_n29526__ = ~pi11 & ~new_new_n29525__;
  assign new_new_n29527__ = new_new_n8477__ & ~new_new_n27029__;
  assign new_new_n29528__ = pi11 & ~new_new_n29527__;
  assign new_new_n29529__ = new_new_n8855__ & ~new_new_n27029__;
  assign new_new_n29530__ = ~new_new_n29528__ & ~new_new_n29529__;
  assign new_new_n29531__ = new_new_n29525__ & ~new_new_n29530__;
  assign new_new_n29532__ = ~new_new_n29526__ & ~new_new_n29531__;
  assign new_new_n29533__ = new_new_n8474__ & ~new_new_n27029__;
  assign new_new_n29534__ = ~new_new_n8479__ & ~new_new_n27021__;
  assign new_new_n29535__ = new_new_n8858__ & ~new_new_n27003__;
  assign new_new_n29536__ = ~new_new_n29533__ & ~new_new_n29534__;
  assign new_new_n29537__ = ~new_new_n29535__ & new_new_n29536__;
  assign new_new_n29538__ = new_new_n8469__ & new_new_n27962__;
  assign new_new_n29539__ = pi11 & ~new_new_n29538__;
  assign new_new_n29540__ = new_new_n11530__ & new_new_n27962__;
  assign new_new_n29541__ = ~new_new_n29539__ & ~new_new_n29540__;
  assign new_new_n29542__ = new_new_n29537__ & ~new_new_n29541__;
  assign new_new_n29543__ = ~pi11 & ~new_new_n29537__;
  assign new_new_n29544__ = ~new_new_n29542__ & ~new_new_n29543__;
  assign new_new_n29545__ = new_new_n29103__ & new_new_n29199__;
  assign new_new_n29546__ = ~new_new_n29200__ & ~new_new_n29545__;
  assign new_new_n29547__ = new_new_n29103__ & new_new_n29205__;
  assign new_new_n29548__ = ~new_new_n29202__ & ~new_new_n29547__;
  assign new_new_n29549__ = new_new_n29546__ & ~new_new_n29548__;
  assign new_new_n29550__ = ~new_new_n29202__ & ~new_new_n29205__;
  assign new_new_n29551__ = ~new_new_n29546__ & new_new_n29550__;
  assign new_new_n29552__ = ~new_new_n29549__ & ~new_new_n29551__;
  assign new_new_n29553__ = new_new_n8474__ & ~new_new_n27033__;
  assign new_new_n29554__ = ~new_new_n8479__ & ~new_new_n27054__;
  assign new_new_n29555__ = ~new_new_n29553__ & ~new_new_n29554__;
  assign new_new_n29556__ = new_new_n8469__ & new_new_n27687__;
  assign new_new_n29557__ = new_new_n29555__ & ~new_new_n29556__;
  assign new_new_n29558__ = pi11 & ~new_new_n29557__;
  assign new_new_n29559__ = new_new_n8469__ & ~new_new_n27691__;
  assign new_new_n29560__ = ~pi11 & ~new_new_n29559__;
  assign new_new_n29561__ = ~pi10 & new_new_n27111__;
  assign new_new_n29562__ = pi10 & ~new_new_n27111__;
  assign new_new_n29563__ = new_new_n8469__ & ~new_new_n29561__;
  assign new_new_n29564__ = ~new_new_n29562__ & new_new_n29563__;
  assign new_new_n29565__ = new_new_n27686__ & new_new_n29564__;
  assign new_new_n29566__ = ~new_new_n29560__ & ~new_new_n29565__;
  assign new_new_n29567__ = new_new_n29555__ & ~new_new_n29566__;
  assign new_new_n29568__ = ~new_new_n29558__ & ~new_new_n29567__;
  assign new_new_n29569__ = ~new_new_n8479__ & new_new_n27041__;
  assign new_new_n29570__ = new_new_n8474__ & ~new_new_n27054__;
  assign new_new_n29571__ = ~new_new_n29569__ & ~new_new_n29570__;
  assign new_new_n29572__ = new_new_n8469__ & new_new_n27545__;
  assign new_new_n29573__ = new_new_n29571__ & ~new_new_n29572__;
  assign new_new_n29574__ = pi11 & ~new_new_n29573__;
  assign new_new_n29575__ = new_new_n8469__ & ~new_new_n27535__;
  assign new_new_n29576__ = ~pi11 & ~new_new_n29575__;
  assign new_new_n29577__ = pi10 & ~new_new_n27033__;
  assign new_new_n29578__ = ~pi10 & new_new_n27033__;
  assign new_new_n29579__ = ~new_new_n29577__ & ~new_new_n29578__;
  assign new_new_n29580__ = new_new_n8469__ & ~new_new_n29579__;
  assign new_new_n29581__ = ~new_new_n27102__ & new_new_n29580__;
  assign new_new_n29582__ = ~new_new_n29576__ & ~new_new_n29581__;
  assign new_new_n29583__ = new_new_n29571__ & ~new_new_n29582__;
  assign new_new_n29584__ = ~new_new_n29574__ & ~new_new_n29583__;
  assign new_new_n29585__ = ~new_new_n29153__ & ~new_new_n29157__;
  assign new_new_n29586__ = ~new_new_n29158__ & ~new_new_n29585__;
  assign new_new_n29587__ = new_new_n8474__ & new_new_n27059__;
  assign new_new_n29588__ = ~new_new_n8468__ & new_new_n28443__;
  assign new_new_n29589__ = ~new_new_n28442__ & ~new_new_n29588__;
  assign new_new_n29590__ = new_new_n8469__ & ~new_new_n29589__;
  assign new_new_n29591__ = new_new_n8858__ & ~new_new_n27071__;
  assign new_new_n29592__ = ~new_new_n29587__ & ~new_new_n29591__;
  assign new_new_n29593__ = ~new_new_n29590__ & new_new_n29592__;
  assign new_new_n29594__ = ~pi11 & ~new_new_n29593__;
  assign new_new_n29595__ = new_new_n8477__ & new_new_n26118__;
  assign new_new_n29596__ = pi11 & ~new_new_n29595__;
  assign new_new_n29597__ = new_new_n8855__ & new_new_n26118__;
  assign new_new_n29598__ = ~new_new_n29596__ & ~new_new_n29597__;
  assign new_new_n29599__ = new_new_n29593__ & ~new_new_n29598__;
  assign new_new_n29600__ = ~new_new_n29594__ & ~new_new_n29599__;
  assign new_new_n29601__ = new_new_n6994__ & ~new_new_n27075__;
  assign new_new_n29602__ = ~new_new_n23470__ & ~new_new_n27577__;
  assign new_new_n29603__ = new_new_n8858__ & new_new_n27059__;
  assign new_new_n29604__ = ~new_new_n8468__ & new_new_n27846__;
  assign new_new_n29605__ = ~new_new_n28718__ & ~new_new_n29604__;
  assign new_new_n29606__ = new_new_n8469__ & ~new_new_n29605__;
  assign new_new_n29607__ = new_new_n8469__ & new_new_n27059__;
  assign new_new_n29608__ = new_new_n8479__ & ~new_new_n29607__;
  assign new_new_n29609__ = ~new_new_n27075__ & ~new_new_n29608__;
  assign new_new_n29610__ = ~new_new_n29603__ & ~new_new_n29609__;
  assign new_new_n29611__ = ~new_new_n29606__ & new_new_n29610__;
  assign new_new_n29612__ = pi11 & ~new_new_n29602__;
  assign new_new_n29613__ = new_new_n29611__ & new_new_n29612__;
  assign new_new_n29614__ = ~new_new_n29601__ & ~new_new_n29613__;
  assign new_new_n29615__ = ~new_new_n29600__ & ~new_new_n29614__;
  assign new_new_n29616__ = new_new_n6982__ & new_new_n27087__;
  assign new_new_n29617__ = ~new_new_n6994__ & new_new_n27582__;
  assign new_new_n29618__ = ~new_new_n6981__ & new_new_n26118__;
  assign new_new_n29619__ = new_new_n6984__ & ~new_new_n29618__;
  assign new_new_n29620__ = ~new_new_n23485__ & ~new_new_n27577__;
  assign new_new_n29621__ = ~new_new_n29616__ & new_new_n29620__;
  assign new_new_n29622__ = ~new_new_n29617__ & ~new_new_n29619__;
  assign new_new_n29623__ = new_new_n29621__ & new_new_n29622__;
  assign new_new_n29624__ = new_new_n29615__ & new_new_n29623__;
  assign new_new_n29625__ = ~new_new_n29615__ & ~new_new_n29623__;
  assign new_new_n29626__ = new_new_n8474__ & ~new_new_n27071__;
  assign new_new_n29627__ = ~new_new_n8479__ & new_new_n27059__;
  assign new_new_n29628__ = new_new_n8858__ & new_new_n27041__;
  assign new_new_n29629__ = ~new_new_n29626__ & ~new_new_n29627__;
  assign new_new_n29630__ = ~new_new_n29628__ & new_new_n29629__;
  assign new_new_n29631__ = new_new_n8470__ & new_new_n27567__;
  assign new_new_n29632__ = new_new_n29630__ & ~new_new_n29631__;
  assign new_new_n29633__ = ~pi11 & ~new_new_n29632__;
  assign new_new_n29634__ = pi11 & new_new_n29632__;
  assign new_new_n29635__ = ~new_new_n29633__ & ~new_new_n29634__;
  assign new_new_n29636__ = ~new_new_n29625__ & ~new_new_n29635__;
  assign new_new_n29637__ = ~new_new_n29624__ & ~new_new_n29636__;
  assign new_new_n29638__ = ~new_new_n29586__ & new_new_n29637__;
  assign new_new_n29639__ = new_new_n29586__ & ~new_new_n29637__;
  assign new_new_n29640__ = new_new_n8858__ & ~new_new_n27054__;
  assign new_new_n29641__ = ~new_new_n8479__ & ~new_new_n27071__;
  assign new_new_n29642__ = new_new_n8474__ & new_new_n27041__;
  assign new_new_n29643__ = new_new_n8470__ & ~new_new_n27094__;
  assign new_new_n29644__ = ~new_new_n29641__ & ~new_new_n29642__;
  assign new_new_n29645__ = ~new_new_n29640__ & new_new_n29644__;
  assign new_new_n29646__ = ~new_new_n29643__ & new_new_n29645__;
  assign new_new_n29647__ = pi11 & ~new_new_n29646__;
  assign new_new_n29648__ = ~pi11 & new_new_n29646__;
  assign new_new_n29649__ = ~new_new_n29647__ & ~new_new_n29648__;
  assign new_new_n29650__ = ~new_new_n29639__ & ~new_new_n29649__;
  assign new_new_n29651__ = ~new_new_n29638__ & ~new_new_n29650__;
  assign new_new_n29652__ = new_new_n29584__ & new_new_n29651__;
  assign new_new_n29653__ = ~new_new_n29584__ & ~new_new_n29651__;
  assign new_new_n29654__ = new_new_n29158__ & new_new_n29159__;
  assign new_new_n29655__ = ~new_new_n29176__ & ~new_new_n29654__;
  assign new_new_n29656__ = new_new_n29160__ & ~new_new_n29655__;
  assign new_new_n29657__ = ~new_new_n29160__ & new_new_n29655__;
  assign new_new_n29658__ = ~new_new_n29656__ & ~new_new_n29657__;
  assign new_new_n29659__ = ~new_new_n29653__ & new_new_n29658__;
  assign new_new_n29660__ = ~new_new_n29652__ & ~new_new_n29659__;
  assign new_new_n29661__ = new_new_n29568__ & ~new_new_n29660__;
  assign new_new_n29662__ = ~new_new_n29568__ & new_new_n29660__;
  assign new_new_n29663__ = ~new_new_n29178__ & ~new_new_n29179__;
  assign new_new_n29664__ = new_new_n29187__ & ~new_new_n29663__;
  assign new_new_n29665__ = ~new_new_n29187__ & new_new_n29663__;
  assign new_new_n29666__ = ~new_new_n29664__ & ~new_new_n29665__;
  assign new_new_n29667__ = ~new_new_n29662__ & ~new_new_n29666__;
  assign new_new_n29668__ = ~new_new_n29661__ & ~new_new_n29667__;
  assign new_new_n29669__ = new_new_n28133__ & ~new_new_n29194__;
  assign new_new_n29670__ = ~new_new_n28133__ & new_new_n29194__;
  assign new_new_n29671__ = ~new_new_n29669__ & ~new_new_n29670__;
  assign new_new_n29672__ = new_new_n29120__ & ~new_new_n29189__;
  assign new_new_n29673__ = ~new_new_n29120__ & new_new_n29189__;
  assign new_new_n29674__ = ~new_new_n29672__ & ~new_new_n29673__;
  assign new_new_n29675__ = new_new_n29671__ & new_new_n29674__;
  assign new_new_n29676__ = ~new_new_n29671__ & ~new_new_n29674__;
  assign new_new_n29677__ = ~new_new_n29675__ & ~new_new_n29676__;
  assign new_new_n29678__ = new_new_n29668__ & new_new_n29677__;
  assign new_new_n29679__ = ~new_new_n29668__ & ~new_new_n29677__;
  assign new_new_n29680__ = new_new_n8470__ & new_new_n27796__;
  assign new_new_n29681__ = new_new_n8474__ & new_new_n27111__;
  assign new_new_n29682__ = ~new_new_n8479__ & ~new_new_n27033__;
  assign new_new_n29683__ = new_new_n8858__ & ~new_new_n27021__;
  assign new_new_n29684__ = ~new_new_n29681__ & ~new_new_n29682__;
  assign new_new_n29685__ = ~new_new_n29683__ & new_new_n29684__;
  assign new_new_n29686__ = ~new_new_n29680__ & new_new_n29685__;
  assign new_new_n29687__ = pi11 & ~new_new_n29686__;
  assign new_new_n29688__ = ~pi11 & new_new_n29686__;
  assign new_new_n29689__ = ~new_new_n29687__ & ~new_new_n29688__;
  assign new_new_n29690__ = ~new_new_n29679__ & ~new_new_n29689__;
  assign new_new_n29691__ = ~new_new_n29678__ & ~new_new_n29690__;
  assign new_new_n29692__ = ~new_new_n29552__ & ~new_new_n29691__;
  assign new_new_n29693__ = new_new_n29552__ & new_new_n29691__;
  assign new_new_n29694__ = new_new_n8858__ & ~new_new_n27029__;
  assign new_new_n29695__ = new_new_n8474__ & ~new_new_n27021__;
  assign new_new_n29696__ = ~new_new_n8479__ & new_new_n27111__;
  assign new_new_n29697__ = new_new_n8470__ & new_new_n27764__;
  assign new_new_n29698__ = ~new_new_n29695__ & ~new_new_n29696__;
  assign new_new_n29699__ = ~new_new_n29694__ & new_new_n29698__;
  assign new_new_n29700__ = ~new_new_n29697__ & new_new_n29699__;
  assign new_new_n29701__ = ~pi11 & ~new_new_n29700__;
  assign new_new_n29702__ = pi11 & new_new_n29700__;
  assign new_new_n29703__ = ~new_new_n29701__ & ~new_new_n29702__;
  assign new_new_n29704__ = ~new_new_n29693__ & new_new_n29703__;
  assign new_new_n29705__ = ~new_new_n29692__ & ~new_new_n29704__;
  assign new_new_n29706__ = new_new_n29544__ & ~new_new_n29705__;
  assign new_new_n29707__ = ~new_new_n29544__ & new_new_n29705__;
  assign new_new_n29708__ = ~new_new_n29209__ & ~new_new_n29210__;
  assign new_new_n29709__ = ~new_new_n29212__ & new_new_n29708__;
  assign new_new_n29710__ = new_new_n29212__ & ~new_new_n29708__;
  assign new_new_n29711__ = ~new_new_n29709__ & ~new_new_n29710__;
  assign new_new_n29712__ = ~new_new_n29707__ & new_new_n29711__;
  assign new_new_n29713__ = ~new_new_n29706__ & ~new_new_n29712__;
  assign new_new_n29714__ = ~new_new_n29532__ & new_new_n29713__;
  assign new_new_n29715__ = new_new_n29532__ & ~new_new_n29713__;
  assign new_new_n29716__ = new_new_n29214__ & ~new_new_n29233__;
  assign new_new_n29717__ = ~new_new_n29214__ & new_new_n29233__;
  assign new_new_n29718__ = ~new_new_n29716__ & ~new_new_n29717__;
  assign new_new_n29719__ = new_new_n29071__ & ~new_new_n29718__;
  assign new_new_n29720__ = ~new_new_n29071__ & new_new_n29718__;
  assign new_new_n29721__ = ~new_new_n29719__ & ~new_new_n29720__;
  assign new_new_n29722__ = ~new_new_n29715__ & ~new_new_n29721__;
  assign new_new_n29723__ = ~new_new_n29714__ & ~new_new_n29722__;
  assign new_new_n29724__ = ~new_new_n29520__ & new_new_n29723__;
  assign new_new_n29725__ = new_new_n29520__ & ~new_new_n29723__;
  assign new_new_n29726__ = ~new_new_n29724__ & ~new_new_n29725__;
  assign new_new_n29727__ = ~new_new_n29238__ & ~new_new_n29239__;
  assign new_new_n29728__ = ~new_new_n29726__ & new_new_n29727__;
  assign new_new_n29729__ = new_new_n29726__ & ~new_new_n29727__;
  assign new_new_n29730__ = ~new_new_n29728__ & ~new_new_n29729__;
  assign new_new_n29731__ = new_new_n29250__ & ~new_new_n29730__;
  assign new_new_n29732__ = ~new_new_n29237__ & ~new_new_n29731__;
  assign new_new_n29733__ = ~new_new_n29250__ & new_new_n29730__;
  assign new_new_n29734__ = new_new_n29237__ & ~new_new_n29733__;
  assign new_new_n29735__ = new_new_n29069__ & ~new_new_n29732__;
  assign new_new_n29736__ = ~new_new_n29734__ & new_new_n29735__;
  assign new_new_n29737__ = ~new_new_n29237__ & ~new_new_n29733__;
  assign new_new_n29738__ = new_new_n29237__ & ~new_new_n29731__;
  assign new_new_n29739__ = ~new_new_n29069__ & ~new_new_n29737__;
  assign new_new_n29740__ = ~new_new_n29738__ & new_new_n29739__;
  assign new_new_n29741__ = ~new_new_n29724__ & ~new_new_n29736__;
  assign new_new_n29742__ = ~new_new_n29740__ & new_new_n29741__;
  assign new_new_n29743__ = new_new_n29508__ & ~new_new_n29742__;
  assign new_new_n29744__ = ~new_new_n29508__ & new_new_n29742__;
  assign new_new_n29745__ = new_new_n8858__ & ~new_new_n26937__;
  assign new_new_n29746__ = ~new_new_n8479__ & ~new_new_n26978__;
  assign new_new_n29747__ = new_new_n8474__ & new_new_n26971__;
  assign new_new_n29748__ = new_new_n8470__ & new_new_n28005__;
  assign new_new_n29749__ = ~new_new_n29746__ & ~new_new_n29747__;
  assign new_new_n29750__ = ~new_new_n29745__ & new_new_n29749__;
  assign new_new_n29751__ = ~new_new_n29748__ & new_new_n29750__;
  assign new_new_n29752__ = pi11 & ~new_new_n29751__;
  assign new_new_n29753__ = ~pi11 & new_new_n29751__;
  assign new_new_n29754__ = ~new_new_n29752__ & ~new_new_n29753__;
  assign new_new_n29755__ = ~new_new_n29744__ & ~new_new_n29754__;
  assign new_new_n29756__ = ~new_new_n29743__ & ~new_new_n29755__;
  assign new_new_n29757__ = ~new_new_n29504__ & ~new_new_n29756__;
  assign new_new_n29758__ = ~new_new_n29503__ & ~new_new_n29757__;
  assign new_new_n29759__ = ~new_new_n29488__ & ~new_new_n29758__;
  assign new_new_n29760__ = new_new_n29488__ & new_new_n29758__;
  assign new_new_n29761__ = ~new_new_n29024__ & ~new_new_n29025__;
  assign new_new_n29762__ = ~new_new_n29258__ & new_new_n29761__;
  assign new_new_n29763__ = new_new_n29258__ & ~new_new_n29761__;
  assign new_new_n29764__ = ~new_new_n29762__ & ~new_new_n29763__;
  assign new_new_n29765__ = ~new_new_n29760__ & ~new_new_n29764__;
  assign new_new_n29766__ = ~new_new_n29759__ & ~new_new_n29765__;
  assign new_new_n29767__ = ~new_new_n29476__ & ~new_new_n29766__;
  assign new_new_n29768__ = new_new_n29476__ & new_new_n29766__;
  assign new_new_n29769__ = new_new_n29002__ & new_new_n29267__;
  assign new_new_n29770__ = ~new_new_n29268__ & ~new_new_n29769__;
  assign new_new_n29771__ = ~new_new_n29768__ & ~new_new_n29770__;
  assign new_new_n29772__ = ~new_new_n29767__ & ~new_new_n29771__;
  assign new_new_n29773__ = ~new_new_n29466__ & new_new_n29772__;
  assign new_new_n29774__ = new_new_n29466__ & ~new_new_n29772__;
  assign new_new_n29775__ = new_new_n8858__ & new_new_n26917__;
  assign new_new_n29776__ = ~new_new_n8479__ & ~new_new_n26941__;
  assign new_new_n29777__ = new_new_n8474__ & new_new_n26928__;
  assign new_new_n29778__ = new_new_n8470__ & ~new_new_n27462__;
  assign new_new_n29779__ = ~new_new_n29776__ & ~new_new_n29777__;
  assign new_new_n29780__ = ~new_new_n29775__ & new_new_n29779__;
  assign new_new_n29781__ = ~new_new_n29778__ & new_new_n29780__;
  assign new_new_n29782__ = pi11 & ~new_new_n29781__;
  assign new_new_n29783__ = ~pi11 & new_new_n29781__;
  assign new_new_n29784__ = ~new_new_n29782__ & ~new_new_n29783__;
  assign new_new_n29785__ = ~new_new_n29774__ & new_new_n29784__;
  assign new_new_n29786__ = ~new_new_n29773__ & ~new_new_n29785__;
  assign new_new_n29787__ = ~new_new_n29462__ & new_new_n29786__;
  assign new_new_n29788__ = new_new_n29462__ & ~new_new_n29786__;
  assign new_new_n29789__ = new_new_n8474__ & new_new_n26917__;
  assign new_new_n29790__ = new_new_n8858__ & ~new_new_n27168__;
  assign new_new_n29791__ = ~new_new_n8479__ & new_new_n26928__;
  assign new_new_n29792__ = new_new_n8470__ & ~new_new_n28799__;
  assign new_new_n29793__ = ~new_new_n29790__ & ~new_new_n29791__;
  assign new_new_n29794__ = ~new_new_n29789__ & new_new_n29793__;
  assign new_new_n29795__ = ~new_new_n29792__ & new_new_n29794__;
  assign new_new_n29796__ = pi11 & ~new_new_n29795__;
  assign new_new_n29797__ = ~pi11 & new_new_n29795__;
  assign new_new_n29798__ = ~new_new_n29796__ & ~new_new_n29797__;
  assign new_new_n29799__ = ~new_new_n29788__ & ~new_new_n29798__;
  assign new_new_n29800__ = ~new_new_n29787__ & ~new_new_n29799__;
  assign new_new_n29801__ = ~new_new_n29458__ & new_new_n29800__;
  assign new_new_n29802__ = new_new_n29458__ & ~new_new_n29800__;
  assign new_new_n29803__ = ~new_new_n29308__ & ~new_new_n29309__;
  assign new_new_n29804__ = new_new_n29326__ & ~new_new_n29803__;
  assign new_new_n29805__ = ~new_new_n29326__ & new_new_n29803__;
  assign new_new_n29806__ = ~new_new_n29804__ & ~new_new_n29805__;
  assign new_new_n29807__ = ~new_new_n29802__ & new_new_n29806__;
  assign new_new_n29808__ = ~new_new_n29801__ & ~new_new_n29807__;
  assign new_new_n29809__ = ~new_new_n28968__ & ~new_new_n28969__;
  assign new_new_n29810__ = new_new_n29328__ & ~new_new_n29809__;
  assign new_new_n29811__ = ~new_new_n29328__ & new_new_n29809__;
  assign new_new_n29812__ = ~new_new_n29810__ & ~new_new_n29811__;
  assign new_new_n29813__ = new_new_n29808__ & ~new_new_n29812__;
  assign new_new_n29814__ = ~new_new_n29808__ & new_new_n29812__;
  assign new_new_n29815__ = new_new_n8474__ & new_new_n26922__;
  assign new_new_n29816__ = ~new_new_n8479__ & ~new_new_n27168__;
  assign new_new_n29817__ = new_new_n8858__ & ~new_new_n26888__;
  assign new_new_n29818__ = ~new_new_n29815__ & ~new_new_n29816__;
  assign new_new_n29819__ = ~new_new_n29817__ & new_new_n29818__;
  assign new_new_n29820__ = new_new_n8469__ & new_new_n27180__;
  assign new_new_n29821__ = ~pi11 & ~new_new_n29820__;
  assign new_new_n29822__ = new_new_n11368__ & new_new_n27180__;
  assign new_new_n29823__ = ~new_new_n29821__ & ~new_new_n29822__;
  assign new_new_n29824__ = new_new_n29819__ & ~new_new_n29823__;
  assign new_new_n29825__ = pi11 & ~new_new_n29819__;
  assign new_new_n29826__ = ~new_new_n29824__ & ~new_new_n29825__;
  assign new_new_n29827__ = ~new_new_n29814__ & ~new_new_n29826__;
  assign new_new_n29828__ = ~new_new_n29813__ & ~new_new_n29827__;
  assign new_new_n29829__ = ~new_new_n29331__ & ~new_new_n29332__;
  assign new_new_n29830__ = new_new_n29349__ & ~new_new_n29829__;
  assign new_new_n29831__ = ~new_new_n29349__ & new_new_n29829__;
  assign new_new_n29832__ = ~new_new_n29830__ & ~new_new_n29831__;
  assign new_new_n29833__ = new_new_n29828__ & new_new_n29832__;
  assign new_new_n29834__ = new_new_n29446__ & ~new_new_n29833__;
  assign new_new_n29835__ = ~new_new_n29828__ & ~new_new_n29832__;
  assign new_new_n29836__ = ~new_new_n29834__ & ~new_new_n29835__;
  assign new_new_n29837__ = ~new_new_n29434__ & ~new_new_n29836__;
  assign new_new_n29838__ = new_new_n29434__ & new_new_n29836__;
  assign new_new_n29839__ = ~new_new_n29356__ & ~new_new_n29357__;
  assign new_new_n29840__ = new_new_n29374__ & ~new_new_n29839__;
  assign new_new_n29841__ = ~new_new_n29374__ & new_new_n29839__;
  assign new_new_n29842__ = ~new_new_n29840__ & ~new_new_n29841__;
  assign new_new_n29843__ = ~new_new_n29838__ & ~new_new_n29842__;
  assign new_new_n29844__ = ~new_new_n29837__ & ~new_new_n29843__;
  assign new_new_n29845__ = ~new_new_n29410__ & new_new_n29844__;
  assign new_new_n29846__ = new_new_n29410__ & ~new_new_n29844__;
  assign new_new_n29847__ = ~new_new_n29377__ & ~new_new_n29378__;
  assign new_new_n29848__ = ~new_new_n29389__ & ~new_new_n29847__;
  assign new_new_n29849__ = new_new_n29389__ & new_new_n29847__;
  assign new_new_n29850__ = ~new_new_n29848__ & ~new_new_n29849__;
  assign new_new_n29851__ = ~new_new_n29846__ & ~new_new_n29850__;
  assign new_new_n29852__ = ~new_new_n29845__ & ~new_new_n29851__;
  assign new_new_n29853__ = new_new_n29394__ & ~new_new_n29852__;
  assign new_new_n29854__ = ~new_new_n29394__ & new_new_n29852__;
  assign new_new_n29855__ = ~new_new_n29853__ & ~new_new_n29854__;
  assign new_new_n29856__ = pi11 & ~new_new_n29855__;
  assign new_new_n29857__ = ~pi11 & new_new_n29855__;
  assign new_new_n29858__ = ~new_new_n29856__ & ~new_new_n29857__;
  assign new_new_n29859__ = new_new_n27415__ & new_new_n29858__;
  assign new_new_n29860__ = ~new_new_n27415__ & ~new_new_n29858__;
  assign new_new_n29861__ = ~new_new_n29859__ & ~new_new_n29860__;
  assign new_new_n29862__ = ~new_new_n27405__ & ~new_new_n29861__;
  assign new_new_n29863__ = new_new_n27405__ & new_new_n29861__;
  assign new_new_n29864__ = ~new_new_n29389__ & new_new_n29410__;
  assign new_new_n29865__ = new_new_n29389__ & ~new_new_n29410__;
  assign new_new_n29866__ = ~new_new_n29864__ & ~new_new_n29865__;
  assign new_new_n29867__ = new_new_n29847__ & ~new_new_n29866__;
  assign new_new_n29868__ = ~new_new_n29847__ & new_new_n29866__;
  assign new_new_n29869__ = ~new_new_n29867__ & ~new_new_n29868__;
  assign new_new_n29870__ = new_new_n29844__ & new_new_n29869__;
  assign new_new_n29871__ = ~new_new_n29844__ & ~new_new_n29869__;
  assign new_new_n29872__ = ~new_new_n29870__ & ~new_new_n29871__;
  assign new_new_n29873__ = ~new_new_n11409__ & ~new_new_n26854__;
  assign new_new_n29874__ = new_new_n10702__ & new_new_n26847__;
  assign new_new_n29875__ = ~new_new_n29873__ & ~new_new_n29874__;
  assign new_new_n29876__ = new_new_n10694__ & ~new_new_n26823__;
  assign new_new_n29877__ = ~new_new_n29400__ & new_new_n29876__;
  assign new_new_n29878__ = new_new_n29875__ & ~new_new_n29877__;
  assign new_new_n29879__ = ~pi08 & ~new_new_n29878__;
  assign new_new_n29880__ = new_new_n26823__ & new_new_n29400__;
  assign new_new_n29881__ = new_new_n10694__ & ~new_new_n29880__;
  assign new_new_n29882__ = ~pi08 & ~new_new_n29881__;
  assign new_new_n29883__ = ~pi07 & new_new_n29400__;
  assign new_new_n29884__ = pi07 & new_new_n26823__;
  assign new_new_n29885__ = new_new_n10694__ & ~new_new_n29884__;
  assign new_new_n29886__ = ~new_new_n29883__ & new_new_n29885__;
  assign new_new_n29887__ = new_new_n29875__ & ~new_new_n29886__;
  assign new_new_n29888__ = ~new_new_n29882__ & new_new_n29887__;
  assign new_new_n29889__ = ~new_new_n29879__ & ~new_new_n29888__;
  assign new_new_n29890__ = ~new_new_n29787__ & ~new_new_n29788__;
  assign new_new_n29891__ = ~new_new_n29798__ & new_new_n29890__;
  assign new_new_n29892__ = new_new_n29798__ & ~new_new_n29890__;
  assign new_new_n29893__ = ~new_new_n29891__ & ~new_new_n29892__;
  assign new_new_n29894__ = new_new_n10698__ & new_new_n26847__;
  assign new_new_n29895__ = new_new_n10702__ & ~new_new_n26854__;
  assign new_new_n29896__ = ~new_new_n11409__ & ~new_new_n26888__;
  assign new_new_n29897__ = new_new_n11378__ & new_new_n29424__;
  assign new_new_n29898__ = ~new_new_n29895__ & ~new_new_n29896__;
  assign new_new_n29899__ = ~new_new_n29894__ & new_new_n29898__;
  assign new_new_n29900__ = ~new_new_n29897__ & new_new_n29899__;
  assign new_new_n29901__ = ~new_new_n29801__ & ~new_new_n29802__;
  assign new_new_n29902__ = new_new_n29806__ & new_new_n29901__;
  assign new_new_n29903__ = ~new_new_n29806__ & ~new_new_n29901__;
  assign new_new_n29904__ = ~new_new_n29902__ & ~new_new_n29903__;
  assign new_new_n29905__ = new_new_n11378__ & ~new_new_n27430__;
  assign new_new_n29906__ = ~new_new_n11409__ & new_new_n26922__;
  assign new_new_n29907__ = new_new_n10702__ & ~new_new_n26888__;
  assign new_new_n29908__ = new_new_n10698__ & ~new_new_n26854__;
  assign new_new_n29909__ = ~new_new_n29906__ & ~new_new_n29907__;
  assign new_new_n29910__ = ~new_new_n29908__ & new_new_n29909__;
  assign new_new_n29911__ = ~new_new_n29905__ & new_new_n29910__;
  assign new_new_n29912__ = ~new_new_n29904__ & new_new_n29911__;
  assign new_new_n29913__ = pi08 & ~new_new_n29911__;
  assign new_new_n29914__ = ~new_new_n29912__ & ~new_new_n29913__;
  assign new_new_n29915__ = ~new_new_n29900__ & new_new_n29914__;
  assign new_new_n29916__ = new_new_n29904__ & ~new_new_n29911__;
  assign new_new_n29917__ = ~new_new_n29773__ & ~new_new_n29774__;
  assign new_new_n29918__ = new_new_n29784__ & new_new_n29917__;
  assign new_new_n29919__ = ~new_new_n29784__ & ~new_new_n29917__;
  assign new_new_n29920__ = ~new_new_n29918__ & ~new_new_n29919__;
  assign new_new_n29921__ = ~new_new_n11409__ & new_new_n26917__;
  assign new_new_n29922__ = new_new_n10702__ & ~new_new_n27168__;
  assign new_new_n29923__ = new_new_n10698__ & new_new_n26922__;
  assign new_new_n29924__ = ~new_new_n29921__ & ~new_new_n29922__;
  assign new_new_n29925__ = ~new_new_n29923__ & new_new_n29924__;
  assign new_new_n29926__ = new_new_n10694__ & ~new_new_n29366__;
  assign new_new_n29927__ = ~pi08 & ~new_new_n29926__;
  assign new_new_n29928__ = new_new_n12121__ & ~new_new_n29366__;
  assign new_new_n29929__ = ~new_new_n29927__ & ~new_new_n29928__;
  assign new_new_n29930__ = new_new_n29925__ & ~new_new_n29929__;
  assign new_new_n29931__ = pi08 & ~new_new_n29925__;
  assign new_new_n29932__ = ~new_new_n29930__ & ~new_new_n29931__;
  assign new_new_n29933__ = new_new_n11378__ & ~new_new_n28799__;
  assign new_new_n29934__ = ~new_new_n11409__ & new_new_n26928__;
  assign new_new_n29935__ = new_new_n10702__ & new_new_n26917__;
  assign new_new_n29936__ = ~new_new_n29934__ & ~new_new_n29935__;
  assign new_new_n29937__ = ~new_new_n29933__ & new_new_n29936__;
  assign new_new_n29938__ = new_new_n10694__ & ~new_new_n27168__;
  assign new_new_n29939__ = ~pi08 & ~new_new_n29938__;
  assign new_new_n29940__ = new_new_n11498__ & ~new_new_n27168__;
  assign new_new_n29941__ = ~new_new_n29939__ & ~new_new_n29940__;
  assign new_new_n29942__ = new_new_n29937__ & ~new_new_n29941__;
  assign new_new_n29943__ = pi08 & ~new_new_n29937__;
  assign new_new_n29944__ = ~new_new_n29942__ & ~new_new_n29943__;
  assign new_new_n29945__ = ~new_new_n29714__ & ~new_new_n29715__;
  assign new_new_n29946__ = new_new_n29721__ & new_new_n29945__;
  assign new_new_n29947__ = ~new_new_n29721__ & ~new_new_n29945__;
  assign new_new_n29948__ = ~new_new_n29946__ & ~new_new_n29947__;
  assign new_new_n29949__ = new_new_n10698__ & new_new_n27152__;
  assign new_new_n29950__ = ~new_new_n11409__ & new_new_n26971__;
  assign new_new_n29951__ = new_new_n10702__ & ~new_new_n26937__;
  assign new_new_n29952__ = ~new_new_n29950__ & ~new_new_n29951__;
  assign new_new_n29953__ = ~new_new_n29949__ & new_new_n29952__;
  assign new_new_n29954__ = new_new_n12408__ & new_new_n29953__;
  assign new_new_n29955__ = new_new_n12415__ & ~new_new_n27152__;
  assign new_new_n29956__ = pi08 & new_new_n27152__;
  assign new_new_n29957__ = new_new_n29953__ & new_new_n29956__;
  assign new_new_n29958__ = ~new_new_n29955__ & ~new_new_n29957__;
  assign new_new_n29959__ = new_new_n27477__ & ~new_new_n29958__;
  assign new_new_n29960__ = new_new_n12415__ & new_new_n27152__;
  assign new_new_n29961__ = pi08 & ~new_new_n27152__;
  assign new_new_n29962__ = new_new_n29953__ & new_new_n29961__;
  assign new_new_n29963__ = ~new_new_n29960__ & ~new_new_n29962__;
  assign new_new_n29964__ = ~new_new_n27477__ & ~new_new_n29963__;
  assign new_new_n29965__ = ~pi08 & ~new_new_n29953__;
  assign new_new_n29966__ = ~new_new_n29954__ & ~new_new_n29965__;
  assign new_new_n29967__ = ~new_new_n29959__ & new_new_n29966__;
  assign new_new_n29968__ = ~new_new_n29964__ & new_new_n29967__;
  assign new_new_n29969__ = ~new_new_n29948__ & ~new_new_n29968__;
  assign new_new_n29970__ = new_new_n29948__ & new_new_n29968__;
  assign new_new_n29971__ = ~new_new_n29706__ & ~new_new_n29707__;
  assign new_new_n29972__ = ~new_new_n29711__ & new_new_n29971__;
  assign new_new_n29973__ = new_new_n29711__ & ~new_new_n29971__;
  assign new_new_n29974__ = ~new_new_n29972__ & ~new_new_n29973__;
  assign new_new_n29975__ = new_new_n10698__ & new_new_n26971__;
  assign new_new_n29976__ = ~new_new_n11409__ & ~new_new_n27003__;
  assign new_new_n29977__ = new_new_n10702__ & ~new_new_n26978__;
  assign new_new_n29978__ = ~new_new_n29976__ & ~new_new_n29977__;
  assign new_new_n29979__ = ~new_new_n29975__ & new_new_n29978__;
  assign new_new_n29980__ = new_new_n10694__ & new_new_n28277__;
  assign new_new_n29981__ = pi08 & ~new_new_n29980__;
  assign new_new_n29982__ = new_new_n11498__ & new_new_n28277__;
  assign new_new_n29983__ = ~new_new_n29981__ & ~new_new_n29982__;
  assign new_new_n29984__ = new_new_n29979__ & ~new_new_n29983__;
  assign new_new_n29985__ = ~pi08 & ~new_new_n29979__;
  assign new_new_n29986__ = ~new_new_n29984__ & ~new_new_n29985__;
  assign new_new_n29987__ = ~new_new_n29678__ & ~new_new_n29679__;
  assign new_new_n29988__ = ~new_new_n29689__ & new_new_n29987__;
  assign new_new_n29989__ = new_new_n29689__ & ~new_new_n29987__;
  assign new_new_n29990__ = ~new_new_n29988__ & ~new_new_n29989__;
  assign new_new_n29991__ = new_new_n10698__ & ~new_new_n27029__;
  assign new_new_n29992__ = new_new_n10702__ & ~new_new_n27021__;
  assign new_new_n29993__ = ~new_new_n11409__ & new_new_n27111__;
  assign new_new_n29994__ = new_new_n11378__ & new_new_n27764__;
  assign new_new_n29995__ = ~new_new_n29992__ & ~new_new_n29993__;
  assign new_new_n29996__ = ~new_new_n29991__ & new_new_n29995__;
  assign new_new_n29997__ = ~new_new_n29994__ & new_new_n29996__;
  assign new_new_n29998__ = pi08 & ~new_new_n29997__;
  assign new_new_n29999__ = ~pi08 & new_new_n29997__;
  assign new_new_n30000__ = ~new_new_n29998__ & ~new_new_n29999__;
  assign new_new_n30001__ = ~new_new_n29638__ & ~new_new_n29639__;
  assign new_new_n30002__ = ~new_new_n29649__ & new_new_n30001__;
  assign new_new_n30003__ = new_new_n29649__ & ~new_new_n30001__;
  assign new_new_n30004__ = ~new_new_n30002__ & ~new_new_n30003__;
  assign new_new_n30005__ = new_new_n10702__ & ~new_new_n27033__;
  assign new_new_n30006__ = ~new_new_n11409__ & ~new_new_n27054__;
  assign new_new_n30007__ = ~new_new_n30005__ & ~new_new_n30006__;
  assign new_new_n30008__ = new_new_n10694__ & new_new_n27687__;
  assign new_new_n30009__ = new_new_n30007__ & ~new_new_n30008__;
  assign new_new_n30010__ = pi08 & ~new_new_n30009__;
  assign new_new_n30011__ = new_new_n10694__ & ~new_new_n27691__;
  assign new_new_n30012__ = ~pi08 & ~new_new_n30011__;
  assign new_new_n30013__ = ~pi07 & new_new_n27111__;
  assign new_new_n30014__ = pi07 & ~new_new_n27111__;
  assign new_new_n30015__ = new_new_n10694__ & ~new_new_n30013__;
  assign new_new_n30016__ = ~new_new_n30014__ & new_new_n30015__;
  assign new_new_n30017__ = new_new_n27686__ & new_new_n30016__;
  assign new_new_n30018__ = ~new_new_n30012__ & ~new_new_n30017__;
  assign new_new_n30019__ = new_new_n30007__ & ~new_new_n30018__;
  assign new_new_n30020__ = ~new_new_n30010__ & ~new_new_n30019__;
  assign new_new_n30021__ = new_new_n8469__ & new_new_n27567__;
  assign new_new_n30022__ = ~pi10 & ~new_new_n29623__;
  assign new_new_n30023__ = pi10 & new_new_n29623__;
  assign new_new_n30024__ = ~new_new_n30022__ & ~new_new_n30023__;
  assign new_new_n30025__ = new_new_n30021__ & ~new_new_n30024__;
  assign new_new_n30026__ = pi11 & ~new_new_n29623__;
  assign new_new_n30027__ = ~pi11 & new_new_n29623__;
  assign new_new_n30028__ = ~new_new_n30026__ & ~new_new_n30027__;
  assign new_new_n30029__ = ~new_new_n30021__ & new_new_n30028__;
  assign new_new_n30030__ = ~new_new_n30025__ & ~new_new_n30029__;
  assign new_new_n30031__ = new_new_n29630__ & ~new_new_n30030__;
  assign new_new_n30032__ = ~new_new_n29630__ & ~new_new_n30028__;
  assign new_new_n30033__ = ~new_new_n30031__ & ~new_new_n30032__;
  assign new_new_n30034__ = ~new_new_n29615__ & ~new_new_n30033__;
  assign new_new_n30035__ = new_new_n30020__ & ~new_new_n30034__;
  assign new_new_n30036__ = ~new_new_n30020__ & new_new_n30034__;
  assign new_new_n30037__ = new_new_n29601__ & new_new_n29613__;
  assign new_new_n30038__ = ~new_new_n29600__ & ~new_new_n30037__;
  assign new_new_n30039__ = new_new_n29614__ & ~new_new_n30038__;
  assign new_new_n30040__ = ~new_new_n29614__ & new_new_n30038__;
  assign new_new_n30041__ = ~new_new_n30039__ & ~new_new_n30040__;
  assign new_new_n30042__ = new_new_n10698__ & ~new_new_n27054__;
  assign new_new_n30043__ = ~new_new_n11409__ & ~new_new_n27071__;
  assign new_new_n30044__ = new_new_n10702__ & new_new_n27041__;
  assign new_new_n30045__ = ~new_new_n30043__ & ~new_new_n30044__;
  assign new_new_n30046__ = ~new_new_n30042__ & new_new_n30045__;
  assign new_new_n30047__ = new_new_n10694__ & ~new_new_n27094__;
  assign new_new_n30048__ = ~pi08 & ~new_new_n30047__;
  assign new_new_n30049__ = new_new_n12121__ & ~new_new_n27094__;
  assign new_new_n30050__ = ~new_new_n30048__ & ~new_new_n30049__;
  assign new_new_n30051__ = new_new_n30046__ & ~new_new_n30050__;
  assign new_new_n30052__ = pi08 & ~new_new_n30046__;
  assign new_new_n30053__ = ~new_new_n30051__ & ~new_new_n30052__;
  assign new_new_n30054__ = new_new_n8469__ & ~new_new_n27075__;
  assign new_new_n30055__ = new_new_n10694__ & new_new_n26118__;
  assign new_new_n30056__ = new_new_n27075__ & ~new_new_n30055__;
  assign new_new_n30057__ = ~new_new_n12276__ & ~new_new_n30056__;
  assign new_new_n30058__ = new_new_n10702__ & new_new_n26118__;
  assign new_new_n30059__ = ~new_new_n11409__ & ~new_new_n27075__;
  assign new_new_n30060__ = ~new_new_n10697__ & new_new_n27582__;
  assign new_new_n30061__ = new_new_n27059__ & new_new_n30060__;
  assign new_new_n30062__ = ~new_new_n27059__ & ~new_new_n30060__;
  assign new_new_n30063__ = new_new_n10694__ & ~new_new_n30061__;
  assign new_new_n30064__ = ~new_new_n30062__ & new_new_n30063__;
  assign new_new_n30065__ = ~new_new_n30058__ & ~new_new_n30059__;
  assign new_new_n30066__ = ~new_new_n30064__ & new_new_n30065__;
  assign new_new_n30067__ = pi08 & ~new_new_n30057__;
  assign new_new_n30068__ = new_new_n30066__ & new_new_n30067__;
  assign new_new_n30069__ = ~new_new_n30054__ & ~new_new_n30068__;
  assign new_new_n30070__ = new_new_n10698__ & ~new_new_n27071__;
  assign new_new_n30071__ = ~new_new_n11409__ & new_new_n26118__;
  assign new_new_n30072__ = new_new_n10702__ & new_new_n27059__;
  assign new_new_n30073__ = ~new_new_n30071__ & ~new_new_n30072__;
  assign new_new_n30074__ = ~new_new_n30070__ & new_new_n30073__;
  assign new_new_n30075__ = new_new_n10694__ & new_new_n27600__;
  assign new_new_n30076__ = pi08 & ~new_new_n30075__;
  assign new_new_n30077__ = new_new_n11498__ & new_new_n27600__;
  assign new_new_n30078__ = ~new_new_n30076__ & ~new_new_n30077__;
  assign new_new_n30079__ = new_new_n30074__ & ~new_new_n30078__;
  assign new_new_n30080__ = ~pi08 & ~new_new_n30074__;
  assign new_new_n30081__ = ~new_new_n30079__ & ~new_new_n30080__;
  assign new_new_n30082__ = ~new_new_n30069__ & ~new_new_n30081__;
  assign new_new_n30083__ = new_new_n8472__ & new_new_n27087__;
  assign new_new_n30084__ = ~new_new_n8469__ & new_new_n27582__;
  assign new_new_n30085__ = ~new_new_n8301__ & new_new_n26118__;
  assign new_new_n30086__ = new_new_n8473__ & ~new_new_n30085__;
  assign new_new_n30087__ = ~new_new_n8855__ & ~new_new_n27577__;
  assign new_new_n30088__ = ~new_new_n30083__ & new_new_n30087__;
  assign new_new_n30089__ = ~new_new_n30084__ & ~new_new_n30086__;
  assign new_new_n30090__ = new_new_n30088__ & new_new_n30089__;
  assign new_new_n30091__ = ~new_new_n30082__ & ~new_new_n30090__;
  assign new_new_n30092__ = new_new_n30082__ & new_new_n30090__;
  assign new_new_n30093__ = new_new_n10698__ & new_new_n27041__;
  assign new_new_n30094__ = new_new_n10702__ & ~new_new_n27071__;
  assign new_new_n30095__ = ~new_new_n11409__ & new_new_n27059__;
  assign new_new_n30096__ = new_new_n11378__ & new_new_n27567__;
  assign new_new_n30097__ = ~new_new_n30093__ & ~new_new_n30095__;
  assign new_new_n30098__ = ~new_new_n30094__ & new_new_n30097__;
  assign new_new_n30099__ = ~new_new_n30096__ & new_new_n30098__;
  assign new_new_n30100__ = pi08 & ~new_new_n30099__;
  assign new_new_n30101__ = ~pi08 & new_new_n30099__;
  assign new_new_n30102__ = ~new_new_n30100__ & ~new_new_n30101__;
  assign new_new_n30103__ = ~new_new_n30092__ & ~new_new_n30102__;
  assign new_new_n30104__ = ~new_new_n30091__ & ~new_new_n30103__;
  assign new_new_n30105__ = ~new_new_n30053__ & ~new_new_n30104__;
  assign new_new_n30106__ = new_new_n30053__ & new_new_n30104__;
  assign new_new_n30107__ = ~pi11 & ~new_new_n26118__;
  assign new_new_n30108__ = new_new_n24042__ & new_new_n27087__;
  assign new_new_n30109__ = ~new_new_n8474__ & ~new_new_n20003__;
  assign new_new_n30110__ = ~new_new_n27577__ & ~new_new_n30109__;
  assign new_new_n30111__ = ~new_new_n30107__ & new_new_n30110__;
  assign new_new_n30112__ = ~new_new_n30108__ & new_new_n30111__;
  assign new_new_n30113__ = new_new_n29611__ & ~new_new_n30112__;
  assign new_new_n30114__ = new_new_n8474__ & ~new_new_n27087__;
  assign new_new_n30115__ = new_new_n20003__ & ~new_new_n27577__;
  assign new_new_n30116__ = ~new_new_n30114__ & new_new_n30115__;
  assign new_new_n30117__ = ~new_new_n29611__ & new_new_n30116__;
  assign new_new_n30118__ = ~new_new_n30113__ & ~new_new_n30117__;
  assign new_new_n30119__ = ~new_new_n30106__ & ~new_new_n30118__;
  assign new_new_n30120__ = ~new_new_n30105__ & ~new_new_n30119__;
  assign new_new_n30121__ = ~new_new_n30041__ & ~new_new_n30120__;
  assign new_new_n30122__ = new_new_n10698__ & ~new_new_n27033__;
  assign new_new_n30123__ = ~new_new_n11409__ & new_new_n27041__;
  assign new_new_n30124__ = new_new_n10702__ & ~new_new_n27054__;
  assign new_new_n30125__ = ~new_new_n30123__ & ~new_new_n30124__;
  assign new_new_n30126__ = ~new_new_n30122__ & new_new_n30125__;
  assign new_new_n30127__ = new_new_n10694__ & ~new_new_n27535__;
  assign new_new_n30128__ = ~new_new_n29095__ & new_new_n30127__;
  assign new_new_n30129__ = pi08 & ~new_new_n30128__;
  assign new_new_n30130__ = pi07 & new_new_n30128__;
  assign new_new_n30131__ = ~new_new_n30129__ & ~new_new_n30130__;
  assign new_new_n30132__ = new_new_n30126__ & ~new_new_n30131__;
  assign new_new_n30133__ = ~pi08 & ~new_new_n30126__;
  assign new_new_n30134__ = ~new_new_n30132__ & ~new_new_n30133__;
  assign new_new_n30135__ = ~new_new_n30121__ & ~new_new_n30134__;
  assign new_new_n30136__ = new_new_n30041__ & new_new_n30120__;
  assign new_new_n30137__ = ~new_new_n30135__ & ~new_new_n30136__;
  assign new_new_n30138__ = ~new_new_n30036__ & ~new_new_n30137__;
  assign new_new_n30139__ = ~new_new_n30035__ & ~new_new_n30138__;
  assign new_new_n30140__ = new_new_n30020__ & new_new_n30135__;
  assign new_new_n30141__ = new_new_n29615__ & new_new_n30033__;
  assign new_new_n30142__ = ~new_new_n30140__ & new_new_n30141__;
  assign new_new_n30143__ = ~new_new_n30139__ & ~new_new_n30142__;
  assign new_new_n30144__ = ~new_new_n30004__ & new_new_n30143__;
  assign new_new_n30145__ = new_new_n30004__ & ~new_new_n30143__;
  assign new_new_n30146__ = new_new_n10698__ & ~new_new_n27021__;
  assign new_new_n30147__ = ~new_new_n11409__ & ~new_new_n27033__;
  assign new_new_n30148__ = new_new_n10702__ & new_new_n27111__;
  assign new_new_n30149__ = ~new_new_n30147__ & ~new_new_n30148__;
  assign new_new_n30150__ = ~new_new_n30146__ & new_new_n30149__;
  assign new_new_n30151__ = new_new_n11378__ & new_new_n27796__;
  assign new_new_n30152__ = new_new_n30150__ & ~new_new_n30151__;
  assign new_new_n30153__ = ~pi08 & ~new_new_n30152__;
  assign new_new_n30154__ = pi08 & new_new_n30152__;
  assign new_new_n30155__ = ~new_new_n30153__ & ~new_new_n30154__;
  assign new_new_n30156__ = ~new_new_n30145__ & ~new_new_n30155__;
  assign new_new_n30157__ = ~new_new_n30144__ & ~new_new_n30156__;
  assign new_new_n30158__ = new_new_n30000__ & ~new_new_n30157__;
  assign new_new_n30159__ = ~new_new_n30000__ & new_new_n30157__;
  assign new_new_n30160__ = ~new_new_n29652__ & ~new_new_n29653__;
  assign new_new_n30161__ = new_new_n29658__ & new_new_n30160__;
  assign new_new_n30162__ = ~new_new_n29658__ & ~new_new_n30160__;
  assign new_new_n30163__ = ~new_new_n30161__ & ~new_new_n30162__;
  assign new_new_n30164__ = ~new_new_n30159__ & new_new_n30163__;
  assign new_new_n30165__ = ~new_new_n30158__ & ~new_new_n30164__;
  assign new_new_n30166__ = ~new_new_n29661__ & ~new_new_n29662__;
  assign new_new_n30167__ = ~new_new_n29666__ & new_new_n30166__;
  assign new_new_n30168__ = new_new_n29666__ & ~new_new_n30166__;
  assign new_new_n30169__ = ~new_new_n30167__ & ~new_new_n30168__;
  assign new_new_n30170__ = new_new_n30165__ & ~new_new_n30169__;
  assign new_new_n30171__ = ~new_new_n30165__ & new_new_n30169__;
  assign new_new_n30172__ = new_new_n10698__ & ~new_new_n27003__;
  assign new_new_n30173__ = ~new_new_n11409__ & ~new_new_n27021__;
  assign new_new_n30174__ = new_new_n10702__ & ~new_new_n27029__;
  assign new_new_n30175__ = ~new_new_n30173__ & ~new_new_n30174__;
  assign new_new_n30176__ = ~new_new_n30172__ & new_new_n30175__;
  assign new_new_n30177__ = new_new_n10694__ & new_new_n27962__;
  assign new_new_n30178__ = pi08 & ~new_new_n30177__;
  assign new_new_n30179__ = new_new_n11498__ & new_new_n27962__;
  assign new_new_n30180__ = ~new_new_n30178__ & ~new_new_n30179__;
  assign new_new_n30181__ = new_new_n30176__ & ~new_new_n30180__;
  assign new_new_n30182__ = ~pi08 & ~new_new_n30176__;
  assign new_new_n30183__ = ~new_new_n30181__ & ~new_new_n30182__;
  assign new_new_n30184__ = ~new_new_n30171__ & new_new_n30183__;
  assign new_new_n30185__ = ~new_new_n30170__ & ~new_new_n30184__;
  assign new_new_n30186__ = new_new_n29990__ & ~new_new_n30185__;
  assign new_new_n30187__ = ~new_new_n29990__ & new_new_n30185__;
  assign new_new_n30188__ = new_new_n10698__ & ~new_new_n26978__;
  assign new_new_n30189__ = ~new_new_n11409__ & ~new_new_n27029__;
  assign new_new_n30190__ = new_new_n10702__ & ~new_new_n27003__;
  assign new_new_n30191__ = new_new_n11378__ & new_new_n27986__;
  assign new_new_n30192__ = ~new_new_n30189__ & ~new_new_n30190__;
  assign new_new_n30193__ = ~new_new_n30188__ & new_new_n30192__;
  assign new_new_n30194__ = ~new_new_n30191__ & new_new_n30193__;
  assign new_new_n30195__ = ~pi08 & ~new_new_n30194__;
  assign new_new_n30196__ = pi08 & new_new_n30194__;
  assign new_new_n30197__ = ~new_new_n30195__ & ~new_new_n30196__;
  assign new_new_n30198__ = ~new_new_n30187__ & new_new_n30197__;
  assign new_new_n30199__ = ~new_new_n30186__ & ~new_new_n30198__;
  assign new_new_n30200__ = ~new_new_n29986__ & new_new_n30199__;
  assign new_new_n30201__ = new_new_n29986__ & ~new_new_n30199__;
  assign new_new_n30202__ = pi11 & ~new_new_n29552__;
  assign new_new_n30203__ = ~pi11 & new_new_n29552__;
  assign new_new_n30204__ = ~new_new_n30202__ & ~new_new_n30203__;
  assign new_new_n30205__ = ~new_new_n29691__ & new_new_n30204__;
  assign new_new_n30206__ = new_new_n29691__ & ~new_new_n30204__;
  assign new_new_n30207__ = ~new_new_n30205__ & ~new_new_n30206__;
  assign new_new_n30208__ = new_new_n29700__ & new_new_n30207__;
  assign new_new_n30209__ = ~new_new_n29700__ & ~new_new_n30207__;
  assign new_new_n30210__ = ~new_new_n30208__ & ~new_new_n30209__;
  assign new_new_n30211__ = ~new_new_n30201__ & ~new_new_n30210__;
  assign new_new_n30212__ = ~new_new_n30200__ & ~new_new_n30211__;
  assign new_new_n30213__ = new_new_n29974__ & ~new_new_n30212__;
  assign new_new_n30214__ = ~new_new_n29974__ & new_new_n30212__;
  assign new_new_n30215__ = new_new_n10702__ & new_new_n26971__;
  assign new_new_n30216__ = ~new_new_n11409__ & ~new_new_n26978__;
  assign new_new_n30217__ = new_new_n10698__ & ~new_new_n26937__;
  assign new_new_n30218__ = ~new_new_n30215__ & ~new_new_n30216__;
  assign new_new_n30219__ = ~new_new_n30217__ & new_new_n30218__;
  assign new_new_n30220__ = new_new_n10694__ & new_new_n28005__;
  assign new_new_n30221__ = pi08 & ~new_new_n30220__;
  assign new_new_n30222__ = new_new_n11498__ & new_new_n28005__;
  assign new_new_n30223__ = ~new_new_n30221__ & ~new_new_n30222__;
  assign new_new_n30224__ = new_new_n30219__ & ~new_new_n30223__;
  assign new_new_n30225__ = ~pi08 & ~new_new_n30219__;
  assign new_new_n30226__ = ~new_new_n30224__ & ~new_new_n30225__;
  assign new_new_n30227__ = ~new_new_n30214__ & ~new_new_n30226__;
  assign new_new_n30228__ = ~new_new_n30213__ & ~new_new_n30227__;
  assign new_new_n30229__ = ~new_new_n29970__ & ~new_new_n30228__;
  assign new_new_n30230__ = ~new_new_n29969__ & ~new_new_n30229__;
  assign new_new_n30231__ = ~new_new_n29731__ & ~new_new_n29733__;
  assign new_new_n30232__ = new_new_n10702__ & new_new_n27152__;
  assign new_new_n30233__ = ~new_new_n11409__ & ~new_new_n26937__;
  assign new_new_n30234__ = new_new_n10698__ & ~new_new_n26941__;
  assign new_new_n30235__ = ~new_new_n30233__ & ~new_new_n30234__;
  assign new_new_n30236__ = ~new_new_n30232__ & new_new_n30235__;
  assign new_new_n30237__ = new_new_n10694__ & ~new_new_n27502__;
  assign new_new_n30238__ = pi08 & ~new_new_n30237__;
  assign new_new_n30239__ = new_new_n11498__ & ~new_new_n27502__;
  assign new_new_n30240__ = ~new_new_n30238__ & ~new_new_n30239__;
  assign new_new_n30241__ = new_new_n30236__ & ~new_new_n30240__;
  assign new_new_n30242__ = ~pi08 & ~new_new_n30236__;
  assign new_new_n30243__ = ~new_new_n30241__ & ~new_new_n30242__;
  assign new_new_n30244__ = new_new_n30231__ & new_new_n30243__;
  assign new_new_n30245__ = ~new_new_n30230__ & ~new_new_n30244__;
  assign new_new_n30246__ = ~new_new_n30231__ & ~new_new_n30243__;
  assign new_new_n30247__ = ~new_new_n30245__ & ~new_new_n30246__;
  assign new_new_n30248__ = ~new_new_n29743__ & ~new_new_n29744__;
  assign new_new_n30249__ = ~new_new_n29754__ & new_new_n30248__;
  assign new_new_n30250__ = new_new_n29754__ & ~new_new_n30248__;
  assign new_new_n30251__ = ~new_new_n30249__ & ~new_new_n30250__;
  assign new_new_n30252__ = ~new_new_n30247__ & ~new_new_n30251__;
  assign new_new_n30253__ = new_new_n30247__ & new_new_n30251__;
  assign new_new_n30254__ = new_new_n10698__ & new_new_n26928__;
  assign new_new_n30255__ = new_new_n10702__ & ~new_new_n26941__;
  assign new_new_n30256__ = ~new_new_n11409__ & new_new_n27152__;
  assign new_new_n30257__ = new_new_n11378__ & new_new_n27488__;
  assign new_new_n30258__ = ~new_new_n30255__ & ~new_new_n30256__;
  assign new_new_n30259__ = ~new_new_n30254__ & new_new_n30258__;
  assign new_new_n30260__ = ~new_new_n30257__ & new_new_n30259__;
  assign new_new_n30261__ = ~pi08 & ~new_new_n30260__;
  assign new_new_n30262__ = pi08 & new_new_n30260__;
  assign new_new_n30263__ = ~new_new_n30261__ & ~new_new_n30262__;
  assign new_new_n30264__ = ~new_new_n30253__ & ~new_new_n30263__;
  assign new_new_n30265__ = ~new_new_n30252__ & ~new_new_n30264__;
  assign new_new_n30266__ = ~new_new_n29503__ & ~new_new_n29504__;
  assign new_new_n30267__ = new_new_n29756__ & new_new_n30266__;
  assign new_new_n30268__ = ~new_new_n29756__ & ~new_new_n30266__;
  assign new_new_n30269__ = ~new_new_n30267__ & ~new_new_n30268__;
  assign new_new_n30270__ = new_new_n30265__ & ~new_new_n30269__;
  assign new_new_n30271__ = ~new_new_n30265__ & new_new_n30269__;
  assign new_new_n30272__ = new_new_n10698__ & new_new_n26917__;
  assign new_new_n30273__ = new_new_n10702__ & new_new_n26928__;
  assign new_new_n30274__ = ~new_new_n11409__ & ~new_new_n26941__;
  assign new_new_n30275__ = new_new_n11378__ & ~new_new_n27462__;
  assign new_new_n30276__ = ~new_new_n30273__ & ~new_new_n30274__;
  assign new_new_n30277__ = ~new_new_n30272__ & new_new_n30276__;
  assign new_new_n30278__ = ~new_new_n30275__ & new_new_n30277__;
  assign new_new_n30279__ = pi08 & ~new_new_n30278__;
  assign new_new_n30280__ = ~pi08 & new_new_n30278__;
  assign new_new_n30281__ = ~new_new_n30279__ & ~new_new_n30280__;
  assign new_new_n30282__ = ~new_new_n30271__ & ~new_new_n30281__;
  assign new_new_n30283__ = ~new_new_n30270__ & ~new_new_n30282__;
  assign new_new_n30284__ = ~new_new_n29944__ & ~new_new_n30283__;
  assign new_new_n30285__ = new_new_n29944__ & new_new_n30283__;
  assign new_new_n30286__ = ~new_new_n29759__ & ~new_new_n29760__;
  assign new_new_n30287__ = ~new_new_n29764__ & new_new_n30286__;
  assign new_new_n30288__ = new_new_n29764__ & ~new_new_n30286__;
  assign new_new_n30289__ = ~new_new_n30287__ & ~new_new_n30288__;
  assign new_new_n30290__ = ~new_new_n30285__ & new_new_n30289__;
  assign new_new_n30291__ = ~new_new_n30284__ & ~new_new_n30290__;
  assign new_new_n30292__ = new_new_n29932__ & new_new_n30291__;
  assign new_new_n30293__ = ~new_new_n29932__ & ~new_new_n30291__;
  assign new_new_n30294__ = ~new_new_n29476__ & ~new_new_n29770__;
  assign new_new_n30295__ = new_new_n29476__ & new_new_n29770__;
  assign new_new_n30296__ = ~new_new_n30294__ & ~new_new_n30295__;
  assign new_new_n30297__ = ~new_new_n29766__ & new_new_n30296__;
  assign new_new_n30298__ = new_new_n29766__ & ~new_new_n30296__;
  assign new_new_n30299__ = ~new_new_n30297__ & ~new_new_n30298__;
  assign new_new_n30300__ = ~new_new_n30293__ & ~new_new_n30299__;
  assign new_new_n30301__ = ~new_new_n30292__ & ~new_new_n30300__;
  assign new_new_n30302__ = new_new_n29920__ & ~new_new_n30301__;
  assign new_new_n30303__ = ~new_new_n29920__ & new_new_n30301__;
  assign new_new_n30304__ = new_new_n10698__ & ~new_new_n26888__;
  assign new_new_n30305__ = new_new_n10702__ & new_new_n26922__;
  assign new_new_n30306__ = ~new_new_n11409__ & ~new_new_n27168__;
  assign new_new_n30307__ = new_new_n11378__ & new_new_n27180__;
  assign new_new_n30308__ = ~new_new_n30305__ & ~new_new_n30306__;
  assign new_new_n30309__ = ~new_new_n30304__ & new_new_n30308__;
  assign new_new_n30310__ = ~new_new_n30307__ & new_new_n30309__;
  assign new_new_n30311__ = pi08 & ~new_new_n30310__;
  assign new_new_n30312__ = ~pi08 & new_new_n30310__;
  assign new_new_n30313__ = ~new_new_n30311__ & ~new_new_n30312__;
  assign new_new_n30314__ = ~new_new_n30303__ & new_new_n30313__;
  assign new_new_n30315__ = ~new_new_n30302__ & ~new_new_n30314__;
  assign new_new_n30316__ = ~new_new_n29911__ & new_new_n30315__;
  assign new_new_n30317__ = pi08 & ~new_new_n30316__;
  assign new_new_n30318__ = ~new_new_n29916__ & ~new_new_n30317__;
  assign new_new_n30319__ = new_new_n29900__ & ~new_new_n30318__;
  assign new_new_n30320__ = ~pi08 & ~new_new_n29900__;
  assign new_new_n30321__ = ~new_new_n29904__ & ~new_new_n30320__;
  assign new_new_n30322__ = ~new_new_n30315__ & ~new_new_n30321__;
  assign new_new_n30323__ = ~new_new_n29915__ & ~new_new_n30322__;
  assign new_new_n30324__ = ~new_new_n30319__ & new_new_n30323__;
  assign new_new_n30325__ = ~new_new_n29893__ & ~new_new_n30324__;
  assign new_new_n30326__ = pi08 & new_new_n29904__;
  assign new_new_n30327__ = pi08 & new_new_n29911__;
  assign new_new_n30328__ = ~new_new_n29916__ & ~new_new_n30327__;
  assign new_new_n30329__ = ~new_new_n30315__ & ~new_new_n30328__;
  assign new_new_n30330__ = ~new_new_n30326__ & ~new_new_n30329__;
  assign new_new_n30331__ = new_new_n29900__ & ~new_new_n30330__;
  assign new_new_n30332__ = ~pi08 & new_new_n29904__;
  assign new_new_n30333__ = new_new_n29914__ & ~new_new_n30315__;
  assign new_new_n30334__ = ~new_new_n30332__ & ~new_new_n30333__;
  assign new_new_n30335__ = ~new_new_n29900__ & ~new_new_n30334__;
  assign new_new_n30336__ = ~new_new_n30331__ & ~new_new_n30335__;
  assign new_new_n30337__ = ~new_new_n30325__ & new_new_n30336__;
  assign new_new_n30338__ = ~new_new_n29889__ & ~new_new_n30337__;
  assign new_new_n30339__ = new_new_n29889__ & new_new_n30337__;
  assign new_new_n30340__ = ~new_new_n29813__ & ~new_new_n29814__;
  assign new_new_n30341__ = new_new_n29826__ & new_new_n30340__;
  assign new_new_n30342__ = ~new_new_n29826__ & ~new_new_n30340__;
  assign new_new_n30343__ = ~new_new_n30341__ & ~new_new_n30342__;
  assign new_new_n30344__ = ~new_new_n30339__ & new_new_n30343__;
  assign new_new_n30345__ = ~new_new_n30338__ & ~new_new_n30344__;
  assign new_new_n30346__ = ~new_new_n29446__ & new_new_n29828__;
  assign new_new_n30347__ = new_new_n29446__ & ~new_new_n29828__;
  assign new_new_n30348__ = ~new_new_n30346__ & ~new_new_n30347__;
  assign new_new_n30349__ = ~new_new_n29832__ & new_new_n30345__;
  assign new_new_n30350__ = new_new_n29832__ & ~new_new_n30345__;
  assign new_new_n30351__ = ~new_new_n30349__ & ~new_new_n30350__;
  assign new_new_n30352__ = new_new_n30348__ & new_new_n30351__;
  assign new_new_n30353__ = ~new_new_n30348__ & ~new_new_n30351__;
  assign new_new_n30354__ = ~new_new_n30352__ & ~new_new_n30353__;
  assign new_new_n30355__ = ~new_new_n30345__ & ~new_new_n30354__;
  assign new_new_n30356__ = new_new_n10698__ & ~new_new_n27221__;
  assign new_new_n30357__ = ~new_new_n11409__ & new_new_n26847__;
  assign new_new_n30358__ = new_new_n10702__ & ~new_new_n26823__;
  assign new_new_n30359__ = ~new_new_n30357__ & ~new_new_n30358__;
  assign new_new_n30360__ = ~new_new_n30356__ & new_new_n30359__;
  assign new_new_n30361__ = new_new_n10694__ & new_new_n27411__;
  assign new_new_n30362__ = pi08 & ~new_new_n30361__;
  assign new_new_n30363__ = new_new_n11498__ & new_new_n27411__;
  assign new_new_n30364__ = ~new_new_n30362__ & ~new_new_n30363__;
  assign new_new_n30365__ = new_new_n30360__ & ~new_new_n30364__;
  assign new_new_n30366__ = ~pi08 & ~new_new_n30360__;
  assign new_new_n30367__ = ~new_new_n30365__ & ~new_new_n30366__;
  assign new_new_n30368__ = new_new_n30354__ & ~new_new_n30367__;
  assign new_new_n30369__ = ~new_new_n30355__ & ~new_new_n30368__;
  assign new_new_n30370__ = new_new_n29351__ & ~new_new_n29836__;
  assign new_new_n30371__ = ~new_new_n29351__ & new_new_n29836__;
  assign new_new_n30372__ = ~new_new_n30370__ & ~new_new_n30371__;
  assign new_new_n30373__ = ~new_new_n29374__ & new_new_n29434__;
  assign new_new_n30374__ = new_new_n29374__ & ~new_new_n29434__;
  assign new_new_n30375__ = ~new_new_n30373__ & ~new_new_n30374__;
  assign new_new_n30376__ = new_new_n30372__ & ~new_new_n30375__;
  assign new_new_n30377__ = ~new_new_n30372__ & new_new_n30375__;
  assign new_new_n30378__ = ~new_new_n30376__ & ~new_new_n30377__;
  assign new_new_n30379__ = new_new_n29355__ & new_new_n30378__;
  assign new_new_n30380__ = ~new_new_n29355__ & ~new_new_n30378__;
  assign new_new_n30381__ = ~new_new_n30379__ & ~new_new_n30380__;
  assign new_new_n30382__ = ~new_new_n30369__ & new_new_n30381__;
  assign new_new_n30383__ = new_new_n30369__ & ~new_new_n30381__;
  assign new_new_n30384__ = new_new_n10698__ & ~new_new_n26741__;
  assign new_new_n30385__ = ~new_new_n11409__ & ~new_new_n26823__;
  assign new_new_n30386__ = new_new_n10702__ & ~new_new_n27221__;
  assign new_new_n30387__ = ~new_new_n26823__ & new_new_n27221__;
  assign new_new_n30388__ = new_new_n26823__ & ~new_new_n27221__;
  assign new_new_n30389__ = ~new_new_n30387__ & ~new_new_n30388__;
  assign new_new_n30390__ = new_new_n27191__ & ~new_new_n30389__;
  assign new_new_n30391__ = ~new_new_n26741__ & new_new_n30390__;
  assign new_new_n30392__ = new_new_n26741__ & ~new_new_n30390__;
  assign new_new_n30393__ = ~new_new_n30391__ & ~new_new_n30392__;
  assign new_new_n30394__ = new_new_n11378__ & new_new_n30393__;
  assign new_new_n30395__ = ~new_new_n30385__ & ~new_new_n30386__;
  assign new_new_n30396__ = ~new_new_n30384__ & new_new_n30395__;
  assign new_new_n30397__ = ~new_new_n30394__ & new_new_n30396__;
  assign new_new_n30398__ = pi08 & ~new_new_n30397__;
  assign new_new_n30399__ = ~pi08 & new_new_n30397__;
  assign new_new_n30400__ = ~new_new_n30398__ & ~new_new_n30399__;
  assign new_new_n30401__ = ~new_new_n30383__ & new_new_n30400__;
  assign new_new_n30402__ = ~new_new_n30382__ & ~new_new_n30401__;
  assign new_new_n30403__ = new_new_n29872__ & ~new_new_n30402__;
  assign new_new_n30404__ = ~new_new_n29872__ & new_new_n30402__;
  assign new_new_n30405__ = new_new_n10698__ & ~new_new_n26802__;
  assign new_new_n30406__ = ~new_new_n11409__ & ~new_new_n27221__;
  assign new_new_n30407__ = new_new_n10702__ & ~new_new_n26741__;
  assign new_new_n30408__ = ~new_new_n30406__ & ~new_new_n30407__;
  assign new_new_n30409__ = ~new_new_n30405__ & new_new_n30408__;
  assign new_new_n30410__ = ~new_new_n26802__ & new_new_n27390__;
  assign new_new_n30411__ = ~new_new_n27391__ & ~new_new_n30410__;
  assign new_new_n30412__ = new_new_n10694__ & new_new_n30411__;
  assign new_new_n30413__ = pi08 & ~new_new_n30412__;
  assign new_new_n30414__ = new_new_n11498__ & new_new_n30411__;
  assign new_new_n30415__ = ~new_new_n30413__ & ~new_new_n30414__;
  assign new_new_n30416__ = new_new_n30409__ & ~new_new_n30415__;
  assign new_new_n30417__ = ~pi08 & ~new_new_n30409__;
  assign new_new_n30418__ = ~new_new_n30416__ & ~new_new_n30417__;
  assign new_new_n30419__ = ~new_new_n30404__ & ~new_new_n30418__;
  assign new_new_n30420__ = ~new_new_n30403__ & ~new_new_n30419__;
  assign new_new_n30421__ = ~new_new_n29863__ & new_new_n30420__;
  assign new_new_n30422__ = ~new_new_n29862__ & ~new_new_n30421__;
  assign new_new_n30423__ = new_new_n27385__ & ~new_new_n30422__;
  assign new_new_n30424__ = ~new_new_n27385__ & new_new_n30422__;
  assign new_new_n30425__ = ~new_new_n30423__ & ~new_new_n30424__;
  assign new_new_n30426__ = new_new_n8474__ & ~new_new_n27221__;
  assign new_new_n30427__ = ~new_new_n8479__ & ~new_new_n26823__;
  assign new_new_n30428__ = new_new_n8858__ & ~new_new_n26741__;
  assign new_new_n30429__ = ~new_new_n30426__ & ~new_new_n30427__;
  assign new_new_n30430__ = ~new_new_n30428__ & new_new_n30429__;
  assign new_new_n30431__ = new_new_n8469__ & new_new_n30393__;
  assign new_new_n30432__ = pi11 & ~new_new_n30431__;
  assign new_new_n30433__ = new_new_n11530__ & new_new_n30393__;
  assign new_new_n30434__ = ~new_new_n30432__ & ~new_new_n30433__;
  assign new_new_n30435__ = new_new_n30430__ & ~new_new_n30434__;
  assign new_new_n30436__ = ~pi11 & ~new_new_n30430__;
  assign new_new_n30437__ = ~new_new_n30435__ & ~new_new_n30436__;
  assign new_new_n30438__ = ~new_new_n28939__ & ~new_new_n29391__;
  assign new_new_n30439__ = ~new_new_n28938__ & ~new_new_n30438__;
  assign new_new_n30440__ = new_new_n6991__ & ~new_new_n26888__;
  assign new_new_n30441__ = new_new_n6985__ & ~new_new_n26854__;
  assign new_new_n30442__ = ~new_new_n30440__ & ~new_new_n30441__;
  assign new_new_n30443__ = new_new_n6994__ & new_new_n26847__;
  assign new_new_n30444__ = new_new_n29424__ & new_new_n30443__;
  assign new_new_n30445__ = new_new_n30442__ & ~new_new_n30444__;
  assign new_new_n30446__ = ~pi14 & ~new_new_n30445__;
  assign new_new_n30447__ = ~new_new_n26847__ & ~new_new_n29423__;
  assign new_new_n30448__ = new_new_n6994__ & ~new_new_n30447__;
  assign new_new_n30449__ = ~pi13 & new_new_n29424__;
  assign new_new_n30450__ = pi13 & new_new_n26847__;
  assign new_new_n30451__ = new_new_n30448__ & ~new_new_n30450__;
  assign new_new_n30452__ = ~new_new_n30449__ & new_new_n30451__;
  assign new_new_n30453__ = pi14 & new_new_n30442__;
  assign new_new_n30454__ = ~new_new_n30448__ & new_new_n30453__;
  assign new_new_n30455__ = ~new_new_n30446__ & ~new_new_n30454__;
  assign new_new_n30456__ = ~new_new_n30452__ & new_new_n30455__;
  assign new_new_n30457__ = new_new_n7935__ & new_new_n26922__;
  assign new_new_n30458__ = new_new_n6968__ & ~new_new_n27168__;
  assign new_new_n30459__ = new_new_n6964__ & new_new_n26917__;
  assign new_new_n30460__ = new_new_n6959__ & ~new_new_n29366__;
  assign new_new_n30461__ = ~new_new_n30458__ & ~new_new_n30459__;
  assign new_new_n30462__ = ~new_new_n30457__ & new_new_n30461__;
  assign new_new_n30463__ = ~new_new_n30460__ & new_new_n30462__;
  assign new_new_n30464__ = ~new_new_n28807__ & new_new_n28934__;
  assign new_new_n30465__ = ~new_new_n28808__ & ~new_new_n30464__;
  assign new_new_n30466__ = new_new_n6634__ & new_new_n26928__;
  assign new_new_n30467__ = new_new_n6629__ & ~new_new_n26941__;
  assign new_new_n30468__ = ~new_new_n6625__ & new_new_n27152__;
  assign new_new_n30469__ = ~new_new_n30467__ & ~new_new_n30468__;
  assign new_new_n30470__ = ~new_new_n30466__ & new_new_n30469__;
  assign new_new_n30471__ = new_new_n6631__ & new_new_n27488__;
  assign new_new_n30472__ = pi20 & ~new_new_n30471__;
  assign new_new_n30473__ = new_new_n6640__ & new_new_n27488__;
  assign new_new_n30474__ = ~new_new_n30472__ & ~new_new_n30473__;
  assign new_new_n30475__ = new_new_n30470__ & ~new_new_n30474__;
  assign new_new_n30476__ = ~pi20 & ~new_new_n30470__;
  assign new_new_n30477__ = ~new_new_n30475__ & ~new_new_n30476__;
  assign new_new_n30478__ = new_new_n3311__ & ~new_new_n27003__;
  assign new_new_n30479__ = ~new_new_n333__ & ~new_new_n27021__;
  assign new_new_n30480__ = new_new_n873__ & ~new_new_n27029__;
  assign new_new_n30481__ = ~new_new_n30479__ & ~new_new_n30480__;
  assign new_new_n30482__ = ~new_new_n30478__ & new_new_n30481__;
  assign new_new_n30483__ = ~pi26 & ~new_new_n30482__;
  assign new_new_n30484__ = new_new_n512__ & new_new_n27962__;
  assign new_new_n30485__ = new_new_n801__ & new_new_n27962__;
  assign new_new_n30486__ = pi26 & ~new_new_n30485__;
  assign new_new_n30487__ = ~new_new_n30484__ & ~new_new_n30486__;
  assign new_new_n30488__ = new_new_n30482__ & ~new_new_n30487__;
  assign new_new_n30489__ = ~new_new_n30483__ & ~new_new_n30488__;
  assign new_new_n30490__ = ~new_new_n28834__ & ~new_new_n28903__;
  assign new_new_n30491__ = ~new_new_n28833__ & ~new_new_n30490__;
  assign new_new_n30492__ = ~new_new_n30489__ & ~new_new_n30491__;
  assign new_new_n30493__ = new_new_n30489__ & new_new_n30491__;
  assign new_new_n30494__ = ~new_new_n30492__ & ~new_new_n30493__;
  assign new_new_n30495__ = new_new_n4212__ & ~new_new_n27033__;
  assign new_new_n30496__ = ~new_new_n4818__ & ~new_new_n27054__;
  assign new_new_n30497__ = ~new_new_n30495__ & ~new_new_n30496__;
  assign new_new_n30498__ = new_new_n4214__ & new_new_n27687__;
  assign new_new_n30499__ = new_new_n30497__ & ~new_new_n30498__;
  assign new_new_n30500__ = pi29 & ~new_new_n30499__;
  assign new_new_n30501__ = new_new_n4214__ & ~new_new_n27691__;
  assign new_new_n30502__ = ~pi29 & ~new_new_n30501__;
  assign new_new_n30503__ = ~pi28 & new_new_n27111__;
  assign new_new_n30504__ = pi28 & ~new_new_n27111__;
  assign new_new_n30505__ = new_new_n4214__ & ~new_new_n30503__;
  assign new_new_n30506__ = ~new_new_n30504__ & new_new_n30505__;
  assign new_new_n30507__ = new_new_n27686__ & new_new_n30506__;
  assign new_new_n30508__ = ~new_new_n30502__ & ~new_new_n30507__;
  assign new_new_n30509__ = new_new_n30497__ & ~new_new_n30508__;
  assign new_new_n30510__ = ~new_new_n30500__ & ~new_new_n30509__;
  assign new_new_n30511__ = new_new_n161__ & ~new_new_n27071__;
  assign new_new_n30512__ = new_new_n765__ & new_new_n27041__;
  assign new_new_n30513__ = ~new_new_n30511__ & ~new_new_n30512__;
  assign new_new_n30514__ = ~pi31 & ~new_new_n30513__;
  assign new_new_n30515__ = new_new_n71__ & new_new_n27071__;
  assign new_new_n30516__ = ~new_new_n27071__ & new_new_n27559__;
  assign new_new_n30517__ = ~new_new_n27565__ & ~new_new_n30516__;
  assign new_new_n30518__ = ~new_new_n15853__ & ~new_new_n30517__;
  assign new_new_n30519__ = ~new_new_n161__ & ~new_new_n27083__;
  assign new_new_n30520__ = ~new_new_n27560__ & new_new_n30519__;
  assign new_new_n30521__ = ~new_new_n71__ & ~new_new_n27059__;
  assign new_new_n30522__ = ~new_new_n30520__ & new_new_n30521__;
  assign new_new_n30523__ = pi31 & ~new_new_n30515__;
  assign new_new_n30524__ = ~new_new_n30522__ & new_new_n30523__;
  assign new_new_n30525__ = ~new_new_n30518__ & new_new_n30524__;
  assign new_new_n30526__ = ~new_new_n30514__ & ~new_new_n30525__;
  assign new_new_n30527__ = ~new_new_n212__ & ~new_new_n692__;
  assign new_new_n30528__ = ~new_new_n311__ & new_new_n30527__;
  assign new_new_n30529__ = new_new_n4343__ & new_new_n5383__;
  assign new_new_n30530__ = new_new_n30528__ & new_new_n30529__;
  assign new_new_n30531__ = new_new_n743__ & new_new_n1508__;
  assign new_new_n30532__ = new_new_n4228__ & new_new_n7126__;
  assign new_new_n30533__ = new_new_n16812__ & new_new_n30532__;
  assign new_new_n30534__ = new_new_n30530__ & new_new_n30531__;
  assign new_new_n30535__ = new_new_n30533__ & new_new_n30534__;
  assign new_new_n30536__ = new_new_n16166__ & new_new_n30535__;
  assign new_new_n30537__ = new_new_n16234__ & new_new_n30536__;
  assign new_new_n30538__ = new_new_n16146__ & new_new_n30537__;
  assign new_new_n30539__ = new_new_n19399__ & new_new_n30538__;
  assign new_new_n30540__ = new_new_n30526__ & new_new_n30539__;
  assign new_new_n30541__ = ~new_new_n30526__ & ~new_new_n30539__;
  assign new_new_n30542__ = ~new_new_n30540__ & ~new_new_n30541__;
  assign new_new_n30543__ = ~new_new_n28875__ & ~new_new_n28892__;
  assign new_new_n30544__ = ~new_new_n28874__ & ~new_new_n30543__;
  assign new_new_n30545__ = ~new_new_n30542__ & new_new_n30544__;
  assign new_new_n30546__ = ~new_new_n30540__ & ~new_new_n30544__;
  assign new_new_n30547__ = ~new_new_n30541__ & new_new_n30546__;
  assign new_new_n30548__ = ~new_new_n30545__ & ~new_new_n30547__;
  assign new_new_n30549__ = ~new_new_n30510__ & ~new_new_n30548__;
  assign new_new_n30550__ = new_new_n30510__ & new_new_n30548__;
  assign new_new_n30551__ = ~new_new_n30549__ & ~new_new_n30550__;
  assign new_new_n30552__ = ~new_new_n28851__ & ~new_new_n28899__;
  assign new_new_n30553__ = ~new_new_n28898__ & ~new_new_n30552__;
  assign new_new_n30554__ = new_new_n30551__ & ~new_new_n30553__;
  assign new_new_n30555__ = ~new_new_n30551__ & new_new_n30553__;
  assign new_new_n30556__ = ~new_new_n30554__ & ~new_new_n30555__;
  assign new_new_n30557__ = ~new_new_n30494__ & ~new_new_n30556__;
  assign new_new_n30558__ = ~new_new_n30493__ & new_new_n30556__;
  assign new_new_n30559__ = ~new_new_n30492__ & new_new_n30558__;
  assign new_new_n30560__ = ~new_new_n30557__ & ~new_new_n30559__;
  assign new_new_n30561__ = new_new_n5215__ & new_new_n28005__;
  assign new_new_n30562__ = new_new_n5191__ & ~new_new_n26978__;
  assign new_new_n30563__ = new_new_n5183__ & new_new_n26971__;
  assign new_new_n30564__ = ~new_new_n30562__ & ~new_new_n30563__;
  assign new_new_n30565__ = ~new_new_n30561__ & new_new_n30564__;
  assign new_new_n30566__ = new_new_n5195__ & ~new_new_n26937__;
  assign new_new_n30567__ = ~pi23 & ~new_new_n30566__;
  assign new_new_n30568__ = new_new_n7878__ & ~new_new_n26937__;
  assign new_new_n30569__ = ~new_new_n30567__ & ~new_new_n30568__;
  assign new_new_n30570__ = new_new_n30565__ & ~new_new_n30569__;
  assign new_new_n30571__ = pi23 & ~new_new_n30565__;
  assign new_new_n30572__ = ~new_new_n30570__ & ~new_new_n30571__;
  assign new_new_n30573__ = ~new_new_n28907__ & ~new_new_n28911__;
  assign new_new_n30574__ = ~new_new_n28908__ & ~new_new_n30573__;
  assign new_new_n30575__ = ~new_new_n30572__ & new_new_n30574__;
  assign new_new_n30576__ = new_new_n30572__ & ~new_new_n30574__;
  assign new_new_n30577__ = ~new_new_n30575__ & ~new_new_n30576__;
  assign new_new_n30578__ = ~new_new_n30560__ & new_new_n30577__;
  assign new_new_n30579__ = new_new_n30560__ & ~new_new_n30577__;
  assign new_new_n30580__ = ~new_new_n30578__ & ~new_new_n30579__;
  assign new_new_n30581__ = ~new_new_n30477__ & ~new_new_n30580__;
  assign new_new_n30582__ = new_new_n30477__ & new_new_n30580__;
  assign new_new_n30583__ = ~new_new_n30581__ & ~new_new_n30582__;
  assign new_new_n30584__ = ~new_new_n28917__ & ~new_new_n28931__;
  assign new_new_n30585__ = ~new_new_n28918__ & ~new_new_n30584__;
  assign new_new_n30586__ = new_new_n30583__ & ~new_new_n30585__;
  assign new_new_n30587__ = ~new_new_n30583__ & new_new_n30585__;
  assign new_new_n30588__ = ~new_new_n30586__ & ~new_new_n30587__;
  assign new_new_n30589__ = pi17 & ~new_new_n30588__;
  assign new_new_n30590__ = ~pi17 & new_new_n30588__;
  assign new_new_n30591__ = ~new_new_n30589__ & ~new_new_n30590__;
  assign new_new_n30592__ = new_new_n30465__ & ~new_new_n30591__;
  assign new_new_n30593__ = ~new_new_n30465__ & new_new_n30591__;
  assign new_new_n30594__ = ~new_new_n30592__ & ~new_new_n30593__;
  assign new_new_n30595__ = new_new_n30463__ & new_new_n30594__;
  assign new_new_n30596__ = ~new_new_n30463__ & ~new_new_n30594__;
  assign new_new_n30597__ = ~new_new_n30595__ & ~new_new_n30596__;
  assign new_new_n30598__ = ~new_new_n30456__ & new_new_n30597__;
  assign new_new_n30599__ = new_new_n30456__ & ~new_new_n30597__;
  assign new_new_n30600__ = ~new_new_n30598__ & ~new_new_n30599__;
  assign new_new_n30601__ = new_new_n30439__ & new_new_n30600__;
  assign new_new_n30602__ = ~new_new_n30439__ & ~new_new_n30600__;
  assign new_new_n30603__ = ~new_new_n30601__ & ~new_new_n30602__;
  assign new_new_n30604__ = new_new_n30437__ & new_new_n30603__;
  assign new_new_n30605__ = ~new_new_n30437__ & ~new_new_n30603__;
  assign new_new_n30606__ = ~new_new_n30604__ & ~new_new_n30605__;
  assign new_new_n30607__ = ~new_new_n29854__ & ~new_new_n29861__;
  assign new_new_n30608__ = ~new_new_n29853__ & ~new_new_n30607__;
  assign new_new_n30609__ = ~new_new_n30606__ & new_new_n30608__;
  assign new_new_n30610__ = new_new_n30606__ & ~new_new_n30608__;
  assign new_new_n30611__ = ~new_new_n30609__ & ~new_new_n30610__;
  assign new_new_n30612__ = new_new_n30425__ & new_new_n30611__;
  assign new_new_n30613__ = ~new_new_n30425__ & ~new_new_n30611__;
  assign new_new_n30614__ = ~new_new_n30612__ & ~new_new_n30613__;
  assign new_new_n30615__ = ~new_new_n27367__ & ~new_new_n30614__;
  assign new_new_n30616__ = new_new_n27367__ & new_new_n30614__;
  assign new_new_n30617__ = new_new_n11475__ & new_new_n26774__;
  assign new_new_n30618__ = new_new_n11471__ & new_new_n26810__;
  assign new_new_n30619__ = new_new_n12850__ & new_new_n26729__;
  assign new_new_n30620__ = ~new_new_n30617__ & ~new_new_n30618__;
  assign new_new_n30621__ = ~new_new_n30619__ & new_new_n30620__;
  assign new_new_n30622__ = pi05 & ~new_new_n30621__;
  assign new_new_n30623__ = ~new_new_n26729__ & new_new_n27370__;
  assign new_new_n30624__ = ~new_new_n26729__ & new_new_n26810__;
  assign new_new_n30625__ = new_new_n26802__ & new_new_n30624__;
  assign new_new_n30626__ = new_new_n26729__ & new_new_n27368__;
  assign new_new_n30627__ = ~new_new_n27226__ & new_new_n30626__;
  assign new_new_n30628__ = ~new_new_n30625__ & ~new_new_n30627__;
  assign new_new_n30629__ = new_new_n26741__ & ~new_new_n30628__;
  assign new_new_n30630__ = ~new_new_n26802__ & new_new_n26811__;
  assign new_new_n30631__ = ~new_new_n26774__ & new_new_n27230__;
  assign new_new_n30632__ = new_new_n27226__ & new_new_n30631__;
  assign new_new_n30633__ = ~new_new_n30630__ & ~new_new_n30632__;
  assign new_new_n30634__ = ~new_new_n26741__ & ~new_new_n30633__;
  assign new_new_n30635__ = new_new_n26811__ & new_new_n27226__;
  assign new_new_n30636__ = ~new_new_n30631__ & ~new_new_n30635__;
  assign new_new_n30637__ = ~new_new_n26802__ & ~new_new_n30636__;
  assign new_new_n30638__ = ~new_new_n27226__ & new_new_n30624__;
  assign new_new_n30639__ = ~new_new_n30626__ & ~new_new_n30638__;
  assign new_new_n30640__ = new_new_n26802__ & ~new_new_n30639__;
  assign new_new_n30641__ = ~new_new_n30637__ & ~new_new_n30640__;
  assign new_new_n30642__ = ~new_new_n30629__ & new_new_n30641__;
  assign new_new_n30643__ = ~new_new_n30634__ & new_new_n30642__;
  assign new_new_n30644__ = ~new_new_n30623__ & new_new_n30643__;
  assign new_new_n30645__ = new_new_n12856__ & new_new_n30644__;
  assign new_new_n30646__ = new_new_n11469__ & new_new_n30644__;
  assign new_new_n30647__ = ~pi05 & ~new_new_n30646__;
  assign new_new_n30648__ = ~new_new_n30645__ & ~new_new_n30647__;
  assign new_new_n30649__ = new_new_n30621__ & ~new_new_n30648__;
  assign new_new_n30650__ = ~new_new_n30622__ & ~new_new_n30649__;
  assign new_new_n30651__ = new_new_n13111__ & ~new_new_n26802__;
  assign new_new_n30652__ = new_new_n11469__ & ~new_new_n27373__;
  assign new_new_n30653__ = ~new_new_n30651__ & ~new_new_n30652__;
  assign new_new_n30654__ = new_new_n11478__ & ~new_new_n30653__;
  assign new_new_n30655__ = new_new_n11475__ & new_new_n26810__;
  assign new_new_n30656__ = ~new_new_n30654__ & ~new_new_n30655__;
  assign new_new_n30657__ = pi05 & ~new_new_n30656__;
  assign new_new_n30658__ = new_new_n12873__ & new_new_n26774__;
  assign new_new_n30659__ = new_new_n11469__ & new_new_n26774__;
  assign new_new_n30660__ = ~pi05 & ~new_new_n30659__;
  assign new_new_n30661__ = ~new_new_n30658__ & ~new_new_n30660__;
  assign new_new_n30662__ = new_new_n30656__ & ~new_new_n30661__;
  assign new_new_n30663__ = ~new_new_n30657__ & ~new_new_n30662__;
  assign new_new_n30664__ = ~new_new_n30382__ & ~new_new_n30383__;
  assign new_new_n30665__ = ~new_new_n30400__ & ~new_new_n30664__;
  assign new_new_n30666__ = new_new_n30400__ & new_new_n30664__;
  assign new_new_n30667__ = ~new_new_n30665__ & ~new_new_n30666__;
  assign new_new_n30668__ = new_new_n30663__ & new_new_n30667__;
  assign new_new_n30669__ = ~new_new_n30663__ & ~new_new_n30667__;
  assign new_new_n30670__ = new_new_n11475__ & ~new_new_n26802__;
  assign new_new_n30671__ = ~new_new_n11478__ & ~new_new_n26810__;
  assign new_new_n30672__ = new_new_n11478__ & ~new_new_n27395__;
  assign new_new_n30673__ = ~new_new_n11482__ & ~new_new_n30671__;
  assign new_new_n30674__ = ~new_new_n30672__ & new_new_n30673__;
  assign new_new_n30675__ = ~new_new_n30670__ & ~new_new_n30674__;
  assign new_new_n30676__ = ~pi05 & ~new_new_n30675__;
  assign new_new_n30677__ = new_new_n12830__ & ~new_new_n26741__;
  assign new_new_n30678__ = pi05 & ~new_new_n30677__;
  assign new_new_n30679__ = new_new_n12828__ & ~new_new_n26741__;
  assign new_new_n30680__ = ~new_new_n30678__ & ~new_new_n30679__;
  assign new_new_n30681__ = new_new_n30675__ & ~new_new_n30680__;
  assign new_new_n30682__ = ~new_new_n30676__ & ~new_new_n30681__;
  assign new_new_n30683__ = new_new_n12832__ & ~new_new_n27221__;
  assign new_new_n30684__ = new_new_n11475__ & ~new_new_n26741__;
  assign new_new_n30685__ = ~new_new_n30683__ & ~new_new_n30684__;
  assign new_new_n30686__ = ~new_new_n11482__ & ~new_new_n26802__;
  assign new_new_n30687__ = new_new_n30411__ & new_new_n30686__;
  assign new_new_n30688__ = new_new_n30685__ & ~new_new_n30687__;
  assign new_new_n30689__ = pi05 & ~new_new_n30688__;
  assign new_new_n30690__ = new_new_n11469__ & ~new_new_n27391__;
  assign new_new_n30691__ = ~pi05 & ~new_new_n30690__;
  assign new_new_n30692__ = new_new_n26802__ & new_new_n27390__;
  assign new_new_n30693__ = ~pi04 & ~new_new_n30692__;
  assign new_new_n30694__ = pi04 & ~new_new_n30410__;
  assign new_new_n30695__ = ~new_new_n11482__ & ~new_new_n30693__;
  assign new_new_n30696__ = ~new_new_n30694__ & new_new_n30695__;
  assign new_new_n30697__ = ~new_new_n30691__ & ~new_new_n30696__;
  assign new_new_n30698__ = new_new_n30685__ & ~new_new_n30697__;
  assign new_new_n30699__ = ~new_new_n30689__ & ~new_new_n30698__;
  assign new_new_n30700__ = ~new_new_n29893__ & ~new_new_n30315__;
  assign new_new_n30701__ = new_new_n29893__ & new_new_n30315__;
  assign new_new_n30702__ = ~new_new_n30700__ & ~new_new_n30701__;
  assign new_new_n30703__ = ~pi08 & new_new_n29911__;
  assign new_new_n30704__ = ~new_new_n29913__ & ~new_new_n30703__;
  assign new_new_n30705__ = new_new_n30702__ & new_new_n30704__;
  assign new_new_n30706__ = ~new_new_n30702__ & ~new_new_n30704__;
  assign new_new_n30707__ = ~new_new_n30705__ & ~new_new_n30706__;
  assign new_new_n30708__ = ~new_new_n30302__ & ~new_new_n30303__;
  assign new_new_n30709__ = new_new_n30313__ & new_new_n30708__;
  assign new_new_n30710__ = ~new_new_n30313__ & ~new_new_n30708__;
  assign new_new_n30711__ = ~new_new_n30709__ & ~new_new_n30710__;
  assign new_new_n30712__ = ~new_new_n30284__ & ~new_new_n30285__;
  assign new_new_n30713__ = ~new_new_n30289__ & new_new_n30712__;
  assign new_new_n30714__ = new_new_n30289__ & ~new_new_n30712__;
  assign new_new_n30715__ = ~new_new_n30713__ & ~new_new_n30714__;
  assign new_new_n30716__ = ~new_new_n30252__ & ~new_new_n30253__;
  assign new_new_n30717__ = ~new_new_n30263__ & new_new_n30716__;
  assign new_new_n30718__ = new_new_n30263__ & ~new_new_n30716__;
  assign new_new_n30719__ = ~new_new_n30717__ & ~new_new_n30718__;
  assign new_new_n30720__ = new_new_n11475__ & new_new_n26917__;
  assign new_new_n30721__ = new_new_n11471__ & new_new_n26928__;
  assign new_new_n30722__ = new_new_n12850__ & ~new_new_n27168__;
  assign new_new_n30723__ = ~new_new_n30721__ & ~new_new_n30722__;
  assign new_new_n30724__ = ~new_new_n30720__ & new_new_n30723__;
  assign new_new_n30725__ = pi05 & ~new_new_n30724__;
  assign new_new_n30726__ = new_new_n12856__ & ~new_new_n28799__;
  assign new_new_n30727__ = new_new_n11469__ & ~new_new_n28799__;
  assign new_new_n30728__ = ~pi05 & ~new_new_n30727__;
  assign new_new_n30729__ = ~new_new_n30726__ & ~new_new_n30728__;
  assign new_new_n30730__ = new_new_n30724__ & ~new_new_n30729__;
  assign new_new_n30731__ = ~new_new_n30725__ & ~new_new_n30730__;
  assign new_new_n30732__ = new_new_n13069__ & ~new_new_n27462__;
  assign new_new_n30733__ = new_new_n11475__ & new_new_n26928__;
  assign new_new_n30734__ = ~new_new_n30732__ & ~new_new_n30733__;
  assign new_new_n30735__ = new_new_n11471__ & ~new_new_n26941__;
  assign new_new_n30736__ = new_new_n12850__ & new_new_n26917__;
  assign new_new_n30737__ = ~new_new_n30735__ & ~new_new_n30736__;
  assign new_new_n30738__ = new_new_n30734__ & new_new_n30737__;
  assign new_new_n30739__ = pi05 & ~new_new_n30738__;
  assign new_new_n30740__ = ~new_new_n11471__ & ~new_new_n26917__;
  assign new_new_n30741__ = new_new_n12850__ & ~new_new_n30740__;
  assign new_new_n30742__ = ~pi05 & ~new_new_n30735__;
  assign new_new_n30743__ = ~new_new_n30741__ & new_new_n30742__;
  assign new_new_n30744__ = new_new_n30734__ & new_new_n30743__;
  assign new_new_n30745__ = ~new_new_n30739__ & ~new_new_n30744__;
  assign new_new_n30746__ = ~new_new_n29969__ & ~new_new_n29970__;
  assign new_new_n30747__ = ~new_new_n30228__ & new_new_n30746__;
  assign new_new_n30748__ = new_new_n30228__ & ~new_new_n30746__;
  assign new_new_n30749__ = ~new_new_n30747__ & ~new_new_n30748__;
  assign new_new_n30750__ = new_new_n30745__ & new_new_n30749__;
  assign new_new_n30751__ = ~new_new_n30745__ & ~new_new_n30749__;
  assign new_new_n30752__ = new_new_n11471__ & new_new_n27152__;
  assign new_new_n30753__ = new_new_n11475__ & ~new_new_n26941__;
  assign new_new_n30754__ = new_new_n12850__ & new_new_n26928__;
  assign new_new_n30755__ = ~new_new_n30752__ & ~new_new_n30753__;
  assign new_new_n30756__ = ~new_new_n30754__ & new_new_n30755__;
  assign new_new_n30757__ = pi05 & ~new_new_n30756__;
  assign new_new_n30758__ = new_new_n12856__ & new_new_n27488__;
  assign new_new_n30759__ = new_new_n11469__ & new_new_n27488__;
  assign new_new_n30760__ = ~pi05 & ~new_new_n30759__;
  assign new_new_n30761__ = ~new_new_n30758__ & ~new_new_n30760__;
  assign new_new_n30762__ = new_new_n30756__ & ~new_new_n30761__;
  assign new_new_n30763__ = ~new_new_n30757__ & ~new_new_n30762__;
  assign new_new_n30764__ = ~pi05 & new_new_n12873__;
  assign new_new_n30765__ = new_new_n27152__ & new_new_n30764__;
  assign new_new_n30766__ = new_new_n12850__ & new_new_n27152__;
  assign new_new_n30767__ = new_new_n11471__ & new_new_n26971__;
  assign new_new_n30768__ = new_new_n11475__ & ~new_new_n26937__;
  assign new_new_n30769__ = ~new_new_n30767__ & ~new_new_n30768__;
  assign new_new_n30770__ = ~new_new_n30766__ & new_new_n30769__;
  assign new_new_n30771__ = pi05 & ~new_new_n27152__;
  assign new_new_n30772__ = new_new_n30770__ & new_new_n30771__;
  assign new_new_n30773__ = ~new_new_n30765__ & ~new_new_n30772__;
  assign new_new_n30774__ = ~new_new_n27477__ & ~new_new_n30773__;
  assign new_new_n30775__ = ~new_new_n27152__ & new_new_n30764__;
  assign new_new_n30776__ = pi05 & new_new_n27152__;
  assign new_new_n30777__ = new_new_n30770__ & new_new_n30776__;
  assign new_new_n30778__ = ~new_new_n30775__ & ~new_new_n30777__;
  assign new_new_n30779__ = new_new_n27477__ & ~new_new_n30778__;
  assign new_new_n30780__ = ~pi05 & ~new_new_n30770__;
  assign new_new_n30781__ = pi05 & ~new_new_n12856__;
  assign new_new_n30782__ = new_new_n30770__ & new_new_n30781__;
  assign new_new_n30783__ = ~new_new_n30780__ & ~new_new_n30782__;
  assign new_new_n30784__ = ~new_new_n30774__ & new_new_n30783__;
  assign new_new_n30785__ = ~new_new_n30779__ & new_new_n30784__;
  assign new_new_n30786__ = ~new_new_n30186__ & ~new_new_n30187__;
  assign new_new_n30787__ = pi08 & ~new_new_n30194__;
  assign new_new_n30788__ = ~pi08 & new_new_n30194__;
  assign new_new_n30789__ = ~new_new_n30787__ & ~new_new_n30788__;
  assign new_new_n30790__ = new_new_n30786__ & new_new_n30789__;
  assign new_new_n30791__ = ~new_new_n30786__ & ~new_new_n30789__;
  assign new_new_n30792__ = ~new_new_n30790__ & ~new_new_n30791__;
  assign new_new_n30793__ = new_new_n30785__ & ~new_new_n30792__;
  assign new_new_n30794__ = ~new_new_n30785__ & new_new_n30792__;
  assign new_new_n30795__ = ~new_new_n30170__ & ~new_new_n30171__;
  assign new_new_n30796__ = new_new_n30183__ & new_new_n30795__;
  assign new_new_n30797__ = ~new_new_n30183__ & ~new_new_n30795__;
  assign new_new_n30798__ = ~new_new_n30796__ & ~new_new_n30797__;
  assign new_new_n30799__ = new_new_n12850__ & new_new_n26971__;
  assign new_new_n30800__ = new_new_n11471__ & ~new_new_n27003__;
  assign new_new_n30801__ = new_new_n11475__ & ~new_new_n26978__;
  assign new_new_n30802__ = ~new_new_n30800__ & ~new_new_n30801__;
  assign new_new_n30803__ = ~new_new_n30799__ & new_new_n30802__;
  assign new_new_n30804__ = ~pi05 & ~new_new_n30803__;
  assign new_new_n30805__ = new_new_n12873__ & new_new_n28277__;
  assign new_new_n30806__ = new_new_n11469__ & new_new_n28277__;
  assign new_new_n30807__ = pi05 & ~new_new_n30806__;
  assign new_new_n30808__ = ~new_new_n30805__ & ~new_new_n30807__;
  assign new_new_n30809__ = new_new_n30803__ & ~new_new_n30808__;
  assign new_new_n30810__ = ~new_new_n30804__ & ~new_new_n30809__;
  assign new_new_n30811__ = ~new_new_n30158__ & ~new_new_n30159__;
  assign new_new_n30812__ = new_new_n30163__ & new_new_n30811__;
  assign new_new_n30813__ = ~new_new_n30163__ & ~new_new_n30811__;
  assign new_new_n30814__ = ~new_new_n30812__ & ~new_new_n30813__;
  assign new_new_n30815__ = new_new_n30810__ & ~new_new_n30814__;
  assign new_new_n30816__ = ~new_new_n30810__ & new_new_n30814__;
  assign new_new_n30817__ = new_new_n12832__ & ~new_new_n27029__;
  assign new_new_n30818__ = new_new_n11475__ & ~new_new_n27003__;
  assign new_new_n30819__ = ~new_new_n30817__ & ~new_new_n30818__;
  assign new_new_n30820__ = new_new_n11469__ & new_new_n27992__;
  assign new_new_n30821__ = new_new_n30819__ & ~new_new_n30820__;
  assign new_new_n30822__ = pi05 & ~new_new_n30821__;
  assign new_new_n30823__ = new_new_n11469__ & ~new_new_n27996__;
  assign new_new_n30824__ = ~pi05 & ~new_new_n30823__;
  assign new_new_n30825__ = ~pi04 & ~new_new_n29034__;
  assign new_new_n30826__ = pi04 & ~new_new_n29032__;
  assign new_new_n30827__ = ~new_new_n11482__ & ~new_new_n30825__;
  assign new_new_n30828__ = ~new_new_n30826__ & new_new_n30827__;
  assign new_new_n30829__ = ~new_new_n30824__ & ~new_new_n30828__;
  assign new_new_n30830__ = new_new_n30819__ & ~new_new_n30829__;
  assign new_new_n30831__ = ~new_new_n30822__ & ~new_new_n30830__;
  assign new_new_n30832__ = ~new_new_n30020__ & new_new_n30033__;
  assign new_new_n30833__ = new_new_n30020__ & ~new_new_n30033__;
  assign new_new_n30834__ = ~new_new_n30832__ & ~new_new_n30833__;
  assign new_new_n30835__ = new_new_n29615__ & ~new_new_n30135__;
  assign new_new_n30836__ = ~new_new_n29615__ & ~new_new_n30137__;
  assign new_new_n30837__ = ~new_new_n30835__ & ~new_new_n30836__;
  assign new_new_n30838__ = ~new_new_n30033__ & new_new_n30136__;
  assign new_new_n30839__ = new_new_n30837__ & ~new_new_n30838__;
  assign new_new_n30840__ = new_new_n30834__ & ~new_new_n30839__;
  assign new_new_n30841__ = ~new_new_n30834__ & new_new_n30837__;
  assign new_new_n30842__ = ~new_new_n30840__ & ~new_new_n30841__;
  assign new_new_n30843__ = new_new_n12832__ & ~new_new_n27033__;
  assign new_new_n30844__ = new_new_n11475__ & new_new_n27111__;
  assign new_new_n30845__ = ~new_new_n30843__ & ~new_new_n30844__;
  assign new_new_n30846__ = ~new_new_n11482__ & ~new_new_n27021__;
  assign new_new_n30847__ = new_new_n27796__ & new_new_n30846__;
  assign new_new_n30848__ = new_new_n30845__ & ~new_new_n30847__;
  assign new_new_n30849__ = pi05 & ~new_new_n30848__;
  assign new_new_n30850__ = new_new_n11469__ & ~new_new_n29228__;
  assign new_new_n30851__ = ~pi05 & ~new_new_n30850__;
  assign new_new_n30852__ = ~pi04 & ~new_new_n29224__;
  assign new_new_n30853__ = pi04 & ~new_new_n29222__;
  assign new_new_n30854__ = ~new_new_n11482__ & ~new_new_n30853__;
  assign new_new_n30855__ = ~new_new_n30852__ & new_new_n30854__;
  assign new_new_n30856__ = ~new_new_n30851__ & ~new_new_n30855__;
  assign new_new_n30857__ = new_new_n30845__ & ~new_new_n30856__;
  assign new_new_n30858__ = ~new_new_n30849__ & ~new_new_n30857__;
  assign new_new_n30859__ = new_new_n12832__ & ~new_new_n27054__;
  assign new_new_n30860__ = new_new_n11475__ & ~new_new_n27033__;
  assign new_new_n30861__ = ~new_new_n30859__ & ~new_new_n30860__;
  assign new_new_n30862__ = new_new_n11469__ & ~new_new_n27691__;
  assign new_new_n30863__ = pi05 & ~new_new_n30862__;
  assign new_new_n30864__ = pi04 & new_new_n27111__;
  assign new_new_n30865__ = ~pi04 & ~new_new_n27111__;
  assign new_new_n30866__ = ~new_new_n11482__ & ~new_new_n30864__;
  assign new_new_n30867__ = ~new_new_n30865__ & new_new_n30866__;
  assign new_new_n30868__ = new_new_n27686__ & new_new_n30867__;
  assign new_new_n30869__ = ~new_new_n30863__ & ~new_new_n30868__;
  assign new_new_n30870__ = new_new_n30861__ & ~new_new_n30869__;
  assign new_new_n30871__ = new_new_n11469__ & new_new_n27687__;
  assign new_new_n30872__ = new_new_n30861__ & ~new_new_n30871__;
  assign new_new_n30873__ = ~pi05 & ~new_new_n30872__;
  assign new_new_n30874__ = ~new_new_n30870__ & ~new_new_n30873__;
  assign new_new_n30875__ = ~new_new_n30091__ & ~new_new_n30092__;
  assign new_new_n30876__ = ~new_new_n30102__ & new_new_n30875__;
  assign new_new_n30877__ = new_new_n30102__ & ~new_new_n30875__;
  assign new_new_n30878__ = ~new_new_n30876__ & ~new_new_n30877__;
  assign new_new_n30879__ = ~new_new_n30874__ & ~new_new_n30878__;
  assign new_new_n30880__ = new_new_n30874__ & new_new_n30878__;
  assign new_new_n30881__ = new_new_n12832__ & new_new_n27041__;
  assign new_new_n30882__ = new_new_n11475__ & ~new_new_n27054__;
  assign new_new_n30883__ = ~new_new_n30881__ & ~new_new_n30882__;
  assign new_new_n30884__ = new_new_n11469__ & ~new_new_n27535__;
  assign new_new_n30885__ = pi05 & ~new_new_n30884__;
  assign new_new_n30886__ = ~pi04 & new_new_n27033__;
  assign new_new_n30887__ = pi04 & ~new_new_n27033__;
  assign new_new_n30888__ = ~new_new_n11482__ & ~new_new_n30886__;
  assign new_new_n30889__ = ~new_new_n30887__ & new_new_n30888__;
  assign new_new_n30890__ = ~new_new_n27102__ & new_new_n30889__;
  assign new_new_n30891__ = ~new_new_n30885__ & ~new_new_n30890__;
  assign new_new_n30892__ = new_new_n30883__ & ~new_new_n30891__;
  assign new_new_n30893__ = new_new_n11469__ & new_new_n27545__;
  assign new_new_n30894__ = new_new_n30883__ & ~new_new_n30893__;
  assign new_new_n30895__ = ~pi05 & ~new_new_n30894__;
  assign new_new_n30896__ = ~new_new_n30892__ & ~new_new_n30895__;
  assign new_new_n30897__ = ~new_new_n30054__ & ~new_new_n30081__;
  assign new_new_n30898__ = new_new_n30068__ & ~new_new_n30897__;
  assign new_new_n30899__ = new_new_n12850__ & new_new_n27041__;
  assign new_new_n30900__ = new_new_n11471__ & new_new_n27059__;
  assign new_new_n30901__ = new_new_n11475__ & ~new_new_n27071__;
  assign new_new_n30902__ = ~new_new_n30899__ & ~new_new_n30900__;
  assign new_new_n30903__ = ~new_new_n30901__ & new_new_n30902__;
  assign new_new_n30904__ = pi05 & ~new_new_n30903__;
  assign new_new_n30905__ = new_new_n12856__ & new_new_n27567__;
  assign new_new_n30906__ = new_new_n11469__ & new_new_n27567__;
  assign new_new_n30907__ = ~pi05 & ~new_new_n30906__;
  assign new_new_n30908__ = ~new_new_n30905__ & ~new_new_n30907__;
  assign new_new_n30909__ = new_new_n30903__ & ~new_new_n30908__;
  assign new_new_n30910__ = ~new_new_n30904__ & ~new_new_n30909__;
  assign new_new_n30911__ = new_new_n11475__ & new_new_n27059__;
  assign new_new_n30912__ = new_new_n11478__ & new_new_n28441__;
  assign new_new_n30913__ = new_new_n27071__ & ~new_new_n30912__;
  assign new_new_n30914__ = ~new_new_n27071__ & new_new_n30912__;
  assign new_new_n30915__ = new_new_n11469__ & ~new_new_n30913__;
  assign new_new_n30916__ = ~new_new_n30914__ & new_new_n30915__;
  assign new_new_n30917__ = ~new_new_n30911__ & ~new_new_n30916__;
  assign new_new_n30918__ = ~pi05 & ~new_new_n30917__;
  assign new_new_n30919__ = new_new_n12830__ & new_new_n26118__;
  assign new_new_n30920__ = pi05 & ~new_new_n30919__;
  assign new_new_n30921__ = new_new_n12828__ & new_new_n26118__;
  assign new_new_n30922__ = ~new_new_n30920__ & ~new_new_n30921__;
  assign new_new_n30923__ = new_new_n30917__ & ~new_new_n30922__;
  assign new_new_n30924__ = ~new_new_n30918__ & ~new_new_n30923__;
  assign new_new_n30925__ = new_new_n10694__ & ~new_new_n27075__;
  assign new_new_n30926__ = new_new_n11469__ & new_new_n26118__;
  assign new_new_n30927__ = new_new_n27075__ & ~new_new_n30926__;
  assign new_new_n30928__ = ~new_new_n13111__ & ~new_new_n30927__;
  assign new_new_n30929__ = new_new_n13069__ & new_new_n27553__;
  assign new_new_n30930__ = new_new_n13082__ & ~new_new_n30929__;
  assign new_new_n30931__ = new_new_n26118__ & ~new_new_n30930__;
  assign new_new_n30932__ = ~new_new_n11482__ & new_new_n27059__;
  assign new_new_n30933__ = new_new_n11471__ & ~new_new_n27075__;
  assign new_new_n30934__ = ~new_new_n30932__ & ~new_new_n30933__;
  assign new_new_n30935__ = new_new_n11478__ & new_new_n27075__;
  assign new_new_n30936__ = new_new_n26118__ & new_new_n30935__;
  assign new_new_n30937__ = ~new_new_n30934__ & ~new_new_n30936__;
  assign new_new_n30938__ = ~new_new_n30931__ & ~new_new_n30937__;
  assign new_new_n30939__ = pi05 & ~new_new_n30928__;
  assign new_new_n30940__ = new_new_n30938__ & new_new_n30939__;
  assign new_new_n30941__ = ~new_new_n30925__ & ~new_new_n30940__;
  assign new_new_n30942__ = ~new_new_n30924__ & ~new_new_n30941__;
  assign new_new_n30943__ = ~new_new_n30910__ & ~new_new_n30942__;
  assign new_new_n30944__ = new_new_n30910__ & new_new_n30942__;
  assign new_new_n30945__ = new_new_n10700__ & new_new_n27087__;
  assign new_new_n30946__ = ~new_new_n10694__ & new_new_n27582__;
  assign new_new_n30947__ = ~new_new_n9697__ & new_new_n26118__;
  assign new_new_n30948__ = new_new_n10701__ & ~new_new_n30947__;
  assign new_new_n30949__ = ~new_new_n17566__ & ~new_new_n27577__;
  assign new_new_n30950__ = ~new_new_n30945__ & new_new_n30949__;
  assign new_new_n30951__ = ~new_new_n30946__ & ~new_new_n30948__;
  assign new_new_n30952__ = new_new_n30950__ & new_new_n30951__;
  assign new_new_n30953__ = ~new_new_n30944__ & ~new_new_n30952__;
  assign new_new_n30954__ = ~new_new_n30943__ & ~new_new_n30953__;
  assign new_new_n30955__ = new_new_n13064__ & ~new_new_n30056__;
  assign new_new_n30956__ = new_new_n30066__ & ~new_new_n30955__;
  assign new_new_n30957__ = pi08 & new_new_n30057__;
  assign new_new_n30958__ = ~new_new_n30066__ & new_new_n30957__;
  assign new_new_n30959__ = ~new_new_n30956__ & ~new_new_n30958__;
  assign new_new_n30960__ = ~new_new_n30954__ & ~new_new_n30959__;
  assign new_new_n30961__ = new_new_n30954__ & new_new_n30959__;
  assign new_new_n30962__ = new_new_n13069__ & ~new_new_n27094__;
  assign new_new_n30963__ = new_new_n12850__ & ~new_new_n27054__;
  assign new_new_n30964__ = new_new_n11471__ & ~new_new_n27071__;
  assign new_new_n30965__ = new_new_n11475__ & new_new_n27041__;
  assign new_new_n30966__ = ~new_new_n30964__ & ~new_new_n30965__;
  assign new_new_n30967__ = ~new_new_n30963__ & new_new_n30966__;
  assign new_new_n30968__ = ~new_new_n30962__ & new_new_n30967__;
  assign new_new_n30969__ = pi05 & ~new_new_n30968__;
  assign new_new_n30970__ = ~pi05 & new_new_n30968__;
  assign new_new_n30971__ = ~new_new_n30969__ & ~new_new_n30970__;
  assign new_new_n30972__ = ~new_new_n30961__ & ~new_new_n30971__;
  assign new_new_n30973__ = ~new_new_n30960__ & ~new_new_n30972__;
  assign new_new_n30974__ = ~new_new_n30898__ & ~new_new_n30973__;
  assign new_new_n30975__ = ~new_new_n30896__ & ~new_new_n30974__;
  assign new_new_n30976__ = new_new_n30896__ & ~new_new_n30973__;
  assign new_new_n30977__ = ~new_new_n30054__ & new_new_n30081__;
  assign new_new_n30978__ = ~new_new_n30082__ & ~new_new_n30977__;
  assign new_new_n30979__ = ~new_new_n30976__ & new_new_n30978__;
  assign new_new_n30980__ = ~new_new_n30975__ & ~new_new_n30979__;
  assign new_new_n30981__ = ~new_new_n30880__ & ~new_new_n30980__;
  assign new_new_n30982__ = ~new_new_n30879__ & ~new_new_n30981__;
  assign new_new_n30983__ = ~new_new_n30858__ & new_new_n30982__;
  assign new_new_n30984__ = new_new_n30858__ & ~new_new_n30982__;
  assign new_new_n30985__ = ~new_new_n30105__ & ~new_new_n30106__;
  assign new_new_n30986__ = new_new_n30118__ & ~new_new_n30985__;
  assign new_new_n30987__ = ~new_new_n30118__ & new_new_n30985__;
  assign new_new_n30988__ = ~new_new_n30986__ & ~new_new_n30987__;
  assign new_new_n30989__ = ~new_new_n30984__ & new_new_n30988__;
  assign new_new_n30990__ = ~new_new_n30983__ & ~new_new_n30989__;
  assign new_new_n30991__ = ~new_new_n30121__ & ~new_new_n30136__;
  assign new_new_n30992__ = new_new_n30134__ & ~new_new_n30991__;
  assign new_new_n30993__ = ~new_new_n30134__ & new_new_n30991__;
  assign new_new_n30994__ = ~new_new_n30992__ & ~new_new_n30993__;
  assign new_new_n30995__ = new_new_n30990__ & new_new_n30994__;
  assign new_new_n30996__ = ~new_new_n30990__ & ~new_new_n30994__;
  assign new_new_n30997__ = new_new_n11471__ & new_new_n27111__;
  assign new_new_n30998__ = new_new_n11475__ & ~new_new_n27021__;
  assign new_new_n30999__ = ~new_new_n11478__ & new_new_n27029__;
  assign new_new_n31000__ = new_new_n11478__ & ~new_new_n27764__;
  assign new_new_n31001__ = ~new_new_n11482__ & ~new_new_n30999__;
  assign new_new_n31002__ = ~new_new_n31000__ & new_new_n31001__;
  assign new_new_n31003__ = ~new_new_n30997__ & ~new_new_n30998__;
  assign new_new_n31004__ = ~new_new_n31002__ & new_new_n31003__;
  assign new_new_n31005__ = pi05 & ~new_new_n31004__;
  assign new_new_n31006__ = ~pi05 & new_new_n31004__;
  assign new_new_n31007__ = ~new_new_n31005__ & ~new_new_n31006__;
  assign new_new_n31008__ = ~new_new_n30996__ & new_new_n31007__;
  assign new_new_n31009__ = ~new_new_n30995__ & ~new_new_n31008__;
  assign new_new_n31010__ = ~new_new_n30842__ & ~new_new_n31009__;
  assign new_new_n31011__ = new_new_n30842__ & new_new_n31009__;
  assign new_new_n31012__ = new_new_n12850__ & ~new_new_n27003__;
  assign new_new_n31013__ = new_new_n11475__ & ~new_new_n27029__;
  assign new_new_n31014__ = new_new_n11471__ & ~new_new_n27021__;
  assign new_new_n31015__ = new_new_n13069__ & new_new_n27962__;
  assign new_new_n31016__ = ~new_new_n31013__ & ~new_new_n31014__;
  assign new_new_n31017__ = ~new_new_n31012__ & new_new_n31016__;
  assign new_new_n31018__ = ~new_new_n31015__ & new_new_n31017__;
  assign new_new_n31019__ = pi05 & ~new_new_n31018__;
  assign new_new_n31020__ = ~pi05 & new_new_n31018__;
  assign new_new_n31021__ = ~new_new_n31019__ & ~new_new_n31020__;
  assign new_new_n31022__ = ~new_new_n31011__ & new_new_n31021__;
  assign new_new_n31023__ = ~new_new_n31010__ & ~new_new_n31022__;
  assign new_new_n31024__ = new_new_n30831__ & ~new_new_n31023__;
  assign new_new_n31025__ = ~new_new_n30831__ & new_new_n31023__;
  assign new_new_n31026__ = new_new_n10694__ & new_new_n27796__;
  assign new_new_n31027__ = pi07 & ~new_new_n30004__;
  assign new_new_n31028__ = ~pi07 & new_new_n30004__;
  assign new_new_n31029__ = ~new_new_n31027__ & ~new_new_n31028__;
  assign new_new_n31030__ = new_new_n31026__ & ~new_new_n31029__;
  assign new_new_n31031__ = pi08 & new_new_n30004__;
  assign new_new_n31032__ = ~pi08 & ~new_new_n30004__;
  assign new_new_n31033__ = ~new_new_n31031__ & ~new_new_n31032__;
  assign new_new_n31034__ = ~new_new_n31026__ & new_new_n31033__;
  assign new_new_n31035__ = ~new_new_n31030__ & ~new_new_n31034__;
  assign new_new_n31036__ = new_new_n30150__ & ~new_new_n31035__;
  assign new_new_n31037__ = ~new_new_n30150__ & ~new_new_n31033__;
  assign new_new_n31038__ = ~new_new_n31036__ & ~new_new_n31037__;
  assign new_new_n31039__ = new_new_n30143__ & ~new_new_n31038__;
  assign new_new_n31040__ = ~new_new_n30143__ & new_new_n31038__;
  assign new_new_n31041__ = ~new_new_n31039__ & ~new_new_n31040__;
  assign new_new_n31042__ = ~new_new_n31025__ & ~new_new_n31041__;
  assign new_new_n31043__ = ~new_new_n31024__ & ~new_new_n31042__;
  assign new_new_n31044__ = ~new_new_n30816__ & new_new_n31043__;
  assign new_new_n31045__ = ~new_new_n30815__ & ~new_new_n31044__;
  assign new_new_n31046__ = new_new_n30798__ & ~new_new_n31045__;
  assign new_new_n31047__ = ~new_new_n30798__ & new_new_n31045__;
  assign new_new_n31048__ = new_new_n11475__ & new_new_n26971__;
  assign new_new_n31049__ = new_new_n11471__ & ~new_new_n26978__;
  assign new_new_n31050__ = new_new_n12850__ & ~new_new_n26937__;
  assign new_new_n31051__ = ~new_new_n31048__ & ~new_new_n31049__;
  assign new_new_n31052__ = ~new_new_n31050__ & new_new_n31051__;
  assign new_new_n31053__ = ~pi05 & ~new_new_n31052__;
  assign new_new_n31054__ = new_new_n12873__ & new_new_n28005__;
  assign new_new_n31055__ = new_new_n11469__ & new_new_n28005__;
  assign new_new_n31056__ = pi05 & ~new_new_n31055__;
  assign new_new_n31057__ = ~new_new_n31054__ & ~new_new_n31056__;
  assign new_new_n31058__ = new_new_n31052__ & ~new_new_n31057__;
  assign new_new_n31059__ = ~new_new_n31053__ & ~new_new_n31058__;
  assign new_new_n31060__ = ~new_new_n31047__ & new_new_n31059__;
  assign new_new_n31061__ = ~new_new_n31046__ & ~new_new_n31060__;
  assign new_new_n31062__ = ~new_new_n30794__ & ~new_new_n31061__;
  assign new_new_n31063__ = ~new_new_n30793__ & ~new_new_n31062__;
  assign new_new_n31064__ = new_new_n29700__ & ~new_new_n30199__;
  assign new_new_n31065__ = ~new_new_n29700__ & new_new_n30199__;
  assign new_new_n31066__ = ~new_new_n31064__ & ~new_new_n31065__;
  assign new_new_n31067__ = new_new_n29691__ & new_new_n31066__;
  assign new_new_n31068__ = ~new_new_n29691__ & ~new_new_n31066__;
  assign new_new_n31069__ = ~new_new_n31067__ & ~new_new_n31068__;
  assign new_new_n31070__ = new_new_n29986__ & ~new_new_n31069__;
  assign new_new_n31071__ = ~new_new_n29986__ & new_new_n31069__;
  assign new_new_n31072__ = ~new_new_n31070__ & ~new_new_n31071__;
  assign new_new_n31073__ = new_new_n30204__ & new_new_n31072__;
  assign new_new_n31074__ = ~new_new_n30204__ & ~new_new_n31072__;
  assign new_new_n31075__ = ~new_new_n31073__ & ~new_new_n31074__;
  assign new_new_n31076__ = new_new_n31063__ & ~new_new_n31075__;
  assign new_new_n31077__ = ~new_new_n31063__ & new_new_n31075__;
  assign new_new_n31078__ = new_new_n12850__ & ~new_new_n26941__;
  assign new_new_n31079__ = new_new_n13111__ & ~new_new_n26937__;
  assign new_new_n31080__ = new_new_n11469__ & ~new_new_n27502__;
  assign new_new_n31081__ = ~new_new_n31079__ & ~new_new_n31080__;
  assign new_new_n31082__ = new_new_n11478__ & ~new_new_n31081__;
  assign new_new_n31083__ = new_new_n11475__ & new_new_n27152__;
  assign new_new_n31084__ = ~new_new_n31078__ & ~new_new_n31083__;
  assign new_new_n31085__ = ~new_new_n31082__ & new_new_n31084__;
  assign new_new_n31086__ = pi05 & ~new_new_n31085__;
  assign new_new_n31087__ = ~pi05 & new_new_n31085__;
  assign new_new_n31088__ = ~new_new_n31086__ & ~new_new_n31087__;
  assign new_new_n31089__ = ~new_new_n31077__ & new_new_n31088__;
  assign new_new_n31090__ = ~new_new_n31076__ & ~new_new_n31089__;
  assign new_new_n31091__ = new_new_n30763__ & ~new_new_n31090__;
  assign new_new_n31092__ = ~new_new_n30763__ & new_new_n31090__;
  assign new_new_n31093__ = ~new_new_n30213__ & ~new_new_n30214__;
  assign new_new_n31094__ = ~new_new_n30226__ & new_new_n31093__;
  assign new_new_n31095__ = new_new_n30226__ & ~new_new_n31093__;
  assign new_new_n31096__ = ~new_new_n31094__ & ~new_new_n31095__;
  assign new_new_n31097__ = ~new_new_n31092__ & new_new_n31096__;
  assign new_new_n31098__ = ~new_new_n31091__ & ~new_new_n31097__;
  assign new_new_n31099__ = ~new_new_n30751__ & ~new_new_n31098__;
  assign new_new_n31100__ = ~new_new_n30750__ & ~new_new_n31099__;
  assign new_new_n31101__ = ~new_new_n30731__ & new_new_n31100__;
  assign new_new_n31102__ = new_new_n30731__ & ~new_new_n31100__;
  assign new_new_n31103__ = new_new_n30231__ & ~new_new_n30243__;
  assign new_new_n31104__ = ~new_new_n30231__ & new_new_n30243__;
  assign new_new_n31105__ = ~new_new_n31103__ & ~new_new_n31104__;
  assign new_new_n31106__ = new_new_n30230__ & new_new_n31105__;
  assign new_new_n31107__ = ~new_new_n30230__ & ~new_new_n31105__;
  assign new_new_n31108__ = ~new_new_n31106__ & ~new_new_n31107__;
  assign new_new_n31109__ = ~new_new_n31102__ & ~new_new_n31108__;
  assign new_new_n31110__ = ~new_new_n31101__ & ~new_new_n31109__;
  assign new_new_n31111__ = ~new_new_n30719__ & ~new_new_n31110__;
  assign new_new_n31112__ = new_new_n30719__ & new_new_n31110__;
  assign new_new_n31113__ = new_new_n12850__ & new_new_n26922__;
  assign new_new_n31114__ = new_new_n11475__ & ~new_new_n27168__;
  assign new_new_n31115__ = new_new_n11471__ & new_new_n26917__;
  assign new_new_n31116__ = new_new_n13069__ & ~new_new_n29366__;
  assign new_new_n31117__ = ~new_new_n31114__ & ~new_new_n31115__;
  assign new_new_n31118__ = ~new_new_n31113__ & new_new_n31117__;
  assign new_new_n31119__ = ~new_new_n31116__ & new_new_n31118__;
  assign new_new_n31120__ = ~pi05 & ~new_new_n31119__;
  assign new_new_n31121__ = pi05 & new_new_n31119__;
  assign new_new_n31122__ = ~new_new_n31120__ & ~new_new_n31121__;
  assign new_new_n31123__ = ~new_new_n31112__ & new_new_n31122__;
  assign new_new_n31124__ = ~new_new_n31111__ & ~new_new_n31123__;
  assign new_new_n31125__ = ~new_new_n30270__ & ~new_new_n30271__;
  assign new_new_n31126__ = ~new_new_n30281__ & new_new_n31125__;
  assign new_new_n31127__ = new_new_n30281__ & ~new_new_n31125__;
  assign new_new_n31128__ = ~new_new_n31126__ & ~new_new_n31127__;
  assign new_new_n31129__ = ~new_new_n31124__ & new_new_n31128__;
  assign new_new_n31130__ = new_new_n31124__ & ~new_new_n31128__;
  assign new_new_n31131__ = new_new_n11471__ & ~new_new_n27168__;
  assign new_new_n31132__ = new_new_n11475__ & new_new_n26922__;
  assign new_new_n31133__ = ~new_new_n11478__ & new_new_n26888__;
  assign new_new_n31134__ = new_new_n11478__ & ~new_new_n27180__;
  assign new_new_n31135__ = ~new_new_n11482__ & ~new_new_n31133__;
  assign new_new_n31136__ = ~new_new_n31134__ & new_new_n31135__;
  assign new_new_n31137__ = ~new_new_n31131__ & ~new_new_n31132__;
  assign new_new_n31138__ = ~new_new_n31136__ & new_new_n31137__;
  assign new_new_n31139__ = pi05 & ~new_new_n31138__;
  assign new_new_n31140__ = ~pi05 & new_new_n31138__;
  assign new_new_n31141__ = ~new_new_n31139__ & ~new_new_n31140__;
  assign new_new_n31142__ = ~new_new_n31130__ & ~new_new_n31141__;
  assign new_new_n31143__ = ~new_new_n31129__ & ~new_new_n31142__;
  assign new_new_n31144__ = ~new_new_n30715__ & ~new_new_n31143__;
  assign new_new_n31145__ = new_new_n30715__ & new_new_n31143__;
  assign new_new_n31146__ = new_new_n12850__ & ~new_new_n26854__;
  assign new_new_n31147__ = new_new_n13111__ & new_new_n26922__;
  assign new_new_n31148__ = new_new_n11469__ & ~new_new_n27430__;
  assign new_new_n31149__ = ~new_new_n31147__ & ~new_new_n31148__;
  assign new_new_n31150__ = new_new_n11478__ & ~new_new_n31149__;
  assign new_new_n31151__ = new_new_n11475__ & ~new_new_n26888__;
  assign new_new_n31152__ = ~new_new_n31146__ & ~new_new_n31151__;
  assign new_new_n31153__ = ~new_new_n31150__ & new_new_n31152__;
  assign new_new_n31154__ = ~pi05 & ~new_new_n31153__;
  assign new_new_n31155__ = pi05 & new_new_n31153__;
  assign new_new_n31156__ = ~new_new_n31154__ & ~new_new_n31155__;
  assign new_new_n31157__ = ~new_new_n31145__ & new_new_n31156__;
  assign new_new_n31158__ = ~new_new_n31144__ & ~new_new_n31157__;
  assign new_new_n31159__ = new_new_n29932__ & ~new_new_n30291__;
  assign new_new_n31160__ = ~new_new_n29932__ & new_new_n30291__;
  assign new_new_n31161__ = ~new_new_n31159__ & ~new_new_n31160__;
  assign new_new_n31162__ = new_new_n30299__ & new_new_n31161__;
  assign new_new_n31163__ = ~new_new_n30299__ & ~new_new_n31161__;
  assign new_new_n31164__ = ~new_new_n31162__ & ~new_new_n31163__;
  assign new_new_n31165__ = new_new_n31158__ & new_new_n31164__;
  assign new_new_n31166__ = ~new_new_n31158__ & ~new_new_n31164__;
  assign new_new_n31167__ = new_new_n11471__ & ~new_new_n26888__;
  assign new_new_n31168__ = new_new_n11475__ & ~new_new_n26854__;
  assign new_new_n31169__ = ~new_new_n11478__ & ~new_new_n26847__;
  assign new_new_n31170__ = new_new_n11478__ & ~new_new_n29424__;
  assign new_new_n31171__ = ~new_new_n11482__ & ~new_new_n31169__;
  assign new_new_n31172__ = ~new_new_n31170__ & new_new_n31171__;
  assign new_new_n31173__ = ~new_new_n31167__ & ~new_new_n31168__;
  assign new_new_n31174__ = ~new_new_n31172__ & new_new_n31173__;
  assign new_new_n31175__ = ~pi05 & ~new_new_n31174__;
  assign new_new_n31176__ = pi05 & new_new_n31174__;
  assign new_new_n31177__ = ~new_new_n31175__ & ~new_new_n31176__;
  assign new_new_n31178__ = ~new_new_n31166__ & ~new_new_n31177__;
  assign new_new_n31179__ = ~new_new_n31165__ & ~new_new_n31178__;
  assign new_new_n31180__ = new_new_n30711__ & ~new_new_n31179__;
  assign new_new_n31181__ = ~new_new_n30711__ & new_new_n31179__;
  assign new_new_n31182__ = new_new_n12850__ & ~new_new_n26823__;
  assign new_new_n31183__ = new_new_n13111__ & ~new_new_n26854__;
  assign new_new_n31184__ = new_new_n11469__ & ~new_new_n29400__;
  assign new_new_n31185__ = ~new_new_n31183__ & ~new_new_n31184__;
  assign new_new_n31186__ = new_new_n11478__ & ~new_new_n31185__;
  assign new_new_n31187__ = new_new_n11475__ & new_new_n26847__;
  assign new_new_n31188__ = ~new_new_n31182__ & ~new_new_n31187__;
  assign new_new_n31189__ = ~new_new_n31186__ & new_new_n31188__;
  assign new_new_n31190__ = pi05 & ~new_new_n31189__;
  assign new_new_n31191__ = ~pi05 & new_new_n31189__;
  assign new_new_n31192__ = ~new_new_n31190__ & ~new_new_n31191__;
  assign new_new_n31193__ = ~new_new_n31181__ & new_new_n31192__;
  assign new_new_n31194__ = ~new_new_n31180__ & ~new_new_n31193__;
  assign new_new_n31195__ = new_new_n30707__ & ~new_new_n31194__;
  assign new_new_n31196__ = ~new_new_n30707__ & new_new_n31194__;
  assign new_new_n31197__ = new_new_n12850__ & ~new_new_n27221__;
  assign new_new_n31198__ = new_new_n11475__ & ~new_new_n26823__;
  assign new_new_n31199__ = new_new_n11471__ & new_new_n26847__;
  assign new_new_n31200__ = new_new_n13069__ & new_new_n27411__;
  assign new_new_n31201__ = ~new_new_n31198__ & ~new_new_n31199__;
  assign new_new_n31202__ = ~new_new_n31197__ & new_new_n31201__;
  assign new_new_n31203__ = ~new_new_n31200__ & new_new_n31202__;
  assign new_new_n31204__ = pi05 & ~new_new_n31203__;
  assign new_new_n31205__ = ~pi05 & new_new_n31203__;
  assign new_new_n31206__ = ~new_new_n31204__ & ~new_new_n31205__;
  assign new_new_n31207__ = ~new_new_n31196__ & new_new_n31206__;
  assign new_new_n31208__ = ~new_new_n31195__ & ~new_new_n31207__;
  assign new_new_n31209__ = pi08 & ~new_new_n29904__;
  assign new_new_n31210__ = ~new_new_n30332__ & ~new_new_n31209__;
  assign new_new_n31211__ = new_new_n29900__ & new_new_n31210__;
  assign new_new_n31212__ = ~new_new_n29900__ & ~new_new_n31210__;
  assign new_new_n31213__ = ~new_new_n31211__ & ~new_new_n31212__;
  assign new_new_n31214__ = new_new_n30701__ & ~new_new_n31213__;
  assign new_new_n31215__ = new_new_n30700__ & new_new_n31213__;
  assign new_new_n31216__ = ~new_new_n29912__ & ~new_new_n29916__;
  assign new_new_n31217__ = new_new_n29900__ & new_new_n31216__;
  assign new_new_n31218__ = ~new_new_n29900__ & ~new_new_n31216__;
  assign new_new_n31219__ = new_new_n30702__ & ~new_new_n31217__;
  assign new_new_n31220__ = ~new_new_n31218__ & new_new_n31219__;
  assign new_new_n31221__ = ~new_new_n31214__ & ~new_new_n31215__;
  assign new_new_n31222__ = ~new_new_n31220__ & new_new_n31221__;
  assign new_new_n31223__ = ~new_new_n31208__ & new_new_n31222__;
  assign new_new_n31224__ = new_new_n31208__ & ~new_new_n31222__;
  assign new_new_n31225__ = new_new_n11475__ & ~new_new_n27221__;
  assign new_new_n31226__ = new_new_n11471__ & ~new_new_n26823__;
  assign new_new_n31227__ = new_new_n12850__ & ~new_new_n26741__;
  assign new_new_n31228__ = ~new_new_n31225__ & ~new_new_n31226__;
  assign new_new_n31229__ = ~new_new_n31227__ & new_new_n31228__;
  assign new_new_n31230__ = pi05 & ~new_new_n31229__;
  assign new_new_n31231__ = new_new_n12856__ & new_new_n30393__;
  assign new_new_n31232__ = new_new_n11469__ & new_new_n30393__;
  assign new_new_n31233__ = ~pi05 & ~new_new_n31232__;
  assign new_new_n31234__ = ~new_new_n31231__ & ~new_new_n31233__;
  assign new_new_n31235__ = new_new_n31229__ & ~new_new_n31234__;
  assign new_new_n31236__ = ~new_new_n31230__ & ~new_new_n31235__;
  assign new_new_n31237__ = ~new_new_n31224__ & new_new_n31236__;
  assign new_new_n31238__ = ~new_new_n31223__ & ~new_new_n31237__;
  assign new_new_n31239__ = new_new_n30699__ & ~new_new_n31238__;
  assign new_new_n31240__ = ~new_new_n30699__ & new_new_n31238__;
  assign new_new_n31241__ = ~new_new_n30338__ & ~new_new_n30339__;
  assign new_new_n31242__ = new_new_n30343__ & ~new_new_n31241__;
  assign new_new_n31243__ = ~new_new_n30343__ & new_new_n31241__;
  assign new_new_n31244__ = ~new_new_n31242__ & ~new_new_n31243__;
  assign new_new_n31245__ = ~new_new_n31240__ & ~new_new_n31244__;
  assign new_new_n31246__ = ~new_new_n31239__ & ~new_new_n31245__;
  assign new_new_n31247__ = ~new_new_n30682__ & ~new_new_n31246__;
  assign new_new_n31248__ = new_new_n30682__ & new_new_n31246__;
  assign new_new_n31249__ = ~new_new_n30354__ & new_new_n30367__;
  assign new_new_n31250__ = ~new_new_n30368__ & ~new_new_n31249__;
  assign new_new_n31251__ = ~new_new_n31248__ & new_new_n31250__;
  assign new_new_n31252__ = ~new_new_n31247__ & ~new_new_n31251__;
  assign new_new_n31253__ = ~new_new_n30669__ & ~new_new_n31252__;
  assign new_new_n31254__ = ~new_new_n30668__ & ~new_new_n31253__;
  assign new_new_n31255__ = ~new_new_n30650__ & new_new_n31254__;
  assign new_new_n31256__ = new_new_n30650__ & ~new_new_n31254__;
  assign new_new_n31257__ = ~new_new_n30403__ & ~new_new_n30404__;
  assign new_new_n31258__ = new_new_n30418__ & ~new_new_n31257__;
  assign new_new_n31259__ = ~new_new_n30418__ & new_new_n31257__;
  assign new_new_n31260__ = ~new_new_n31258__ & ~new_new_n31259__;
  assign new_new_n31261__ = ~new_new_n31256__ & ~new_new_n31260__;
  assign new_new_n31262__ = ~new_new_n31255__ & ~new_new_n31261__;
  assign new_new_n31263__ = ~new_new_n29862__ & ~new_new_n29863__;
  assign new_new_n31264__ = new_new_n30420__ & new_new_n31263__;
  assign new_new_n31265__ = ~new_new_n30420__ & ~new_new_n31263__;
  assign new_new_n31266__ = ~new_new_n31264__ & ~new_new_n31265__;
  assign new_new_n31267__ = ~new_new_n31262__ & new_new_n31266__;
  assign new_new_n31268__ = new_new_n31262__ & ~new_new_n31266__;
  assign new_new_n31269__ = new_new_n11475__ & new_new_n26729__;
  assign new_new_n31270__ = ~new_new_n11478__ & ~new_new_n26722__;
  assign new_new_n31271__ = new_new_n11478__ & new_new_n27348__;
  assign new_new_n31272__ = ~new_new_n11482__ & ~new_new_n31270__;
  assign new_new_n31273__ = ~new_new_n31271__ & new_new_n31272__;
  assign new_new_n31274__ = ~new_new_n31269__ & ~new_new_n31273__;
  assign new_new_n31275__ = new_new_n11466__ & new_new_n26774__;
  assign new_new_n31276__ = pi05 & ~new_new_n31275__;
  assign new_new_n31277__ = new_new_n11467__ & new_new_n26774__;
  assign new_new_n31278__ = ~pi05 & ~new_new_n31277__;
  assign new_new_n31279__ = pi02 & ~new_new_n31278__;
  assign new_new_n31280__ = ~new_new_n31276__ & ~new_new_n31279__;
  assign new_new_n31281__ = new_new_n31274__ & ~new_new_n31280__;
  assign new_new_n31282__ = ~pi05 & ~new_new_n31274__;
  assign new_new_n31283__ = ~new_new_n31281__ & ~new_new_n31282__;
  assign new_new_n31284__ = ~new_new_n31268__ & new_new_n31283__;
  assign new_new_n31285__ = ~new_new_n31267__ & ~new_new_n31284__;
  assign new_new_n31286__ = ~new_new_n30616__ & ~new_new_n31285__;
  assign new_new_n31287__ = ~new_new_n30615__ & ~new_new_n31286__;
  assign new_new_n31288__ = new_new_n27317__ & ~new_new_n31287__;
  assign new_new_n31289__ = ~new_new_n27317__ & new_new_n31287__;
  assign new_new_n31290__ = ~new_new_n31288__ & ~new_new_n31289__;
  assign new_new_n31291__ = new_new_n10702__ & new_new_n26774__;
  assign new_new_n31292__ = ~new_new_n11409__ & new_new_n26810__;
  assign new_new_n31293__ = new_new_n10698__ & new_new_n26729__;
  assign new_new_n31294__ = ~new_new_n31291__ & ~new_new_n31292__;
  assign new_new_n31295__ = ~new_new_n31293__ & new_new_n31294__;
  assign new_new_n31296__ = new_new_n10694__ & new_new_n30644__;
  assign new_new_n31297__ = new_new_n8474__ & ~new_new_n26741__;
  assign new_new_n31298__ = ~new_new_n8479__ & ~new_new_n27221__;
  assign new_new_n31299__ = ~new_new_n31297__ & ~new_new_n31298__;
  assign new_new_n31300__ = new_new_n8469__ & ~new_new_n26802__;
  assign new_new_n31301__ = new_new_n30411__ & new_new_n31300__;
  assign new_new_n31302__ = new_new_n31299__ & ~new_new_n31301__;
  assign new_new_n31303__ = pi11 & ~new_new_n31302__;
  assign new_new_n31304__ = new_new_n8469__ & ~new_new_n27391__;
  assign new_new_n31305__ = ~pi11 & ~new_new_n31304__;
  assign new_new_n31306__ = ~pi10 & ~new_new_n30692__;
  assign new_new_n31307__ = pi10 & ~new_new_n30410__;
  assign new_new_n31308__ = new_new_n8469__ & ~new_new_n31306__;
  assign new_new_n31309__ = ~new_new_n31307__ & new_new_n31308__;
  assign new_new_n31310__ = ~new_new_n31305__ & ~new_new_n31309__;
  assign new_new_n31311__ = new_new_n31299__ & ~new_new_n31310__;
  assign new_new_n31312__ = ~new_new_n31303__ & ~new_new_n31311__;
  assign new_new_n31313__ = new_new_n30439__ & ~new_new_n30598__;
  assign new_new_n31314__ = ~new_new_n30599__ & ~new_new_n31313__;
  assign new_new_n31315__ = ~new_new_n31312__ & new_new_n31314__;
  assign new_new_n31316__ = new_new_n31312__ & ~new_new_n31314__;
  assign new_new_n31317__ = ~new_new_n31315__ & ~new_new_n31316__;
  assign new_new_n31318__ = new_new_n5213__ & new_new_n27152__;
  assign new_new_n31319__ = new_new_n5183__ & ~new_new_n26937__;
  assign new_new_n31320__ = new_new_n5191__ & new_new_n26971__;
  assign new_new_n31321__ = new_new_n5215__ & ~new_new_n28666__;
  assign new_new_n31322__ = ~new_new_n31319__ & ~new_new_n31320__;
  assign new_new_n31323__ = ~new_new_n31318__ & new_new_n31322__;
  assign new_new_n31324__ = ~new_new_n31321__ & new_new_n31323__;
  assign new_new_n31325__ = ~new_new_n4900__ & new_new_n27986__;
  assign new_new_n31326__ = new_new_n873__ & ~new_new_n27003__;
  assign new_new_n31327__ = ~new_new_n333__ & ~new_new_n27029__;
  assign new_new_n31328__ = new_new_n3311__ & ~new_new_n26978__;
  assign new_new_n31329__ = ~new_new_n31326__ & ~new_new_n31327__;
  assign new_new_n31330__ = ~new_new_n31328__ & new_new_n31329__;
  assign new_new_n31331__ = ~new_new_n31325__ & new_new_n31330__;
  assign new_new_n31332__ = ~pi26 & ~new_new_n31331__;
  assign new_new_n31333__ = pi26 & new_new_n31331__;
  assign new_new_n31334__ = ~new_new_n31332__ & ~new_new_n31333__;
  assign new_new_n31335__ = ~new_new_n30550__ & new_new_n30553__;
  assign new_new_n31336__ = ~new_new_n30549__ & ~new_new_n31335__;
  assign new_new_n31337__ = ~new_new_n31334__ & new_new_n31336__;
  assign new_new_n31338__ = new_new_n31334__ & ~new_new_n31336__;
  assign new_new_n31339__ = ~new_new_n31337__ & ~new_new_n31338__;
  assign new_new_n31340__ = ~new_new_n30541__ & ~new_new_n30546__;
  assign new_new_n31341__ = new_new_n31339__ & ~new_new_n31340__;
  assign new_new_n31342__ = ~new_new_n31339__ & new_new_n31340__;
  assign new_new_n31343__ = ~new_new_n31341__ & ~new_new_n31342__;
  assign new_new_n31344__ = new_new_n161__ & new_new_n27041__;
  assign new_new_n31345__ = new_new_n765__ & ~new_new_n27054__;
  assign new_new_n31346__ = ~new_new_n31344__ & ~new_new_n31345__;
  assign new_new_n31347__ = ~pi31 & ~new_new_n31346__;
  assign new_new_n31348__ = new_new_n71__ & new_new_n27041__;
  assign new_new_n31349__ = new_new_n765__ & ~new_new_n27094__;
  assign new_new_n31350__ = ~new_new_n30511__ & ~new_new_n31348__;
  assign new_new_n31351__ = ~new_new_n31349__ & new_new_n31350__;
  assign new_new_n31352__ = pi31 & ~new_new_n31351__;
  assign new_new_n31353__ = ~new_new_n31347__ & ~new_new_n31352__;
  assign new_new_n31354__ = new_new_n135__ & ~new_new_n752__;
  assign new_new_n31355__ = ~new_new_n749__ & ~new_new_n877__;
  assign new_new_n31356__ = ~new_new_n306__ & new_new_n31355__;
  assign new_new_n31357__ = new_new_n2516__ & new_new_n6758__;
  assign new_new_n31358__ = new_new_n18568__ & ~new_new_n31354__;
  assign new_new_n31359__ = new_new_n31357__ & new_new_n31358__;
  assign new_new_n31360__ = new_new_n830__ & new_new_n31356__;
  assign new_new_n31361__ = new_new_n1705__ & new_new_n31360__;
  assign new_new_n31362__ = new_new_n2028__ & new_new_n31359__;
  assign new_new_n31363__ = new_new_n2543__ & new_new_n31362__;
  assign new_new_n31364__ = new_new_n5565__ & new_new_n31361__;
  assign new_new_n31365__ = new_new_n16816__ & new_new_n31364__;
  assign new_new_n31366__ = new_new_n4373__ & new_new_n31363__;
  assign new_new_n31367__ = new_new_n31365__ & new_new_n31366__;
  assign new_new_n31368__ = new_new_n5429__ & new_new_n31367__;
  assign new_new_n31369__ = new_new_n16792__ & new_new_n31368__;
  assign new_new_n31370__ = new_new_n31353__ & new_new_n31369__;
  assign new_new_n31371__ = ~new_new_n31353__ & ~new_new_n31369__;
  assign new_new_n31372__ = ~new_new_n31370__ & ~new_new_n31371__;
  assign new_new_n31373__ = new_new_n4815__ & ~new_new_n27021__;
  assign new_new_n31374__ = ~new_new_n4818__ & ~new_new_n27033__;
  assign new_new_n31375__ = new_new_n4212__ & new_new_n27111__;
  assign new_new_n31376__ = ~new_new_n31374__ & ~new_new_n31375__;
  assign new_new_n31377__ = ~new_new_n31373__ & new_new_n31376__;
  assign new_new_n31378__ = new_new_n4214__ & new_new_n27796__;
  assign new_new_n31379__ = ~pi29 & ~new_new_n31378__;
  assign new_new_n31380__ = new_new_n5732__ & new_new_n27796__;
  assign new_new_n31381__ = ~new_new_n31379__ & ~new_new_n31380__;
  assign new_new_n31382__ = new_new_n31377__ & ~new_new_n31381__;
  assign new_new_n31383__ = pi29 & ~new_new_n31377__;
  assign new_new_n31384__ = ~new_new_n31382__ & ~new_new_n31383__;
  assign new_new_n31385__ = new_new_n31372__ & ~new_new_n31384__;
  assign new_new_n31386__ = ~new_new_n31372__ & new_new_n31384__;
  assign new_new_n31387__ = ~new_new_n31385__ & ~new_new_n31386__;
  assign new_new_n31388__ = new_new_n31343__ & new_new_n31387__;
  assign new_new_n31389__ = ~new_new_n31343__ & ~new_new_n31387__;
  assign new_new_n31390__ = ~new_new_n31388__ & ~new_new_n31389__;
  assign new_new_n31391__ = new_new_n30492__ & ~new_new_n31390__;
  assign new_new_n31392__ = new_new_n30493__ & new_new_n31390__;
  assign new_new_n31393__ = ~new_new_n31391__ & ~new_new_n31392__;
  assign new_new_n31394__ = ~new_new_n30556__ & ~new_new_n31393__;
  assign new_new_n31395__ = new_new_n30559__ & ~new_new_n31390__;
  assign new_new_n31396__ = ~new_new_n31394__ & ~new_new_n31395__;
  assign new_new_n31397__ = ~new_new_n30576__ & ~new_new_n31396__;
  assign new_new_n31398__ = ~new_new_n30492__ & ~new_new_n30558__;
  assign new_new_n31399__ = new_new_n31390__ & new_new_n31398__;
  assign new_new_n31400__ = ~new_new_n31391__ & ~new_new_n31399__;
  assign new_new_n31401__ = new_new_n30575__ & ~new_new_n31400__;
  assign new_new_n31402__ = ~new_new_n31397__ & ~new_new_n31401__;
  assign new_new_n31403__ = ~new_new_n30492__ & new_new_n31390__;
  assign new_new_n31404__ = ~new_new_n31391__ & ~new_new_n31403__;
  assign new_new_n31405__ = new_new_n30560__ & new_new_n31404__;
  assign new_new_n31406__ = ~new_new_n30575__ & new_new_n31405__;
  assign new_new_n31407__ = ~new_new_n30493__ & ~new_new_n31390__;
  assign new_new_n31408__ = ~new_new_n31399__ & ~new_new_n31407__;
  assign new_new_n31409__ = new_new_n30576__ & new_new_n31408__;
  assign new_new_n31410__ = ~new_new_n31406__ & ~new_new_n31409__;
  assign new_new_n31411__ = new_new_n31402__ & new_new_n31410__;
  assign new_new_n31412__ = pi23 & ~new_new_n31411__;
  assign new_new_n31413__ = ~pi23 & new_new_n31411__;
  assign new_new_n31414__ = ~new_new_n31412__ & ~new_new_n31413__;
  assign new_new_n31415__ = new_new_n31324__ & new_new_n31414__;
  assign new_new_n31416__ = ~new_new_n31324__ & ~new_new_n31414__;
  assign new_new_n31417__ = ~new_new_n31415__ & ~new_new_n31416__;
  assign new_new_n31418__ = ~new_new_n30581__ & ~new_new_n30585__;
  assign new_new_n31419__ = ~new_new_n30582__ & ~new_new_n31418__;
  assign new_new_n31420__ = new_new_n31417__ & new_new_n31419__;
  assign new_new_n31421__ = ~new_new_n31417__ & ~new_new_n31419__;
  assign new_new_n31422__ = ~new_new_n31420__ & ~new_new_n31421__;
  assign new_new_n31423__ = new_new_n6629__ & new_new_n26928__;
  assign new_new_n31424__ = ~new_new_n6625__ & ~new_new_n26941__;
  assign new_new_n31425__ = new_new_n6634__ & new_new_n26917__;
  assign new_new_n31426__ = ~new_new_n31423__ & ~new_new_n31424__;
  assign new_new_n31427__ = ~new_new_n31425__ & new_new_n31426__;
  assign new_new_n31428__ = new_new_n6631__ & ~new_new_n27462__;
  assign new_new_n31429__ = pi20 & ~new_new_n31428__;
  assign new_new_n31430__ = new_new_n6640__ & ~new_new_n27462__;
  assign new_new_n31431__ = ~new_new_n31429__ & ~new_new_n31430__;
  assign new_new_n31432__ = new_new_n31427__ & ~new_new_n31431__;
  assign new_new_n31433__ = ~pi20 & ~new_new_n31427__;
  assign new_new_n31434__ = ~new_new_n31432__ & ~new_new_n31433__;
  assign new_new_n31435__ = new_new_n31422__ & ~new_new_n31434__;
  assign new_new_n31436__ = ~new_new_n31422__ & new_new_n31434__;
  assign new_new_n31437__ = ~new_new_n31435__ & ~new_new_n31436__;
  assign new_new_n31438__ = new_new_n7935__ & ~new_new_n26888__;
  assign new_new_n31439__ = new_new_n6964__ & ~new_new_n27168__;
  assign new_new_n31440__ = new_new_n6968__ & new_new_n26922__;
  assign new_new_n31441__ = ~new_new_n31439__ & ~new_new_n31440__;
  assign new_new_n31442__ = ~new_new_n31438__ & new_new_n31441__;
  assign new_new_n31443__ = new_new_n6958__ & new_new_n27180__;
  assign new_new_n31444__ = pi17 & ~new_new_n31443__;
  assign new_new_n31445__ = new_new_n7942__ & new_new_n27180__;
  assign new_new_n31446__ = ~new_new_n31444__ & ~new_new_n31445__;
  assign new_new_n31447__ = new_new_n31442__ & ~new_new_n31446__;
  assign new_new_n31448__ = ~pi17 & ~new_new_n31442__;
  assign new_new_n31449__ = ~new_new_n31447__ & ~new_new_n31448__;
  assign new_new_n31450__ = new_new_n30588__ & new_new_n30597__;
  assign new_new_n31451__ = ~new_new_n30588__ & ~new_new_n30597__;
  assign new_new_n31452__ = ~new_new_n30465__ & ~new_new_n31451__;
  assign new_new_n31453__ = ~new_new_n31450__ & ~new_new_n31452__;
  assign new_new_n31454__ = new_new_n31449__ & ~new_new_n31453__;
  assign new_new_n31455__ = ~new_new_n31449__ & new_new_n31453__;
  assign new_new_n31456__ = ~new_new_n31454__ & ~new_new_n31455__;
  assign new_new_n31457__ = new_new_n31437__ & new_new_n31456__;
  assign new_new_n31458__ = ~new_new_n31437__ & ~new_new_n31456__;
  assign new_new_n31459__ = ~new_new_n31457__ & ~new_new_n31458__;
  assign new_new_n31460__ = new_new_n31317__ & ~new_new_n31459__;
  assign new_new_n31461__ = ~new_new_n31317__ & new_new_n31459__;
  assign new_new_n31462__ = ~new_new_n31460__ & ~new_new_n31461__;
  assign new_new_n31463__ = new_new_n6985__ & ~new_new_n26847__;
  assign new_new_n31464__ = ~new_new_n10772__ & ~new_new_n26823__;
  assign new_new_n31465__ = new_new_n10772__ & ~new_new_n29400__;
  assign new_new_n31466__ = new_new_n6994__ & ~new_new_n31464__;
  assign new_new_n31467__ = ~new_new_n31465__ & new_new_n31466__;
  assign new_new_n31468__ = ~new_new_n10998__ & new_new_n26854__;
  assign new_new_n31469__ = ~new_new_n20015__ & ~new_new_n31468__;
  assign new_new_n31470__ = ~new_new_n31463__ & new_new_n31469__;
  assign new_new_n31471__ = ~new_new_n31467__ & new_new_n31470__;
  assign new_new_n31472__ = ~pi14 & ~new_new_n31471__;
  assign new_new_n31473__ = pi14 & new_new_n31471__;
  assign new_new_n31474__ = ~new_new_n31472__ & ~new_new_n31473__;
  assign new_new_n31475__ = ~new_new_n30604__ & ~new_new_n30608__;
  assign new_new_n31476__ = ~new_new_n30605__ & ~new_new_n31475__;
  assign new_new_n31477__ = new_new_n31474__ & ~new_new_n31476__;
  assign new_new_n31478__ = ~new_new_n31474__ & new_new_n31476__;
  assign new_new_n31479__ = ~new_new_n31477__ & ~new_new_n31478__;
  assign new_new_n31480__ = new_new_n31462__ & new_new_n31479__;
  assign new_new_n31481__ = ~new_new_n31462__ & ~new_new_n31479__;
  assign new_new_n31482__ = ~new_new_n31480__ & ~new_new_n31481__;
  assign new_new_n31483__ = pi07 & ~new_new_n31482__;
  assign new_new_n31484__ = ~pi07 & new_new_n31482__;
  assign new_new_n31485__ = ~new_new_n31483__ & ~new_new_n31484__;
  assign new_new_n31486__ = new_new_n31296__ & ~new_new_n31485__;
  assign new_new_n31487__ = pi08 & new_new_n31482__;
  assign new_new_n31488__ = ~pi08 & ~new_new_n31482__;
  assign new_new_n31489__ = ~new_new_n31487__ & ~new_new_n31488__;
  assign new_new_n31490__ = ~new_new_n31296__ & new_new_n31489__;
  assign new_new_n31491__ = ~new_new_n31486__ & ~new_new_n31490__;
  assign new_new_n31492__ = new_new_n31295__ & ~new_new_n31491__;
  assign new_new_n31493__ = ~new_new_n31295__ & ~new_new_n31489__;
  assign new_new_n31494__ = ~new_new_n31492__ & ~new_new_n31493__;
  assign new_new_n31495__ = ~new_new_n30423__ & new_new_n30611__;
  assign new_new_n31496__ = ~new_new_n30424__ & ~new_new_n31495__;
  assign new_new_n31497__ = new_new_n31494__ & ~new_new_n31496__;
  assign new_new_n31498__ = ~new_new_n31494__ & new_new_n31496__;
  assign new_new_n31499__ = ~new_new_n31497__ & ~new_new_n31498__;
  assign new_new_n31500__ = new_new_n31290__ & new_new_n31499__;
  assign new_new_n31501__ = ~new_new_n31290__ & ~new_new_n31499__;
  assign new_new_n31502__ = ~new_new_n31500__ & ~new_new_n31501__;
  assign new_new_n31503__ = ~new_new_n27305__ & ~new_new_n31502__;
  assign new_new_n31504__ = new_new_n27305__ & new_new_n31502__;
  assign new_new_n31505__ = ~new_new_n31503__ & ~new_new_n31504__;
  assign new_new_n31506__ = pi01 & new_new_n27250__;
  assign new_new_n31507__ = ~pi00 & ~new_new_n31506__;
  assign new_new_n31508__ = ~new_new_n27277__ & ~new_new_n27279__;
  assign new_new_n31509__ = new_new_n26698__ & ~new_new_n31508__;
  assign new_new_n31510__ = ~new_new_n27277__ & new_new_n27280__;
  assign new_new_n31511__ = ~new_new_n31509__ & ~new_new_n31510__;
  assign new_new_n31512__ = pi00 & ~new_new_n26698__;
  assign new_new_n31513__ = ~new_new_n31511__ & new_new_n31512__;
  assign new_new_n31514__ = ~new_new_n31507__ & ~new_new_n31513__;
  assign new_new_n31515__ = ~pi02 & ~new_new_n31514__;
  assign new_new_n31516__ = ~pi01 & ~new_new_n27242__;
  assign new_new_n31517__ = new_new_n31507__ & ~new_new_n31516__;
  assign new_new_n31518__ = pi00 & ~new_new_n31511__;
  assign new_new_n31519__ = pi02 & ~new_new_n31517__;
  assign new_new_n31520__ = ~new_new_n31512__ & new_new_n31519__;
  assign new_new_n31521__ = ~new_new_n31518__ & new_new_n31520__;
  assign new_new_n31522__ = pi01 & new_new_n26698__;
  assign new_new_n31523__ = ~new_new_n27299__ & ~new_new_n31522__;
  assign new_new_n31524__ = pi00 & ~new_new_n31523__;
  assign new_new_n31525__ = ~new_new_n31508__ & new_new_n31524__;
  assign new_new_n31526__ = ~new_new_n31521__ & ~new_new_n31525__;
  assign new_new_n31527__ = ~new_new_n31515__ & new_new_n31526__;
  assign new_new_n31528__ = ~pi01 & ~new_new_n27250__;
  assign new_new_n31529__ = pi02 & new_new_n27250__;
  assign new_new_n31530__ = ~new_new_n31528__ & ~new_new_n31529__;
  assign new_new_n31531__ = ~new_new_n27271__ & new_new_n31530__;
  assign new_new_n31532__ = ~pi02 & ~new_new_n27250__;
  assign new_new_n31533__ = ~new_new_n31506__ & ~new_new_n31532__;
  assign new_new_n31534__ = new_new_n27271__ & new_new_n31533__;
  assign new_new_n31535__ = pi00 & ~new_new_n31531__;
  assign new_new_n31536__ = ~new_new_n31534__ & new_new_n31535__;
  assign new_new_n31537__ = pi02 & ~new_new_n27242__;
  assign new_new_n31538__ = ~pi02 & new_new_n27242__;
  assign new_new_n31539__ = pi01 & ~new_new_n31537__;
  assign new_new_n31540__ = ~new_new_n31538__ & new_new_n31539__;
  assign new_new_n31541__ = new_new_n12798__ & ~new_new_n26722__;
  assign new_new_n31542__ = ~pi00 & ~new_new_n31540__;
  assign new_new_n31543__ = ~new_new_n31541__ & new_new_n31542__;
  assign new_new_n31544__ = ~new_new_n31536__ & ~new_new_n31543__;
  assign new_new_n31545__ = ~new_new_n31255__ & ~new_new_n31256__;
  assign new_new_n31546__ = ~new_new_n31260__ & new_new_n31545__;
  assign new_new_n31547__ = new_new_n31260__ & ~new_new_n31545__;
  assign new_new_n31548__ = ~new_new_n31546__ & ~new_new_n31547__;
  assign new_new_n31549__ = ~new_new_n31544__ & new_new_n31548__;
  assign new_new_n31550__ = new_new_n31544__ & ~new_new_n31548__;
  assign new_new_n31551__ = pi02 & ~new_new_n27352__;
  assign new_new_n31552__ = pi01 & new_new_n27352__;
  assign new_new_n31553__ = ~new_new_n31551__ & ~new_new_n31552__;
  assign new_new_n31554__ = ~new_new_n27242__ & new_new_n31553__;
  assign new_new_n31555__ = new_new_n27242__ & ~new_new_n31553__;
  assign new_new_n31556__ = pi00 & ~new_new_n31554__;
  assign new_new_n31557__ = ~new_new_n31555__ & new_new_n31556__;
  assign new_new_n31558__ = new_new_n13508__ & new_new_n26722__;
  assign new_new_n31559__ = ~pi01 & ~new_new_n26729__;
  assign new_new_n31560__ = pi01 & ~new_new_n26722__;
  assign new_new_n31561__ = ~new_new_n31559__ & ~new_new_n31560__;
  assign new_new_n31562__ = pi02 & ~new_new_n31561__;
  assign new_new_n31563__ = ~pi00 & ~new_new_n31558__;
  assign new_new_n31564__ = ~new_new_n31562__ & new_new_n31563__;
  assign new_new_n31565__ = ~new_new_n31557__ & ~new_new_n31564__;
  assign new_new_n31566__ = ~new_new_n30668__ & ~new_new_n30669__;
  assign new_new_n31567__ = ~new_new_n31252__ & new_new_n31566__;
  assign new_new_n31568__ = new_new_n31252__ & ~new_new_n31566__;
  assign new_new_n31569__ = ~new_new_n31567__ & ~new_new_n31568__;
  assign new_new_n31570__ = ~new_new_n31565__ & ~new_new_n31569__;
  assign new_new_n31571__ = new_new_n31565__ & new_new_n31569__;
  assign new_new_n31572__ = pi01 & new_new_n26774__;
  assign new_new_n31573__ = ~pi01 & new_new_n26810__;
  assign new_new_n31574__ = pi02 & ~new_new_n31573__;
  assign new_new_n31575__ = ~new_new_n31572__ & ~new_new_n31574__;
  assign new_new_n31576__ = pi02 & new_new_n31572__;
  assign new_new_n31577__ = ~pi00 & ~new_new_n31575__;
  assign new_new_n31578__ = ~new_new_n31576__ & new_new_n31577__;
  assign new_new_n31579__ = ~new_new_n26774__ & new_new_n27330__;
  assign new_new_n31580__ = new_new_n26774__ & ~new_new_n27330__;
  assign new_new_n31581__ = ~new_new_n31579__ & ~new_new_n31580__;
  assign new_new_n31582__ = ~new_new_n27370__ & new_new_n31581__;
  assign new_new_n31583__ = pi01 & new_new_n26729__;
  assign new_new_n31584__ = ~new_new_n31559__ & ~new_new_n31583__;
  assign new_new_n31585__ = new_new_n31582__ & ~new_new_n31584__;
  assign new_new_n31586__ = pi02 & new_new_n26729__;
  assign new_new_n31587__ = ~pi02 & ~new_new_n26729__;
  assign new_new_n31588__ = ~new_new_n31586__ & ~new_new_n31587__;
  assign new_new_n31589__ = ~new_new_n31582__ & ~new_new_n31588__;
  assign new_new_n31590__ = pi00 & ~new_new_n31585__;
  assign new_new_n31591__ = ~new_new_n31589__ & new_new_n31590__;
  assign new_new_n31592__ = ~new_new_n31578__ & ~new_new_n31591__;
  assign new_new_n31593__ = new_new_n13508__ & new_new_n26810__;
  assign new_new_n31594__ = ~pi01 & new_new_n26802__;
  assign new_new_n31595__ = pi01 & ~new_new_n26810__;
  assign new_new_n31596__ = ~new_new_n31594__ & ~new_new_n31595__;
  assign new_new_n31597__ = pi02 & ~new_new_n31596__;
  assign new_new_n31598__ = ~new_new_n31593__ & ~new_new_n31597__;
  assign new_new_n31599__ = ~pi00 & ~new_new_n31598__;
  assign new_new_n31600__ = pi01 & new_new_n27373__;
  assign new_new_n31601__ = pi02 & ~new_new_n27373__;
  assign new_new_n31602__ = new_new_n26774__ & ~new_new_n31600__;
  assign new_new_n31603__ = ~new_new_n31601__ & new_new_n31602__;
  assign new_new_n31604__ = ~pi01 & ~new_new_n27373__;
  assign new_new_n31605__ = ~pi02 & new_new_n27373__;
  assign new_new_n31606__ = ~new_new_n26774__ & ~new_new_n31604__;
  assign new_new_n31607__ = ~new_new_n31605__ & new_new_n31606__;
  assign new_new_n31608__ = ~new_new_n31603__ & ~new_new_n31607__;
  assign new_new_n31609__ = pi00 & ~new_new_n31608__;
  assign new_new_n31610__ = ~new_new_n31599__ & ~new_new_n31609__;
  assign new_new_n31611__ = ~pi01 & ~new_new_n26741__;
  assign new_new_n31612__ = pi01 & ~new_new_n26802__;
  assign new_new_n31613__ = pi02 & ~new_new_n31611__;
  assign new_new_n31614__ = ~new_new_n31612__ & new_new_n31613__;
  assign new_new_n31615__ = new_new_n13508__ & ~new_new_n26802__;
  assign new_new_n31616__ = ~new_new_n31614__ & ~new_new_n31615__;
  assign new_new_n31617__ = ~pi00 & ~new_new_n31616__;
  assign new_new_n31618__ = pi02 & new_new_n27395__;
  assign new_new_n31619__ = pi01 & ~new_new_n27395__;
  assign new_new_n31620__ = new_new_n26810__ & ~new_new_n31618__;
  assign new_new_n31621__ = ~new_new_n31619__ & new_new_n31620__;
  assign new_new_n31622__ = ~pi02 & ~new_new_n27395__;
  assign new_new_n31623__ = ~pi01 & new_new_n27395__;
  assign new_new_n31624__ = ~new_new_n26810__ & ~new_new_n31622__;
  assign new_new_n31625__ = ~new_new_n31623__ & new_new_n31624__;
  assign new_new_n31626__ = ~new_new_n31621__ & ~new_new_n31625__;
  assign new_new_n31627__ = pi00 & ~new_new_n31626__;
  assign new_new_n31628__ = ~new_new_n31617__ & ~new_new_n31627__;
  assign new_new_n31629__ = ~new_new_n31195__ & ~new_new_n31196__;
  assign new_new_n31630__ = new_new_n31206__ & new_new_n31629__;
  assign new_new_n31631__ = ~new_new_n31206__ & ~new_new_n31629__;
  assign new_new_n31632__ = ~new_new_n31630__ & ~new_new_n31631__;
  assign new_new_n31633__ = ~new_new_n31628__ & new_new_n31632__;
  assign new_new_n31634__ = new_new_n31628__ & ~new_new_n31632__;
  assign new_new_n31635__ = pi01 & ~new_new_n26741__;
  assign new_new_n31636__ = ~pi01 & ~new_new_n27221__;
  assign new_new_n31637__ = pi02 & new_new_n31636__;
  assign new_new_n31638__ = ~new_new_n31635__ & ~new_new_n31637__;
  assign new_new_n31639__ = ~pi00 & ~new_new_n31638__;
  assign new_new_n31640__ = pi00 & ~new_new_n26802__;
  assign new_new_n31641__ = new_new_n30411__ & new_new_n31640__;
  assign new_new_n31642__ = ~new_new_n31639__ & ~new_new_n31641__;
  assign new_new_n31643__ = ~pi02 & ~new_new_n31642__;
  assign new_new_n31644__ = pi00 & ~new_new_n31594__;
  assign new_new_n31645__ = ~new_new_n31612__ & new_new_n31644__;
  assign new_new_n31646__ = new_new_n27390__ & new_new_n31645__;
  assign new_new_n31647__ = pi00 & ~new_new_n27391__;
  assign new_new_n31648__ = pi02 & ~new_new_n31639__;
  assign new_new_n31649__ = ~new_new_n31647__ & new_new_n31648__;
  assign new_new_n31650__ = ~new_new_n31646__ & ~new_new_n31649__;
  assign new_new_n31651__ = ~new_new_n31643__ & new_new_n31650__;
  assign new_new_n31652__ = pi02 & ~new_new_n30390__;
  assign new_new_n31653__ = pi01 & new_new_n30390__;
  assign new_new_n31654__ = ~new_new_n31652__ & ~new_new_n31653__;
  assign new_new_n31655__ = ~new_new_n26741__ & ~new_new_n31654__;
  assign new_new_n31656__ = new_new_n26741__ & new_new_n31654__;
  assign new_new_n31657__ = pi00 & ~new_new_n31655__;
  assign new_new_n31658__ = ~new_new_n31656__ & new_new_n31657__;
  assign new_new_n31659__ = ~pi02 & new_new_n27221__;
  assign new_new_n31660__ = pi01 & new_new_n27221__;
  assign new_new_n31661__ = ~pi01 & new_new_n26823__;
  assign new_new_n31662__ = pi02 & ~new_new_n31661__;
  assign new_new_n31663__ = ~new_new_n31660__ & new_new_n31662__;
  assign new_new_n31664__ = new_new_n25566__ & ~new_new_n31659__;
  assign new_new_n31665__ = ~new_new_n31663__ & new_new_n31664__;
  assign new_new_n31666__ = ~new_new_n31658__ & ~new_new_n31665__;
  assign new_new_n31667__ = ~new_new_n31165__ & ~new_new_n31166__;
  assign new_new_n31668__ = new_new_n31177__ & ~new_new_n31667__;
  assign new_new_n31669__ = ~new_new_n31177__ & new_new_n31667__;
  assign new_new_n31670__ = ~new_new_n31668__ & ~new_new_n31669__;
  assign new_new_n31671__ = ~new_new_n31666__ & new_new_n31670__;
  assign new_new_n31672__ = new_new_n31666__ & ~new_new_n31670__;
  assign new_new_n31673__ = ~new_new_n31144__ & ~new_new_n31145__;
  assign new_new_n31674__ = new_new_n31156__ & new_new_n31673__;
  assign new_new_n31675__ = ~new_new_n31156__ & ~new_new_n31673__;
  assign new_new_n31676__ = ~new_new_n31674__ & ~new_new_n31675__;
  assign new_new_n31677__ = ~pi02 & ~new_new_n29424__;
  assign new_new_n31678__ = ~pi01 & new_new_n29424__;
  assign new_new_n31679__ = ~new_new_n26847__ & ~new_new_n31677__;
  assign new_new_n31680__ = ~new_new_n31678__ & new_new_n31679__;
  assign new_new_n31681__ = pi02 & new_new_n29424__;
  assign new_new_n31682__ = pi01 & ~new_new_n29424__;
  assign new_new_n31683__ = new_new_n26847__ & ~new_new_n31681__;
  assign new_new_n31684__ = ~new_new_n31682__ & new_new_n31683__;
  assign new_new_n31685__ = ~new_new_n31680__ & ~new_new_n31684__;
  assign new_new_n31686__ = pi00 & ~new_new_n31685__;
  assign new_new_n31687__ = pi02 & new_new_n26854__;
  assign new_new_n31688__ = ~pi02 & ~new_new_n26854__;
  assign new_new_n31689__ = ~new_new_n31687__ & ~new_new_n31688__;
  assign new_new_n31690__ = pi01 & ~new_new_n31689__;
  assign new_new_n31691__ = new_new_n12798__ & new_new_n26888__;
  assign new_new_n31692__ = ~new_new_n31690__ & ~new_new_n31691__;
  assign new_new_n31693__ = ~pi00 & ~new_new_n31692__;
  assign new_new_n31694__ = ~new_new_n31686__ & ~new_new_n31693__;
  assign new_new_n31695__ = pi01 & ~new_new_n26888__;
  assign new_new_n31696__ = ~pi01 & new_new_n26922__;
  assign new_new_n31697__ = ~new_new_n31695__ & ~new_new_n31696__;
  assign new_new_n31698__ = pi02 & ~new_new_n31697__;
  assign new_new_n31699__ = ~pi02 & ~new_new_n31695__;
  assign new_new_n31700__ = ~pi00 & ~new_new_n31699__;
  assign new_new_n31701__ = ~new_new_n31698__ & new_new_n31700__;
  assign new_new_n31702__ = pi01 & ~new_new_n26854__;
  assign new_new_n31703__ = ~pi01 & new_new_n26854__;
  assign new_new_n31704__ = ~new_new_n31702__ & ~new_new_n31703__;
  assign new_new_n31705__ = new_new_n27421__ & ~new_new_n31704__;
  assign new_new_n31706__ = ~new_new_n27421__ & new_new_n31689__;
  assign new_new_n31707__ = pi00 & ~new_new_n31705__;
  assign new_new_n31708__ = ~new_new_n31706__ & new_new_n31707__;
  assign new_new_n31709__ = ~new_new_n31701__ & ~new_new_n31708__;
  assign new_new_n31710__ = ~new_new_n31101__ & ~new_new_n31102__;
  assign new_new_n31711__ = ~new_new_n31108__ & new_new_n31710__;
  assign new_new_n31712__ = new_new_n31108__ & ~new_new_n31710__;
  assign new_new_n31713__ = ~new_new_n31711__ & ~new_new_n31712__;
  assign new_new_n31714__ = ~new_new_n31709__ & ~new_new_n31713__;
  assign new_new_n31715__ = new_new_n31709__ & new_new_n31713__;
  assign new_new_n31716__ = pi02 & ~new_new_n27177__;
  assign new_new_n31717__ = pi01 & new_new_n27177__;
  assign new_new_n31718__ = ~new_new_n31716__ & ~new_new_n31717__;
  assign new_new_n31719__ = ~new_new_n26888__ & new_new_n31718__;
  assign new_new_n31720__ = new_new_n26888__ & ~new_new_n31718__;
  assign new_new_n31721__ = pi00 & ~new_new_n31719__;
  assign new_new_n31722__ = ~new_new_n31720__ & new_new_n31721__;
  assign new_new_n31723__ = new_new_n13508__ & new_new_n26922__;
  assign new_new_n31724__ = pi01 & new_new_n26922__;
  assign new_new_n31725__ = ~pi01 & ~new_new_n27168__;
  assign new_new_n31726__ = pi02 & ~new_new_n31725__;
  assign new_new_n31727__ = ~new_new_n31724__ & new_new_n31726__;
  assign new_new_n31728__ = ~pi00 & ~new_new_n31723__;
  assign new_new_n31729__ = ~new_new_n31727__ & new_new_n31728__;
  assign new_new_n31730__ = ~new_new_n31722__ & ~new_new_n31729__;
  assign new_new_n31731__ = new_new_n13508__ & ~new_new_n27168__;
  assign new_new_n31732__ = pi01 & new_new_n27168__;
  assign new_new_n31733__ = ~pi01 & ~new_new_n26917__;
  assign new_new_n31734__ = ~new_new_n31732__ & ~new_new_n31733__;
  assign new_new_n31735__ = pi02 & ~new_new_n31734__;
  assign new_new_n31736__ = ~new_new_n31731__ & ~new_new_n31735__;
  assign new_new_n31737__ = ~pi00 & ~new_new_n31736__;
  assign new_new_n31738__ = pi01 & new_new_n29366__;
  assign new_new_n31739__ = pi02 & ~new_new_n29366__;
  assign new_new_n31740__ = new_new_n26922__ & ~new_new_n31738__;
  assign new_new_n31741__ = ~new_new_n31739__ & new_new_n31740__;
  assign new_new_n31742__ = ~pi01 & ~new_new_n29366__;
  assign new_new_n31743__ = ~pi02 & new_new_n29366__;
  assign new_new_n31744__ = ~new_new_n26922__ & ~new_new_n31742__;
  assign new_new_n31745__ = ~new_new_n31743__ & new_new_n31744__;
  assign new_new_n31746__ = ~new_new_n31741__ & ~new_new_n31745__;
  assign new_new_n31747__ = pi00 & ~new_new_n31746__;
  assign new_new_n31748__ = ~new_new_n31737__ & ~new_new_n31747__;
  assign new_new_n31749__ = ~pi02 & ~new_new_n28799__;
  assign new_new_n31750__ = ~pi01 & new_new_n28799__;
  assign new_new_n31751__ = ~new_new_n27168__ & ~new_new_n31749__;
  assign new_new_n31752__ = ~new_new_n31750__ & new_new_n31751__;
  assign new_new_n31753__ = pi02 & new_new_n28799__;
  assign new_new_n31754__ = pi01 & ~new_new_n28799__;
  assign new_new_n31755__ = new_new_n27168__ & ~new_new_n31753__;
  assign new_new_n31756__ = ~new_new_n31754__ & new_new_n31755__;
  assign new_new_n31757__ = ~new_new_n31752__ & ~new_new_n31756__;
  assign new_new_n31758__ = pi00 & ~new_new_n31757__;
  assign new_new_n31759__ = new_new_n13508__ & new_new_n26917__;
  assign new_new_n31760__ = ~pi01 & new_new_n26928__;
  assign new_new_n31761__ = pi01 & new_new_n26917__;
  assign new_new_n31762__ = pi02 & ~new_new_n31760__;
  assign new_new_n31763__ = ~new_new_n31761__ & new_new_n31762__;
  assign new_new_n31764__ = ~pi00 & ~new_new_n31759__;
  assign new_new_n31765__ = ~new_new_n31763__ & new_new_n31764__;
  assign new_new_n31766__ = ~new_new_n31758__ & ~new_new_n31765__;
  assign new_new_n31767__ = ~new_new_n31076__ & ~new_new_n31077__;
  assign new_new_n31768__ = new_new_n31088__ & new_new_n31767__;
  assign new_new_n31769__ = ~new_new_n31088__ & ~new_new_n31767__;
  assign new_new_n31770__ = ~new_new_n31768__ & ~new_new_n31769__;
  assign new_new_n31771__ = ~new_new_n31766__ & ~new_new_n31770__;
  assign new_new_n31772__ = new_new_n31766__ & new_new_n31770__;
  assign new_new_n31773__ = pi02 & new_new_n26941__;
  assign new_new_n31774__ = ~pi02 & ~new_new_n26941__;
  assign new_new_n31775__ = ~new_new_n31773__ & ~new_new_n31774__;
  assign new_new_n31776__ = pi01 & ~new_new_n31775__;
  assign new_new_n31777__ = new_new_n12798__ & ~new_new_n27152__;
  assign new_new_n31778__ = ~new_new_n31776__ & ~new_new_n31777__;
  assign new_new_n31779__ = ~pi00 & ~new_new_n31778__;
  assign new_new_n31780__ = pi02 & ~new_new_n26928__;
  assign new_new_n31781__ = ~new_new_n31760__ & ~new_new_n31780__;
  assign new_new_n31782__ = ~new_new_n27488__ & new_new_n31781__;
  assign new_new_n31783__ = pi01 & ~new_new_n26928__;
  assign new_new_n31784__ = ~pi02 & new_new_n26928__;
  assign new_new_n31785__ = ~new_new_n31783__ & ~new_new_n31784__;
  assign new_new_n31786__ = new_new_n27488__ & new_new_n31785__;
  assign new_new_n31787__ = pi00 & ~new_new_n31782__;
  assign new_new_n31788__ = ~new_new_n31786__ & new_new_n31787__;
  assign new_new_n31789__ = ~new_new_n31779__ & ~new_new_n31788__;
  assign new_new_n31790__ = new_new_n13508__ & new_new_n27152__;
  assign new_new_n31791__ = ~pi01 & new_new_n26937__;
  assign new_new_n31792__ = pi01 & ~new_new_n27152__;
  assign new_new_n31793__ = ~new_new_n31791__ & ~new_new_n31792__;
  assign new_new_n31794__ = pi02 & ~new_new_n31793__;
  assign new_new_n31795__ = ~new_new_n31790__ & ~new_new_n31794__;
  assign new_new_n31796__ = ~pi00 & ~new_new_n31795__;
  assign new_new_n31797__ = ~pi01 & new_new_n26941__;
  assign new_new_n31798__ = pi01 & ~new_new_n26941__;
  assign new_new_n31799__ = ~new_new_n31797__ & ~new_new_n31798__;
  assign new_new_n31800__ = new_new_n27481__ & ~new_new_n31799__;
  assign new_new_n31801__ = ~new_new_n27481__ & new_new_n31775__;
  assign new_new_n31802__ = pi00 & ~new_new_n31800__;
  assign new_new_n31803__ = ~new_new_n31801__ & new_new_n31802__;
  assign new_new_n31804__ = ~new_new_n31796__ & ~new_new_n31803__;
  assign new_new_n31805__ = ~new_new_n30815__ & ~new_new_n30816__;
  assign new_new_n31806__ = ~new_new_n31043__ & new_new_n31805__;
  assign new_new_n31807__ = new_new_n31043__ & ~new_new_n31805__;
  assign new_new_n31808__ = ~new_new_n31806__ & ~new_new_n31807__;
  assign new_new_n31809__ = new_new_n31804__ & ~new_new_n31808__;
  assign new_new_n31810__ = ~new_new_n31804__ & new_new_n31808__;
  assign new_new_n31811__ = pi02 & ~new_new_n27477__;
  assign new_new_n31812__ = pi01 & new_new_n27477__;
  assign new_new_n31813__ = ~new_new_n31811__ & ~new_new_n31812__;
  assign new_new_n31814__ = new_new_n27152__ & new_new_n31813__;
  assign new_new_n31815__ = ~new_new_n27152__ & ~new_new_n31813__;
  assign new_new_n31816__ = pi00 & ~new_new_n31814__;
  assign new_new_n31817__ = ~new_new_n31815__ & new_new_n31816__;
  assign new_new_n31818__ = new_new_n13508__ & ~new_new_n26937__;
  assign new_new_n31819__ = ~pi01 & new_new_n26971__;
  assign new_new_n31820__ = pi01 & ~new_new_n26937__;
  assign new_new_n31821__ = pi02 & ~new_new_n31819__;
  assign new_new_n31822__ = ~new_new_n31820__ & new_new_n31821__;
  assign new_new_n31823__ = ~pi00 & ~new_new_n31818__;
  assign new_new_n31824__ = ~new_new_n31822__ & new_new_n31823__;
  assign new_new_n31825__ = ~new_new_n31817__ & ~new_new_n31824__;
  assign new_new_n31826__ = ~pi01 & ~new_new_n27003__;
  assign new_new_n31827__ = pi01 & ~new_new_n26978__;
  assign new_new_n31828__ = pi02 & ~new_new_n31826__;
  assign new_new_n31829__ = ~new_new_n31827__ & new_new_n31828__;
  assign new_new_n31830__ = new_new_n13508__ & ~new_new_n26978__;
  assign new_new_n31831__ = ~new_new_n31829__ & ~new_new_n31830__;
  assign new_new_n31832__ = ~pi00 & ~new_new_n31831__;
  assign new_new_n31833__ = pi02 & ~new_new_n26971__;
  assign new_new_n31834__ = ~new_new_n31819__ & ~new_new_n31833__;
  assign new_new_n31835__ = ~new_new_n28277__ & new_new_n31834__;
  assign new_new_n31836__ = pi01 & ~new_new_n26971__;
  assign new_new_n31837__ = ~pi02 & new_new_n26971__;
  assign new_new_n31838__ = ~new_new_n31836__ & ~new_new_n31837__;
  assign new_new_n31839__ = new_new_n28277__ & new_new_n31838__;
  assign new_new_n31840__ = pi00 & ~new_new_n31835__;
  assign new_new_n31841__ = ~new_new_n31839__ & new_new_n31840__;
  assign new_new_n31842__ = ~new_new_n31832__ & ~new_new_n31841__;
  assign new_new_n31843__ = ~new_new_n30995__ & ~new_new_n30996__;
  assign new_new_n31844__ = new_new_n31007__ & new_new_n31843__;
  assign new_new_n31845__ = ~new_new_n31007__ & ~new_new_n31843__;
  assign new_new_n31846__ = ~new_new_n31844__ & ~new_new_n31845__;
  assign new_new_n31847__ = ~new_new_n31842__ & new_new_n31846__;
  assign new_new_n31848__ = new_new_n31842__ & ~new_new_n31846__;
  assign new_new_n31849__ = new_new_n13508__ & ~new_new_n27003__;
  assign new_new_n31850__ = ~pi01 & ~new_new_n27029__;
  assign new_new_n31851__ = pi01 & ~new_new_n27003__;
  assign new_new_n31852__ = pi02 & ~new_new_n31850__;
  assign new_new_n31853__ = ~new_new_n31851__ & new_new_n31852__;
  assign new_new_n31854__ = ~pi00 & ~new_new_n31849__;
  assign new_new_n31855__ = ~new_new_n31853__ & new_new_n31854__;
  assign new_new_n31856__ = ~pi02 & new_new_n26978__;
  assign new_new_n31857__ = ~new_new_n31827__ & ~new_new_n31856__;
  assign new_new_n31858__ = ~new_new_n27986__ & new_new_n31857__;
  assign new_new_n31859__ = ~pi01 & new_new_n26978__;
  assign new_new_n31860__ = pi02 & ~new_new_n26978__;
  assign new_new_n31861__ = ~new_new_n31859__ & ~new_new_n31860__;
  assign new_new_n31862__ = new_new_n27986__ & new_new_n31861__;
  assign new_new_n31863__ = pi00 & ~new_new_n31858__;
  assign new_new_n31864__ = ~new_new_n31862__ & new_new_n31863__;
  assign new_new_n31865__ = ~new_new_n31855__ & ~new_new_n31864__;
  assign new_new_n31866__ = ~new_new_n30983__ & ~new_new_n30984__;
  assign new_new_n31867__ = new_new_n30988__ & new_new_n31866__;
  assign new_new_n31868__ = ~new_new_n30988__ & ~new_new_n31866__;
  assign new_new_n31869__ = ~new_new_n31867__ & ~new_new_n31868__;
  assign new_new_n31870__ = new_new_n31865__ & ~new_new_n31869__;
  assign new_new_n31871__ = ~new_new_n31865__ & new_new_n31869__;
  assign new_new_n31872__ = ~pi02 & ~new_new_n27003__;
  assign new_new_n31873__ = pi01 & new_new_n27003__;
  assign new_new_n31874__ = ~new_new_n31872__ & ~new_new_n31873__;
  assign new_new_n31875__ = new_new_n27962__ & new_new_n31874__;
  assign new_new_n31876__ = pi02 & new_new_n27003__;
  assign new_new_n31877__ = ~new_new_n31826__ & ~new_new_n31876__;
  assign new_new_n31878__ = ~new_new_n27962__ & new_new_n31877__;
  assign new_new_n31879__ = ~new_new_n31875__ & ~new_new_n31878__;
  assign new_new_n31880__ = pi00 & ~new_new_n31879__;
  assign new_new_n31881__ = new_new_n13508__ & ~new_new_n27029__;
  assign new_new_n31882__ = ~pi01 & new_new_n27021__;
  assign new_new_n31883__ = pi01 & new_new_n27029__;
  assign new_new_n31884__ = ~new_new_n31882__ & ~new_new_n31883__;
  assign new_new_n31885__ = pi02 & ~new_new_n31884__;
  assign new_new_n31886__ = ~pi00 & ~new_new_n31881__;
  assign new_new_n31887__ = ~new_new_n31885__ & new_new_n31886__;
  assign new_new_n31888__ = ~new_new_n31880__ & ~new_new_n31887__;
  assign new_new_n31889__ = ~pi02 & ~new_new_n27021__;
  assign new_new_n31890__ = pi02 & new_new_n27021__;
  assign new_new_n31891__ = ~new_new_n31889__ & ~new_new_n31890__;
  assign new_new_n31892__ = pi01 & ~new_new_n31891__;
  assign new_new_n31893__ = new_new_n12798__ & ~new_new_n27111__;
  assign new_new_n31894__ = ~new_new_n31892__ & ~new_new_n31893__;
  assign new_new_n31895__ = ~pi00 & ~new_new_n31894__;
  assign new_new_n31896__ = pi02 & new_new_n27029__;
  assign new_new_n31897__ = ~new_new_n31850__ & ~new_new_n31896__;
  assign new_new_n31898__ = ~new_new_n27764__ & new_new_n31897__;
  assign new_new_n31899__ = ~pi02 & ~new_new_n27029__;
  assign new_new_n31900__ = ~new_new_n31883__ & ~new_new_n31899__;
  assign new_new_n31901__ = new_new_n27764__ & new_new_n31900__;
  assign new_new_n31902__ = pi00 & ~new_new_n31898__;
  assign new_new_n31903__ = ~new_new_n31901__ & new_new_n31902__;
  assign new_new_n31904__ = ~new_new_n31895__ & ~new_new_n31903__;
  assign new_new_n31905__ = new_new_n30068__ & new_new_n30896__;
  assign new_new_n31906__ = ~new_new_n30896__ & new_new_n30973__;
  assign new_new_n31907__ = ~new_new_n30976__ & ~new_new_n31906__;
  assign new_new_n31908__ = new_new_n30069__ & new_new_n31907__;
  assign new_new_n31909__ = ~new_new_n30069__ & ~new_new_n31907__;
  assign new_new_n31910__ = ~new_new_n31908__ & ~new_new_n31909__;
  assign new_new_n31911__ = new_new_n30081__ & ~new_new_n31905__;
  assign new_new_n31912__ = new_new_n31910__ & new_new_n31911__;
  assign new_new_n31913__ = new_new_n30054__ & new_new_n30068__;
  assign new_new_n31914__ = ~new_new_n30896__ & new_new_n31913__;
  assign new_new_n31915__ = ~new_new_n30973__ & new_new_n31914__;
  assign new_new_n31916__ = ~new_new_n30081__ & ~new_new_n31913__;
  assign new_new_n31917__ = ~new_new_n31910__ & new_new_n31916__;
  assign new_new_n31918__ = ~new_new_n31912__ & ~new_new_n31915__;
  assign new_new_n31919__ = ~new_new_n31917__ & new_new_n31918__;
  assign new_new_n31920__ = ~new_new_n31904__ & new_new_n31919__;
  assign new_new_n31921__ = new_new_n31904__ & ~new_new_n31919__;
  assign new_new_n31922__ = ~new_new_n30924__ & ~new_new_n30925__;
  assign new_new_n31923__ = new_new_n30924__ & new_new_n30925__;
  assign new_new_n31924__ = ~new_new_n31922__ & ~new_new_n31923__;
  assign new_new_n31925__ = pi02 & new_new_n27102__;
  assign new_new_n31926__ = pi01 & ~new_new_n27102__;
  assign new_new_n31927__ = ~new_new_n31925__ & ~new_new_n31926__;
  assign new_new_n31928__ = ~new_new_n27033__ & ~new_new_n31927__;
  assign new_new_n31929__ = new_new_n27033__ & new_new_n31927__;
  assign new_new_n31930__ = pi00 & ~new_new_n31928__;
  assign new_new_n31931__ = ~new_new_n31929__ & new_new_n31930__;
  assign new_new_n31932__ = pi01 & ~new_new_n27054__;
  assign new_new_n31933__ = ~pi02 & ~new_new_n31932__;
  assign new_new_n31934__ = ~pi01 & new_new_n27038__;
  assign new_new_n31935__ = ~new_new_n31932__ & ~new_new_n31934__;
  assign new_new_n31936__ = pi02 & ~new_new_n31935__;
  assign new_new_n31937__ = ~pi00 & ~new_new_n31933__;
  assign new_new_n31938__ = ~new_new_n31936__ & new_new_n31937__;
  assign new_new_n31939__ = ~new_new_n31931__ & ~new_new_n31938__;
  assign new_new_n31940__ = new_new_n31922__ & ~new_new_n31939__;
  assign new_new_n31941__ = new_new_n12798__ & ~new_new_n27071__;
  assign new_new_n31942__ = pi01 & new_new_n27041__;
  assign new_new_n31943__ = ~pi00 & ~new_new_n31941__;
  assign new_new_n31944__ = ~new_new_n31942__ & new_new_n31943__;
  assign new_new_n31945__ = new_new_n25294__ & ~new_new_n27054__;
  assign new_new_n31946__ = ~new_new_n25294__ & ~new_new_n27094__;
  assign new_new_n31947__ = pi00 & ~new_new_n31945__;
  assign new_new_n31948__ = ~new_new_n31946__ & new_new_n31947__;
  assign new_new_n31949__ = ~new_new_n31944__ & ~new_new_n31948__;
  assign new_new_n31950__ = new_new_n12798__ & new_new_n27059__;
  assign new_new_n31951__ = pi01 & ~new_new_n27071__;
  assign new_new_n31952__ = ~pi00 & ~new_new_n31950__;
  assign new_new_n31953__ = ~new_new_n31951__ & new_new_n31952__;
  assign new_new_n31954__ = ~new_new_n25294__ & new_new_n27567__;
  assign new_new_n31955__ = new_new_n25294__ & new_new_n27041__;
  assign new_new_n31956__ = pi00 & ~new_new_n31955__;
  assign new_new_n31957__ = ~new_new_n31954__ & new_new_n31956__;
  assign new_new_n31958__ = ~new_new_n31953__ & ~new_new_n31957__;
  assign new_new_n31959__ = new_new_n14117__ & ~new_new_n30927__;
  assign new_new_n31960__ = new_new_n30938__ & ~new_new_n31959__;
  assign new_new_n31961__ = pi05 & new_new_n30928__;
  assign new_new_n31962__ = ~new_new_n30938__ & new_new_n31961__;
  assign new_new_n31963__ = ~new_new_n31960__ & ~new_new_n31962__;
  assign new_new_n31964__ = new_new_n31958__ & new_new_n31963__;
  assign new_new_n31965__ = pi02 & ~new_new_n31958__;
  assign new_new_n31966__ = ~new_new_n31964__ & ~new_new_n31965__;
  assign new_new_n31967__ = ~new_new_n31949__ & ~new_new_n31966__;
  assign new_new_n31968__ = pi02 & new_new_n31958__;
  assign new_new_n31969__ = ~new_new_n31958__ & ~new_new_n31963__;
  assign new_new_n31970__ = new_new_n31949__ & ~new_new_n31968__;
  assign new_new_n31971__ = ~new_new_n31969__ & new_new_n31970__;
  assign new_new_n31972__ = ~new_new_n31967__ & ~new_new_n31971__;
  assign new_new_n31973__ = ~new_new_n25294__ & new_new_n28441__;
  assign new_new_n31974__ = new_new_n27071__ & ~new_new_n31973__;
  assign new_new_n31975__ = ~new_new_n27071__ & new_new_n31973__;
  assign new_new_n31976__ = pi00 & ~new_new_n31974__;
  assign new_new_n31977__ = ~new_new_n31975__ & new_new_n31976__;
  assign new_new_n31978__ = pi02 & new_new_n27577__;
  assign new_new_n31979__ = ~new_new_n27059__ & new_new_n31978__;
  assign new_new_n31980__ = new_new_n25581__ & new_new_n26118__;
  assign new_new_n31981__ = new_new_n25583__ & new_new_n27059__;
  assign new_new_n31982__ = ~new_new_n31980__ & ~new_new_n31981__;
  assign new_new_n31983__ = new_new_n11481__ & ~new_new_n27075__;
  assign new_new_n31984__ = new_new_n31982__ & new_new_n31983__;
  assign new_new_n31985__ = ~new_new_n31979__ & ~new_new_n31984__;
  assign new_new_n31986__ = ~new_new_n31977__ & ~new_new_n31985__;
  assign new_new_n31987__ = ~new_new_n31977__ & new_new_n31982__;
  assign new_new_n31988__ = new_new_n11480__ & ~new_new_n27075__;
  assign new_new_n31989__ = ~new_new_n31987__ & new_new_n31988__;
  assign new_new_n31990__ = ~new_new_n31986__ & ~new_new_n31989__;
  assign new_new_n31991__ = ~new_new_n31972__ & ~new_new_n31990__;
  assign new_new_n31992__ = ~pi02 & new_new_n31949__;
  assign new_new_n31993__ = pi02 & ~new_new_n31949__;
  assign new_new_n31994__ = ~new_new_n31992__ & ~new_new_n31993__;
  assign new_new_n31995__ = new_new_n31963__ & ~new_new_n31994__;
  assign new_new_n31996__ = new_new_n11474__ & new_new_n27087__;
  assign new_new_n31997__ = ~new_new_n10726__ & new_new_n26118__;
  assign new_new_n31998__ = new_new_n11473__ & ~new_new_n31997__;
  assign new_new_n31999__ = new_new_n31958__ & new_new_n31990__;
  assign new_new_n32000__ = pi02 & ~new_new_n31999__;
  assign new_new_n32001__ = ~new_new_n31964__ & ~new_new_n32000__;
  assign new_new_n32002__ = ~new_new_n31949__ & ~new_new_n32001__;
  assign new_new_n32003__ = ~new_new_n31963__ & ~new_new_n31992__;
  assign new_new_n32004__ = ~new_new_n31990__ & ~new_new_n32003__;
  assign new_new_n32005__ = ~new_new_n31971__ & ~new_new_n32002__;
  assign new_new_n32006__ = ~new_new_n32004__ & new_new_n32005__;
  assign new_new_n32007__ = ~new_new_n12828__ & ~new_new_n30927__;
  assign new_new_n32008__ = ~new_new_n31996__ & ~new_new_n31998__;
  assign new_new_n32009__ = new_new_n32007__ & new_new_n32008__;
  assign new_new_n32010__ = ~new_new_n32006__ & new_new_n32009__;
  assign new_new_n32011__ = ~new_new_n31991__ & ~new_new_n31995__;
  assign new_new_n32012__ = ~new_new_n32010__ & new_new_n32011__;
  assign new_new_n32013__ = ~new_new_n31940__ & new_new_n32012__;
  assign new_new_n32014__ = ~new_new_n30940__ & ~new_new_n31924__;
  assign new_new_n32015__ = ~new_new_n32013__ & new_new_n32014__;
  assign new_new_n32016__ = new_new_n30940__ & ~new_new_n31922__;
  assign new_new_n32017__ = ~new_new_n31923__ & ~new_new_n32016__;
  assign new_new_n32018__ = new_new_n32012__ & new_new_n32017__;
  assign new_new_n32019__ = ~new_new_n31939__ & ~new_new_n32018__;
  assign new_new_n32020__ = ~new_new_n32015__ & ~new_new_n32019__;
  assign new_new_n32021__ = new_new_n13508__ & ~new_new_n27033__;
  assign new_new_n32022__ = ~pi01 & ~new_new_n27054__;
  assign new_new_n32023__ = pi01 & ~new_new_n27033__;
  assign new_new_n32024__ = pi02 & ~new_new_n32022__;
  assign new_new_n32025__ = ~new_new_n32023__ & new_new_n32024__;
  assign new_new_n32026__ = ~pi00 & ~new_new_n32021__;
  assign new_new_n32027__ = ~new_new_n32025__ & new_new_n32026__;
  assign new_new_n32028__ = pi02 & ~new_new_n27686__;
  assign new_new_n32029__ = pi01 & new_new_n27686__;
  assign new_new_n32030__ = ~new_new_n32028__ & ~new_new_n32029__;
  assign new_new_n32031__ = new_new_n27111__ & new_new_n32030__;
  assign new_new_n32032__ = ~new_new_n27111__ & ~new_new_n32030__;
  assign new_new_n32033__ = pi00 & ~new_new_n32031__;
  assign new_new_n32034__ = ~new_new_n32032__ & new_new_n32033__;
  assign new_new_n32035__ = ~new_new_n32027__ & ~new_new_n32034__;
  assign new_new_n32036__ = new_new_n32020__ & ~new_new_n32035__;
  assign new_new_n32037__ = ~new_new_n32020__ & new_new_n32035__;
  assign new_new_n32038__ = ~new_new_n30943__ & ~new_new_n30944__;
  assign new_new_n32039__ = new_new_n30952__ & ~new_new_n32038__;
  assign new_new_n32040__ = ~new_new_n30952__ & new_new_n32038__;
  assign new_new_n32041__ = ~new_new_n32039__ & ~new_new_n32040__;
  assign new_new_n32042__ = ~new_new_n32037__ & new_new_n32041__;
  assign new_new_n32043__ = ~pi01 & ~new_new_n27033__;
  assign new_new_n32044__ = pi02 & ~new_new_n32043__;
  assign new_new_n32045__ = pi01 & new_new_n27111__;
  assign new_new_n32046__ = ~new_new_n32044__ & ~new_new_n32045__;
  assign new_new_n32047__ = pi02 & new_new_n32045__;
  assign new_new_n32048__ = ~pi00 & ~new_new_n32046__;
  assign new_new_n32049__ = ~new_new_n32047__ & new_new_n32048__;
  assign new_new_n32050__ = ~new_new_n27686__ & ~new_new_n27743__;
  assign new_new_n32051__ = new_new_n31891__ & ~new_new_n32050__;
  assign new_new_n32052__ = pi01 & ~new_new_n27020__;
  assign new_new_n32053__ = ~new_new_n31882__ & ~new_new_n32052__;
  assign new_new_n32054__ = new_new_n32050__ & ~new_new_n32053__;
  assign new_new_n32055__ = pi00 & ~new_new_n32051__;
  assign new_new_n32056__ = ~new_new_n32054__ & new_new_n32055__;
  assign new_new_n32057__ = ~new_new_n32049__ & ~new_new_n32056__;
  assign new_new_n32058__ = ~new_new_n30960__ & ~new_new_n30961__;
  assign new_new_n32059__ = ~new_new_n30971__ & new_new_n32058__;
  assign new_new_n32060__ = new_new_n30971__ & ~new_new_n32058__;
  assign new_new_n32061__ = ~new_new_n32059__ & ~new_new_n32060__;
  assign new_new_n32062__ = new_new_n32057__ & new_new_n32061__;
  assign new_new_n32063__ = ~new_new_n32036__ & ~new_new_n32062__;
  assign new_new_n32064__ = ~new_new_n32042__ & new_new_n32063__;
  assign new_new_n32065__ = ~new_new_n32057__ & ~new_new_n32061__;
  assign new_new_n32066__ = ~new_new_n32064__ & ~new_new_n32065__;
  assign new_new_n32067__ = ~new_new_n31921__ & ~new_new_n32066__;
  assign new_new_n32068__ = ~new_new_n31920__ & ~new_new_n32067__;
  assign new_new_n32069__ = new_new_n31888__ & ~new_new_n32068__;
  assign new_new_n32070__ = ~new_new_n31888__ & new_new_n32068__;
  assign new_new_n32071__ = ~new_new_n30879__ & ~new_new_n30880__;
  assign new_new_n32072__ = new_new_n30980__ & ~new_new_n32071__;
  assign new_new_n32073__ = ~new_new_n30980__ & new_new_n32071__;
  assign new_new_n32074__ = ~new_new_n32072__ & ~new_new_n32073__;
  assign new_new_n32075__ = ~new_new_n32070__ & new_new_n32074__;
  assign new_new_n32076__ = ~new_new_n32069__ & ~new_new_n32075__;
  assign new_new_n32077__ = ~new_new_n31871__ & ~new_new_n32076__;
  assign new_new_n32078__ = ~new_new_n31870__ & ~new_new_n32077__;
  assign new_new_n32079__ = ~new_new_n31848__ & ~new_new_n32078__;
  assign new_new_n32080__ = new_new_n13508__ & new_new_n26971__;
  assign new_new_n32081__ = ~new_new_n31836__ & ~new_new_n31859__;
  assign new_new_n32082__ = pi02 & ~new_new_n32081__;
  assign new_new_n32083__ = ~pi00 & ~new_new_n32080__;
  assign new_new_n32084__ = ~new_new_n32082__ & new_new_n32083__;
  assign new_new_n32085__ = ~pi02 & new_new_n26937__;
  assign new_new_n32086__ = ~new_new_n31820__ & ~new_new_n32085__;
  assign new_new_n32087__ = ~new_new_n28005__ & new_new_n32086__;
  assign new_new_n32088__ = pi02 & ~new_new_n26937__;
  assign new_new_n32089__ = ~new_new_n31791__ & ~new_new_n32088__;
  assign new_new_n32090__ = new_new_n28005__ & new_new_n32089__;
  assign new_new_n32091__ = pi00 & ~new_new_n32087__;
  assign new_new_n32092__ = ~new_new_n32090__ & new_new_n32091__;
  assign new_new_n32093__ = ~new_new_n32084__ & ~new_new_n32092__;
  assign new_new_n32094__ = ~new_new_n31010__ & ~new_new_n31011__;
  assign new_new_n32095__ = ~new_new_n31021__ & new_new_n32094__;
  assign new_new_n32096__ = new_new_n31021__ & ~new_new_n32094__;
  assign new_new_n32097__ = ~new_new_n32095__ & ~new_new_n32096__;
  assign new_new_n32098__ = new_new_n32093__ & ~new_new_n32097__;
  assign new_new_n32099__ = ~new_new_n31847__ & ~new_new_n32079__;
  assign new_new_n32100__ = ~new_new_n32098__ & new_new_n32099__;
  assign new_new_n32101__ = ~new_new_n32093__ & new_new_n32097__;
  assign new_new_n32102__ = ~new_new_n32100__ & ~new_new_n32101__;
  assign new_new_n32103__ = ~new_new_n31825__ & ~new_new_n32102__;
  assign new_new_n32104__ = new_new_n31825__ & new_new_n32102__;
  assign new_new_n32105__ = ~new_new_n31024__ & ~new_new_n31025__;
  assign new_new_n32106__ = new_new_n31041__ & new_new_n32105__;
  assign new_new_n32107__ = ~new_new_n31041__ & ~new_new_n32105__;
  assign new_new_n32108__ = ~new_new_n32106__ & ~new_new_n32107__;
  assign new_new_n32109__ = ~new_new_n32104__ & new_new_n32108__;
  assign new_new_n32110__ = ~new_new_n32103__ & ~new_new_n32109__;
  assign new_new_n32111__ = ~new_new_n31810__ & ~new_new_n32110__;
  assign new_new_n32112__ = ~new_new_n31809__ & ~new_new_n32111__;
  assign new_new_n32113__ = new_new_n31789__ & ~new_new_n32112__;
  assign new_new_n32114__ = ~new_new_n31789__ & new_new_n32112__;
  assign new_new_n32115__ = ~new_new_n31046__ & ~new_new_n31047__;
  assign new_new_n32116__ = new_new_n31059__ & ~new_new_n32115__;
  assign new_new_n32117__ = ~new_new_n31059__ & new_new_n32115__;
  assign new_new_n32118__ = ~new_new_n32116__ & ~new_new_n32117__;
  assign new_new_n32119__ = ~new_new_n32114__ & ~new_new_n32118__;
  assign new_new_n32120__ = ~new_new_n32113__ & ~new_new_n32119__;
  assign new_new_n32121__ = ~new_new_n30793__ & ~new_new_n30794__;
  assign new_new_n32122__ = ~new_new_n31061__ & new_new_n32121__;
  assign new_new_n32123__ = new_new_n31061__ & ~new_new_n32121__;
  assign new_new_n32124__ = ~new_new_n32122__ & ~new_new_n32123__;
  assign new_new_n32125__ = ~new_new_n32120__ & new_new_n32124__;
  assign new_new_n32126__ = new_new_n32120__ & ~new_new_n32124__;
  assign new_new_n32127__ = new_new_n13508__ & new_new_n26928__;
  assign new_new_n32128__ = ~new_new_n31783__ & ~new_new_n31797__;
  assign new_new_n32129__ = pi02 & ~new_new_n32128__;
  assign new_new_n32130__ = ~pi00 & ~new_new_n32127__;
  assign new_new_n32131__ = ~new_new_n32129__ & new_new_n32130__;
  assign new_new_n32132__ = pi02 & new_new_n26917__;
  assign new_new_n32133__ = ~new_new_n31733__ & ~new_new_n32132__;
  assign new_new_n32134__ = ~new_new_n27462__ & new_new_n32133__;
  assign new_new_n32135__ = ~pi02 & ~new_new_n26917__;
  assign new_new_n32136__ = ~new_new_n31761__ & ~new_new_n32135__;
  assign new_new_n32137__ = new_new_n27462__ & new_new_n32136__;
  assign new_new_n32138__ = pi00 & ~new_new_n32134__;
  assign new_new_n32139__ = ~new_new_n32137__ & new_new_n32138__;
  assign new_new_n32140__ = ~new_new_n32131__ & ~new_new_n32139__;
  assign new_new_n32141__ = ~new_new_n32126__ & ~new_new_n32140__;
  assign new_new_n32142__ = ~new_new_n32125__ & ~new_new_n32141__;
  assign new_new_n32143__ = ~new_new_n31772__ & ~new_new_n32142__;
  assign new_new_n32144__ = ~new_new_n31771__ & ~new_new_n32143__;
  assign new_new_n32145__ = ~new_new_n31748__ & new_new_n32144__;
  assign new_new_n32146__ = new_new_n31748__ & ~new_new_n32144__;
  assign new_new_n32147__ = ~new_new_n31091__ & ~new_new_n31092__;
  assign new_new_n32148__ = new_new_n31096__ & new_new_n32147__;
  assign new_new_n32149__ = ~new_new_n31096__ & ~new_new_n32147__;
  assign new_new_n32150__ = ~new_new_n32148__ & ~new_new_n32149__;
  assign new_new_n32151__ = ~new_new_n32146__ & new_new_n32150__;
  assign new_new_n32152__ = ~new_new_n32145__ & ~new_new_n32151__;
  assign new_new_n32153__ = new_new_n31730__ & ~new_new_n32152__;
  assign new_new_n32154__ = ~new_new_n31730__ & new_new_n32152__;
  assign new_new_n32155__ = ~new_new_n30750__ & ~new_new_n30751__;
  assign new_new_n32156__ = ~new_new_n31098__ & ~new_new_n32155__;
  assign new_new_n32157__ = new_new_n31098__ & new_new_n32155__;
  assign new_new_n32158__ = ~new_new_n32156__ & ~new_new_n32157__;
  assign new_new_n32159__ = ~new_new_n32154__ & ~new_new_n32158__;
  assign new_new_n32160__ = ~new_new_n32153__ & ~new_new_n32159__;
  assign new_new_n32161__ = ~new_new_n31715__ & ~new_new_n32160__;
  assign new_new_n32162__ = ~new_new_n31714__ & ~new_new_n32161__;
  assign new_new_n32163__ = ~new_new_n31694__ & ~new_new_n32162__;
  assign new_new_n32164__ = new_new_n31694__ & new_new_n32162__;
  assign new_new_n32165__ = ~new_new_n31111__ & ~new_new_n31112__;
  assign new_new_n32166__ = ~new_new_n31122__ & new_new_n32165__;
  assign new_new_n32167__ = new_new_n31122__ & ~new_new_n32165__;
  assign new_new_n32168__ = ~new_new_n32166__ & ~new_new_n32167__;
  assign new_new_n32169__ = ~new_new_n32164__ & new_new_n32168__;
  assign new_new_n32170__ = ~new_new_n32163__ & ~new_new_n32169__;
  assign new_new_n32171__ = new_new_n13508__ & new_new_n26847__;
  assign new_new_n32172__ = pi01 & ~new_new_n26847__;
  assign new_new_n32173__ = ~new_new_n31703__ & ~new_new_n32172__;
  assign new_new_n32174__ = pi02 & ~new_new_n32173__;
  assign new_new_n32175__ = ~new_new_n32171__ & ~new_new_n32174__;
  assign new_new_n32176__ = ~pi00 & ~new_new_n32175__;
  assign new_new_n32177__ = pi02 & ~new_new_n26823__;
  assign new_new_n32178__ = ~new_new_n31661__ & ~new_new_n32177__;
  assign new_new_n32179__ = ~new_new_n29400__ & ~new_new_n32178__;
  assign new_new_n32180__ = pi01 & ~new_new_n26823__;
  assign new_new_n32181__ = ~pi02 & new_new_n26823__;
  assign new_new_n32182__ = ~new_new_n32180__ & ~new_new_n32181__;
  assign new_new_n32183__ = new_new_n29400__ & ~new_new_n32182__;
  assign new_new_n32184__ = pi00 & ~new_new_n32179__;
  assign new_new_n32185__ = ~new_new_n32183__ & new_new_n32184__;
  assign new_new_n32186__ = ~new_new_n32176__ & ~new_new_n32185__;
  assign new_new_n32187__ = ~new_new_n31129__ & ~new_new_n31130__;
  assign new_new_n32188__ = ~new_new_n31141__ & new_new_n32187__;
  assign new_new_n32189__ = new_new_n31141__ & ~new_new_n32187__;
  assign new_new_n32190__ = ~new_new_n32188__ & ~new_new_n32189__;
  assign new_new_n32191__ = new_new_n32186__ & new_new_n32190__;
  assign new_new_n32192__ = ~new_new_n32170__ & ~new_new_n32191__;
  assign new_new_n32193__ = ~new_new_n32186__ & ~new_new_n32190__;
  assign new_new_n32194__ = ~new_new_n32192__ & ~new_new_n32193__;
  assign new_new_n32195__ = ~new_new_n31676__ & ~new_new_n32194__;
  assign new_new_n32196__ = new_new_n31676__ & new_new_n32194__;
  assign new_new_n32197__ = ~pi01 & new_new_n26847__;
  assign new_new_n32198__ = pi02 & ~new_new_n32197__;
  assign new_new_n32199__ = ~new_new_n32180__ & new_new_n32198__;
  assign new_new_n32200__ = new_new_n13508__ & ~new_new_n26823__;
  assign new_new_n32201__ = ~new_new_n32199__ & ~new_new_n32200__;
  assign new_new_n32202__ = ~pi00 & ~new_new_n32201__;
  assign new_new_n32203__ = ~new_new_n31636__ & ~new_new_n31660__;
  assign new_new_n32204__ = ~new_new_n27191__ & new_new_n32203__;
  assign new_new_n32205__ = pi02 & ~new_new_n27221__;
  assign new_new_n32206__ = ~new_new_n31659__ & ~new_new_n32205__;
  assign new_new_n32207__ = new_new_n27191__ & ~new_new_n32206__;
  assign new_new_n32208__ = pi00 & ~new_new_n32204__;
  assign new_new_n32209__ = ~new_new_n32207__ & new_new_n32208__;
  assign new_new_n32210__ = ~new_new_n32202__ & ~new_new_n32209__;
  assign new_new_n32211__ = ~new_new_n32196__ & ~new_new_n32210__;
  assign new_new_n32212__ = ~new_new_n32195__ & ~new_new_n32211__;
  assign new_new_n32213__ = ~new_new_n31672__ & ~new_new_n32212__;
  assign new_new_n32214__ = ~new_new_n31671__ & ~new_new_n32213__;
  assign new_new_n32215__ = ~new_new_n31651__ & ~new_new_n32214__;
  assign new_new_n32216__ = new_new_n31651__ & new_new_n32214__;
  assign new_new_n32217__ = ~new_new_n31180__ & ~new_new_n31181__;
  assign new_new_n32218__ = new_new_n31192__ & ~new_new_n32217__;
  assign new_new_n32219__ = ~new_new_n31192__ & new_new_n32217__;
  assign new_new_n32220__ = ~new_new_n32218__ & ~new_new_n32219__;
  assign new_new_n32221__ = ~new_new_n32216__ & ~new_new_n32220__;
  assign new_new_n32222__ = ~new_new_n32215__ & ~new_new_n32221__;
  assign new_new_n32223__ = ~new_new_n31634__ & ~new_new_n32222__;
  assign new_new_n32224__ = ~new_new_n31633__ & ~new_new_n32223__;
  assign new_new_n32225__ = ~new_new_n31610__ & ~new_new_n32224__;
  assign new_new_n32226__ = new_new_n31610__ & new_new_n32224__;
  assign new_new_n32227__ = ~new_new_n31223__ & ~new_new_n31224__;
  assign new_new_n32228__ = new_new_n31236__ & ~new_new_n32227__;
  assign new_new_n32229__ = ~new_new_n31236__ & new_new_n32227__;
  assign new_new_n32230__ = ~new_new_n32228__ & ~new_new_n32229__;
  assign new_new_n32231__ = ~new_new_n32226__ & ~new_new_n32230__;
  assign new_new_n32232__ = ~new_new_n32225__ & ~new_new_n32231__;
  assign new_new_n32233__ = ~new_new_n31592__ & ~new_new_n32232__;
  assign new_new_n32234__ = new_new_n31592__ & new_new_n32232__;
  assign new_new_n32235__ = new_new_n29826__ & ~new_new_n30699__;
  assign new_new_n32236__ = ~new_new_n29826__ & new_new_n30699__;
  assign new_new_n32237__ = ~new_new_n32235__ & ~new_new_n32236__;
  assign new_new_n32238__ = new_new_n29889__ & ~new_new_n30337__;
  assign new_new_n32239__ = ~new_new_n29889__ & new_new_n30337__;
  assign new_new_n32240__ = ~new_new_n32238__ & ~new_new_n32239__;
  assign new_new_n32241__ = new_new_n31238__ & ~new_new_n32240__;
  assign new_new_n32242__ = ~new_new_n31238__ & new_new_n32240__;
  assign new_new_n32243__ = ~new_new_n32241__ & ~new_new_n32242__;
  assign new_new_n32244__ = ~new_new_n32237__ & new_new_n32243__;
  assign new_new_n32245__ = new_new_n32237__ & ~new_new_n32243__;
  assign new_new_n32246__ = ~new_new_n32244__ & ~new_new_n32245__;
  assign new_new_n32247__ = new_new_n30340__ & new_new_n32246__;
  assign new_new_n32248__ = ~new_new_n30340__ & ~new_new_n32246__;
  assign new_new_n32249__ = ~new_new_n32247__ & ~new_new_n32248__;
  assign new_new_n32250__ = ~new_new_n32234__ & ~new_new_n32249__;
  assign new_new_n32251__ = pi01 & new_new_n31588__;
  assign new_new_n32252__ = new_new_n12798__ & ~new_new_n26774__;
  assign new_new_n32253__ = ~new_new_n32251__ & ~new_new_n32252__;
  assign new_new_n32254__ = ~pi00 & ~new_new_n32253__;
  assign new_new_n32255__ = pi01 & new_new_n27348__;
  assign new_new_n32256__ = pi02 & ~new_new_n27348__;
  assign new_new_n32257__ = new_new_n26722__ & ~new_new_n32255__;
  assign new_new_n32258__ = ~new_new_n32256__ & new_new_n32257__;
  assign new_new_n32259__ = ~pi01 & ~new_new_n27348__;
  assign new_new_n32260__ = ~pi02 & new_new_n27348__;
  assign new_new_n32261__ = ~new_new_n26722__ & ~new_new_n32259__;
  assign new_new_n32262__ = ~new_new_n32260__ & new_new_n32261__;
  assign new_new_n32263__ = ~new_new_n32258__ & ~new_new_n32262__;
  assign new_new_n32264__ = pi00 & ~new_new_n32263__;
  assign new_new_n32265__ = ~new_new_n32254__ & ~new_new_n32264__;
  assign new_new_n32266__ = ~new_new_n31247__ & ~new_new_n31248__;
  assign new_new_n32267__ = new_new_n31250__ & ~new_new_n32266__;
  assign new_new_n32268__ = ~new_new_n31250__ & new_new_n32266__;
  assign new_new_n32269__ = ~new_new_n32267__ & ~new_new_n32268__;
  assign new_new_n32270__ = ~new_new_n32265__ & ~new_new_n32269__;
  assign new_new_n32271__ = ~new_new_n32233__ & ~new_new_n32250__;
  assign new_new_n32272__ = ~new_new_n32270__ & new_new_n32271__;
  assign new_new_n32273__ = new_new_n32265__ & new_new_n32269__;
  assign new_new_n32274__ = ~new_new_n32272__ & ~new_new_n32273__;
  assign new_new_n32275__ = ~new_new_n31571__ & ~new_new_n32274__;
  assign new_new_n32276__ = ~new_new_n31570__ & ~new_new_n32275__;
  assign new_new_n32277__ = ~new_new_n31550__ & ~new_new_n32276__;
  assign new_new_n32278__ = ~new_new_n31549__ & ~new_new_n32277__;
  assign new_new_n32279__ = new_new_n31527__ & new_new_n32278__;
  assign new_new_n32280__ = ~new_new_n30615__ & ~new_new_n30616__;
  assign new_new_n32281__ = new_new_n31267__ & new_new_n32280__;
  assign new_new_n32282__ = new_new_n31285__ & ~new_new_n32280__;
  assign new_new_n32283__ = ~new_new_n32281__ & ~new_new_n32282__;
  assign new_new_n32284__ = new_new_n32279__ & ~new_new_n32283__;
  assign new_new_n32285__ = ~new_new_n31527__ & ~new_new_n32278__;
  assign new_new_n32286__ = new_new_n31268__ & ~new_new_n31283__;
  assign new_new_n32287__ = ~new_new_n32280__ & ~new_new_n32286__;
  assign new_new_n32288__ = new_new_n31267__ & new_new_n31283__;
  assign new_new_n32289__ = ~new_new_n31285__ & ~new_new_n32288__;
  assign new_new_n32290__ = new_new_n32280__ & ~new_new_n32289__;
  assign new_new_n32291__ = ~new_new_n32285__ & ~new_new_n32287__;
  assign new_new_n32292__ = ~new_new_n32290__ & new_new_n32291__;
  assign new_new_n32293__ = ~new_new_n32284__ & ~new_new_n32292__;
  assign new_new_n32294__ = ~new_new_n31505__ & ~new_new_n32293__;
  assign new_new_n32295__ = new_new_n31505__ & new_new_n32293__;
  assign new_new_n32296__ = ~new_new_n32294__ & ~new_new_n32295__;
  assign new_new_n32297__ = new_new_n26698__ & ~new_new_n27273__;
  assign new_new_n32298__ = ~new_new_n26698__ & new_new_n27273__;
  assign new_new_n32299__ = ~new_new_n32297__ & ~new_new_n32298__;
  assign new_new_n32300__ = new_new_n31508__ & ~new_new_n32299__;
  assign new_new_n32301__ = ~new_new_n25294__ & new_new_n32300__;
  assign new_new_n32302__ = ~new_new_n26674__ & ~new_new_n32301__;
  assign new_new_n32303__ = new_new_n26674__ & new_new_n32301__;
  assign new_new_n32304__ = ~new_new_n32302__ & ~new_new_n32303__;
  assign new_new_n32305__ = pi00 & ~new_new_n32304__;
  assign new_new_n32306__ = ~pi01 & new_new_n31529__;
  assign new_new_n32307__ = ~new_new_n31522__ & ~new_new_n32306__;
  assign new_new_n32308__ = ~pi00 & ~new_new_n32307__;
  assign new_new_n32309__ = ~new_new_n32305__ & ~new_new_n32308__;
  assign new_new_n32310__ = pi02 & ~new_new_n32309__;
  assign new_new_n32311__ = ~pi02 & new_new_n32309__;
  assign new_new_n32312__ = ~new_new_n32310__ & ~new_new_n32311__;
  assign new_new_n32313__ = ~new_new_n32296__ & new_new_n32312__;
  assign new_new_n32314__ = ~new_new_n31267__ & ~new_new_n32280__;
  assign new_new_n32315__ = ~new_new_n32286__ & ~new_new_n32289__;
  assign new_new_n32316__ = ~new_new_n32279__ & new_new_n32315__;
  assign new_new_n32317__ = ~new_new_n32281__ & ~new_new_n32314__;
  assign new_new_n32318__ = new_new_n32316__ & new_new_n32317__;
  assign new_new_n32319__ = ~new_new_n31268__ & new_new_n32280__;
  assign new_new_n32320__ = ~new_new_n32282__ & new_new_n32285__;
  assign new_new_n32321__ = ~new_new_n32319__ & new_new_n32320__;
  assign new_new_n32322__ = ~new_new_n32318__ & ~new_new_n32321__;
  assign new_new_n32323__ = ~new_new_n31505__ & new_new_n32322__;
  assign new_new_n32324__ = new_new_n31505__ & ~new_new_n32322__;
  assign new_new_n32325__ = ~new_new_n32312__ & ~new_new_n32323__;
  assign new_new_n32326__ = ~new_new_n32324__ & new_new_n32325__;
  assign po00 = ~new_new_n32313__ & ~new_new_n32326__;
  assign new_new_n32328__ = new_new_n32293__ & new_new_n32322__;
  assign new_new_n32329__ = new_new_n26667__ & new_new_n26674__;
  assign new_new_n32330__ = ~new_new_n26667__ & ~new_new_n27284__;
  assign new_new_n32331__ = new_new_n26667__ & new_new_n27284__;
  assign new_new_n32332__ = ~new_new_n32330__ & ~new_new_n32331__;
  assign new_new_n32333__ = ~new_new_n26698__ & ~new_new_n32329__;
  assign new_new_n32334__ = ~new_new_n32332__ & new_new_n32333__;
  assign new_new_n32335__ = new_new_n26698__ & ~new_new_n27288__;
  assign new_new_n32336__ = new_new_n32332__ & new_new_n32335__;
  assign new_new_n32337__ = ~new_new_n32334__ & ~new_new_n32336__;
  assign new_new_n32338__ = new_new_n26667__ & ~new_new_n32337__;
  assign new_new_n32339__ = ~new_new_n26667__ & new_new_n32300__;
  assign new_new_n32340__ = new_new_n32337__ & ~new_new_n32339__;
  assign new_new_n32341__ = ~new_new_n26667__ & new_new_n32340__;
  assign new_new_n32342__ = ~new_new_n26667__ & ~new_new_n26674__;
  assign new_new_n32343__ = ~new_new_n32329__ & ~new_new_n32342__;
  assign new_new_n32344__ = ~new_new_n32338__ & new_new_n32343__;
  assign new_new_n32345__ = ~new_new_n32341__ & new_new_n32344__;
  assign new_new_n32346__ = pi02 & ~new_new_n32345__;
  assign new_new_n32347__ = pi01 & new_new_n32345__;
  assign new_new_n32348__ = ~new_new_n32346__ & ~new_new_n32347__;
  assign new_new_n32349__ = ~new_new_n15968__ & ~new_new_n16041__;
  assign new_new_n32350__ = ~new_new_n15969__ & ~new_new_n32349__;
  assign new_new_n32351__ = ~pi30 & new_new_n16056__;
  assign new_new_n32352__ = ~new_new_n15853__ & ~new_new_n32351__;
  assign new_new_n32353__ = ~new_new_n16051__ & new_new_n32352__;
  assign new_new_n32354__ = ~new_new_n4876__ & ~new_new_n15971__;
  assign new_new_n32355__ = ~new_new_n32353__ & new_new_n32354__;
  assign new_new_n32356__ = ~new_new_n70__ & ~new_new_n32355__;
  assign new_new_n32357__ = new_new_n70__ & new_new_n32355__;
  assign new_new_n32358__ = ~new_new_n32356__ & ~new_new_n32357__;
  assign new_new_n32359__ = new_new_n16044__ & new_new_n26585__;
  assign new_new_n32360__ = ~new_new_n16044__ & ~new_new_n26585__;
  assign new_new_n32361__ = ~new_new_n26639__ & ~new_new_n32360__;
  assign new_new_n32362__ = new_new_n16044__ & ~new_new_n26641__;
  assign new_new_n32363__ = ~new_new_n26644__ & ~new_new_n32362__;
  assign new_new_n32364__ = ~new_new_n26642__ & ~new_new_n32363__;
  assign new_new_n32365__ = ~new_new_n32359__ & ~new_new_n32364__;
  assign new_new_n32366__ = ~new_new_n32361__ & new_new_n32365__;
  assign new_new_n32367__ = new_new_n465__ & new_new_n3764__;
  assign new_new_n32368__ = new_new_n16035__ & new_new_n16038__;
  assign new_new_n32369__ = new_new_n16034__ & ~new_new_n16038__;
  assign new_new_n32370__ = ~new_new_n32368__ & ~new_new_n32369__;
  assign new_new_n32371__ = new_new_n32367__ & ~new_new_n32370__;
  assign new_new_n32372__ = ~new_new_n32367__ & new_new_n32370__;
  assign new_new_n32373__ = ~new_new_n32371__ & ~new_new_n32372__;
  assign new_new_n32374__ = ~new_new_n32366__ & ~new_new_n32373__;
  assign new_new_n32375__ = new_new_n32366__ & new_new_n32373__;
  assign new_new_n32376__ = ~new_new_n32374__ & ~new_new_n32375__;
  assign new_new_n32377__ = new_new_n32358__ & ~new_new_n32376__;
  assign new_new_n32378__ = ~new_new_n32358__ & new_new_n32376__;
  assign new_new_n32379__ = ~new_new_n32377__ & ~new_new_n32378__;
  assign new_new_n32380__ = new_new_n32350__ & new_new_n32379__;
  assign new_new_n32381__ = ~new_new_n32350__ & ~new_new_n32379__;
  assign new_new_n32382__ = ~new_new_n32380__ & ~new_new_n32381__;
  assign new_new_n32383__ = new_new_n32348__ & ~new_new_n32382__;
  assign new_new_n32384__ = ~new_new_n32348__ & new_new_n32382__;
  assign new_new_n32385__ = pi00 & ~new_new_n32383__;
  assign new_new_n32386__ = ~new_new_n32384__ & new_new_n32385__;
  assign new_new_n32387__ = pi01 & ~new_new_n26667__;
  assign new_new_n32388__ = ~pi01 & ~new_new_n26674__;
  assign new_new_n32389__ = pi02 & ~new_new_n32388__;
  assign new_new_n32390__ = ~new_new_n32387__ & ~new_new_n32389__;
  assign new_new_n32391__ = pi02 & new_new_n32387__;
  assign new_new_n32392__ = ~pi00 & ~new_new_n32390__;
  assign new_new_n32393__ = ~new_new_n32391__ & new_new_n32392__;
  assign new_new_n32394__ = ~new_new_n32386__ & ~new_new_n32393__;
  assign new_new_n32395__ = new_new_n13111__ & ~new_new_n27242__;
  assign new_new_n32396__ = new_new_n11469__ & new_new_n31511__;
  assign new_new_n32397__ = ~new_new_n32395__ & ~new_new_n32396__;
  assign new_new_n32398__ = new_new_n11478__ & ~new_new_n32397__;
  assign new_new_n32399__ = new_new_n11475__ & new_new_n27250__;
  assign new_new_n32400__ = ~new_new_n32398__ & ~new_new_n32399__;
  assign new_new_n32401__ = pi05 & ~new_new_n32400__;
  assign new_new_n32402__ = new_new_n12873__ & new_new_n26698__;
  assign new_new_n32403__ = new_new_n11469__ & new_new_n26698__;
  assign new_new_n32404__ = ~pi05 & ~new_new_n32403__;
  assign new_new_n32405__ = ~new_new_n32402__ & ~new_new_n32404__;
  assign new_new_n32406__ = new_new_n32400__ & ~new_new_n32405__;
  assign new_new_n32407__ = ~new_new_n32401__ & ~new_new_n32406__;
  assign new_new_n32408__ = new_new_n10698__ & new_new_n26722__;
  assign new_new_n32409__ = ~new_new_n11409__ & new_new_n26774__;
  assign new_new_n32410__ = new_new_n10702__ & new_new_n26729__;
  assign new_new_n32411__ = ~new_new_n32409__ & ~new_new_n32410__;
  assign new_new_n32412__ = ~new_new_n32408__ & new_new_n32411__;
  assign new_new_n32413__ = new_new_n10694__ & ~new_new_n27348__;
  assign new_new_n32414__ = ~pi08 & ~new_new_n32413__;
  assign new_new_n32415__ = new_new_n12121__ & ~new_new_n27348__;
  assign new_new_n32416__ = ~new_new_n32414__ & ~new_new_n32415__;
  assign new_new_n32417__ = new_new_n32412__ & ~new_new_n32416__;
  assign new_new_n32418__ = pi08 & ~new_new_n32412__;
  assign new_new_n32419__ = ~new_new_n32417__ & ~new_new_n32418__;
  assign new_new_n32420__ = new_new_n6968__ & ~new_new_n26888__;
  assign new_new_n32421__ = new_new_n6964__ & new_new_n26922__;
  assign new_new_n32422__ = new_new_n7935__ & ~new_new_n26854__;
  assign new_new_n32423__ = ~new_new_n32420__ & ~new_new_n32421__;
  assign new_new_n32424__ = ~new_new_n32422__ & new_new_n32423__;
  assign new_new_n32425__ = new_new_n6958__ & ~new_new_n27430__;
  assign new_new_n32426__ = ~pi17 & ~new_new_n32425__;
  assign new_new_n32427__ = new_new_n8160__ & ~new_new_n27430__;
  assign new_new_n32428__ = ~new_new_n32426__ & ~new_new_n32427__;
  assign new_new_n32429__ = new_new_n32424__ & ~new_new_n32428__;
  assign new_new_n32430__ = pi17 & ~new_new_n32424__;
  assign new_new_n32431__ = ~new_new_n32429__ & ~new_new_n32430__;
  assign new_new_n32432__ = pi23 & ~new_new_n31402__;
  assign new_new_n32433__ = new_new_n31410__ & new_new_n32432__;
  assign new_new_n32434__ = ~new_new_n31324__ & new_new_n31410__;
  assign new_new_n32435__ = ~pi23 & ~new_new_n31410__;
  assign new_new_n32436__ = ~new_new_n32434__ & ~new_new_n32435__;
  assign new_new_n32437__ = new_new_n31402__ & ~new_new_n32436__;
  assign new_new_n32438__ = ~new_new_n32433__ & ~new_new_n32437__;
  assign new_new_n32439__ = new_new_n3311__ & new_new_n26971__;
  assign new_new_n32440__ = new_new_n873__ & ~new_new_n26978__;
  assign new_new_n32441__ = ~new_new_n333__ & ~new_new_n27003__;
  assign new_new_n32442__ = ~new_new_n4900__ & new_new_n28277__;
  assign new_new_n32443__ = ~new_new_n32440__ & ~new_new_n32441__;
  assign new_new_n32444__ = ~new_new_n32439__ & new_new_n32443__;
  assign new_new_n32445__ = ~new_new_n32442__ & new_new_n32444__;
  assign new_new_n32446__ = ~pi26 & ~new_new_n32445__;
  assign new_new_n32447__ = pi26 & new_new_n32445__;
  assign new_new_n32448__ = ~new_new_n32446__ & ~new_new_n32447__;
  assign new_new_n32449__ = new_new_n31334__ & new_new_n31390__;
  assign new_new_n32450__ = ~new_new_n31390__ & new_new_n31398__;
  assign new_new_n32451__ = ~new_new_n32449__ & ~new_new_n32450__;
  assign new_new_n32452__ = new_new_n32448__ & ~new_new_n32451__;
  assign new_new_n32453__ = ~new_new_n32448__ & new_new_n32451__;
  assign new_new_n32454__ = ~new_new_n32452__ & ~new_new_n32453__;
  assign new_new_n32455__ = new_new_n4815__ & ~new_new_n27029__;
  assign new_new_n32456__ = new_new_n4212__ & ~new_new_n27021__;
  assign new_new_n32457__ = ~new_new_n4818__ & new_new_n27111__;
  assign new_new_n32458__ = new_new_n4813__ & new_new_n27764__;
  assign new_new_n32459__ = ~new_new_n32456__ & ~new_new_n32457__;
  assign new_new_n32460__ = ~new_new_n32455__ & new_new_n32459__;
  assign new_new_n32461__ = ~new_new_n32458__ & new_new_n32460__;
  assign new_new_n32462__ = pi29 & ~new_new_n32461__;
  assign new_new_n32463__ = ~pi29 & new_new_n32461__;
  assign new_new_n32464__ = ~new_new_n32462__ & ~new_new_n32463__;
  assign new_new_n32465__ = ~new_new_n27054__ & ~new_new_n27097__;
  assign new_new_n32466__ = ~new_new_n15853__ & ~new_new_n27100__;
  assign new_new_n32467__ = ~new_new_n32465__ & new_new_n32466__;
  assign new_new_n32468__ = ~new_new_n27055__ & ~new_new_n32467__;
  assign new_new_n32469__ = ~new_new_n27033__ & ~new_new_n32468__;
  assign new_new_n32470__ = new_new_n27033__ & new_new_n27098__;
  assign new_new_n32471__ = ~new_new_n71__ & ~new_new_n32470__;
  assign new_new_n32472__ = ~new_new_n161__ & ~new_new_n27054__;
  assign new_new_n32473__ = ~new_new_n32471__ & new_new_n32472__;
  assign new_new_n32474__ = new_new_n27097__ & new_new_n27683__;
  assign new_new_n32475__ = ~new_new_n161__ & ~new_new_n32474__;
  assign new_new_n32476__ = ~new_new_n71__ & new_new_n27041__;
  assign new_new_n32477__ = ~new_new_n32475__ & new_new_n32476__;
  assign new_new_n32478__ = ~new_new_n32469__ & ~new_new_n32473__;
  assign new_new_n32479__ = ~new_new_n32477__ & new_new_n32478__;
  assign new_new_n32480__ = pi31 & ~new_new_n32479__;
  assign new_new_n32481__ = new_new_n161__ & ~new_new_n27054__;
  assign new_new_n32482__ = new_new_n765__ & ~new_new_n27033__;
  assign new_new_n32483__ = ~new_new_n32481__ & ~new_new_n32482__;
  assign new_new_n32484__ = ~pi31 & ~new_new_n32483__;
  assign new_new_n32485__ = ~new_new_n32480__ & ~new_new_n32484__;
  assign new_new_n32486__ = ~new_new_n31340__ & ~new_new_n31370__;
  assign new_new_n32487__ = ~new_new_n31371__ & ~new_new_n32486__;
  assign new_new_n32488__ = new_new_n32485__ & new_new_n32487__;
  assign new_new_n32489__ = ~new_new_n32485__ & ~new_new_n32487__;
  assign new_new_n32490__ = ~new_new_n32488__ & ~new_new_n32489__;
  assign new_new_n32491__ = ~new_new_n921__ & new_new_n2908__;
  assign new_new_n32492__ = new_new_n91__ & ~new_new_n355__;
  assign new_new_n32493__ = ~new_new_n88__ & ~new_new_n130__;
  assign new_new_n32494__ = ~new_new_n247__ & ~new_new_n309__;
  assign new_new_n32495__ = ~new_new_n385__ & ~new_new_n597__;
  assign new_new_n32496__ = ~new_new_n1081__ & ~new_new_n2170__;
  assign new_new_n32497__ = new_new_n32495__ & new_new_n32496__;
  assign new_new_n32498__ = new_new_n32493__ & new_new_n32494__;
  assign new_new_n32499__ = ~new_new_n322__ & new_new_n1522__;
  assign new_new_n32500__ = new_new_n2158__ & new_new_n2590__;
  assign new_new_n32501__ = new_new_n4459__ & ~new_new_n32492__;
  assign new_new_n32502__ = new_new_n32500__ & new_new_n32501__;
  assign new_new_n32503__ = new_new_n32498__ & new_new_n32499__;
  assign new_new_n32504__ = new_new_n17256__ & new_new_n32497__;
  assign new_new_n32505__ = new_new_n32503__ & new_new_n32504__;
  assign new_new_n32506__ = new_new_n2028__ & new_new_n32502__;
  assign new_new_n32507__ = new_new_n32505__ & new_new_n32506__;
  assign new_new_n32508__ = new_new_n669__ & new_new_n7492__;
  assign new_new_n32509__ = new_new_n7656__ & new_new_n32508__;
  assign new_new_n32510__ = new_new_n32507__ & new_new_n32509__;
  assign new_new_n32511__ = new_new_n17536__ & new_new_n32510__;
  assign new_new_n32512__ = new_new_n983__ & new_new_n32491__;
  assign new_new_n32513__ = new_new_n32511__ & new_new_n32512__;
  assign new_new_n32514__ = ~new_new_n32490__ & new_new_n32513__;
  assign new_new_n32515__ = new_new_n32490__ & ~new_new_n32513__;
  assign new_new_n32516__ = ~new_new_n32514__ & ~new_new_n32515__;
  assign new_new_n32517__ = new_new_n31336__ & new_new_n31384__;
  assign new_new_n32518__ = ~new_new_n31336__ & ~new_new_n31384__;
  assign new_new_n32519__ = ~new_new_n31340__ & ~new_new_n31372__;
  assign new_new_n32520__ = new_new_n31340__ & new_new_n31372__;
  assign new_new_n32521__ = ~new_new_n32519__ & ~new_new_n32520__;
  assign new_new_n32522__ = ~new_new_n32518__ & ~new_new_n32521__;
  assign new_new_n32523__ = ~new_new_n32517__ & ~new_new_n32522__;
  assign new_new_n32524__ = ~new_new_n32516__ & new_new_n32523__;
  assign new_new_n32525__ = new_new_n32516__ & ~new_new_n32523__;
  assign new_new_n32526__ = ~new_new_n32524__ & ~new_new_n32525__;
  assign new_new_n32527__ = ~new_new_n32464__ & ~new_new_n32526__;
  assign new_new_n32528__ = new_new_n32464__ & new_new_n32526__;
  assign new_new_n32529__ = ~new_new_n32527__ & ~new_new_n32528__;
  assign new_new_n32530__ = new_new_n32454__ & ~new_new_n32529__;
  assign new_new_n32531__ = ~new_new_n32454__ & new_new_n32529__;
  assign new_new_n32532__ = ~new_new_n32530__ & ~new_new_n32531__;
  assign new_new_n32533__ = new_new_n5183__ & new_new_n27152__;
  assign new_new_n32534__ = new_new_n5191__ & ~new_new_n26937__;
  assign new_new_n32535__ = new_new_n5213__ & ~new_new_n26941__;
  assign new_new_n32536__ = new_new_n5215__ & ~new_new_n27502__;
  assign new_new_n32537__ = ~new_new_n32534__ & ~new_new_n32535__;
  assign new_new_n32538__ = ~new_new_n32533__ & new_new_n32537__;
  assign new_new_n32539__ = ~new_new_n32536__ & new_new_n32538__;
  assign new_new_n32540__ = new_new_n32532__ & new_new_n32539__;
  assign new_new_n32541__ = ~new_new_n32532__ & ~new_new_n32539__;
  assign new_new_n32542__ = ~new_new_n32540__ & ~new_new_n32541__;
  assign new_new_n32543__ = ~new_new_n32438__ & new_new_n32542__;
  assign new_new_n32544__ = new_new_n31402__ & new_new_n32434__;
  assign new_new_n32545__ = ~new_new_n32432__ & ~new_new_n32542__;
  assign new_new_n32546__ = ~new_new_n32435__ & new_new_n32545__;
  assign new_new_n32547__ = ~new_new_n32544__ & new_new_n32546__;
  assign new_new_n32548__ = ~new_new_n32543__ & ~new_new_n32547__;
  assign new_new_n32549__ = ~new_new_n31420__ & new_new_n31434__;
  assign new_new_n32550__ = ~new_new_n31421__ & ~new_new_n32549__;
  assign new_new_n32551__ = new_new_n6629__ & new_new_n26917__;
  assign new_new_n32552__ = ~new_new_n6625__ & new_new_n26928__;
  assign new_new_n32553__ = new_new_n6634__ & ~new_new_n27168__;
  assign new_new_n32554__ = ~new_new_n32552__ & ~new_new_n32553__;
  assign new_new_n32555__ = ~new_new_n32551__ & new_new_n32554__;
  assign new_new_n32556__ = new_new_n6631__ & ~new_new_n28799__;
  assign new_new_n32557__ = ~pi20 & ~new_new_n32556__;
  assign new_new_n32558__ = new_new_n7015__ & ~new_new_n28799__;
  assign new_new_n32559__ = ~new_new_n32557__ & ~new_new_n32558__;
  assign new_new_n32560__ = new_new_n32555__ & ~new_new_n32559__;
  assign new_new_n32561__ = pi20 & ~new_new_n32555__;
  assign new_new_n32562__ = ~new_new_n32560__ & ~new_new_n32561__;
  assign new_new_n32563__ = new_new_n32550__ & ~new_new_n32562__;
  assign new_new_n32564__ = ~new_new_n32550__ & new_new_n32562__;
  assign new_new_n32565__ = ~new_new_n32563__ & ~new_new_n32564__;
  assign new_new_n32566__ = new_new_n32548__ & ~new_new_n32565__;
  assign new_new_n32567__ = ~new_new_n32548__ & new_new_n32565__;
  assign new_new_n32568__ = ~new_new_n32566__ & ~new_new_n32567__;
  assign new_new_n32569__ = new_new_n31437__ & ~new_new_n31454__;
  assign new_new_n32570__ = ~new_new_n31455__ & ~new_new_n32569__;
  assign new_new_n32571__ = new_new_n32568__ & ~new_new_n32570__;
  assign new_new_n32572__ = ~new_new_n32568__ & new_new_n32570__;
  assign new_new_n32573__ = ~new_new_n32571__ & ~new_new_n32572__;
  assign new_new_n32574__ = new_new_n6985__ & ~new_new_n26823__;
  assign new_new_n32575__ = new_new_n6991__ & new_new_n26847__;
  assign new_new_n32576__ = ~new_new_n32574__ & ~new_new_n32575__;
  assign new_new_n32577__ = new_new_n6994__ & ~new_new_n27221__;
  assign new_new_n32578__ = new_new_n27411__ & new_new_n32577__;
  assign new_new_n32579__ = new_new_n32576__ & ~new_new_n32578__;
  assign new_new_n32580__ = pi14 & ~new_new_n32579__;
  assign new_new_n32581__ = pi13 & new_new_n27221__;
  assign new_new_n32582__ = ~pi13 & ~new_new_n27221__;
  assign new_new_n32583__ = new_new_n6994__ & ~new_new_n32581__;
  assign new_new_n32584__ = ~new_new_n32582__ & new_new_n32583__;
  assign new_new_n32585__ = ~new_new_n27191__ & new_new_n32584__;
  assign new_new_n32586__ = new_new_n6994__ & ~new_new_n27410__;
  assign new_new_n32587__ = ~pi14 & new_new_n32576__;
  assign new_new_n32588__ = ~new_new_n32586__ & new_new_n32587__;
  assign new_new_n32589__ = ~new_new_n32585__ & ~new_new_n32588__;
  assign new_new_n32590__ = ~new_new_n32580__ & new_new_n32589__;
  assign new_new_n32591__ = new_new_n32573__ & ~new_new_n32590__;
  assign new_new_n32592__ = ~new_new_n32573__ & new_new_n32590__;
  assign new_new_n32593__ = ~new_new_n32591__ & ~new_new_n32592__;
  assign new_new_n32594__ = new_new_n32431__ & new_new_n32593__;
  assign new_new_n32595__ = ~new_new_n32431__ & ~new_new_n32593__;
  assign new_new_n32596__ = ~new_new_n32594__ & ~new_new_n32595__;
  assign new_new_n32597__ = ~new_new_n31314__ & ~new_new_n31459__;
  assign new_new_n32598__ = new_new_n31314__ & new_new_n31459__;
  assign new_new_n32599__ = ~new_new_n31474__ & ~new_new_n32598__;
  assign new_new_n32600__ = ~new_new_n32597__ & ~new_new_n32599__;
  assign new_new_n32601__ = ~new_new_n32596__ & new_new_n32600__;
  assign new_new_n32602__ = new_new_n32596__ & ~new_new_n32600__;
  assign new_new_n32603__ = ~new_new_n32601__ & ~new_new_n32602__;
  assign new_new_n32604__ = ~new_new_n31312__ & new_new_n31476__;
  assign new_new_n32605__ = new_new_n31312__ & ~new_new_n31476__;
  assign new_new_n32606__ = ~new_new_n32597__ & ~new_new_n32598__;
  assign new_new_n32607__ = ~new_new_n31474__ & ~new_new_n32606__;
  assign new_new_n32608__ = new_new_n31474__ & new_new_n32606__;
  assign new_new_n32609__ = ~new_new_n32607__ & ~new_new_n32608__;
  assign new_new_n32610__ = ~new_new_n32605__ & ~new_new_n32609__;
  assign new_new_n32611__ = ~new_new_n32604__ & ~new_new_n32610__;
  assign new_new_n32612__ = new_new_n8474__ & ~new_new_n26802__;
  assign new_new_n32613__ = ~new_new_n8479__ & ~new_new_n26741__;
  assign new_new_n32614__ = new_new_n8468__ & ~new_new_n26810__;
  assign new_new_n32615__ = ~new_new_n8468__ & ~new_new_n27395__;
  assign new_new_n32616__ = new_new_n8469__ & ~new_new_n32614__;
  assign new_new_n32617__ = ~new_new_n32615__ & new_new_n32616__;
  assign new_new_n32618__ = ~new_new_n32612__ & ~new_new_n32613__;
  assign new_new_n32619__ = ~new_new_n32617__ & new_new_n32618__;
  assign new_new_n32620__ = new_new_n8474__ & ~new_new_n8479__;
  assign new_new_n32621__ = pi11 & ~new_new_n32620__;
  assign new_new_n32622__ = new_new_n32619__ & ~new_new_n32621__;
  assign new_new_n32623__ = pi11 & ~new_new_n32619__;
  assign new_new_n32624__ = ~new_new_n32622__ & ~new_new_n32623__;
  assign new_new_n32625__ = new_new_n31482__ & ~new_new_n31496__;
  assign new_new_n32626__ = ~new_new_n31482__ & new_new_n31496__;
  assign new_new_n32627__ = new_new_n11378__ & new_new_n30644__;
  assign new_new_n32628__ = new_new_n31295__ & ~new_new_n32627__;
  assign new_new_n32629__ = ~pi08 & ~new_new_n32628__;
  assign new_new_n32630__ = pi08 & new_new_n32628__;
  assign new_new_n32631__ = ~new_new_n32629__ & ~new_new_n32630__;
  assign new_new_n32632__ = ~new_new_n32626__ & ~new_new_n32631__;
  assign new_new_n32633__ = ~new_new_n32625__ & ~new_new_n32632__;
  assign new_new_n32634__ = new_new_n32624__ & ~new_new_n32633__;
  assign new_new_n32635__ = ~new_new_n32624__ & new_new_n32633__;
  assign new_new_n32636__ = ~new_new_n32634__ & ~new_new_n32635__;
  assign new_new_n32637__ = new_new_n32611__ & new_new_n32636__;
  assign new_new_n32638__ = ~new_new_n32611__ & ~new_new_n32636__;
  assign new_new_n32639__ = ~new_new_n32637__ & ~new_new_n32638__;
  assign new_new_n32640__ = new_new_n32603__ & ~new_new_n32639__;
  assign new_new_n32641__ = ~new_new_n32603__ & new_new_n32639__;
  assign new_new_n32642__ = ~new_new_n32640__ & ~new_new_n32641__;
  assign new_new_n32643__ = new_new_n32419__ & new_new_n32642__;
  assign new_new_n32644__ = ~new_new_n32419__ & ~new_new_n32642__;
  assign new_new_n32645__ = ~new_new_n32643__ & ~new_new_n32644__;
  assign new_new_n32646__ = new_new_n32407__ & ~new_new_n32645__;
  assign new_new_n32647__ = ~new_new_n32407__ & new_new_n32645__;
  assign new_new_n32648__ = ~new_new_n32646__ & ~new_new_n32647__;
  assign new_new_n32649__ = new_new_n27317__ & new_new_n31287__;
  assign new_new_n32650__ = ~new_new_n27317__ & ~new_new_n31287__;
  assign new_new_n32651__ = ~new_new_n31499__ & ~new_new_n32650__;
  assign new_new_n32652__ = ~new_new_n32649__ & ~new_new_n32651__;
  assign new_new_n32653__ = new_new_n32648__ & new_new_n32652__;
  assign new_new_n32654__ = ~new_new_n32648__ & ~new_new_n32652__;
  assign new_new_n32655__ = ~new_new_n32653__ & ~new_new_n32654__;
  assign new_new_n32656__ = new_new_n32293__ & ~new_new_n32312__;
  assign new_new_n32657__ = new_new_n32322__ & ~new_new_n32656__;
  assign new_new_n32658__ = ~new_new_n31503__ & new_new_n32657__;
  assign new_new_n32659__ = ~new_new_n31504__ & ~new_new_n32658__;
  assign new_new_n32660__ = new_new_n32655__ & new_new_n32659__;
  assign new_new_n32661__ = ~new_new_n32655__ & ~new_new_n32659__;
  assign new_new_n32662__ = ~new_new_n32660__ & ~new_new_n32661__;
  assign new_new_n32663__ = ~new_new_n32394__ & new_new_n32662__;
  assign new_new_n32664__ = new_new_n32394__ & ~new_new_n32662__;
  assign new_new_n32665__ = ~new_new_n32663__ & ~new_new_n32664__;
  assign new_new_n32666__ = ~new_new_n32328__ & new_new_n32665__;
  assign new_new_n32667__ = new_new_n32295__ & new_new_n32322__;
  assign new_new_n32668__ = ~new_new_n32665__ & new_new_n32667__;
  assign new_new_n32669__ = ~new_new_n32666__ & ~new_new_n32668__;
  assign new_new_n32670__ = ~new_new_n32312__ & ~new_new_n32669__;
  assign new_new_n32671__ = new_new_n32296__ & new_new_n32665__;
  assign new_new_n32672__ = ~new_new_n32294__ & ~new_new_n32324__;
  assign new_new_n32673__ = ~new_new_n32665__ & new_new_n32672__;
  assign new_new_n32674__ = new_new_n32312__ & ~new_new_n32666__;
  assign new_new_n32675__ = ~new_new_n32673__ & new_new_n32674__;
  assign new_new_n32676__ = ~new_new_n32670__ & ~new_new_n32671__;
  assign po01 = new_new_n32675__ | ~new_new_n32676__;
  assign new_new_n32678__ = ~pi31 & new_new_n71__;
  assign new_new_n32679__ = ~new_new_n66__ & ~new_new_n32678__;
  assign new_new_n32680__ = ~new_new_n69__ & ~new_new_n32679__;
  assign new_new_n32681__ = ~pi30 & ~pi31;
  assign new_new_n32682__ = new_new_n69__ & ~new_new_n32681__;
  assign new_new_n32683__ = ~new_new_n32680__ & ~new_new_n32682__;
  assign new_new_n32684__ = ~new_new_n421__ & new_new_n16035__;
  assign new_new_n32685__ = new_new_n421__ & ~new_new_n16035__;
  assign new_new_n32686__ = new_new_n16038__ & new_new_n32685__;
  assign new_new_n32687__ = ~new_new_n16033__ & ~new_new_n32367__;
  assign new_new_n32688__ = ~new_new_n16038__ & ~new_new_n32687__;
  assign new_new_n32689__ = ~new_new_n32684__ & ~new_new_n32688__;
  assign new_new_n32690__ = ~new_new_n32686__ & new_new_n32689__;
  assign new_new_n32691__ = new_new_n32683__ & ~new_new_n32690__;
  assign new_new_n32692__ = ~new_new_n16031__ & new_new_n32683__;
  assign new_new_n32693__ = ~new_new_n32369__ & ~new_new_n32683__;
  assign new_new_n32694__ = ~new_new_n32367__ & ~new_new_n32692__;
  assign new_new_n32695__ = ~new_new_n32693__ & new_new_n32694__;
  assign new_new_n32696__ = new_new_n16038__ & ~new_new_n32683__;
  assign new_new_n32697__ = new_new_n32367__ & new_new_n32696__;
  assign new_new_n32698__ = ~new_new_n32684__ & new_new_n32697__;
  assign new_new_n32699__ = ~new_new_n32685__ & new_new_n32698__;
  assign new_new_n32700__ = ~new_new_n32695__ & ~new_new_n32699__;
  assign new_new_n32701__ = ~new_new_n32691__ & new_new_n32700__;
  assign new_new_n32702__ = new_new_n32350__ & new_new_n32373__;
  assign new_new_n32703__ = ~new_new_n32357__ & ~new_new_n32702__;
  assign new_new_n32704__ = ~new_new_n32350__ & ~new_new_n32373__;
  assign new_new_n32705__ = new_new_n32366__ & ~new_new_n32704__;
  assign new_new_n32706__ = ~new_new_n32703__ & new_new_n32705__;
  assign new_new_n32707__ = new_new_n70__ & new_new_n32702__;
  assign new_new_n32708__ = new_new_n32355__ & new_new_n32707__;
  assign new_new_n32709__ = ~new_new_n32350__ & ~new_new_n32357__;
  assign new_new_n32710__ = new_new_n32374__ & new_new_n32709__;
  assign new_new_n32711__ = ~new_new_n32356__ & ~new_new_n32708__;
  assign new_new_n32712__ = ~new_new_n32706__ & new_new_n32711__;
  assign new_new_n32713__ = ~new_new_n32710__ & new_new_n32712__;
  assign new_new_n32714__ = ~new_new_n32701__ & ~new_new_n32713__;
  assign new_new_n32715__ = ~new_new_n70__ & ~new_new_n32702__;
  assign new_new_n32716__ = new_new_n32355__ & ~new_new_n32715__;
  assign new_new_n32717__ = new_new_n32705__ & new_new_n32716__;
  assign new_new_n32718__ = new_new_n32356__ & new_new_n32704__;
  assign new_new_n32719__ = ~new_new_n32350__ & ~new_new_n32355__;
  assign new_new_n32720__ = new_new_n32350__ & new_new_n32355__;
  assign new_new_n32721__ = ~new_new_n70__ & ~new_new_n32373__;
  assign new_new_n32722__ = ~new_new_n32720__ & new_new_n32721__;
  assign new_new_n32723__ = ~new_new_n32707__ & ~new_new_n32719__;
  assign new_new_n32724__ = ~new_new_n32722__ & new_new_n32723__;
  assign new_new_n32725__ = ~new_new_n32366__ & ~new_new_n32724__;
  assign new_new_n32726__ = new_new_n32701__ & ~new_new_n32718__;
  assign new_new_n32727__ = ~new_new_n32725__ & new_new_n32726__;
  assign new_new_n32728__ = ~new_new_n32717__ & new_new_n32727__;
  assign new_new_n32729__ = ~new_new_n32714__ & ~new_new_n32728__;
  assign new_new_n32730__ = new_new_n32382__ & ~new_new_n32729__;
  assign new_new_n32731__ = ~new_new_n27284__ & new_new_n32730__;
  assign new_new_n32732__ = ~new_new_n32382__ & new_new_n32729__;
  assign new_new_n32733__ = ~new_new_n26667__ & new_new_n32732__;
  assign new_new_n32734__ = ~new_new_n32731__ & ~new_new_n32733__;
  assign new_new_n32735__ = ~new_new_n26674__ & ~new_new_n32734__;
  assign new_new_n32736__ = ~new_new_n26667__ & new_new_n32382__;
  assign new_new_n32737__ = new_new_n26667__ & ~new_new_n32382__;
  assign new_new_n32738__ = ~new_new_n32736__ & ~new_new_n32737__;
  assign new_new_n32739__ = ~new_new_n32729__ & ~new_new_n32738__;
  assign new_new_n32740__ = ~new_new_n32382__ & ~new_new_n32729__;
  assign new_new_n32741__ = new_new_n27284__ & new_new_n32740__;
  assign new_new_n32742__ = new_new_n26667__ & new_new_n32382__;
  assign new_new_n32743__ = new_new_n32729__ & new_new_n32742__;
  assign new_new_n32744__ = ~new_new_n32741__ & ~new_new_n32743__;
  assign new_new_n32745__ = new_new_n26674__ & ~new_new_n32744__;
  assign new_new_n32746__ = new_new_n27284__ & new_new_n32743__;
  assign new_new_n32747__ = new_new_n26674__ & ~new_new_n32382__;
  assign new_new_n32748__ = ~new_new_n32729__ & new_new_n32747__;
  assign new_new_n32749__ = ~new_new_n32746__ & ~new_new_n32748__;
  assign new_new_n32750__ = ~new_new_n26698__ & ~new_new_n32749__;
  assign new_new_n32751__ = ~new_new_n26674__ & new_new_n32730__;
  assign new_new_n32752__ = new_new_n32330__ & new_new_n32732__;
  assign new_new_n32753__ = ~new_new_n32751__ & ~new_new_n32752__;
  assign new_new_n32754__ = new_new_n26698__ & ~new_new_n32753__;
  assign new_new_n32755__ = ~new_new_n32735__ & ~new_new_n32739__;
  assign new_new_n32756__ = ~new_new_n32745__ & ~new_new_n32750__;
  assign new_new_n32757__ = new_new_n32755__ & new_new_n32756__;
  assign new_new_n32758__ = ~new_new_n32754__ & new_new_n32757__;
  assign new_new_n32759__ = pi02 & ~new_new_n32729__;
  assign new_new_n32760__ = ~pi01 & new_new_n32729__;
  assign new_new_n32761__ = ~new_new_n32759__ & ~new_new_n32760__;
  assign new_new_n32762__ = ~new_new_n32758__ & ~new_new_n32761__;
  assign new_new_n32763__ = ~pi01 & ~new_new_n32729__;
  assign new_new_n32764__ = pi02 & new_new_n32729__;
  assign new_new_n32765__ = ~new_new_n32763__ & ~new_new_n32764__;
  assign new_new_n32766__ = new_new_n32758__ & new_new_n32765__;
  assign new_new_n32767__ = ~new_new_n32762__ & ~new_new_n32766__;
  assign new_new_n32768__ = pi00 & ~new_new_n32767__;
  assign new_new_n32769__ = pi01 & new_new_n32382__;
  assign new_new_n32770__ = ~pi02 & ~new_new_n32769__;
  assign new_new_n32771__ = ~pi01 & ~new_new_n26667__;
  assign new_new_n32772__ = ~new_new_n32769__ & ~new_new_n32771__;
  assign new_new_n32773__ = pi02 & ~new_new_n32772__;
  assign new_new_n32774__ = ~pi00 & ~new_new_n32770__;
  assign new_new_n32775__ = ~new_new_n32773__ & new_new_n32774__;
  assign new_new_n32776__ = ~new_new_n32768__ & ~new_new_n32775__;
  assign new_new_n32777__ = new_new_n13111__ & new_new_n27250__;
  assign new_new_n32778__ = new_new_n11469__ & new_new_n27284__;
  assign new_new_n32779__ = ~new_new_n32777__ & ~new_new_n32778__;
  assign new_new_n32780__ = new_new_n11478__ & ~new_new_n32779__;
  assign new_new_n32781__ = new_new_n11475__ & new_new_n26698__;
  assign new_new_n32782__ = ~new_new_n32780__ & ~new_new_n32781__;
  assign new_new_n32783__ = pi05 & ~new_new_n32782__;
  assign new_new_n32784__ = new_new_n12873__ & ~new_new_n26674__;
  assign new_new_n32785__ = new_new_n11469__ & ~new_new_n26674__;
  assign new_new_n32786__ = ~pi05 & ~new_new_n32785__;
  assign new_new_n32787__ = ~new_new_n32784__ & ~new_new_n32786__;
  assign new_new_n32788__ = new_new_n32782__ & ~new_new_n32787__;
  assign new_new_n32789__ = ~new_new_n32783__ & ~new_new_n32788__;
  assign new_new_n32790__ = ~new_new_n32647__ & ~new_new_n32652__;
  assign new_new_n32791__ = ~new_new_n32646__ & ~new_new_n32790__;
  assign new_new_n32792__ = new_new_n32789__ & ~new_new_n32791__;
  assign new_new_n32793__ = ~new_new_n32789__ & new_new_n32791__;
  assign new_new_n32794__ = ~new_new_n32792__ & ~new_new_n32793__;
  assign new_new_n32795__ = new_new_n10702__ & new_new_n26722__;
  assign new_new_n32796__ = ~new_new_n10697__ & new_new_n27352__;
  assign new_new_n32797__ = new_new_n27242__ & ~new_new_n32796__;
  assign new_new_n32798__ = ~new_new_n27242__ & new_new_n32796__;
  assign new_new_n32799__ = new_new_n10694__ & ~new_new_n32797__;
  assign new_new_n32800__ = ~new_new_n32798__ & new_new_n32799__;
  assign new_new_n32801__ = ~new_new_n32795__ & ~new_new_n32800__;
  assign new_new_n32802__ = new_new_n10709__ & new_new_n26729__;
  assign new_new_n32803__ = pi08 & ~new_new_n32802__;
  assign new_new_n32804__ = new_new_n10712__ & new_new_n26729__;
  assign new_new_n32805__ = ~pi08 & ~new_new_n32804__;
  assign new_new_n32806__ = pi05 & ~new_new_n32805__;
  assign new_new_n32807__ = ~new_new_n32803__ & ~new_new_n32806__;
  assign new_new_n32808__ = new_new_n32801__ & ~new_new_n32807__;
  assign new_new_n32809__ = ~pi08 & ~new_new_n32801__;
  assign new_new_n32810__ = ~new_new_n32808__ & ~new_new_n32809__;
  assign new_new_n32811__ = new_new_n8474__ & new_new_n26810__;
  assign new_new_n32812__ = ~new_new_n8479__ & ~new_new_n26802__;
  assign new_new_n32813__ = new_new_n8858__ & new_new_n26774__;
  assign new_new_n32814__ = ~new_new_n32811__ & ~new_new_n32812__;
  assign new_new_n32815__ = ~new_new_n32813__ & new_new_n32814__;
  assign new_new_n32816__ = new_new_n8469__ & ~new_new_n27373__;
  assign new_new_n32817__ = pi11 & ~new_new_n32816__;
  assign new_new_n32818__ = new_new_n11530__ & ~new_new_n27373__;
  assign new_new_n32819__ = ~new_new_n32817__ & ~new_new_n32818__;
  assign new_new_n32820__ = new_new_n32815__ & ~new_new_n32819__;
  assign new_new_n32821__ = ~pi11 & ~new_new_n32815__;
  assign new_new_n32822__ = ~new_new_n32820__ & ~new_new_n32821__;
  assign new_new_n32823__ = ~new_new_n32603__ & ~new_new_n32611__;
  assign new_new_n32824__ = new_new_n32603__ & new_new_n32611__;
  assign new_new_n32825__ = ~new_new_n32624__ & ~new_new_n32824__;
  assign new_new_n32826__ = ~new_new_n32823__ & ~new_new_n32825__;
  assign new_new_n32827__ = ~new_new_n32822__ & new_new_n32826__;
  assign new_new_n32828__ = new_new_n32822__ & ~new_new_n32826__;
  assign new_new_n32829__ = ~new_new_n32827__ & ~new_new_n32828__;
  assign new_new_n32830__ = new_new_n6985__ & ~new_new_n27221__;
  assign new_new_n32831__ = new_new_n6991__ & ~new_new_n26823__;
  assign new_new_n32832__ = ~new_new_n32830__ & ~new_new_n32831__;
  assign new_new_n32833__ = new_new_n6994__ & ~new_new_n26741__;
  assign new_new_n32834__ = new_new_n30393__ & new_new_n32833__;
  assign new_new_n32835__ = new_new_n32832__ & ~new_new_n32834__;
  assign new_new_n32836__ = ~pi14 & ~new_new_n32835__;
  assign new_new_n32837__ = ~pi13 & new_new_n26741__;
  assign new_new_n32838__ = pi13 & ~new_new_n26741__;
  assign new_new_n32839__ = new_new_n6994__ & new_new_n30390__;
  assign new_new_n32840__ = ~new_new_n32837__ & new_new_n32839__;
  assign new_new_n32841__ = ~new_new_n32838__ & new_new_n32840__;
  assign new_new_n32842__ = new_new_n6994__ & ~new_new_n30392__;
  assign new_new_n32843__ = pi14 & new_new_n32832__;
  assign new_new_n32844__ = ~new_new_n32842__ & new_new_n32843__;
  assign new_new_n32845__ = ~new_new_n32841__ & ~new_new_n32844__;
  assign new_new_n32846__ = ~new_new_n32836__ & new_new_n32845__;
  assign new_new_n32847__ = new_new_n32590__ & new_new_n32596__;
  assign new_new_n32848__ = ~new_new_n32601__ & ~new_new_n32847__;
  assign new_new_n32849__ = new_new_n32431__ & ~new_new_n32572__;
  assign new_new_n32850__ = ~new_new_n32571__ & ~new_new_n32849__;
  assign new_new_n32851__ = new_new_n6634__ & new_new_n26922__;
  assign new_new_n32852__ = ~new_new_n6625__ & new_new_n26917__;
  assign new_new_n32853__ = new_new_n6629__ & ~new_new_n27168__;
  assign new_new_n32854__ = new_new_n6936__ & ~new_new_n29366__;
  assign new_new_n32855__ = ~new_new_n32852__ & ~new_new_n32853__;
  assign new_new_n32856__ = ~new_new_n32851__ & new_new_n32855__;
  assign new_new_n32857__ = ~new_new_n32854__ & new_new_n32856__;
  assign new_new_n32858__ = ~pi20 & ~new_new_n32857__;
  assign new_new_n32859__ = pi20 & new_new_n32857__;
  assign new_new_n32860__ = ~new_new_n32858__ & ~new_new_n32859__;
  assign new_new_n32861__ = new_new_n7935__ & new_new_n26847__;
  assign new_new_n32862__ = new_new_n6964__ & ~new_new_n26888__;
  assign new_new_n32863__ = new_new_n6968__ & ~new_new_n26854__;
  assign new_new_n32864__ = ~new_new_n32862__ & ~new_new_n32863__;
  assign new_new_n32865__ = ~new_new_n32861__ & new_new_n32864__;
  assign new_new_n32866__ = new_new_n6958__ & new_new_n29424__;
  assign new_new_n32867__ = pi17 & ~new_new_n32866__;
  assign new_new_n32868__ = new_new_n7942__ & new_new_n29424__;
  assign new_new_n32869__ = ~new_new_n32867__ & ~new_new_n32868__;
  assign new_new_n32870__ = new_new_n32865__ & ~new_new_n32869__;
  assign new_new_n32871__ = ~pi17 & ~new_new_n32865__;
  assign new_new_n32872__ = ~new_new_n32870__ & ~new_new_n32871__;
  assign new_new_n32873__ = ~new_new_n32860__ & new_new_n32872__;
  assign new_new_n32874__ = new_new_n32860__ & ~new_new_n32872__;
  assign new_new_n32875__ = ~new_new_n32873__ & ~new_new_n32874__;
  assign new_new_n32876__ = new_new_n32550__ & new_new_n32562__;
  assign new_new_n32877__ = ~new_new_n32566__ & ~new_new_n32876__;
  assign new_new_n32878__ = new_new_n5191__ & new_new_n27152__;
  assign new_new_n32879__ = new_new_n5183__ & ~new_new_n26941__;
  assign new_new_n32880__ = new_new_n5213__ & new_new_n26928__;
  assign new_new_n32881__ = ~new_new_n32878__ & ~new_new_n32879__;
  assign new_new_n32882__ = ~new_new_n32880__ & new_new_n32881__;
  assign new_new_n32883__ = new_new_n5195__ & new_new_n27488__;
  assign new_new_n32884__ = pi23 & ~new_new_n32883__;
  assign new_new_n32885__ = new_new_n7878__ & new_new_n27488__;
  assign new_new_n32886__ = ~new_new_n32884__ & ~new_new_n32885__;
  assign new_new_n32887__ = new_new_n32882__ & ~new_new_n32886__;
  assign new_new_n32888__ = ~pi23 & ~new_new_n32882__;
  assign new_new_n32889__ = ~new_new_n32887__ & ~new_new_n32888__;
  assign new_new_n32890__ = ~pi23 & new_new_n32539__;
  assign new_new_n32891__ = pi23 & ~new_new_n32539__;
  assign new_new_n32892__ = ~new_new_n32890__ & ~new_new_n32891__;
  assign new_new_n32893__ = new_new_n32532__ & ~new_new_n32892__;
  assign new_new_n32894__ = ~new_new_n32532__ & new_new_n32892__;
  assign new_new_n32895__ = pi23 & new_new_n32539__;
  assign new_new_n32896__ = ~new_new_n32541__ & ~new_new_n32895__;
  assign new_new_n32897__ = new_new_n31324__ & ~new_new_n32896__;
  assign new_new_n32898__ = ~new_new_n31324__ & ~new_new_n32891__;
  assign new_new_n32899__ = ~new_new_n32540__ & new_new_n32898__;
  assign new_new_n32900__ = ~new_new_n32897__ & ~new_new_n32899__;
  assign new_new_n32901__ = new_new_n31410__ & new_new_n32900__;
  assign new_new_n32902__ = new_new_n31402__ & ~new_new_n32901__;
  assign new_new_n32903__ = ~new_new_n32894__ & ~new_new_n32902__;
  assign new_new_n32904__ = ~new_new_n32893__ & ~new_new_n32903__;
  assign new_new_n32905__ = new_new_n32889__ & ~new_new_n32904__;
  assign new_new_n32906__ = ~new_new_n32889__ & new_new_n32904__;
  assign new_new_n32907__ = ~new_new_n32905__ & ~new_new_n32906__;
  assign new_new_n32908__ = ~new_new_n4900__ & new_new_n28005__;
  assign new_new_n32909__ = ~new_new_n333__ & ~new_new_n26978__;
  assign new_new_n32910__ = new_new_n873__ & new_new_n26971__;
  assign new_new_n32911__ = ~new_new_n32909__ & ~new_new_n32910__;
  assign new_new_n32912__ = ~new_new_n32908__ & new_new_n32911__;
  assign new_new_n32913__ = pi26 & ~new_new_n32912__;
  assign new_new_n32914__ = new_new_n512__ & ~new_new_n26937__;
  assign new_new_n32915__ = new_new_n801__ & ~new_new_n26937__;
  assign new_new_n32916__ = ~pi26 & ~new_new_n32915__;
  assign new_new_n32917__ = ~new_new_n32914__ & ~new_new_n32916__;
  assign new_new_n32918__ = new_new_n32912__ & ~new_new_n32917__;
  assign new_new_n32919__ = ~new_new_n32913__ & ~new_new_n32918__;
  assign new_new_n32920__ = ~new_new_n32453__ & ~new_new_n32529__;
  assign new_new_n32921__ = ~new_new_n32452__ & ~new_new_n32920__;
  assign new_new_n32922__ = ~new_new_n32919__ & ~new_new_n32921__;
  assign new_new_n32923__ = new_new_n32919__ & new_new_n32921__;
  assign new_new_n32924__ = ~new_new_n32922__ & ~new_new_n32923__;
  assign new_new_n32925__ = new_new_n4815__ & ~new_new_n27003__;
  assign new_new_n32926__ = new_new_n4212__ & ~new_new_n27029__;
  assign new_new_n32927__ = ~new_new_n4818__ & ~new_new_n27021__;
  assign new_new_n32928__ = new_new_n4813__ & new_new_n27962__;
  assign new_new_n32929__ = ~new_new_n32926__ & ~new_new_n32927__;
  assign new_new_n32930__ = ~new_new_n32925__ & new_new_n32929__;
  assign new_new_n32931__ = ~new_new_n32928__ & new_new_n32930__;
  assign new_new_n32932__ = pi29 & ~new_new_n32931__;
  assign new_new_n32933__ = ~pi29 & new_new_n32931__;
  assign new_new_n32934__ = ~new_new_n32932__ & ~new_new_n32933__;
  assign new_new_n32935__ = ~new_new_n32464__ & ~new_new_n32525__;
  assign new_new_n32936__ = ~new_new_n32524__ & ~new_new_n32935__;
  assign new_new_n32937__ = ~new_new_n32934__ & ~new_new_n32936__;
  assign new_new_n32938__ = new_new_n32934__ & new_new_n32936__;
  assign new_new_n32939__ = ~new_new_n32937__ & ~new_new_n32938__;
  assign new_new_n32940__ = ~new_new_n32488__ & ~new_new_n32513__;
  assign new_new_n32941__ = ~new_new_n32489__ & ~new_new_n32940__;
  assign new_new_n32942__ = pi31 & new_new_n32481__;
  assign new_new_n32943__ = new_new_n5053__ & ~new_new_n27033__;
  assign new_new_n32944__ = pi31 & new_new_n27686__;
  assign new_new_n32945__ = new_new_n27111__ & new_new_n32944__;
  assign new_new_n32946__ = ~new_new_n27111__ & ~new_new_n32944__;
  assign new_new_n32947__ = ~new_new_n15853__ & ~new_new_n32945__;
  assign new_new_n32948__ = ~new_new_n32946__ & new_new_n32947__;
  assign new_new_n32949__ = ~new_new_n32942__ & ~new_new_n32943__;
  assign new_new_n32950__ = ~new_new_n32948__ & new_new_n32949__;
  assign new_new_n32951__ = new_new_n32941__ & new_new_n32950__;
  assign new_new_n32952__ = ~new_new_n32941__ & ~new_new_n32950__;
  assign new_new_n32953__ = new_new_n91__ & new_new_n16850__;
  assign new_new_n32954__ = ~new_new_n106__ & ~new_new_n692__;
  assign new_new_n32955__ = new_new_n28575__ & new_new_n32954__;
  assign new_new_n32956__ = ~new_new_n270__ & ~new_new_n311__;
  assign new_new_n32957__ = ~new_new_n871__ & ~new_new_n945__;
  assign new_new_n32958__ = new_new_n1382__ & new_new_n1741__;
  assign new_new_n32959__ = new_new_n2100__ & new_new_n28558__;
  assign new_new_n32960__ = ~new_new_n32953__ & new_new_n32959__;
  assign new_new_n32961__ = new_new_n32957__ & new_new_n32958__;
  assign new_new_n32962__ = new_new_n32955__ & new_new_n32956__;
  assign new_new_n32963__ = new_new_n1114__ & new_new_n1399__;
  assign new_new_n32964__ = new_new_n16852__ & new_new_n32963__;
  assign new_new_n32965__ = new_new_n32961__ & new_new_n32962__;
  assign new_new_n32966__ = new_new_n1381__ & new_new_n32960__;
  assign new_new_n32967__ = ~new_new_n1539__ & new_new_n32966__;
  assign new_new_n32968__ = new_new_n32964__ & new_new_n32965__;
  assign new_new_n32969__ = new_new_n2232__ & new_new_n32968__;
  assign new_new_n32970__ = new_new_n32967__ & new_new_n32969__;
  assign new_new_n32971__ = new_new_n4353__ & new_new_n32970__;
  assign new_new_n32972__ = new_new_n2157__ & new_new_n4340__;
  assign new_new_n32973__ = new_new_n32971__ & new_new_n32972__;
  assign new_new_n32974__ = ~new_new_n32951__ & ~new_new_n32973__;
  assign new_new_n32975__ = ~new_new_n32952__ & ~new_new_n32974__;
  assign new_new_n32976__ = ~new_new_n32951__ & new_new_n32975__;
  assign new_new_n32977__ = ~new_new_n32952__ & new_new_n32974__;
  assign new_new_n32978__ = ~new_new_n32973__ & ~new_new_n32977__;
  assign new_new_n32979__ = ~new_new_n32976__ & ~new_new_n32978__;
  assign new_new_n32980__ = new_new_n32939__ & ~new_new_n32979__;
  assign new_new_n32981__ = ~new_new_n32939__ & new_new_n32979__;
  assign new_new_n32982__ = ~new_new_n32980__ & ~new_new_n32981__;
  assign new_new_n32983__ = new_new_n32924__ & ~new_new_n32982__;
  assign new_new_n32984__ = ~new_new_n32924__ & new_new_n32982__;
  assign new_new_n32985__ = ~new_new_n32983__ & ~new_new_n32984__;
  assign new_new_n32986__ = new_new_n32907__ & ~new_new_n32985__;
  assign new_new_n32987__ = ~new_new_n32907__ & new_new_n32985__;
  assign new_new_n32988__ = ~new_new_n32986__ & ~new_new_n32987__;
  assign new_new_n32989__ = ~new_new_n32877__ & new_new_n32988__;
  assign new_new_n32990__ = new_new_n32877__ & ~new_new_n32988__;
  assign new_new_n32991__ = ~new_new_n32989__ & ~new_new_n32990__;
  assign new_new_n32992__ = new_new_n32875__ & ~new_new_n32991__;
  assign new_new_n32993__ = ~new_new_n32875__ & new_new_n32991__;
  assign new_new_n32994__ = ~new_new_n32992__ & ~new_new_n32993__;
  assign new_new_n32995__ = new_new_n32850__ & new_new_n32994__;
  assign new_new_n32996__ = ~new_new_n32850__ & ~new_new_n32994__;
  assign new_new_n32997__ = ~new_new_n32995__ & ~new_new_n32996__;
  assign new_new_n32998__ = ~new_new_n32848__ & ~new_new_n32997__;
  assign new_new_n32999__ = new_new_n32848__ & new_new_n32997__;
  assign new_new_n33000__ = ~new_new_n32998__ & ~new_new_n32999__;
  assign new_new_n33001__ = ~new_new_n32846__ & new_new_n33000__;
  assign new_new_n33002__ = new_new_n32846__ & ~new_new_n33000__;
  assign new_new_n33003__ = ~new_new_n33001__ & ~new_new_n33002__;
  assign new_new_n33004__ = new_new_n32829__ & ~new_new_n33003__;
  assign new_new_n33005__ = ~new_new_n32829__ & new_new_n33003__;
  assign new_new_n33006__ = ~new_new_n33004__ & ~new_new_n33005__;
  assign new_new_n33007__ = new_new_n32419__ & ~new_new_n32633__;
  assign new_new_n33008__ = ~new_new_n32419__ & new_new_n32633__;
  assign new_new_n33009__ = ~new_new_n32823__ & ~new_new_n32824__;
  assign new_new_n33010__ = new_new_n32624__ & new_new_n33009__;
  assign new_new_n33011__ = ~new_new_n32624__ & ~new_new_n33009__;
  assign new_new_n33012__ = ~new_new_n33010__ & ~new_new_n33011__;
  assign new_new_n33013__ = ~new_new_n33008__ & new_new_n33012__;
  assign new_new_n33014__ = ~new_new_n33007__ & ~new_new_n33013__;
  assign new_new_n33015__ = ~new_new_n33006__ & ~new_new_n33014__;
  assign new_new_n33016__ = new_new_n33006__ & new_new_n33014__;
  assign new_new_n33017__ = ~new_new_n33015__ & ~new_new_n33016__;
  assign new_new_n33018__ = new_new_n32810__ & ~new_new_n33017__;
  assign new_new_n33019__ = ~new_new_n32810__ & new_new_n33017__;
  assign new_new_n33020__ = ~new_new_n33018__ & ~new_new_n33019__;
  assign new_new_n33021__ = new_new_n32794__ & new_new_n33020__;
  assign new_new_n33022__ = ~new_new_n32794__ & ~new_new_n33020__;
  assign new_new_n33023__ = ~new_new_n33021__ & ~new_new_n33022__;
  assign new_new_n33024__ = new_new_n32776__ & ~new_new_n33023__;
  assign new_new_n33025__ = ~new_new_n32776__ & new_new_n33023__;
  assign new_new_n33026__ = ~new_new_n33024__ & ~new_new_n33025__;
  assign new_new_n33027__ = ~new_new_n32394__ & ~new_new_n32660__;
  assign new_new_n33028__ = ~new_new_n32661__ & ~new_new_n33027__;
  assign new_new_n33029__ = ~new_new_n32312__ & ~new_new_n32667__;
  assign new_new_n33030__ = new_new_n32312__ & new_new_n32672__;
  assign new_new_n33031__ = ~new_new_n33029__ & ~new_new_n33030__;
  assign new_new_n33032__ = new_new_n32665__ & new_new_n33031__;
  assign new_new_n33033__ = new_new_n33028__ & ~new_new_n33032__;
  assign new_new_n33034__ = new_new_n32661__ & new_new_n33032__;
  assign new_new_n33035__ = ~new_new_n33033__ & ~new_new_n33034__;
  assign new_new_n33036__ = new_new_n33026__ & ~new_new_n33035__;
  assign new_new_n33037__ = ~new_new_n32394__ & ~new_new_n32659__;
  assign new_new_n33038__ = new_new_n33032__ & new_new_n33037__;
  assign new_new_n33039__ = ~new_new_n33026__ & ~new_new_n33033__;
  assign new_new_n33040__ = ~new_new_n33038__ & new_new_n33039__;
  assign po02 = new_new_n33036__ | new_new_n33040__;
  assign new_new_n33042__ = ~new_new_n32661__ & ~new_new_n33026__;
  assign new_new_n33043__ = new_new_n33026__ & new_new_n33037__;
  assign new_new_n33044__ = new_new_n33032__ & ~new_new_n33042__;
  assign new_new_n33045__ = ~new_new_n33043__ & new_new_n33044__;
  assign new_new_n33046__ = new_new_n27289__ & new_new_n32742__;
  assign new_new_n33047__ = new_new_n27286__ & ~new_new_n32382__;
  assign new_new_n33048__ = new_new_n32729__ & ~new_new_n32737__;
  assign new_new_n33049__ = ~new_new_n33047__ & new_new_n33048__;
  assign new_new_n33050__ = ~new_new_n33046__ & ~new_new_n33049__;
  assign new_new_n33051__ = pi00 & pi02;
  assign new_new_n33052__ = ~new_new_n33050__ & new_new_n33051__;
  assign new_new_n33053__ = new_new_n32382__ & new_new_n32759__;
  assign new_new_n33054__ = pi00 & new_new_n33050__;
  assign new_new_n33055__ = ~new_new_n32740__ & new_new_n33054__;
  assign new_new_n33056__ = new_new_n14382__ & new_new_n32729__;
  assign new_new_n33057__ = ~new_new_n33053__ & ~new_new_n33056__;
  assign new_new_n33058__ = ~new_new_n33055__ & new_new_n33057__;
  assign new_new_n33059__ = pi01 & ~new_new_n33058__;
  assign new_new_n33060__ = ~new_new_n14382__ & ~new_new_n33051__;
  assign new_new_n33061__ = ~new_new_n32729__ & new_new_n33060__;
  assign new_new_n33062__ = ~new_new_n25581__ & ~new_new_n33061__;
  assign new_new_n33063__ = ~new_new_n32382__ & ~new_new_n33062__;
  assign new_new_n33064__ = ~new_new_n33052__ & ~new_new_n33063__;
  assign new_new_n33065__ = ~new_new_n33059__ & new_new_n33064__;
  assign new_new_n33066__ = ~new_new_n33025__ & new_new_n33028__;
  assign new_new_n33067__ = ~new_new_n33024__ & ~new_new_n33066__;
  assign new_new_n33068__ = ~new_new_n33065__ & new_new_n33067__;
  assign new_new_n33069__ = new_new_n33065__ & ~new_new_n33067__;
  assign new_new_n33070__ = ~new_new_n33068__ & ~new_new_n33069__;
  assign new_new_n33071__ = new_new_n13111__ & new_new_n26698__;
  assign new_new_n33072__ = new_new_n11469__ & ~new_new_n32340__;
  assign new_new_n33073__ = ~new_new_n33071__ & ~new_new_n33072__;
  assign new_new_n33074__ = new_new_n11478__ & ~new_new_n33073__;
  assign new_new_n33075__ = new_new_n11475__ & ~new_new_n26674__;
  assign new_new_n33076__ = ~new_new_n33074__ & ~new_new_n33075__;
  assign new_new_n33077__ = pi05 & ~new_new_n33076__;
  assign new_new_n33078__ = new_new_n12873__ & ~new_new_n26667__;
  assign new_new_n33079__ = new_new_n11469__ & ~new_new_n26667__;
  assign new_new_n33080__ = ~pi05 & ~new_new_n33079__;
  assign new_new_n33081__ = ~new_new_n33078__ & ~new_new_n33080__;
  assign new_new_n33082__ = new_new_n33076__ & ~new_new_n33081__;
  assign new_new_n33083__ = ~new_new_n33077__ & ~new_new_n33082__;
  assign new_new_n33084__ = new_new_n10698__ & new_new_n27250__;
  assign new_new_n33085__ = new_new_n10702__ & ~new_new_n27242__;
  assign new_new_n33086__ = ~new_new_n11409__ & new_new_n26722__;
  assign new_new_n33087__ = new_new_n11378__ & ~new_new_n27271__;
  assign new_new_n33088__ = ~new_new_n33085__ & ~new_new_n33086__;
  assign new_new_n33089__ = ~new_new_n33084__ & new_new_n33088__;
  assign new_new_n33090__ = ~new_new_n33087__ & new_new_n33089__;
  assign new_new_n33091__ = pi08 & ~new_new_n33090__;
  assign new_new_n33092__ = ~pi08 & new_new_n33090__;
  assign new_new_n33093__ = ~new_new_n33091__ & ~new_new_n33092__;
  assign new_new_n33094__ = ~new_new_n32810__ & ~new_new_n33016__;
  assign new_new_n33095__ = ~new_new_n33015__ & ~new_new_n33094__;
  assign new_new_n33096__ = new_new_n8858__ & new_new_n26729__;
  assign new_new_n33097__ = ~new_new_n8479__ & new_new_n26810__;
  assign new_new_n33098__ = new_new_n8474__ & new_new_n26774__;
  assign new_new_n33099__ = new_new_n8470__ & new_new_n30644__;
  assign new_new_n33100__ = ~new_new_n33096__ & ~new_new_n33097__;
  assign new_new_n33101__ = ~new_new_n33098__ & new_new_n33100__;
  assign new_new_n33102__ = ~new_new_n33099__ & new_new_n33101__;
  assign new_new_n33103__ = ~new_new_n32827__ & ~new_new_n33003__;
  assign new_new_n33104__ = ~new_new_n32828__ & ~new_new_n33103__;
  assign new_new_n33105__ = new_new_n6991__ & ~new_new_n27221__;
  assign new_new_n33106__ = new_new_n6985__ & ~new_new_n26741__;
  assign new_new_n33107__ = ~new_new_n33105__ & ~new_new_n33106__;
  assign new_new_n33108__ = new_new_n6994__ & ~new_new_n26802__;
  assign new_new_n33109__ = new_new_n30411__ & new_new_n33108__;
  assign new_new_n33110__ = new_new_n33107__ & ~new_new_n33109__;
  assign new_new_n33111__ = pi14 & ~new_new_n33110__;
  assign new_new_n33112__ = ~pi13 & ~new_new_n30692__;
  assign new_new_n33113__ = pi13 & ~new_new_n30410__;
  assign new_new_n33114__ = new_new_n6994__ & ~new_new_n33112__;
  assign new_new_n33115__ = ~new_new_n33113__ & new_new_n33114__;
  assign new_new_n33116__ = new_new_n6994__ & ~new_new_n27391__;
  assign new_new_n33117__ = ~pi14 & new_new_n33107__;
  assign new_new_n33118__ = ~new_new_n33116__ & new_new_n33117__;
  assign new_new_n33119__ = ~new_new_n33115__ & ~new_new_n33118__;
  assign new_new_n33120__ = ~new_new_n33111__ & new_new_n33119__;
  assign new_new_n33121__ = new_new_n6959__ & ~new_new_n29400__;
  assign new_new_n33122__ = new_new_n6964__ & ~new_new_n26854__;
  assign new_new_n33123__ = new_new_n6968__ & new_new_n26847__;
  assign new_new_n33124__ = new_new_n7935__ & ~new_new_n26823__;
  assign new_new_n33125__ = ~new_new_n33122__ & ~new_new_n33123__;
  assign new_new_n33126__ = ~new_new_n33124__ & new_new_n33125__;
  assign new_new_n33127__ = ~new_new_n33121__ & new_new_n33126__;
  assign new_new_n33128__ = pi17 & ~new_new_n33127__;
  assign new_new_n33129__ = ~pi17 & new_new_n33127__;
  assign new_new_n33130__ = ~new_new_n33128__ & ~new_new_n33129__;
  assign new_new_n33131__ = ~new_new_n32906__ & new_new_n32985__;
  assign new_new_n33132__ = ~new_new_n32905__ & ~new_new_n33131__;
  assign new_new_n33133__ = new_new_n4815__ & ~new_new_n26978__;
  assign new_new_n33134__ = new_new_n4212__ & ~new_new_n27003__;
  assign new_new_n33135__ = new_new_n4813__ & new_new_n27986__;
  assign new_new_n33136__ = ~new_new_n33133__ & ~new_new_n33134__;
  assign new_new_n33137__ = ~new_new_n33135__ & new_new_n33136__;
  assign new_new_n33138__ = new_new_n67__ & ~new_new_n27029__;
  assign new_new_n33139__ = pi29 & ~new_new_n33138__;
  assign new_new_n33140__ = new_new_n65__ & ~new_new_n27029__;
  assign new_new_n33141__ = ~pi29 & ~new_new_n33140__;
  assign new_new_n33142__ = pi26 & ~new_new_n33141__;
  assign new_new_n33143__ = ~new_new_n33139__ & ~new_new_n33142__;
  assign new_new_n33144__ = new_new_n33137__ & ~new_new_n33143__;
  assign new_new_n33145__ = ~pi29 & ~new_new_n33137__;
  assign new_new_n33146__ = ~new_new_n33144__ & ~new_new_n33145__;
  assign new_new_n33147__ = ~new_new_n32938__ & new_new_n32979__;
  assign new_new_n33148__ = ~new_new_n32937__ & ~new_new_n33147__;
  assign new_new_n33149__ = new_new_n33146__ & ~new_new_n33148__;
  assign new_new_n33150__ = ~new_new_n33146__ & new_new_n33148__;
  assign new_new_n33151__ = ~new_new_n33149__ & ~new_new_n33150__;
  assign new_new_n33152__ = new_new_n765__ & ~new_new_n27796__;
  assign new_new_n33153__ = new_new_n71__ & ~new_new_n27111__;
  assign new_new_n33154__ = new_new_n161__ & new_new_n27033__;
  assign new_new_n33155__ = pi31 & ~new_new_n33154__;
  assign new_new_n33156__ = ~new_new_n33153__ & new_new_n33155__;
  assign new_new_n33157__ = ~new_new_n33152__ & new_new_n33156__;
  assign new_new_n33158__ = ~new_new_n71__ & ~new_new_n27021__;
  assign new_new_n33159__ = ~new_new_n161__ & ~new_new_n33158__;
  assign new_new_n33160__ = new_new_n161__ & ~new_new_n27111__;
  assign new_new_n33161__ = ~pi31 & ~new_new_n33160__;
  assign new_new_n33162__ = ~new_new_n33159__ & new_new_n33161__;
  assign new_new_n33163__ = ~new_new_n33157__ & ~new_new_n33162__;
  assign new_new_n33164__ = new_new_n32975__ & new_new_n33163__;
  assign new_new_n33165__ = ~new_new_n32975__ & ~new_new_n33163__;
  assign new_new_n33166__ = ~new_new_n33164__ & ~new_new_n33165__;
  assign new_new_n33167__ = new_new_n224__ & ~new_new_n4479__;
  assign new_new_n33168__ = new_new_n744__ & ~new_new_n33167__;
  assign new_new_n33169__ = new_new_n962__ & new_new_n33168__;
  assign new_new_n33170__ = ~new_new_n202__ & ~new_new_n1007__;
  assign new_new_n33171__ = ~new_new_n346__ & new_new_n710__;
  assign new_new_n33172__ = ~new_new_n2329__ & new_new_n4728__;
  assign new_new_n33173__ = new_new_n33171__ & new_new_n33172__;
  assign new_new_n33174__ = new_new_n5313__ & new_new_n33170__;
  assign new_new_n33175__ = new_new_n33173__ & new_new_n33174__;
  assign new_new_n33176__ = new_new_n2315__ & new_new_n2387__;
  assign new_new_n33177__ = new_new_n33175__ & new_new_n33176__;
  assign new_new_n33178__ = new_new_n5569__ & new_new_n19016__;
  assign new_new_n33179__ = new_new_n33169__ & new_new_n33178__;
  assign new_new_n33180__ = new_new_n33177__ & new_new_n33179__;
  assign new_new_n33181__ = new_new_n4594__ & new_new_n33180__;
  assign new_new_n33182__ = new_new_n2790__ & new_new_n7629__;
  assign new_new_n33183__ = new_new_n33181__ & new_new_n33182__;
  assign new_new_n33184__ = ~new_new_n33166__ & new_new_n33183__;
  assign new_new_n33185__ = new_new_n33166__ & ~new_new_n33183__;
  assign new_new_n33186__ = ~new_new_n33184__ & ~new_new_n33185__;
  assign new_new_n33187__ = new_new_n33151__ & new_new_n33186__;
  assign new_new_n33188__ = ~new_new_n33151__ & ~new_new_n33186__;
  assign new_new_n33189__ = ~new_new_n33187__ & ~new_new_n33188__;
  assign new_new_n33190__ = ~new_new_n32923__ & ~new_new_n32982__;
  assign new_new_n33191__ = ~new_new_n32922__ & ~new_new_n33190__;
  assign new_new_n33192__ = new_new_n504__ & ~new_new_n28666__;
  assign new_new_n33193__ = new_new_n3311__ & new_new_n27152__;
  assign new_new_n33194__ = ~new_new_n333__ & new_new_n26971__;
  assign new_new_n33195__ = new_new_n873__ & ~new_new_n26937__;
  assign new_new_n33196__ = ~new_new_n33194__ & ~new_new_n33195__;
  assign new_new_n33197__ = ~new_new_n33193__ & new_new_n33196__;
  assign new_new_n33198__ = ~pi26 & ~new_new_n33197__;
  assign new_new_n33199__ = pi26 & new_new_n33197__;
  assign new_new_n33200__ = ~new_new_n33198__ & ~new_new_n33199__;
  assign new_new_n33201__ = ~new_new_n4899__ & ~new_new_n33200__;
  assign new_new_n33202__ = new_new_n28666__ & new_new_n33199__;
  assign new_new_n33203__ = ~new_new_n33192__ & ~new_new_n33201__;
  assign new_new_n33204__ = ~new_new_n33202__ & new_new_n33203__;
  assign new_new_n33205__ = new_new_n33191__ & ~new_new_n33204__;
  assign new_new_n33206__ = ~new_new_n33191__ & new_new_n33204__;
  assign new_new_n33207__ = ~new_new_n33205__ & ~new_new_n33206__;
  assign new_new_n33208__ = new_new_n33189__ & new_new_n33207__;
  assign new_new_n33209__ = ~new_new_n33189__ & ~new_new_n33207__;
  assign new_new_n33210__ = ~new_new_n33208__ & ~new_new_n33209__;
  assign new_new_n33211__ = new_new_n33132__ & new_new_n33210__;
  assign new_new_n33212__ = ~new_new_n33132__ & ~new_new_n33210__;
  assign new_new_n33213__ = ~new_new_n33211__ & ~new_new_n33212__;
  assign new_new_n33214__ = new_new_n5213__ & new_new_n26917__;
  assign new_new_n33215__ = new_new_n5191__ & ~new_new_n26941__;
  assign new_new_n33216__ = new_new_n5183__ & new_new_n26928__;
  assign new_new_n33217__ = ~new_new_n33215__ & ~new_new_n33216__;
  assign new_new_n33218__ = ~new_new_n33214__ & new_new_n33217__;
  assign new_new_n33219__ = new_new_n5195__ & ~new_new_n27462__;
  assign new_new_n33220__ = ~pi23 & ~new_new_n33219__;
  assign new_new_n33221__ = new_new_n5974__ & ~new_new_n27462__;
  assign new_new_n33222__ = ~new_new_n33220__ & ~new_new_n33221__;
  assign new_new_n33223__ = new_new_n33218__ & ~new_new_n33222__;
  assign new_new_n33224__ = pi23 & ~new_new_n33218__;
  assign new_new_n33225__ = ~new_new_n33223__ & ~new_new_n33224__;
  assign new_new_n33226__ = ~new_new_n33213__ & new_new_n33225__;
  assign new_new_n33227__ = new_new_n33213__ & ~new_new_n33225__;
  assign new_new_n33228__ = ~new_new_n33226__ & ~new_new_n33227__;
  assign new_new_n33229__ = new_new_n6936__ & new_new_n27180__;
  assign new_new_n33230__ = ~new_new_n6625__ & ~new_new_n27168__;
  assign new_new_n33231__ = ~new_new_n33229__ & ~new_new_n33230__;
  assign new_new_n33232__ = new_new_n6629__ & new_new_n26922__;
  assign new_new_n33233__ = new_new_n6634__ & ~new_new_n26888__;
  assign new_new_n33234__ = ~new_new_n33232__ & ~new_new_n33233__;
  assign new_new_n33235__ = new_new_n33231__ & new_new_n33234__;
  assign new_new_n33236__ = pi20 & ~new_new_n33235__;
  assign new_new_n33237__ = ~new_new_n6634__ & ~new_new_n26922__;
  assign new_new_n33238__ = new_new_n6629__ & ~new_new_n33237__;
  assign new_new_n33239__ = ~pi20 & ~new_new_n33238__;
  assign new_new_n33240__ = ~new_new_n33233__ & new_new_n33239__;
  assign new_new_n33241__ = new_new_n33231__ & new_new_n33240__;
  assign new_new_n33242__ = ~new_new_n33236__ & ~new_new_n33241__;
  assign new_new_n33243__ = new_new_n33228__ & ~new_new_n33242__;
  assign new_new_n33244__ = ~new_new_n33228__ & new_new_n33242__;
  assign new_new_n33245__ = ~new_new_n33243__ & ~new_new_n33244__;
  assign new_new_n33246__ = new_new_n32860__ & ~new_new_n32989__;
  assign new_new_n33247__ = ~new_new_n32990__ & ~new_new_n33246__;
  assign new_new_n33248__ = new_new_n33245__ & new_new_n33247__;
  assign new_new_n33249__ = ~new_new_n33245__ & ~new_new_n33247__;
  assign new_new_n33250__ = ~new_new_n33248__ & ~new_new_n33249__;
  assign new_new_n33251__ = new_new_n33130__ & new_new_n33250__;
  assign new_new_n33252__ = ~new_new_n33130__ & ~new_new_n33250__;
  assign new_new_n33253__ = ~new_new_n33251__ & ~new_new_n33252__;
  assign new_new_n33254__ = ~new_new_n32850__ & ~new_new_n32872__;
  assign new_new_n33255__ = new_new_n32850__ & new_new_n32872__;
  assign new_new_n33256__ = new_new_n32860__ & ~new_new_n32991__;
  assign new_new_n33257__ = ~new_new_n32860__ & new_new_n32991__;
  assign new_new_n33258__ = ~new_new_n33256__ & ~new_new_n33257__;
  assign new_new_n33259__ = ~new_new_n33255__ & new_new_n33258__;
  assign new_new_n33260__ = ~new_new_n33254__ & ~new_new_n33259__;
  assign new_new_n33261__ = new_new_n33253__ & ~new_new_n33260__;
  assign new_new_n33262__ = ~new_new_n33253__ & new_new_n33260__;
  assign new_new_n33263__ = ~new_new_n33261__ & ~new_new_n33262__;
  assign new_new_n33264__ = new_new_n33120__ & new_new_n33263__;
  assign new_new_n33265__ = ~new_new_n33120__ & ~new_new_n33263__;
  assign new_new_n33266__ = ~new_new_n33264__ & ~new_new_n33265__;
  assign new_new_n33267__ = ~new_new_n32846__ & ~new_new_n32999__;
  assign new_new_n33268__ = ~new_new_n32998__ & ~new_new_n33267__;
  assign new_new_n33269__ = new_new_n33266__ & new_new_n33268__;
  assign new_new_n33270__ = ~new_new_n33266__ & ~new_new_n33268__;
  assign new_new_n33271__ = ~new_new_n33269__ & ~new_new_n33270__;
  assign new_new_n33272__ = ~new_new_n33104__ & new_new_n33271__;
  assign new_new_n33273__ = new_new_n33104__ & ~new_new_n33271__;
  assign new_new_n33274__ = ~new_new_n33272__ & ~new_new_n33273__;
  assign new_new_n33275__ = pi11 & ~new_new_n33274__;
  assign new_new_n33276__ = ~pi11 & new_new_n33274__;
  assign new_new_n33277__ = ~new_new_n33275__ & ~new_new_n33276__;
  assign new_new_n33278__ = new_new_n33102__ & new_new_n33277__;
  assign new_new_n33279__ = ~new_new_n33102__ & ~new_new_n33277__;
  assign new_new_n33280__ = ~new_new_n33278__ & ~new_new_n33279__;
  assign new_new_n33281__ = new_new_n33095__ & new_new_n33280__;
  assign new_new_n33282__ = ~new_new_n33095__ & ~new_new_n33280__;
  assign new_new_n33283__ = ~new_new_n33281__ & ~new_new_n33282__;
  assign new_new_n33284__ = new_new_n33093__ & ~new_new_n33283__;
  assign new_new_n33285__ = ~new_new_n33093__ & new_new_n33283__;
  assign new_new_n33286__ = ~new_new_n33284__ & ~new_new_n33285__;
  assign new_new_n33287__ = new_new_n32792__ & ~new_new_n33286__;
  assign new_new_n33288__ = new_new_n32793__ & new_new_n33286__;
  assign new_new_n33289__ = ~new_new_n32793__ & ~new_new_n33286__;
  assign new_new_n33290__ = new_new_n32810__ & ~new_new_n33289__;
  assign new_new_n33291__ = ~new_new_n32792__ & new_new_n33286__;
  assign new_new_n33292__ = ~new_new_n32810__ & ~new_new_n33291__;
  assign new_new_n33293__ = new_new_n33017__ & ~new_new_n33290__;
  assign new_new_n33294__ = ~new_new_n33292__ & new_new_n33293__;
  assign new_new_n33295__ = new_new_n32810__ & ~new_new_n33291__;
  assign new_new_n33296__ = ~new_new_n32810__ & ~new_new_n33289__;
  assign new_new_n33297__ = ~new_new_n33017__ & ~new_new_n33295__;
  assign new_new_n33298__ = ~new_new_n33296__ & new_new_n33297__;
  assign new_new_n33299__ = ~new_new_n33288__ & ~new_new_n33294__;
  assign new_new_n33300__ = ~new_new_n33298__ & new_new_n33299__;
  assign new_new_n33301__ = ~new_new_n33287__ & new_new_n33300__;
  assign new_new_n33302__ = new_new_n33083__ & ~new_new_n33301__;
  assign new_new_n33303__ = ~new_new_n33083__ & new_new_n33301__;
  assign new_new_n33304__ = ~new_new_n33302__ & ~new_new_n33303__;
  assign new_new_n33305__ = ~new_new_n33070__ & ~new_new_n33304__;
  assign new_new_n33306__ = new_new_n33070__ & new_new_n33304__;
  assign new_new_n33307__ = ~new_new_n33305__ & ~new_new_n33306__;
  assign new_new_n33308__ = new_new_n33045__ & new_new_n33307__;
  assign new_new_n33309__ = ~new_new_n33045__ & ~new_new_n33307__;
  assign po03 = ~new_new_n33308__ & ~new_new_n33309__;
  assign new_new_n33311__ = pi00 & ~new_new_n33050__;
  assign new_new_n33312__ = ~pi02 & ~new_new_n33311__;
  assign new_new_n33313__ = new_new_n32729__ & ~new_new_n33312__;
  assign new_new_n33314__ = ~new_new_n13986__ & new_new_n32740__;
  assign new_new_n33315__ = ~new_new_n33313__ & ~new_new_n33314__;
  assign new_new_n33316__ = pi01 & ~new_new_n33315__;
  assign new_new_n33317__ = new_new_n32729__ & new_new_n33054__;
  assign new_new_n33318__ = new_new_n14393__ & ~new_new_n32729__;
  assign new_new_n33319__ = ~new_new_n32730__ & ~new_new_n33318__;
  assign new_new_n33320__ = ~new_new_n33317__ & new_new_n33319__;
  assign new_new_n33321__ = pi02 & ~new_new_n33320__;
  assign new_new_n33322__ = ~new_new_n33316__ & ~new_new_n33321__;
  assign new_new_n33323__ = new_new_n33286__ & new_new_n33300__;
  assign new_new_n33324__ = ~new_new_n33302__ & ~new_new_n33323__;
  assign new_new_n33325__ = new_new_n11471__ & ~new_new_n26674__;
  assign new_new_n33326__ = new_new_n11475__ & ~new_new_n26667__;
  assign new_new_n33327__ = ~new_new_n32343__ & new_new_n32382__;
  assign new_new_n33328__ = ~new_new_n26698__ & new_new_n32742__;
  assign new_new_n33329__ = ~new_new_n26667__ & new_new_n32747__;
  assign new_new_n33330__ = ~new_new_n27273__ & new_new_n33329__;
  assign new_new_n33331__ = ~new_new_n33328__ & ~new_new_n33330__;
  assign new_new_n33332__ = ~new_new_n27250__ & ~new_new_n33331__;
  assign new_new_n33333__ = new_new_n26698__ & new_new_n32736__;
  assign new_new_n33334__ = ~new_new_n26674__ & new_new_n32737__;
  assign new_new_n33335__ = new_new_n27273__ & new_new_n33334__;
  assign new_new_n33336__ = ~new_new_n33333__ & ~new_new_n33335__;
  assign new_new_n33337__ = new_new_n27250__ & ~new_new_n33336__;
  assign new_new_n33338__ = new_new_n27273__ & new_new_n32736__;
  assign new_new_n33339__ = ~new_new_n33334__ & ~new_new_n33338__;
  assign new_new_n33340__ = new_new_n26698__ & ~new_new_n33339__;
  assign new_new_n33341__ = ~new_new_n27273__ & new_new_n32742__;
  assign new_new_n33342__ = ~new_new_n33329__ & ~new_new_n33341__;
  assign new_new_n33343__ = ~new_new_n26698__ & ~new_new_n33342__;
  assign new_new_n33344__ = ~new_new_n33340__ & ~new_new_n33343__;
  assign new_new_n33345__ = ~new_new_n33332__ & new_new_n33344__;
  assign new_new_n33346__ = ~new_new_n33337__ & new_new_n33345__;
  assign new_new_n33347__ = ~new_new_n33327__ & new_new_n33346__;
  assign new_new_n33348__ = new_new_n11478__ & new_new_n33347__;
  assign new_new_n33349__ = ~new_new_n11478__ & ~new_new_n32382__;
  assign new_new_n33350__ = ~new_new_n11482__ & ~new_new_n33349__;
  assign new_new_n33351__ = ~new_new_n33348__ & new_new_n33350__;
  assign new_new_n33352__ = ~new_new_n33325__ & ~new_new_n33326__;
  assign new_new_n33353__ = ~new_new_n33351__ & new_new_n33352__;
  assign new_new_n33354__ = pi05 & ~new_new_n33353__;
  assign new_new_n33355__ = ~pi05 & new_new_n33353__;
  assign new_new_n33356__ = ~new_new_n33354__ & ~new_new_n33355__;
  assign new_new_n33357__ = new_new_n7935__ & ~new_new_n27221__;
  assign new_new_n33358__ = new_new_n6964__ & new_new_n26847__;
  assign new_new_n33359__ = new_new_n6968__ & ~new_new_n26823__;
  assign new_new_n33360__ = ~new_new_n33358__ & ~new_new_n33359__;
  assign new_new_n33361__ = ~new_new_n33357__ & new_new_n33360__;
  assign new_new_n33362__ = new_new_n6958__ & new_new_n27411__;
  assign new_new_n33363__ = pi17 & ~new_new_n33362__;
  assign new_new_n33364__ = new_new_n7942__ & new_new_n27411__;
  assign new_new_n33365__ = ~new_new_n33363__ & ~new_new_n33364__;
  assign new_new_n33366__ = new_new_n33361__ & ~new_new_n33365__;
  assign new_new_n33367__ = ~pi17 & ~new_new_n33361__;
  assign new_new_n33368__ = ~new_new_n33366__ & ~new_new_n33367__;
  assign new_new_n33369__ = ~new_new_n33251__ & new_new_n33260__;
  assign new_new_n33370__ = ~new_new_n33252__ & ~new_new_n33369__;
  assign new_new_n33371__ = new_new_n33368__ & ~new_new_n33370__;
  assign new_new_n33372__ = ~new_new_n33368__ & new_new_n33370__;
  assign new_new_n33373__ = ~new_new_n33371__ & ~new_new_n33372__;
  assign new_new_n33374__ = new_new_n5183__ & new_new_n26917__;
  assign new_new_n33375__ = new_new_n5191__ & new_new_n26928__;
  assign new_new_n33376__ = new_new_n5213__ & ~new_new_n27168__;
  assign new_new_n33377__ = ~new_new_n33375__ & ~new_new_n33376__;
  assign new_new_n33378__ = ~new_new_n33374__ & new_new_n33377__;
  assign new_new_n33379__ = new_new_n5195__ & ~new_new_n28799__;
  assign new_new_n33380__ = pi23 & ~new_new_n33379__;
  assign new_new_n33381__ = new_new_n7878__ & ~new_new_n28799__;
  assign new_new_n33382__ = ~new_new_n33380__ & ~new_new_n33381__;
  assign new_new_n33383__ = new_new_n33378__ & ~new_new_n33382__;
  assign new_new_n33384__ = ~pi23 & ~new_new_n33378__;
  assign new_new_n33385__ = ~new_new_n33383__ & ~new_new_n33384__;
  assign new_new_n33386__ = ~new_new_n33211__ & ~new_new_n33225__;
  assign new_new_n33387__ = ~new_new_n33212__ & ~new_new_n33386__;
  assign new_new_n33388__ = ~new_new_n33385__ & new_new_n33387__;
  assign new_new_n33389__ = new_new_n33385__ & ~new_new_n33387__;
  assign new_new_n33390__ = ~new_new_n33388__ & ~new_new_n33389__;
  assign new_new_n33391__ = new_new_n873__ & new_new_n27152__;
  assign new_new_n33392__ = new_new_n3311__ & ~new_new_n26941__;
  assign new_new_n33393__ = ~new_new_n333__ & ~new_new_n26937__;
  assign new_new_n33394__ = ~new_new_n4900__ & ~new_new_n27502__;
  assign new_new_n33395__ = ~new_new_n33392__ & ~new_new_n33393__;
  assign new_new_n33396__ = ~new_new_n33391__ & new_new_n33395__;
  assign new_new_n33397__ = ~new_new_n33394__ & new_new_n33396__;
  assign new_new_n33398__ = new_new_n33189__ & ~new_new_n33206__;
  assign new_new_n33399__ = ~new_new_n33205__ & ~new_new_n33398__;
  assign new_new_n33400__ = ~new_new_n33164__ & ~new_new_n33183__;
  assign new_new_n33401__ = ~new_new_n33165__ & ~new_new_n33400__;
  assign new_new_n33402__ = new_new_n161__ & ~new_new_n27021__;
  assign new_new_n33403__ = new_new_n765__ & ~new_new_n27029__;
  assign new_new_n33404__ = ~new_new_n33402__ & ~new_new_n33403__;
  assign new_new_n33405__ = ~pi31 & ~new_new_n33404__;
  assign new_new_n33406__ = new_new_n765__ & ~new_new_n27764__;
  assign new_new_n33407__ = new_new_n71__ & new_new_n27021__;
  assign new_new_n33408__ = pi31 & ~new_new_n33160__;
  assign new_new_n33409__ = ~new_new_n33407__ & new_new_n33408__;
  assign new_new_n33410__ = ~new_new_n33406__ & new_new_n33409__;
  assign new_new_n33411__ = ~new_new_n33405__ & ~new_new_n33410__;
  assign new_new_n33412__ = ~new_new_n208__ & ~new_new_n247__;
  assign new_new_n33413__ = ~new_new_n312__ & ~new_new_n336__;
  assign new_new_n33414__ = ~new_new_n509__ & ~new_new_n963__;
  assign new_new_n33415__ = new_new_n33413__ & new_new_n33414__;
  assign new_new_n33416__ = ~new_new_n732__ & new_new_n33412__;
  assign new_new_n33417__ = new_new_n5459__ & new_new_n33416__;
  assign new_new_n33418__ = new_new_n7091__ & new_new_n33415__;
  assign new_new_n33419__ = new_new_n16894__ & new_new_n33418__;
  assign new_new_n33420__ = new_new_n3259__ & new_new_n33417__;
  assign new_new_n33421__ = new_new_n33419__ & new_new_n33420__;
  assign new_new_n33422__ = ~new_new_n253__ & ~new_new_n937__;
  assign new_new_n33423__ = ~new_new_n483__ & new_new_n33422__;
  assign new_new_n33424__ = new_new_n1449__ & new_new_n1740__;
  assign new_new_n33425__ = new_new_n2712__ & new_new_n33424__;
  assign new_new_n33426__ = new_new_n1180__ & new_new_n33423__;
  assign new_new_n33427__ = ~new_new_n124__ & ~new_new_n607__;
  assign new_new_n33428__ = new_new_n628__ & new_new_n872__;
  assign new_new_n33429__ = new_new_n2331__ & new_new_n2424__;
  assign new_new_n33430__ = new_new_n3516__ & new_new_n3788__;
  assign new_new_n33431__ = new_new_n33429__ & new_new_n33430__;
  assign new_new_n33432__ = new_new_n33427__ & new_new_n33428__;
  assign new_new_n33433__ = new_new_n33425__ & new_new_n33426__;
  assign new_new_n33434__ = new_new_n2580__ & new_new_n33433__;
  assign new_new_n33435__ = new_new_n33431__ & new_new_n33432__;
  assign new_new_n33436__ = new_new_n33434__ & new_new_n33435__;
  assign new_new_n33437__ = new_new_n33421__ & new_new_n33436__;
  assign new_new_n33438__ = new_new_n4412__ & new_new_n33437__;
  assign new_new_n33439__ = new_new_n5337__ & new_new_n33438__;
  assign new_new_n33440__ = ~new_new_n33411__ & ~new_new_n33439__;
  assign new_new_n33441__ = new_new_n33411__ & new_new_n33439__;
  assign new_new_n33442__ = ~new_new_n33440__ & ~new_new_n33441__;
  assign new_new_n33443__ = ~new_new_n33401__ & new_new_n33442__;
  assign new_new_n33444__ = ~new_new_n5324__ & new_new_n33439__;
  assign new_new_n33445__ = ~new_new_n33442__ & ~new_new_n33444__;
  assign new_new_n33446__ = new_new_n33401__ & new_new_n33445__;
  assign new_new_n33447__ = ~new_new_n33443__ & ~new_new_n33446__;
  assign new_new_n33448__ = new_new_n4815__ & new_new_n26971__;
  assign new_new_n33449__ = new_new_n4212__ & ~new_new_n26978__;
  assign new_new_n33450__ = ~new_new_n4818__ & ~new_new_n27003__;
  assign new_new_n33451__ = new_new_n4813__ & new_new_n28277__;
  assign new_new_n33452__ = ~new_new_n33449__ & ~new_new_n33450__;
  assign new_new_n33453__ = ~new_new_n33448__ & new_new_n33452__;
  assign new_new_n33454__ = ~new_new_n33451__ & new_new_n33453__;
  assign new_new_n33455__ = ~new_new_n33149__ & new_new_n33186__;
  assign new_new_n33456__ = ~new_new_n33150__ & ~new_new_n33455__;
  assign new_new_n33457__ = pi29 & ~new_new_n33456__;
  assign new_new_n33458__ = ~pi29 & new_new_n33456__;
  assign new_new_n33459__ = ~new_new_n33457__ & ~new_new_n33458__;
  assign new_new_n33460__ = new_new_n33454__ & new_new_n33459__;
  assign new_new_n33461__ = ~new_new_n33454__ & ~new_new_n33459__;
  assign new_new_n33462__ = ~new_new_n33460__ & ~new_new_n33461__;
  assign new_new_n33463__ = ~new_new_n33447__ & new_new_n33462__;
  assign new_new_n33464__ = new_new_n33447__ & ~new_new_n33462__;
  assign new_new_n33465__ = ~new_new_n33463__ & ~new_new_n33464__;
  assign new_new_n33466__ = pi26 & ~new_new_n33465__;
  assign new_new_n33467__ = ~pi26 & new_new_n33465__;
  assign new_new_n33468__ = ~new_new_n33466__ & ~new_new_n33467__;
  assign new_new_n33469__ = new_new_n33399__ & ~new_new_n33468__;
  assign new_new_n33470__ = ~new_new_n33399__ & new_new_n33468__;
  assign new_new_n33471__ = ~new_new_n33469__ & ~new_new_n33470__;
  assign new_new_n33472__ = new_new_n33397__ & new_new_n33471__;
  assign new_new_n33473__ = ~new_new_n33397__ & ~new_new_n33471__;
  assign new_new_n33474__ = ~new_new_n33472__ & ~new_new_n33473__;
  assign new_new_n33475__ = new_new_n33390__ & ~new_new_n33474__;
  assign new_new_n33476__ = ~new_new_n33390__ & new_new_n33474__;
  assign new_new_n33477__ = ~new_new_n33475__ & ~new_new_n33476__;
  assign new_new_n33478__ = ~new_new_n33244__ & ~new_new_n33247__;
  assign new_new_n33479__ = ~new_new_n33243__ & ~new_new_n33478__;
  assign new_new_n33480__ = new_new_n33477__ & ~new_new_n33479__;
  assign new_new_n33481__ = ~new_new_n33477__ & new_new_n33479__;
  assign new_new_n33482__ = ~new_new_n33480__ & ~new_new_n33481__;
  assign new_new_n33483__ = new_new_n6634__ & ~new_new_n26854__;
  assign new_new_n33484__ = new_new_n6629__ & ~new_new_n26888__;
  assign new_new_n33485__ = ~new_new_n6625__ & new_new_n26922__;
  assign new_new_n33486__ = new_new_n6936__ & ~new_new_n27430__;
  assign new_new_n33487__ = ~new_new_n33484__ & ~new_new_n33485__;
  assign new_new_n33488__ = ~new_new_n33486__ & new_new_n33487__;
  assign new_new_n33489__ = ~new_new_n33483__ & new_new_n33488__;
  assign new_new_n33490__ = ~pi20 & ~new_new_n33489__;
  assign new_new_n33491__ = ~new_new_n6629__ & new_new_n26854__;
  assign new_new_n33492__ = new_new_n6640__ & ~new_new_n33491__;
  assign new_new_n33493__ = pi20 & ~new_new_n33492__;
  assign new_new_n33494__ = new_new_n33488__ & new_new_n33493__;
  assign new_new_n33495__ = ~new_new_n33490__ & ~new_new_n33494__;
  assign new_new_n33496__ = new_new_n33482__ & new_new_n33495__;
  assign new_new_n33497__ = ~new_new_n33482__ & ~new_new_n33495__;
  assign new_new_n33498__ = ~new_new_n33496__ & ~new_new_n33497__;
  assign new_new_n33499__ = new_new_n33373__ & ~new_new_n33498__;
  assign new_new_n33500__ = ~new_new_n33373__ & new_new_n33498__;
  assign new_new_n33501__ = ~new_new_n33499__ & ~new_new_n33500__;
  assign new_new_n33502__ = ~new_new_n33272__ & ~new_new_n33280__;
  assign new_new_n33503__ = ~new_new_n33273__ & ~new_new_n33502__;
  assign new_new_n33504__ = ~new_new_n33264__ & new_new_n33268__;
  assign new_new_n33505__ = ~new_new_n33265__ & ~new_new_n33504__;
  assign new_new_n33506__ = new_new_n6991__ & ~new_new_n26741__;
  assign new_new_n33507__ = new_new_n6985__ & ~new_new_n26802__;
  assign new_new_n33508__ = ~new_new_n10772__ & ~new_new_n26810__;
  assign new_new_n33509__ = new_new_n10772__ & ~new_new_n27395__;
  assign new_new_n33510__ = new_new_n6994__ & ~new_new_n33508__;
  assign new_new_n33511__ = ~new_new_n33509__ & new_new_n33510__;
  assign new_new_n33512__ = ~new_new_n33506__ & ~new_new_n33507__;
  assign new_new_n33513__ = ~new_new_n33511__ & new_new_n33512__;
  assign new_new_n33514__ = pi14 & ~new_new_n33513__;
  assign new_new_n33515__ = ~pi14 & new_new_n33513__;
  assign new_new_n33516__ = ~new_new_n33514__ & ~new_new_n33515__;
  assign new_new_n33517__ = new_new_n8474__ & new_new_n26729__;
  assign new_new_n33518__ = ~new_new_n8479__ & new_new_n26774__;
  assign new_new_n33519__ = new_new_n8858__ & new_new_n26722__;
  assign new_new_n33520__ = ~new_new_n33517__ & ~new_new_n33518__;
  assign new_new_n33521__ = ~new_new_n33519__ & new_new_n33520__;
  assign new_new_n33522__ = new_new_n8469__ & ~new_new_n27348__;
  assign new_new_n33523__ = pi11 & ~new_new_n33522__;
  assign new_new_n33524__ = new_new_n11530__ & ~new_new_n27348__;
  assign new_new_n33525__ = ~new_new_n33523__ & ~new_new_n33524__;
  assign new_new_n33526__ = new_new_n33521__ & ~new_new_n33525__;
  assign new_new_n33527__ = ~pi11 & ~new_new_n33521__;
  assign new_new_n33528__ = ~new_new_n33526__ & ~new_new_n33527__;
  assign new_new_n33529__ = new_new_n33516__ & ~new_new_n33528__;
  assign new_new_n33530__ = ~new_new_n33516__ & new_new_n33528__;
  assign new_new_n33531__ = ~new_new_n33529__ & ~new_new_n33530__;
  assign new_new_n33532__ = new_new_n33505__ & new_new_n33531__;
  assign new_new_n33533__ = ~new_new_n33505__ & ~new_new_n33531__;
  assign new_new_n33534__ = ~new_new_n33532__ & ~new_new_n33533__;
  assign new_new_n33535__ = new_new_n33503__ & ~new_new_n33534__;
  assign new_new_n33536__ = ~new_new_n33503__ & new_new_n33534__;
  assign new_new_n33537__ = ~new_new_n33535__ & ~new_new_n33536__;
  assign new_new_n33538__ = new_new_n33501__ & new_new_n33537__;
  assign new_new_n33539__ = ~new_new_n33501__ & ~new_new_n33537__;
  assign new_new_n33540__ = ~new_new_n33538__ & ~new_new_n33539__;
  assign new_new_n33541__ = new_new_n33090__ & ~new_new_n33540__;
  assign new_new_n33542__ = ~new_new_n33090__ & new_new_n33540__;
  assign new_new_n33543__ = ~new_new_n33541__ & ~new_new_n33542__;
  assign new_new_n33544__ = new_new_n10702__ & new_new_n27250__;
  assign new_new_n33545__ = ~new_new_n11409__ & ~new_new_n27242__;
  assign new_new_n33546__ = new_new_n10697__ & ~new_new_n26698__;
  assign new_new_n33547__ = ~new_new_n10697__ & ~new_new_n31511__;
  assign new_new_n33548__ = new_new_n10694__ & ~new_new_n33546__;
  assign new_new_n33549__ = ~new_new_n33547__ & new_new_n33548__;
  assign new_new_n33550__ = ~new_new_n33544__ & ~new_new_n33545__;
  assign new_new_n33551__ = ~new_new_n33549__ & new_new_n33550__;
  assign new_new_n33552__ = ~new_new_n33543__ & new_new_n33551__;
  assign new_new_n33553__ = new_new_n33543__ & ~new_new_n33551__;
  assign new_new_n33554__ = ~new_new_n33283__ & ~new_new_n33552__;
  assign new_new_n33555__ = ~new_new_n33553__ & new_new_n33554__;
  assign new_new_n33556__ = ~pi08 & ~new_new_n33551__;
  assign new_new_n33557__ = pi08 & new_new_n33551__;
  assign new_new_n33558__ = ~new_new_n33556__ & ~new_new_n33557__;
  assign new_new_n33559__ = ~new_new_n33095__ & new_new_n33540__;
  assign new_new_n33560__ = ~new_new_n33280__ & ~new_new_n33540__;
  assign new_new_n33561__ = ~new_new_n33559__ & ~new_new_n33560__;
  assign new_new_n33562__ = ~new_new_n33282__ & ~new_new_n33558__;
  assign new_new_n33563__ = ~new_new_n33561__ & new_new_n33562__;
  assign new_new_n33564__ = ~new_new_n33281__ & new_new_n33558__;
  assign new_new_n33565__ = new_new_n33561__ & new_new_n33564__;
  assign new_new_n33566__ = ~new_new_n33563__ & ~new_new_n33565__;
  assign new_new_n33567__ = ~new_new_n33555__ & new_new_n33566__;
  assign new_new_n33568__ = new_new_n33356__ & ~new_new_n33567__;
  assign new_new_n33569__ = ~new_new_n33356__ & new_new_n33567__;
  assign new_new_n33570__ = ~new_new_n33568__ & ~new_new_n33569__;
  assign new_new_n33571__ = ~new_new_n33324__ & new_new_n33570__;
  assign new_new_n33572__ = new_new_n33324__ & ~new_new_n33570__;
  assign new_new_n33573__ = ~new_new_n33571__ & ~new_new_n33572__;
  assign new_new_n33574__ = ~new_new_n33322__ & new_new_n33573__;
  assign new_new_n33575__ = new_new_n33322__ & ~new_new_n33573__;
  assign new_new_n33576__ = ~new_new_n33574__ & ~new_new_n33575__;
  assign new_new_n33577__ = new_new_n33045__ & new_new_n33067__;
  assign new_new_n33578__ = ~new_new_n33576__ & ~new_new_n33577__;
  assign new_new_n33579__ = ~new_new_n33045__ & ~new_new_n33067__;
  assign new_new_n33580__ = new_new_n33576__ & ~new_new_n33579__;
  assign new_new_n33581__ = ~new_new_n33578__ & ~new_new_n33580__;
  assign new_new_n33582__ = new_new_n33065__ & new_new_n33581__;
  assign new_new_n33583__ = new_new_n33578__ & ~new_new_n33579__;
  assign new_new_n33584__ = new_new_n33576__ & ~new_new_n33577__;
  assign new_new_n33585__ = new_new_n33045__ & ~new_new_n33576__;
  assign new_new_n33586__ = ~new_new_n33065__ & ~new_new_n33584__;
  assign new_new_n33587__ = ~new_new_n33585__ & new_new_n33586__;
  assign new_new_n33588__ = ~new_new_n33583__ & ~new_new_n33587__;
  assign new_new_n33589__ = new_new_n33304__ & ~new_new_n33588__;
  assign new_new_n33590__ = new_new_n33065__ & new_new_n33584__;
  assign new_new_n33591__ = ~new_new_n33581__ & ~new_new_n33590__;
  assign new_new_n33592__ = ~new_new_n33304__ & ~new_new_n33591__;
  assign new_new_n33593__ = ~new_new_n33065__ & new_new_n33583__;
  assign new_new_n33594__ = ~new_new_n33582__ & ~new_new_n33593__;
  assign new_new_n33595__ = ~new_new_n33592__ & new_new_n33594__;
  assign po04 = new_new_n33589__ | ~new_new_n33595__;
  assign new_new_n33597__ = ~new_new_n33069__ & new_new_n33304__;
  assign new_new_n33598__ = new_new_n33576__ & new_new_n33597__;
  assign new_new_n33599__ = ~new_new_n33068__ & ~new_new_n33576__;
  assign new_new_n33600__ = new_new_n33045__ & ~new_new_n33305__;
  assign new_new_n33601__ = ~new_new_n33598__ & new_new_n33600__;
  assign new_new_n33602__ = ~new_new_n33599__ & new_new_n33601__;
  assign new_new_n33603__ = new_new_n14393__ & new_new_n32740__;
  assign new_new_n33604__ = pi02 & ~new_new_n33603__;
  assign new_new_n33605__ = ~new_new_n33602__ & ~new_new_n33604__;
  assign new_new_n33606__ = ~new_new_n33568__ & ~new_new_n33571__;
  assign new_new_n33607__ = new_new_n12832__ & ~new_new_n26667__;
  assign new_new_n33608__ = new_new_n11475__ & new_new_n32382__;
  assign new_new_n33609__ = ~new_new_n33607__ & ~new_new_n33608__;
  assign new_new_n33610__ = ~new_new_n11482__ & new_new_n32729__;
  assign new_new_n33611__ = new_new_n32758__ & new_new_n33610__;
  assign new_new_n33612__ = new_new_n33609__ & ~new_new_n33611__;
  assign new_new_n33613__ = pi05 & ~new_new_n33612__;
  assign new_new_n33614__ = ~new_new_n32729__ & ~new_new_n32758__;
  assign new_new_n33615__ = new_new_n11469__ & ~new_new_n33614__;
  assign new_new_n33616__ = ~pi05 & ~new_new_n33615__;
  assign new_new_n33617__ = ~new_new_n32729__ & new_new_n32758__;
  assign new_new_n33618__ = ~pi04 & ~new_new_n33617__;
  assign new_new_n33619__ = new_new_n32729__ & ~new_new_n32758__;
  assign new_new_n33620__ = pi04 & ~new_new_n33619__;
  assign new_new_n33621__ = ~new_new_n11482__ & ~new_new_n33618__;
  assign new_new_n33622__ = ~new_new_n33620__ & new_new_n33621__;
  assign new_new_n33623__ = ~new_new_n33616__ & ~new_new_n33622__;
  assign new_new_n33624__ = new_new_n33609__ & ~new_new_n33623__;
  assign new_new_n33625__ = ~new_new_n33613__ & ~new_new_n33624__;
  assign new_new_n33626__ = new_new_n11378__ & new_new_n27284__;
  assign new_new_n33627__ = ~new_new_n11409__ & new_new_n27250__;
  assign new_new_n33628__ = new_new_n10702__ & new_new_n26698__;
  assign new_new_n33629__ = new_new_n10698__ & ~new_new_n26674__;
  assign new_new_n33630__ = ~new_new_n33627__ & ~new_new_n33628__;
  assign new_new_n33631__ = ~new_new_n33629__ & new_new_n33630__;
  assign new_new_n33632__ = ~new_new_n33626__ & new_new_n33631__;
  assign new_new_n33633__ = pi08 & ~new_new_n33632__;
  assign new_new_n33634__ = ~pi08 & new_new_n33632__;
  assign new_new_n33635__ = ~new_new_n33633__ & ~new_new_n33634__;
  assign new_new_n33636__ = ~new_new_n33091__ & ~new_new_n33541__;
  assign new_new_n33637__ = ~new_new_n33551__ & new_new_n33636__;
  assign new_new_n33638__ = ~new_new_n33090__ & new_new_n33095__;
  assign new_new_n33639__ = pi08 & ~new_new_n33638__;
  assign new_new_n33640__ = ~new_new_n33542__ & ~new_new_n33639__;
  assign new_new_n33641__ = new_new_n33551__ & ~new_new_n33640__;
  assign new_new_n33642__ = ~new_new_n33540__ & ~new_new_n33556__;
  assign new_new_n33643__ = ~new_new_n33095__ & ~new_new_n33642__;
  assign new_new_n33644__ = ~new_new_n33637__ & ~new_new_n33643__;
  assign new_new_n33645__ = ~new_new_n33641__ & new_new_n33644__;
  assign new_new_n33646__ = new_new_n33280__ & ~new_new_n33645__;
  assign new_new_n33647__ = pi08 & new_new_n33540__;
  assign new_new_n33648__ = ~new_new_n33090__ & ~new_new_n33540__;
  assign new_new_n33649__ = ~new_new_n33092__ & ~new_new_n33095__;
  assign new_new_n33650__ = ~new_new_n33648__ & new_new_n33649__;
  assign new_new_n33651__ = ~new_new_n33647__ & ~new_new_n33650__;
  assign new_new_n33652__ = new_new_n33551__ & ~new_new_n33651__;
  assign new_new_n33653__ = ~pi08 & new_new_n33540__;
  assign new_new_n33654__ = ~new_new_n33095__ & new_new_n33636__;
  assign new_new_n33655__ = ~new_new_n33653__ & ~new_new_n33654__;
  assign new_new_n33656__ = ~new_new_n33551__ & ~new_new_n33655__;
  assign new_new_n33657__ = ~new_new_n33652__ & ~new_new_n33656__;
  assign new_new_n33658__ = ~new_new_n33646__ & new_new_n33657__;
  assign new_new_n33659__ = new_new_n8474__ & new_new_n26722__;
  assign new_new_n33660__ = ~new_new_n8479__ & new_new_n26729__;
  assign new_new_n33661__ = ~new_new_n8468__ & new_new_n27352__;
  assign new_new_n33662__ = new_new_n27242__ & ~new_new_n33661__;
  assign new_new_n33663__ = ~new_new_n27242__ & new_new_n33661__;
  assign new_new_n33664__ = new_new_n8469__ & ~new_new_n33662__;
  assign new_new_n33665__ = ~new_new_n33663__ & new_new_n33664__;
  assign new_new_n33666__ = ~new_new_n33659__ & ~new_new_n33660__;
  assign new_new_n33667__ = ~new_new_n33665__ & new_new_n33666__;
  assign new_new_n33668__ = ~pi11 & ~new_new_n33667__;
  assign new_new_n33669__ = pi11 & new_new_n33667__;
  assign new_new_n33670__ = ~new_new_n33668__ & ~new_new_n33669__;
  assign new_new_n33671__ = new_new_n33503__ & new_new_n33528__;
  assign new_new_n33672__ = ~new_new_n33503__ & ~new_new_n33528__;
  assign new_new_n33673__ = new_new_n33501__ & new_new_n33505__;
  assign new_new_n33674__ = ~new_new_n33501__ & ~new_new_n33505__;
  assign new_new_n33675__ = ~new_new_n33673__ & ~new_new_n33674__;
  assign new_new_n33676__ = ~new_new_n33516__ & ~new_new_n33675__;
  assign new_new_n33677__ = new_new_n33516__ & new_new_n33675__;
  assign new_new_n33678__ = ~new_new_n33676__ & ~new_new_n33677__;
  assign new_new_n33679__ = ~new_new_n33672__ & ~new_new_n33678__;
  assign new_new_n33680__ = ~new_new_n33671__ & ~new_new_n33679__;
  assign new_new_n33681__ = ~new_new_n33670__ & new_new_n33680__;
  assign new_new_n33682__ = new_new_n33670__ & ~new_new_n33680__;
  assign new_new_n33683__ = ~new_new_n33681__ & ~new_new_n33682__;
  assign new_new_n33684__ = new_new_n19825__ & new_new_n26810__;
  assign new_new_n33685__ = new_new_n19829__ & ~new_new_n26802__;
  assign new_new_n33686__ = ~new_new_n33684__ & ~new_new_n33685__;
  assign new_new_n33687__ = ~new_new_n6994__ & ~new_new_n33686__;
  assign new_new_n33688__ = new_new_n26774__ & ~new_new_n27373__;
  assign new_new_n33689__ = new_new_n6994__ & new_new_n33688__;
  assign new_new_n33690__ = ~new_new_n33687__ & ~new_new_n33689__;
  assign new_new_n33691__ = ~pi14 & ~new_new_n33690__;
  assign new_new_n33692__ = new_new_n26774__ & new_new_n27373__;
  assign new_new_n33693__ = ~pi13 & ~new_new_n33692__;
  assign new_new_n33694__ = ~new_new_n26774__ & ~new_new_n27373__;
  assign new_new_n33695__ = pi13 & ~new_new_n33694__;
  assign new_new_n33696__ = new_new_n6994__ & ~new_new_n33693__;
  assign new_new_n33697__ = ~new_new_n33695__ & new_new_n33696__;
  assign new_new_n33698__ = ~new_new_n26774__ & new_new_n27373__;
  assign new_new_n33699__ = new_new_n6994__ & ~new_new_n33698__;
  assign new_new_n33700__ = pi14 & ~new_new_n33687__;
  assign new_new_n33701__ = ~new_new_n33699__ & new_new_n33700__;
  assign new_new_n33702__ = ~new_new_n33691__ & ~new_new_n33701__;
  assign new_new_n33703__ = ~new_new_n33697__ & new_new_n33702__;
  assign new_new_n33704__ = ~new_new_n33371__ & ~new_new_n33498__;
  assign new_new_n33705__ = ~new_new_n33372__ & ~new_new_n33704__;
  assign new_new_n33706__ = new_new_n6968__ & ~new_new_n27221__;
  assign new_new_n33707__ = new_new_n6964__ & ~new_new_n26823__;
  assign new_new_n33708__ = new_new_n7935__ & ~new_new_n26741__;
  assign new_new_n33709__ = ~new_new_n33706__ & ~new_new_n33707__;
  assign new_new_n33710__ = ~new_new_n33708__ & new_new_n33709__;
  assign new_new_n33711__ = new_new_n6958__ & new_new_n30393__;
  assign new_new_n33712__ = ~pi17 & ~new_new_n33711__;
  assign new_new_n33713__ = new_new_n8160__ & new_new_n30393__;
  assign new_new_n33714__ = ~new_new_n33712__ & ~new_new_n33713__;
  assign new_new_n33715__ = new_new_n33710__ & ~new_new_n33714__;
  assign new_new_n33716__ = pi17 & ~new_new_n33710__;
  assign new_new_n33717__ = ~new_new_n33715__ & ~new_new_n33716__;
  assign new_new_n33718__ = new_new_n33705__ & ~new_new_n33717__;
  assign new_new_n33719__ = ~new_new_n33705__ & new_new_n33717__;
  assign new_new_n33720__ = ~new_new_n33718__ & ~new_new_n33719__;
  assign new_new_n33721__ = new_new_n6634__ & new_new_n26847__;
  assign new_new_n33722__ = ~new_new_n6625__ & ~new_new_n26888__;
  assign new_new_n33723__ = new_new_n6629__ & ~new_new_n26854__;
  assign new_new_n33724__ = new_new_n6936__ & new_new_n29424__;
  assign new_new_n33725__ = ~new_new_n33722__ & ~new_new_n33723__;
  assign new_new_n33726__ = ~new_new_n33721__ & new_new_n33725__;
  assign new_new_n33727__ = ~new_new_n33724__ & new_new_n33726__;
  assign new_new_n33728__ = ~pi20 & new_new_n33727__;
  assign new_new_n33729__ = pi20 & ~new_new_n33727__;
  assign new_new_n33730__ = ~new_new_n33728__ & ~new_new_n33729__;
  assign new_new_n33731__ = ~new_new_n33389__ & ~new_new_n33475__;
  assign new_new_n33732__ = new_new_n5213__ & new_new_n26922__;
  assign new_new_n33733__ = new_new_n5183__ & ~new_new_n27168__;
  assign new_new_n33734__ = new_new_n5191__ & new_new_n26917__;
  assign new_new_n33735__ = new_new_n5215__ & ~new_new_n29366__;
  assign new_new_n33736__ = ~new_new_n33733__ & ~new_new_n33734__;
  assign new_new_n33737__ = ~new_new_n33732__ & new_new_n33736__;
  assign new_new_n33738__ = ~new_new_n33735__ & new_new_n33737__;
  assign new_new_n33739__ = new_new_n33731__ & ~new_new_n33738__;
  assign new_new_n33740__ = ~new_new_n33731__ & new_new_n33738__;
  assign new_new_n33741__ = ~new_new_n33739__ & ~new_new_n33740__;
  assign new_new_n33742__ = ~new_new_n333__ & new_new_n27152__;
  assign new_new_n33743__ = new_new_n873__ & ~new_new_n26941__;
  assign new_new_n33744__ = new_new_n3311__ & new_new_n26928__;
  assign new_new_n33745__ = ~new_new_n33742__ & ~new_new_n33743__;
  assign new_new_n33746__ = ~new_new_n33744__ & new_new_n33745__;
  assign new_new_n33747__ = ~pi26 & ~new_new_n33746__;
  assign new_new_n33748__ = new_new_n512__ & new_new_n27488__;
  assign new_new_n33749__ = new_new_n801__ & new_new_n27488__;
  assign new_new_n33750__ = pi26 & ~new_new_n33749__;
  assign new_new_n33751__ = ~new_new_n33748__ & ~new_new_n33750__;
  assign new_new_n33752__ = new_new_n33746__ & ~new_new_n33751__;
  assign new_new_n33753__ = ~new_new_n33747__ & ~new_new_n33752__;
  assign new_new_n33754__ = new_new_n4815__ & ~new_new_n26937__;
  assign new_new_n33755__ = new_new_n4212__ & new_new_n26971__;
  assign new_new_n33756__ = ~new_new_n4818__ & ~new_new_n26978__;
  assign new_new_n33757__ = new_new_n4813__ & new_new_n28005__;
  assign new_new_n33758__ = ~new_new_n33755__ & ~new_new_n33756__;
  assign new_new_n33759__ = ~new_new_n33754__ & new_new_n33758__;
  assign new_new_n33760__ = ~new_new_n33757__ & new_new_n33759__;
  assign new_new_n33761__ = new_new_n27021__ & ~new_new_n27764__;
  assign new_new_n33762__ = new_new_n27029__ & new_new_n27762__;
  assign new_new_n33763__ = ~new_new_n33761__ & ~new_new_n33762__;
  assign new_new_n33764__ = new_new_n765__ & ~new_new_n33763__;
  assign new_new_n33765__ = ~new_new_n27118__ & ~new_new_n33764__;
  assign new_new_n33766__ = ~new_new_n27003__ & ~new_new_n33765__;
  assign new_new_n33767__ = new_new_n27003__ & new_new_n27763__;
  assign new_new_n33768__ = ~new_new_n161__ & ~new_new_n33767__;
  assign new_new_n33769__ = new_new_n33158__ & ~new_new_n33768__;
  assign new_new_n33770__ = ~new_new_n71__ & ~new_new_n28270__;
  assign new_new_n33771__ = ~new_new_n27029__ & new_new_n33159__;
  assign new_new_n33772__ = ~new_new_n33770__ & new_new_n33771__;
  assign new_new_n33773__ = ~new_new_n33769__ & ~new_new_n33772__;
  assign new_new_n33774__ = ~new_new_n33766__ & new_new_n33773__;
  assign new_new_n33775__ = pi31 & ~new_new_n33774__;
  assign new_new_n33776__ = ~new_new_n71__ & ~new_new_n27003__;
  assign new_new_n33777__ = ~new_new_n161__ & ~new_new_n33776__;
  assign new_new_n33778__ = new_new_n161__ & new_new_n27029__;
  assign new_new_n33779__ = ~pi31 & ~new_new_n33778__;
  assign new_new_n33780__ = ~new_new_n33777__ & new_new_n33779__;
  assign new_new_n33781__ = ~new_new_n33775__ & ~new_new_n33780__;
  assign new_new_n33782__ = new_new_n33401__ & ~new_new_n33440__;
  assign new_new_n33783__ = ~new_new_n33441__ & ~new_new_n33782__;
  assign new_new_n33784__ = ~new_new_n33781__ & new_new_n33783__;
  assign new_new_n33785__ = new_new_n33781__ & ~new_new_n33783__;
  assign new_new_n33786__ = ~new_new_n33784__ & ~new_new_n33785__;
  assign new_new_n33787__ = ~new_new_n96__ & ~new_new_n208__;
  assign new_new_n33788__ = ~new_new_n472__ & ~new_new_n749__;
  assign new_new_n33789__ = ~new_new_n1031__ & new_new_n33788__;
  assign new_new_n33790__ = new_new_n121__ & new_new_n33787__;
  assign new_new_n33791__ = new_new_n623__ & ~new_new_n842__;
  assign new_new_n33792__ = ~new_new_n1073__ & new_new_n5287__;
  assign new_new_n33793__ = new_new_n33791__ & new_new_n33792__;
  assign new_new_n33794__ = new_new_n33789__ & new_new_n33790__;
  assign new_new_n33795__ = new_new_n2385__ & new_new_n2539__;
  assign new_new_n33796__ = new_new_n33794__ & new_new_n33795__;
  assign new_new_n33797__ = new_new_n33793__ & new_new_n33796__;
  assign new_new_n33798__ = new_new_n714__ & new_new_n4600__;
  assign new_new_n33799__ = new_new_n33797__ & new_new_n33798__;
  assign new_new_n33800__ = new_new_n4464__ & new_new_n33799__;
  assign new_new_n33801__ = new_new_n6181__ & new_new_n33800__;
  assign new_new_n33802__ = new_new_n19340__ & new_new_n33801__;
  assign new_new_n33803__ = ~new_new_n33786__ & new_new_n33802__;
  assign new_new_n33804__ = new_new_n33786__ & ~new_new_n33802__;
  assign new_new_n33805__ = ~new_new_n33803__ & ~new_new_n33804__;
  assign new_new_n33806__ = ~new_new_n33456__ & new_new_n33462__;
  assign new_new_n33807__ = ~new_new_n33464__ & ~new_new_n33806__;
  assign new_new_n33808__ = pi29 & ~new_new_n33807__;
  assign new_new_n33809__ = ~pi29 & new_new_n33807__;
  assign new_new_n33810__ = ~new_new_n33808__ & ~new_new_n33809__;
  assign new_new_n33811__ = new_new_n33805__ & ~new_new_n33810__;
  assign new_new_n33812__ = ~new_new_n33805__ & new_new_n33810__;
  assign new_new_n33813__ = ~new_new_n33811__ & ~new_new_n33812__;
  assign new_new_n33814__ = new_new_n33760__ & new_new_n33813__;
  assign new_new_n33815__ = ~new_new_n33760__ & ~new_new_n33813__;
  assign new_new_n33816__ = ~new_new_n33814__ & ~new_new_n33815__;
  assign new_new_n33817__ = pi23 & ~new_new_n33816__;
  assign new_new_n33818__ = ~pi23 & new_new_n33816__;
  assign new_new_n33819__ = ~new_new_n33817__ & ~new_new_n33818__;
  assign new_new_n33820__ = new_new_n33753__ & new_new_n33819__;
  assign new_new_n33821__ = ~new_new_n33753__ & ~new_new_n33819__;
  assign new_new_n33822__ = ~new_new_n33820__ & ~new_new_n33821__;
  assign new_new_n33823__ = new_new_n33399__ & ~new_new_n33465__;
  assign new_new_n33824__ = ~new_new_n33474__ & ~new_new_n33823__;
  assign new_new_n33825__ = ~new_new_n33399__ & new_new_n33465__;
  assign new_new_n33826__ = ~new_new_n33824__ & ~new_new_n33825__;
  assign new_new_n33827__ = new_new_n33822__ & ~new_new_n33826__;
  assign new_new_n33828__ = ~new_new_n33822__ & new_new_n33826__;
  assign new_new_n33829__ = ~new_new_n33827__ & ~new_new_n33828__;
  assign new_new_n33830__ = new_new_n33741__ & new_new_n33829__;
  assign new_new_n33831__ = ~new_new_n33741__ & ~new_new_n33829__;
  assign new_new_n33832__ = ~new_new_n33830__ & ~new_new_n33831__;
  assign new_new_n33833__ = ~new_new_n33481__ & new_new_n33495__;
  assign new_new_n33834__ = ~new_new_n33480__ & ~new_new_n33833__;
  assign new_new_n33835__ = new_new_n33832__ & ~new_new_n33834__;
  assign new_new_n33836__ = ~new_new_n33832__ & new_new_n33834__;
  assign new_new_n33837__ = ~new_new_n33835__ & ~new_new_n33836__;
  assign new_new_n33838__ = new_new_n33730__ & ~new_new_n33837__;
  assign new_new_n33839__ = ~new_new_n33730__ & new_new_n33837__;
  assign new_new_n33840__ = ~new_new_n33838__ & ~new_new_n33839__;
  assign new_new_n33841__ = new_new_n33720__ & ~new_new_n33840__;
  assign new_new_n33842__ = ~new_new_n33720__ & new_new_n33840__;
  assign new_new_n33843__ = ~new_new_n33841__ & ~new_new_n33842__;
  assign new_new_n33844__ = ~new_new_n33516__ & ~new_new_n33673__;
  assign new_new_n33845__ = ~new_new_n33674__ & ~new_new_n33844__;
  assign new_new_n33846__ = ~new_new_n33843__ & new_new_n33845__;
  assign new_new_n33847__ = new_new_n33843__ & ~new_new_n33845__;
  assign new_new_n33848__ = ~new_new_n33846__ & ~new_new_n33847__;
  assign new_new_n33849__ = new_new_n33703__ & new_new_n33848__;
  assign new_new_n33850__ = ~new_new_n33703__ & ~new_new_n33848__;
  assign new_new_n33851__ = ~new_new_n33849__ & ~new_new_n33850__;
  assign new_new_n33852__ = new_new_n33683__ & new_new_n33851__;
  assign new_new_n33853__ = ~new_new_n33683__ & ~new_new_n33851__;
  assign new_new_n33854__ = ~new_new_n33852__ & ~new_new_n33853__;
  assign new_new_n33855__ = ~new_new_n33658__ & ~new_new_n33854__;
  assign new_new_n33856__ = new_new_n33658__ & new_new_n33854__;
  assign new_new_n33857__ = ~new_new_n33855__ & ~new_new_n33856__;
  assign new_new_n33858__ = new_new_n33635__ & ~new_new_n33857__;
  assign new_new_n33859__ = ~new_new_n33635__ & new_new_n33857__;
  assign new_new_n33860__ = ~new_new_n33858__ & ~new_new_n33859__;
  assign new_new_n33861__ = ~new_new_n33625__ & new_new_n33860__;
  assign new_new_n33862__ = new_new_n33625__ & ~new_new_n33860__;
  assign new_new_n33863__ = ~new_new_n33861__ & ~new_new_n33862__;
  assign new_new_n33864__ = ~new_new_n33606__ & ~new_new_n33863__;
  assign new_new_n33865__ = new_new_n33606__ & new_new_n33863__;
  assign new_new_n33866__ = ~new_new_n33864__ & ~new_new_n33865__;
  assign new_new_n33867__ = ~new_new_n33605__ & new_new_n33866__;
  assign new_new_n33868__ = new_new_n33605__ & ~new_new_n33866__;
  assign new_new_n33869__ = ~new_new_n33867__ & ~new_new_n33868__;
  assign new_new_n33870__ = ~new_new_n33068__ & ~new_new_n33597__;
  assign new_new_n33871__ = ~new_new_n33574__ & new_new_n33870__;
  assign new_new_n33872__ = ~new_new_n33575__ & ~new_new_n33871__;
  assign new_new_n33873__ = ~new_new_n33602__ & ~new_new_n33872__;
  assign new_new_n33874__ = ~new_new_n33604__ & ~new_new_n33872__;
  assign new_new_n33875__ = ~new_new_n33873__ & ~new_new_n33874__;
  assign new_new_n33876__ = new_new_n33869__ & new_new_n33875__;
  assign new_new_n33877__ = ~new_new_n33869__ & ~new_new_n33875__;
  assign po05 = new_new_n33876__ | new_new_n33877__;
  assign new_new_n33879__ = new_new_n12850__ & new_new_n32740__;
  assign new_new_n33880__ = new_new_n13069__ & new_new_n33050__;
  assign new_new_n33881__ = new_new_n12832__ & new_new_n32382__;
  assign new_new_n33882__ = new_new_n11475__ & new_new_n32729__;
  assign new_new_n33883__ = ~new_new_n33881__ & ~new_new_n33882__;
  assign new_new_n33884__ = ~new_new_n33879__ & new_new_n33883__;
  assign new_new_n33885__ = ~new_new_n33880__ & new_new_n33884__;
  assign new_new_n33886__ = pi02 & ~new_new_n33885__;
  assign new_new_n33887__ = ~pi02 & new_new_n33885__;
  assign new_new_n33888__ = ~new_new_n33886__ & ~new_new_n33887__;
  assign new_new_n33889__ = new_new_n10698__ & ~new_new_n26667__;
  assign new_new_n33890__ = new_new_n10702__ & ~new_new_n26674__;
  assign new_new_n33891__ = ~new_new_n11409__ & new_new_n26698__;
  assign new_new_n33892__ = new_new_n11378__ & ~new_new_n32340__;
  assign new_new_n33893__ = ~new_new_n33890__ & ~new_new_n33891__;
  assign new_new_n33894__ = ~new_new_n33889__ & new_new_n33893__;
  assign new_new_n33895__ = ~new_new_n33892__ & new_new_n33894__;
  assign new_new_n33896__ = pi08 & ~new_new_n33895__;
  assign new_new_n33897__ = ~pi08 & new_new_n33895__;
  assign new_new_n33898__ = ~new_new_n33896__ & ~new_new_n33897__;
  assign new_new_n33899__ = new_new_n33635__ & ~new_new_n33856__;
  assign new_new_n33900__ = ~new_new_n33855__ & ~new_new_n33899__;
  assign new_new_n33901__ = ~new_new_n33898__ & new_new_n33900__;
  assign new_new_n33902__ = new_new_n33898__ & ~new_new_n33900__;
  assign new_new_n33903__ = ~new_new_n33901__ & ~new_new_n33902__;
  assign new_new_n33904__ = new_new_n8858__ & new_new_n27250__;
  assign new_new_n33905__ = new_new_n8474__ & ~new_new_n27242__;
  assign new_new_n33906__ = ~new_new_n8479__ & new_new_n26722__;
  assign new_new_n33907__ = new_new_n8470__ & ~new_new_n27271__;
  assign new_new_n33908__ = ~new_new_n33905__ & ~new_new_n33906__;
  assign new_new_n33909__ = ~new_new_n33904__ & new_new_n33908__;
  assign new_new_n33910__ = ~new_new_n33907__ & new_new_n33909__;
  assign new_new_n33911__ = pi11 & ~new_new_n33910__;
  assign new_new_n33912__ = ~pi11 & new_new_n33910__;
  assign new_new_n33913__ = ~new_new_n33911__ & ~new_new_n33912__;
  assign new_new_n33914__ = new_new_n19825__ & new_new_n26774__;
  assign new_new_n33915__ = new_new_n19829__ & new_new_n26810__;
  assign new_new_n33916__ = ~new_new_n6994__ & ~new_new_n33915__;
  assign new_new_n33917__ = ~new_new_n33914__ & new_new_n33916__;
  assign new_new_n33918__ = ~new_new_n26729__ & ~new_new_n30644__;
  assign new_new_n33919__ = new_new_n6994__ & new_new_n33918__;
  assign new_new_n33920__ = ~new_new_n33917__ & ~new_new_n33919__;
  assign new_new_n33921__ = ~pi14 & ~new_new_n33920__;
  assign new_new_n33922__ = new_new_n26729__ & ~new_new_n30643__;
  assign new_new_n33923__ = pi13 & ~new_new_n33922__;
  assign new_new_n33924__ = ~new_new_n26729__ & new_new_n30644__;
  assign new_new_n33925__ = ~pi13 & ~new_new_n33924__;
  assign new_new_n33926__ = new_new_n6994__ & ~new_new_n33923__;
  assign new_new_n33927__ = ~new_new_n33925__ & new_new_n33926__;
  assign new_new_n33928__ = new_new_n6994__ & ~new_new_n30644__;
  assign new_new_n33929__ = new_new_n6994__ & ~new_new_n26729__;
  assign new_new_n33930__ = pi14 & ~new_new_n33929__;
  assign new_new_n33931__ = ~new_new_n33917__ & new_new_n33930__;
  assign new_new_n33932__ = ~new_new_n33928__ & new_new_n33931__;
  assign new_new_n33933__ = ~new_new_n33927__ & ~new_new_n33932__;
  assign new_new_n33934__ = ~new_new_n33921__ & new_new_n33933__;
  assign new_new_n33935__ = ~new_new_n33703__ & ~new_new_n33847__;
  assign new_new_n33936__ = ~new_new_n33846__ & ~new_new_n33935__;
  assign new_new_n33937__ = new_new_n6964__ & ~new_new_n27221__;
  assign new_new_n33938__ = new_new_n6968__ & ~new_new_n26741__;
  assign new_new_n33939__ = ~new_new_n33937__ & ~new_new_n33938__;
  assign new_new_n33940__ = new_new_n6958__ & ~new_new_n26802__;
  assign new_new_n33941__ = new_new_n30411__ & new_new_n33940__;
  assign new_new_n33942__ = new_new_n33939__ & ~new_new_n33941__;
  assign new_new_n33943__ = pi17 & ~new_new_n33942__;
  assign new_new_n33944__ = new_new_n6958__ & ~new_new_n27391__;
  assign new_new_n33945__ = ~pi17 & ~new_new_n33944__;
  assign new_new_n33946__ = ~pi16 & ~new_new_n30692__;
  assign new_new_n33947__ = pi16 & ~new_new_n30410__;
  assign new_new_n33948__ = new_new_n6958__ & ~new_new_n33946__;
  assign new_new_n33949__ = ~new_new_n33947__ & new_new_n33948__;
  assign new_new_n33950__ = ~new_new_n33945__ & ~new_new_n33949__;
  assign new_new_n33951__ = new_new_n33939__ & ~new_new_n33950__;
  assign new_new_n33952__ = ~new_new_n33943__ & ~new_new_n33951__;
  assign new_new_n33953__ = new_new_n33832__ & new_new_n33834__;
  assign new_new_n33954__ = ~new_new_n33832__ & ~new_new_n33834__;
  assign new_new_n33955__ = pi23 & ~new_new_n33738__;
  assign new_new_n33956__ = ~pi23 & new_new_n33738__;
  assign new_new_n33957__ = ~new_new_n33955__ & ~new_new_n33956__;
  assign new_new_n33958__ = ~new_new_n33731__ & ~new_new_n33957__;
  assign new_new_n33959__ = new_new_n33731__ & new_new_n33957__;
  assign new_new_n33960__ = ~new_new_n33816__ & new_new_n33826__;
  assign new_new_n33961__ = new_new_n33816__ & ~new_new_n33826__;
  assign new_new_n33962__ = ~new_new_n33960__ & ~new_new_n33961__;
  assign new_new_n33963__ = new_new_n33753__ & ~new_new_n33962__;
  assign new_new_n33964__ = ~new_new_n33753__ & new_new_n33962__;
  assign new_new_n33965__ = ~new_new_n33963__ & ~new_new_n33964__;
  assign new_new_n33966__ = ~new_new_n33959__ & ~new_new_n33965__;
  assign new_new_n33967__ = ~new_new_n33958__ & ~new_new_n33966__;
  assign new_new_n33968__ = ~new_new_n33753__ & ~new_new_n33960__;
  assign new_new_n33969__ = ~new_new_n33961__ & ~new_new_n33968__;
  assign new_new_n33970__ = ~new_new_n33727__ & new_new_n33969__;
  assign new_new_n33971__ = new_new_n33727__ & ~new_new_n33969__;
  assign new_new_n33972__ = ~new_new_n33970__ & ~new_new_n33971__;
  assign new_new_n33973__ = new_new_n33967__ & new_new_n33972__;
  assign new_new_n33974__ = ~new_new_n33967__ & ~new_new_n33972__;
  assign new_new_n33975__ = ~new_new_n33973__ & ~new_new_n33974__;
  assign new_new_n33976__ = ~new_new_n33953__ & new_new_n33975__;
  assign new_new_n33977__ = ~new_new_n33954__ & new_new_n33976__;
  assign new_new_n33978__ = pi20 & ~new_new_n33969__;
  assign new_new_n33979__ = ~pi20 & new_new_n33969__;
  assign new_new_n33980__ = ~new_new_n33978__ & ~new_new_n33979__;
  assign new_new_n33981__ = ~new_new_n33954__ & ~new_new_n33967__;
  assign new_new_n33982__ = ~new_new_n33953__ & new_new_n33967__;
  assign new_new_n33983__ = ~new_new_n33980__ & ~new_new_n33981__;
  assign new_new_n33984__ = ~new_new_n33982__ & new_new_n33983__;
  assign new_new_n33985__ = ~new_new_n33954__ & new_new_n33967__;
  assign new_new_n33986__ = ~new_new_n33953__ & ~new_new_n33967__;
  assign new_new_n33987__ = new_new_n33980__ & ~new_new_n33985__;
  assign new_new_n33988__ = ~new_new_n33986__ & new_new_n33987__;
  assign new_new_n33989__ = ~new_new_n33977__ & ~new_new_n33984__;
  assign new_new_n33990__ = ~new_new_n33988__ & new_new_n33989__;
  assign new_new_n33991__ = ~new_new_n4818__ & new_new_n26971__;
  assign new_new_n33992__ = new_new_n4212__ & ~new_new_n26937__;
  assign new_new_n33993__ = ~new_new_n4215__ & new_new_n28666__;
  assign new_new_n33994__ = new_new_n4215__ & ~new_new_n27152__;
  assign new_new_n33995__ = new_new_n4214__ & ~new_new_n33994__;
  assign new_new_n33996__ = ~new_new_n33993__ & new_new_n33995__;
  assign new_new_n33997__ = ~new_new_n33991__ & ~new_new_n33992__;
  assign new_new_n33998__ = ~new_new_n33996__ & new_new_n33997__;
  assign new_new_n33999__ = ~new_new_n723__ & ~new_new_n1176__;
  assign new_new_n34000__ = ~new_new_n155__ & new_new_n33999__;
  assign new_new_n34001__ = ~new_new_n939__ & new_new_n34000__;
  assign new_new_n34002__ = new_new_n1310__ & new_new_n6235__;
  assign new_new_n34003__ = new_new_n34001__ & new_new_n34002__;
  assign new_new_n34004__ = new_new_n5312__ & new_new_n34003__;
  assign new_new_n34005__ = ~new_new_n277__ & new_new_n1423__;
  assign new_new_n34006__ = ~new_new_n6184__ & new_new_n34005__;
  assign new_new_n34007__ = new_new_n872__ & new_new_n1164__;
  assign new_new_n34008__ = new_new_n1516__ & new_new_n18149__;
  assign new_new_n34009__ = new_new_n34007__ & new_new_n34008__;
  assign new_new_n34010__ = new_new_n7111__ & new_new_n34006__;
  assign new_new_n34011__ = new_new_n19383__ & new_new_n34010__;
  assign new_new_n34012__ = new_new_n17505__ & new_new_n34009__;
  assign new_new_n34013__ = new_new_n33169__ & new_new_n34012__;
  assign new_new_n34014__ = new_new_n34004__ & new_new_n34011__;
  assign new_new_n34015__ = new_new_n34013__ & new_new_n34014__;
  assign new_new_n34016__ = new_new_n18158__ & new_new_n34015__;
  assign new_new_n34017__ = new_new_n6295__ & new_new_n32491__;
  assign new_new_n34018__ = new_new_n34016__ & new_new_n34017__;
  assign new_new_n34019__ = new_new_n71__ & new_new_n27003__;
  assign new_new_n34020__ = new_new_n765__ & ~new_new_n27986__;
  assign new_new_n34021__ = ~new_new_n33778__ & ~new_new_n34020__;
  assign new_new_n34022__ = pi31 & ~new_new_n34021__;
  assign new_new_n34023__ = new_new_n161__ & new_new_n27003__;
  assign new_new_n34024__ = ~new_new_n161__ & new_new_n26978__;
  assign new_new_n34025__ = ~new_new_n71__ & ~new_new_n34023__;
  assign new_new_n34026__ = ~new_new_n34024__ & new_new_n34025__;
  assign new_new_n34027__ = ~pi31 & ~new_new_n34026__;
  assign new_new_n34028__ = ~new_new_n34019__ & ~new_new_n34027__;
  assign new_new_n34029__ = ~new_new_n34022__ & new_new_n34028__;
  assign new_new_n34030__ = new_new_n34018__ & ~new_new_n34029__;
  assign new_new_n34031__ = ~new_new_n34018__ & new_new_n34029__;
  assign new_new_n34032__ = ~new_new_n34030__ & ~new_new_n34031__;
  assign new_new_n34033__ = ~new_new_n33784__ & new_new_n33802__;
  assign new_new_n34034__ = ~new_new_n33785__ & ~new_new_n34033__;
  assign new_new_n34035__ = new_new_n34032__ & new_new_n34034__;
  assign new_new_n34036__ = ~new_new_n34032__ & ~new_new_n34034__;
  assign new_new_n34037__ = ~new_new_n34035__ & ~new_new_n34036__;
  assign new_new_n34038__ = new_new_n33807__ & new_new_n33816__;
  assign new_new_n34039__ = ~new_new_n33807__ & ~new_new_n33816__;
  assign new_new_n34040__ = ~new_new_n33805__ & ~new_new_n34039__;
  assign new_new_n34041__ = ~new_new_n34038__ & ~new_new_n34040__;
  assign new_new_n34042__ = new_new_n34037__ & new_new_n34041__;
  assign new_new_n34043__ = ~new_new_n34037__ & ~new_new_n34041__;
  assign new_new_n34044__ = ~new_new_n34042__ & ~new_new_n34043__;
  assign new_new_n34045__ = pi29 & ~new_new_n34044__;
  assign new_new_n34046__ = ~pi29 & new_new_n34044__;
  assign new_new_n34047__ = ~new_new_n34045__ & ~new_new_n34046__;
  assign new_new_n34048__ = new_new_n33998__ & new_new_n34047__;
  assign new_new_n34049__ = ~new_new_n33998__ & ~new_new_n34047__;
  assign new_new_n34050__ = ~new_new_n34048__ & ~new_new_n34049__;
  assign new_new_n34051__ = new_new_n33990__ & ~new_new_n34050__;
  assign new_new_n34052__ = ~new_new_n33990__ & new_new_n34050__;
  assign new_new_n34053__ = ~new_new_n34051__ & ~new_new_n34052__;
  assign new_new_n34054__ = new_new_n3311__ & new_new_n26917__;
  assign new_new_n34055__ = ~new_new_n333__ & ~new_new_n26941__;
  assign new_new_n34056__ = new_new_n873__ & new_new_n26928__;
  assign new_new_n34057__ = ~new_new_n34055__ & ~new_new_n34056__;
  assign new_new_n34058__ = ~new_new_n34054__ & new_new_n34057__;
  assign new_new_n34059__ = ~pi26 & ~new_new_n34058__;
  assign new_new_n34060__ = new_new_n512__ & ~new_new_n27462__;
  assign new_new_n34061__ = new_new_n801__ & ~new_new_n27462__;
  assign new_new_n34062__ = pi26 & ~new_new_n34061__;
  assign new_new_n34063__ = ~new_new_n34060__ & ~new_new_n34062__;
  assign new_new_n34064__ = new_new_n34058__ & ~new_new_n34063__;
  assign new_new_n34065__ = ~new_new_n34059__ & ~new_new_n34064__;
  assign new_new_n34066__ = new_new_n5215__ & new_new_n27180__;
  assign new_new_n34067__ = new_new_n5191__ & ~new_new_n27168__;
  assign new_new_n34068__ = new_new_n5183__ & new_new_n26922__;
  assign new_new_n34069__ = ~new_new_n34067__ & ~new_new_n34068__;
  assign new_new_n34070__ = ~new_new_n34066__ & new_new_n34069__;
  assign new_new_n34071__ = new_new_n5195__ & ~new_new_n26888__;
  assign new_new_n34072__ = pi23 & ~new_new_n34071__;
  assign new_new_n34073__ = new_new_n5974__ & ~new_new_n26888__;
  assign new_new_n34074__ = ~new_new_n34072__ & ~new_new_n34073__;
  assign new_new_n34075__ = new_new_n34070__ & ~new_new_n34074__;
  assign new_new_n34076__ = ~pi23 & ~new_new_n34070__;
  assign new_new_n34077__ = ~new_new_n34075__ & ~new_new_n34076__;
  assign new_new_n34078__ = ~new_new_n34065__ & new_new_n34077__;
  assign new_new_n34079__ = new_new_n34065__ & ~new_new_n34077__;
  assign new_new_n34080__ = ~new_new_n34078__ & ~new_new_n34079__;
  assign new_new_n34081__ = new_new_n6936__ & ~new_new_n29400__;
  assign new_new_n34082__ = new_new_n6629__ & new_new_n26847__;
  assign new_new_n34083__ = ~new_new_n6625__ & ~new_new_n26854__;
  assign new_new_n34084__ = new_new_n6634__ & ~new_new_n26823__;
  assign new_new_n34085__ = ~new_new_n34082__ & ~new_new_n34083__;
  assign new_new_n34086__ = ~new_new_n34084__ & new_new_n34085__;
  assign new_new_n34087__ = ~new_new_n34081__ & new_new_n34086__;
  assign new_new_n34088__ = new_new_n34080__ & ~new_new_n34087__;
  assign new_new_n34089__ = ~new_new_n34080__ & new_new_n34087__;
  assign new_new_n34090__ = ~new_new_n34088__ & ~new_new_n34089__;
  assign new_new_n34091__ = new_new_n34053__ & new_new_n34090__;
  assign new_new_n34092__ = ~new_new_n34053__ & ~new_new_n34090__;
  assign new_new_n34093__ = ~new_new_n34091__ & ~new_new_n34092__;
  assign new_new_n34094__ = ~new_new_n33718__ & new_new_n33840__;
  assign new_new_n34095__ = ~new_new_n33719__ & ~new_new_n34094__;
  assign new_new_n34096__ = ~new_new_n34093__ & new_new_n34095__;
  assign new_new_n34097__ = new_new_n34093__ & ~new_new_n34095__;
  assign new_new_n34098__ = ~new_new_n34096__ & ~new_new_n34097__;
  assign new_new_n34099__ = new_new_n33952__ & ~new_new_n34098__;
  assign new_new_n34100__ = ~new_new_n33952__ & new_new_n34098__;
  assign new_new_n34101__ = ~new_new_n34099__ & ~new_new_n34100__;
  assign new_new_n34102__ = ~new_new_n33936__ & ~new_new_n34101__;
  assign new_new_n34103__ = new_new_n33936__ & new_new_n34101__;
  assign new_new_n34104__ = ~new_new_n34102__ & ~new_new_n34103__;
  assign new_new_n34105__ = new_new_n33934__ & new_new_n34104__;
  assign new_new_n34106__ = ~new_new_n33934__ & ~new_new_n34104__;
  assign new_new_n34107__ = ~new_new_n34105__ & ~new_new_n34106__;
  assign new_new_n34108__ = ~new_new_n33682__ & ~new_new_n33851__;
  assign new_new_n34109__ = ~new_new_n33681__ & ~new_new_n34108__;
  assign new_new_n34110__ = new_new_n34107__ & ~new_new_n34109__;
  assign new_new_n34111__ = ~new_new_n34107__ & new_new_n34109__;
  assign new_new_n34112__ = ~new_new_n34110__ & ~new_new_n34111__;
  assign new_new_n34113__ = new_new_n33913__ & new_new_n34112__;
  assign new_new_n34114__ = ~new_new_n33913__ & ~new_new_n34112__;
  assign new_new_n34115__ = ~new_new_n34113__ & ~new_new_n34114__;
  assign new_new_n34116__ = new_new_n33903__ & new_new_n34115__;
  assign new_new_n34117__ = ~new_new_n33903__ & ~new_new_n34115__;
  assign new_new_n34118__ = ~new_new_n34116__ & ~new_new_n34117__;
  assign new_new_n34119__ = pi05 & new_new_n34118__;
  assign new_new_n34120__ = ~pi05 & ~new_new_n34118__;
  assign new_new_n34121__ = ~new_new_n34119__ & ~new_new_n34120__;
  assign new_new_n34122__ = pi02 & ~new_new_n33883__;
  assign new_new_n34123__ = new_new_n33888__ & ~new_new_n34122__;
  assign new_new_n34124__ = new_new_n34121__ & new_new_n34123__;
  assign new_new_n34125__ = ~new_new_n33888__ & ~new_new_n34121__;
  assign new_new_n34126__ = ~new_new_n34124__ & ~new_new_n34125__;
  assign new_new_n34127__ = ~new_new_n33862__ & ~new_new_n34126__;
  assign new_new_n34128__ = ~new_new_n33606__ & ~new_new_n33861__;
  assign new_new_n34129__ = new_new_n34127__ & ~new_new_n34128__;
  assign new_new_n34130__ = ~new_new_n33861__ & new_new_n34126__;
  assign new_new_n34131__ = new_new_n33606__ & ~new_new_n33862__;
  assign new_new_n34132__ = new_new_n34130__ & ~new_new_n34131__;
  assign new_new_n34133__ = ~new_new_n34129__ & ~new_new_n34132__;
  assign new_new_n34134__ = ~new_new_n33866__ & ~new_new_n33874__;
  assign new_new_n34135__ = ~new_new_n33873__ & ~po05;
  assign new_new_n34136__ = ~new_new_n34134__ & ~new_new_n34135__;
  assign new_new_n34137__ = ~new_new_n34133__ & ~new_new_n34136__;
  assign new_new_n34138__ = new_new_n33602__ & ~po05;
  assign new_new_n34139__ = new_new_n33866__ & ~new_new_n33872__;
  assign new_new_n34140__ = new_new_n33605__ & po05;
  assign new_new_n34141__ = ~new_new_n34139__ & ~new_new_n34140__;
  assign new_new_n34142__ = new_new_n34133__ & ~new_new_n34138__;
  assign new_new_n34143__ = ~new_new_n34141__ & new_new_n34142__;
  assign po06 = new_new_n34137__ | new_new_n34143__;
  assign new_new_n34145__ = new_new_n33604__ & ~new_new_n33861__;
  assign new_new_n34146__ = ~new_new_n33862__ & ~new_new_n34145__;
  assign new_new_n34147__ = new_new_n34126__ & ~new_new_n34146__;
  assign new_new_n34148__ = ~new_new_n34126__ & new_new_n34146__;
  assign new_new_n34149__ = ~new_new_n33606__ & new_new_n33872__;
  assign new_new_n34150__ = ~new_new_n34148__ & new_new_n34149__;
  assign new_new_n34151__ = new_new_n33606__ & ~new_new_n33872__;
  assign new_new_n34152__ = ~new_new_n33604__ & ~new_new_n34130__;
  assign new_new_n34153__ = ~new_new_n34127__ & ~new_new_n34151__;
  assign new_new_n34154__ = ~new_new_n34152__ & new_new_n34153__;
  assign new_new_n34155__ = ~new_new_n34147__ & ~new_new_n34150__;
  assign new_new_n34156__ = ~new_new_n34154__ & new_new_n34155__;
  assign new_new_n34157__ = ~new_new_n33602__ & new_new_n34156__;
  assign new_new_n34158__ = new_new_n34133__ & new_new_n34138__;
  assign new_new_n34159__ = ~new_new_n34156__ & new_new_n34158__;
  assign new_new_n34160__ = new_new_n34156__ & ~new_new_n34158__;
  assign new_new_n34161__ = ~new_new_n34159__ & ~new_new_n34160__;
  assign new_new_n34162__ = ~new_new_n7191__ & new_new_n34121__;
  assign new_new_n34163__ = new_new_n33885__ & new_new_n34118__;
  assign new_new_n34164__ = ~new_new_n33886__ & ~new_new_n34163__;
  assign new_new_n34165__ = ~new_new_n34162__ & new_new_n34164__;
  assign new_new_n34166__ = new_new_n34162__ & ~new_new_n34164__;
  assign new_new_n34167__ = ~new_new_n34165__ & ~new_new_n34166__;
  assign new_new_n34168__ = ~new_new_n33901__ & new_new_n34115__;
  assign new_new_n34169__ = ~new_new_n33902__ & ~new_new_n34168__;
  assign new_new_n34170__ = new_new_n34167__ & new_new_n34169__;
  assign new_new_n34171__ = ~new_new_n34167__ & ~new_new_n34169__;
  assign new_new_n34172__ = ~new_new_n34170__ & ~new_new_n34171__;
  assign new_new_n34173__ = new_new_n12832__ & new_new_n32729__;
  assign new_new_n34174__ = new_new_n11475__ & new_new_n32740__;
  assign new_new_n34175__ = ~new_new_n34173__ & ~new_new_n34174__;
  assign new_new_n34176__ = pi05 & ~new_new_n34175__;
  assign new_new_n34177__ = new_new_n32729__ & ~new_new_n33050__;
  assign new_new_n34178__ = ~new_new_n32740__ & ~new_new_n34177__;
  assign new_new_n34179__ = new_new_n12856__ & ~new_new_n34178__;
  assign new_new_n34180__ = new_new_n11469__ & ~new_new_n34178__;
  assign new_new_n34181__ = ~pi05 & ~new_new_n34180__;
  assign new_new_n34182__ = ~new_new_n34179__ & ~new_new_n34181__;
  assign new_new_n34183__ = new_new_n34175__ & ~new_new_n34182__;
  assign new_new_n34184__ = ~new_new_n34176__ & ~new_new_n34183__;
  assign new_new_n34185__ = new_new_n10698__ & new_new_n32382__;
  assign new_new_n34186__ = ~new_new_n11409__ & ~new_new_n26674__;
  assign new_new_n34187__ = new_new_n10702__ & ~new_new_n26667__;
  assign new_new_n34188__ = new_new_n11378__ & ~new_new_n33347__;
  assign new_new_n34189__ = ~new_new_n34186__ & ~new_new_n34187__;
  assign new_new_n34190__ = ~new_new_n34185__ & new_new_n34189__;
  assign new_new_n34191__ = ~new_new_n34188__ & new_new_n34190__;
  assign new_new_n34192__ = ~pi08 & ~new_new_n34191__;
  assign new_new_n34193__ = pi08 & new_new_n34191__;
  assign new_new_n34194__ = ~new_new_n34192__ & ~new_new_n34193__;
  assign new_new_n34195__ = new_new_n8474__ & new_new_n27250__;
  assign new_new_n34196__ = ~new_new_n8479__ & ~new_new_n27242__;
  assign new_new_n34197__ = ~new_new_n34195__ & ~new_new_n34196__;
  assign new_new_n34198__ = new_new_n8469__ & new_new_n26698__;
  assign new_new_n34199__ = new_new_n31511__ & new_new_n34198__;
  assign new_new_n34200__ = new_new_n34197__ & ~new_new_n34199__;
  assign new_new_n34201__ = pi11 & ~new_new_n34200__;
  assign new_new_n34202__ = new_new_n8469__ & ~new_new_n31510__;
  assign new_new_n34203__ = ~pi11 & ~new_new_n34202__;
  assign new_new_n34204__ = ~new_new_n26698__ & ~new_new_n31508__;
  assign new_new_n34205__ = ~pi10 & ~new_new_n34204__;
  assign new_new_n34206__ = pi10 & ~new_new_n31509__;
  assign new_new_n34207__ = new_new_n8469__ & ~new_new_n34205__;
  assign new_new_n34208__ = ~new_new_n34206__ & new_new_n34207__;
  assign new_new_n34209__ = ~new_new_n34203__ & ~new_new_n34208__;
  assign new_new_n34210__ = new_new_n34197__ & ~new_new_n34209__;
  assign new_new_n34211__ = ~new_new_n34201__ & ~new_new_n34210__;
  assign new_new_n34212__ = new_new_n6991__ & new_new_n26774__;
  assign new_new_n34213__ = new_new_n6985__ & new_new_n26729__;
  assign new_new_n34214__ = ~new_new_n34212__ & ~new_new_n34213__;
  assign new_new_n34215__ = new_new_n6994__ & new_new_n27349__;
  assign new_new_n34216__ = new_new_n34214__ & ~new_new_n34215__;
  assign new_new_n34217__ = pi14 & ~new_new_n34216__;
  assign new_new_n34218__ = ~pi13 & new_new_n26722__;
  assign new_new_n34219__ = new_new_n6994__ & ~new_new_n27350__;
  assign new_new_n34220__ = pi13 & ~new_new_n27348__;
  assign new_new_n34221__ = ~new_new_n34218__ & ~new_new_n34220__;
  assign new_new_n34222__ = new_new_n34219__ & new_new_n34221__;
  assign new_new_n34223__ = ~pi14 & new_new_n34214__;
  assign new_new_n34224__ = ~new_new_n34219__ & new_new_n34223__;
  assign new_new_n34225__ = ~new_new_n34222__ & ~new_new_n34224__;
  assign new_new_n34226__ = ~new_new_n34217__ & new_new_n34225__;
  assign new_new_n34227__ = new_new_n6634__ & ~new_new_n27221__;
  assign new_new_n34228__ = new_new_n6629__ & ~new_new_n26823__;
  assign new_new_n34229__ = ~new_new_n6625__ & new_new_n26847__;
  assign new_new_n34230__ = new_new_n6936__ & new_new_n27411__;
  assign new_new_n34231__ = ~new_new_n34228__ & ~new_new_n34229__;
  assign new_new_n34232__ = ~new_new_n34227__ & new_new_n34231__;
  assign new_new_n34233__ = ~new_new_n34230__ & new_new_n34232__;
  assign new_new_n34234__ = pi20 & ~new_new_n34233__;
  assign new_new_n34235__ = ~pi20 & new_new_n34233__;
  assign new_new_n34236__ = ~new_new_n34234__ & ~new_new_n34235__;
  assign new_new_n34237__ = new_new_n5215__ & ~new_new_n27430__;
  assign new_new_n34238__ = new_new_n5191__ & new_new_n26922__;
  assign new_new_n34239__ = new_new_n5183__ & ~new_new_n26888__;
  assign new_new_n34240__ = ~new_new_n34238__ & ~new_new_n34239__;
  assign new_new_n34241__ = ~new_new_n34237__ & new_new_n34240__;
  assign new_new_n34242__ = new_new_n5195__ & ~new_new_n26854__;
  assign new_new_n34243__ = pi23 & ~new_new_n34242__;
  assign new_new_n34244__ = new_new_n5974__ & ~new_new_n26854__;
  assign new_new_n34245__ = ~new_new_n34243__ & ~new_new_n34244__;
  assign new_new_n34246__ = new_new_n34241__ & ~new_new_n34245__;
  assign new_new_n34247__ = ~pi23 & ~new_new_n34241__;
  assign new_new_n34248__ = ~new_new_n34246__ & ~new_new_n34247__;
  assign new_new_n34249__ = new_new_n33969__ & new_new_n34065__;
  assign new_new_n34250__ = ~new_new_n33969__ & ~new_new_n34065__;
  assign new_new_n34251__ = ~new_new_n34050__ & ~new_new_n34250__;
  assign new_new_n34252__ = ~new_new_n34249__ & ~new_new_n34251__;
  assign new_new_n34253__ = ~new_new_n34248__ & new_new_n34252__;
  assign new_new_n34254__ = new_new_n34248__ & ~new_new_n34252__;
  assign new_new_n34255__ = ~new_new_n34253__ & ~new_new_n34254__;
  assign new_new_n34256__ = new_new_n873__ & new_new_n26917__;
  assign new_new_n34257__ = ~new_new_n333__ & new_new_n26928__;
  assign new_new_n34258__ = new_new_n3311__ & ~new_new_n27168__;
  assign new_new_n34259__ = ~new_new_n34257__ & ~new_new_n34258__;
  assign new_new_n34260__ = ~new_new_n34256__ & new_new_n34259__;
  assign new_new_n34261__ = ~pi26 & ~new_new_n34260__;
  assign new_new_n34262__ = new_new_n512__ & ~new_new_n28799__;
  assign new_new_n34263__ = new_new_n801__ & ~new_new_n28799__;
  assign new_new_n34264__ = pi26 & ~new_new_n34263__;
  assign new_new_n34265__ = ~new_new_n34262__ & ~new_new_n34264__;
  assign new_new_n34266__ = new_new_n34260__ & ~new_new_n34265__;
  assign new_new_n34267__ = ~new_new_n34261__ & ~new_new_n34266__;
  assign new_new_n34268__ = new_new_n4212__ & new_new_n27152__;
  assign new_new_n34269__ = new_new_n4815__ & ~new_new_n26941__;
  assign new_new_n34270__ = ~new_new_n4818__ & ~new_new_n26937__;
  assign new_new_n34271__ = new_new_n4813__ & ~new_new_n27502__;
  assign new_new_n34272__ = ~new_new_n34269__ & ~new_new_n34270__;
  assign new_new_n34273__ = ~new_new_n34268__ & new_new_n34272__;
  assign new_new_n34274__ = ~new_new_n34271__ & new_new_n34273__;
  assign new_new_n34275__ = new_new_n26978__ & ~new_new_n27121__;
  assign new_new_n34276__ = ~new_new_n15853__ & ~new_new_n27122__;
  assign new_new_n34277__ = ~new_new_n34275__ & new_new_n34276__;
  assign new_new_n34278__ = ~new_new_n27981__ & ~new_new_n34277__;
  assign new_new_n34279__ = ~new_new_n26971__ & ~new_new_n34278__;
  assign new_new_n34280__ = new_new_n27121__ & new_new_n28265__;
  assign new_new_n34281__ = ~new_new_n161__ & ~new_new_n34280__;
  assign new_new_n34282__ = ~new_new_n71__ & new_new_n27003__;
  assign new_new_n34283__ = ~new_new_n34281__ & new_new_n34282__;
  assign new_new_n34284__ = ~new_new_n27121__ & new_new_n28255__;
  assign new_new_n34285__ = ~new_new_n71__ & ~new_new_n34284__;
  assign new_new_n34286__ = new_new_n34024__ & ~new_new_n34285__;
  assign new_new_n34287__ = pi31 & ~new_new_n34279__;
  assign new_new_n34288__ = ~new_new_n34283__ & ~new_new_n34286__;
  assign new_new_n34289__ = new_new_n34287__ & new_new_n34288__;
  assign new_new_n34290__ = new_new_n161__ & ~new_new_n26978__;
  assign new_new_n34291__ = new_new_n765__ & new_new_n26971__;
  assign new_new_n34292__ = ~new_new_n34290__ & ~new_new_n34291__;
  assign new_new_n34293__ = ~pi31 & ~new_new_n34292__;
  assign new_new_n34294__ = ~new_new_n34289__ & ~new_new_n34293__;
  assign new_new_n34295__ = ~pi02 & new_new_n34294__;
  assign new_new_n34296__ = pi02 & ~new_new_n34294__;
  assign new_new_n34297__ = ~new_new_n34295__ & ~new_new_n34296__;
  assign new_new_n34298__ = ~new_new_n76__ & ~new_new_n138__;
  assign new_new_n34299__ = ~new_new_n496__ & new_new_n34298__;
  assign new_new_n34300__ = ~new_new_n774__ & new_new_n777__;
  assign new_new_n34301__ = ~new_new_n1009__ & new_new_n4577__;
  assign new_new_n34302__ = new_new_n7648__ & new_new_n34301__;
  assign new_new_n34303__ = new_new_n34299__ & new_new_n34300__;
  assign new_new_n34304__ = new_new_n177__ & new_new_n484__;
  assign new_new_n34305__ = new_new_n897__ & new_new_n4989__;
  assign new_new_n34306__ = new_new_n34304__ & new_new_n34305__;
  assign new_new_n34307__ = new_new_n34302__ & new_new_n34303__;
  assign new_new_n34308__ = new_new_n936__ & new_new_n1627__;
  assign new_new_n34309__ = new_new_n3393__ & new_new_n16896__;
  assign new_new_n34310__ = new_new_n34308__ & new_new_n34309__;
  assign new_new_n34311__ = new_new_n34306__ & new_new_n34307__;
  assign new_new_n34312__ = new_new_n34310__ & new_new_n34311__;
  assign new_new_n34313__ = new_new_n2554__ & new_new_n16127__;
  assign new_new_n34314__ = new_new_n34312__ & new_new_n34313__;
  assign new_new_n34315__ = new_new_n3075__ & new_new_n34314__;
  assign new_new_n34316__ = new_new_n370__ & new_new_n34315__;
  assign new_new_n34317__ = ~new_new_n34297__ & new_new_n34316__;
  assign new_new_n34318__ = new_new_n34297__ & ~new_new_n34316__;
  assign new_new_n34319__ = ~new_new_n34317__ & ~new_new_n34318__;
  assign new_new_n34320__ = ~new_new_n34030__ & new_new_n34034__;
  assign new_new_n34321__ = ~new_new_n34031__ & ~new_new_n34320__;
  assign new_new_n34322__ = new_new_n34319__ & ~new_new_n34321__;
  assign new_new_n34323__ = ~new_new_n34319__ & new_new_n34321__;
  assign new_new_n34324__ = ~new_new_n34322__ & ~new_new_n34323__;
  assign new_new_n34325__ = pi29 & ~new_new_n34324__;
  assign new_new_n34326__ = ~pi29 & new_new_n34324__;
  assign new_new_n34327__ = ~new_new_n34325__ & ~new_new_n34326__;
  assign new_new_n34328__ = new_new_n34274__ & new_new_n34327__;
  assign new_new_n34329__ = ~new_new_n34274__ & ~new_new_n34327__;
  assign new_new_n34330__ = ~new_new_n34328__ & ~new_new_n34329__;
  assign new_new_n34331__ = ~new_new_n34043__ & ~new_new_n34050__;
  assign new_new_n34332__ = ~new_new_n34042__ & ~new_new_n34331__;
  assign new_new_n34333__ = ~new_new_n34330__ & new_new_n34332__;
  assign new_new_n34334__ = new_new_n34330__ & ~new_new_n34332__;
  assign new_new_n34335__ = ~new_new_n34333__ & ~new_new_n34334__;
  assign new_new_n34336__ = new_new_n34267__ & new_new_n34335__;
  assign new_new_n34337__ = ~new_new_n34267__ & ~new_new_n34335__;
  assign new_new_n34338__ = ~new_new_n34336__ & ~new_new_n34337__;
  assign new_new_n34339__ = new_new_n34255__ & new_new_n34338__;
  assign new_new_n34340__ = ~new_new_n34255__ & ~new_new_n34338__;
  assign new_new_n34341__ = ~new_new_n34339__ & ~new_new_n34340__;
  assign new_new_n34342__ = ~new_new_n34236__ & new_new_n34341__;
  assign new_new_n34343__ = new_new_n34236__ & ~new_new_n34341__;
  assign new_new_n34344__ = ~new_new_n34342__ & ~new_new_n34343__;
  assign new_new_n34345__ = new_new_n6964__ & ~new_new_n26741__;
  assign new_new_n34346__ = new_new_n6968__ & ~new_new_n26802__;
  assign new_new_n34347__ = ~new_new_n34345__ & ~new_new_n34346__;
  assign new_new_n34348__ = new_new_n6958__ & new_new_n26810__;
  assign new_new_n34349__ = new_new_n27395__ & new_new_n34348__;
  assign new_new_n34350__ = new_new_n34347__ & ~new_new_n34349__;
  assign new_new_n34351__ = ~pi17 & ~new_new_n34350__;
  assign new_new_n34352__ = ~new_new_n26810__ & ~new_new_n27395__;
  assign new_new_n34353__ = new_new_n6958__ & ~new_new_n34352__;
  assign new_new_n34354__ = ~pi17 & ~new_new_n34353__;
  assign new_new_n34355__ = ~pi16 & ~new_new_n27395__;
  assign new_new_n34356__ = pi16 & ~new_new_n26810__;
  assign new_new_n34357__ = new_new_n6958__ & ~new_new_n34356__;
  assign new_new_n34358__ = ~new_new_n34355__ & new_new_n34357__;
  assign new_new_n34359__ = new_new_n34347__ & ~new_new_n34358__;
  assign new_new_n34360__ = ~new_new_n34354__ & new_new_n34359__;
  assign new_new_n34361__ = ~new_new_n34351__ & ~new_new_n34360__;
  assign new_new_n34362__ = new_new_n33967__ & ~new_new_n33969__;
  assign new_new_n34363__ = ~new_new_n33967__ & new_new_n33969__;
  assign new_new_n34364__ = ~new_new_n34362__ & ~new_new_n34363__;
  assign new_new_n34365__ = ~new_new_n34050__ & new_new_n34080__;
  assign new_new_n34366__ = new_new_n34050__ & ~new_new_n34080__;
  assign new_new_n34367__ = ~new_new_n34365__ & ~new_new_n34366__;
  assign new_new_n34368__ = new_new_n34364__ & new_new_n34367__;
  assign new_new_n34369__ = ~new_new_n34364__ & ~new_new_n34367__;
  assign new_new_n34370__ = ~new_new_n34368__ & ~new_new_n34369__;
  assign new_new_n34371__ = new_new_n33727__ & ~new_new_n34370__;
  assign new_new_n34372__ = ~new_new_n33729__ & ~new_new_n34371__;
  assign new_new_n34373__ = ~new_new_n34087__ & new_new_n34372__;
  assign new_new_n34374__ = ~new_new_n33727__ & new_new_n34370__;
  assign new_new_n34375__ = ~new_new_n33727__ & ~new_new_n33834__;
  assign new_new_n34376__ = pi20 & ~new_new_n34375__;
  assign new_new_n34377__ = ~new_new_n34374__ & ~new_new_n34376__;
  assign new_new_n34378__ = new_new_n34087__ & ~new_new_n34377__;
  assign new_new_n34379__ = ~pi20 & ~new_new_n34087__;
  assign new_new_n34380__ = ~new_new_n34370__ & ~new_new_n34379__;
  assign new_new_n34381__ = new_new_n33834__ & ~new_new_n34380__;
  assign new_new_n34382__ = ~new_new_n34373__ & ~new_new_n34381__;
  assign new_new_n34383__ = ~new_new_n34378__ & new_new_n34382__;
  assign new_new_n34384__ = new_new_n33832__ & ~new_new_n34383__;
  assign new_new_n34385__ = pi20 & new_new_n34370__;
  assign new_new_n34386__ = ~new_new_n33727__ & ~new_new_n34370__;
  assign new_new_n34387__ = ~new_new_n33728__ & new_new_n33834__;
  assign new_new_n34388__ = ~new_new_n34386__ & new_new_n34387__;
  assign new_new_n34389__ = ~new_new_n34385__ & ~new_new_n34388__;
  assign new_new_n34390__ = new_new_n34087__ & ~new_new_n34389__;
  assign new_new_n34391__ = ~pi20 & new_new_n34370__;
  assign new_new_n34392__ = new_new_n33834__ & new_new_n34372__;
  assign new_new_n34393__ = ~new_new_n34391__ & ~new_new_n34392__;
  assign new_new_n34394__ = ~new_new_n34087__ & ~new_new_n34393__;
  assign new_new_n34395__ = ~new_new_n34390__ & ~new_new_n34394__;
  assign new_new_n34396__ = ~new_new_n34384__ & new_new_n34395__;
  assign new_new_n34397__ = ~new_new_n34361__ & ~new_new_n34396__;
  assign new_new_n34398__ = new_new_n34361__ & new_new_n34396__;
  assign new_new_n34399__ = ~new_new_n34397__ & ~new_new_n34398__;
  assign new_new_n34400__ = ~new_new_n33967__ & new_new_n34077__;
  assign new_new_n34401__ = new_new_n33967__ & ~new_new_n34077__;
  assign new_new_n34402__ = ~new_new_n34249__ & ~new_new_n34250__;
  assign new_new_n34403__ = ~new_new_n34050__ & new_new_n34402__;
  assign new_new_n34404__ = new_new_n34050__ & ~new_new_n34402__;
  assign new_new_n34405__ = ~new_new_n34403__ & ~new_new_n34404__;
  assign new_new_n34406__ = ~new_new_n34401__ & new_new_n34405__;
  assign new_new_n34407__ = ~new_new_n34400__ & ~new_new_n34406__;
  assign new_new_n34408__ = new_new_n34399__ & ~new_new_n34407__;
  assign new_new_n34409__ = ~new_new_n34399__ & new_new_n34407__;
  assign new_new_n34410__ = ~new_new_n34408__ & ~new_new_n34409__;
  assign new_new_n34411__ = new_new_n34344__ & new_new_n34410__;
  assign new_new_n34412__ = ~new_new_n34344__ & ~new_new_n34410__;
  assign new_new_n34413__ = ~new_new_n34411__ & ~new_new_n34412__;
  assign new_new_n34414__ = new_new_n34226__ & ~new_new_n34413__;
  assign new_new_n34415__ = ~new_new_n34226__ & new_new_n34413__;
  assign new_new_n34416__ = ~new_new_n34414__ & ~new_new_n34415__;
  assign new_new_n34417__ = new_new_n33952__ & ~new_new_n34096__;
  assign new_new_n34418__ = ~new_new_n34097__ & ~new_new_n34417__;
  assign new_new_n34419__ = new_new_n34416__ & new_new_n34418__;
  assign new_new_n34420__ = ~new_new_n34416__ & ~new_new_n34418__;
  assign new_new_n34421__ = ~new_new_n34419__ & ~new_new_n34420__;
  assign new_new_n34422__ = new_new_n34211__ & ~new_new_n34421__;
  assign new_new_n34423__ = ~new_new_n33934__ & ~new_new_n34102__;
  assign new_new_n34424__ = ~new_new_n34211__ & new_new_n34421__;
  assign new_new_n34425__ = ~new_new_n34103__ & ~new_new_n34424__;
  assign new_new_n34426__ = ~new_new_n34423__ & new_new_n34425__;
  assign new_new_n34427__ = ~new_new_n34422__ & new_new_n34426__;
  assign new_new_n34428__ = ~new_new_n33934__ & new_new_n34422__;
  assign new_new_n34429__ = new_new_n33936__ & new_new_n34424__;
  assign new_new_n34430__ = ~new_new_n34428__ & ~new_new_n34429__;
  assign new_new_n34431__ = new_new_n34101__ & ~new_new_n34430__;
  assign new_new_n34432__ = new_new_n33936__ & new_new_n34422__;
  assign new_new_n34433__ = new_new_n34104__ & new_new_n34424__;
  assign new_new_n34434__ = ~new_new_n34432__ & ~new_new_n34433__;
  assign new_new_n34435__ = new_new_n34107__ & ~new_new_n34434__;
  assign new_new_n34436__ = ~new_new_n34427__ & ~new_new_n34431__;
  assign new_new_n34437__ = ~new_new_n34435__ & new_new_n34436__;
  assign new_new_n34438__ = ~new_new_n33913__ & ~new_new_n34110__;
  assign new_new_n34439__ = ~new_new_n34111__ & ~new_new_n34438__;
  assign new_new_n34440__ = new_new_n34437__ & new_new_n34439__;
  assign new_new_n34441__ = ~new_new_n34437__ & ~new_new_n34439__;
  assign new_new_n34442__ = ~new_new_n34440__ & ~new_new_n34441__;
  assign new_new_n34443__ = new_new_n34194__ & ~new_new_n34442__;
  assign new_new_n34444__ = ~new_new_n34194__ & new_new_n34442__;
  assign new_new_n34445__ = ~new_new_n34443__ & ~new_new_n34444__;
  assign new_new_n34446__ = ~new_new_n34184__ & new_new_n34445__;
  assign new_new_n34447__ = new_new_n34184__ & ~new_new_n34445__;
  assign new_new_n34448__ = ~new_new_n34446__ & ~new_new_n34447__;
  assign new_new_n34449__ = new_new_n34172__ & ~new_new_n34448__;
  assign new_new_n34450__ = ~new_new_n34172__ & new_new_n34448__;
  assign new_new_n34451__ = ~new_new_n34449__ & ~new_new_n34450__;
  assign new_new_n34452__ = ~new_new_n34157__ & new_new_n34451__;
  assign new_new_n34453__ = new_new_n34161__ & new_new_n34452__;
  assign new_new_n34454__ = ~new_new_n34161__ & ~new_new_n34451__;
  assign po07 = new_new_n34453__ | new_new_n34454__;
  assign new_new_n34456__ = new_new_n34158__ & ~po07;
  assign new_new_n34457__ = ~new_new_n34156__ & new_new_n34167__;
  assign new_new_n34458__ = ~new_new_n34169__ & new_new_n34445__;
  assign new_new_n34459__ = new_new_n34169__ & ~new_new_n34445__;
  assign new_new_n34460__ = new_new_n34184__ & ~new_new_n34459__;
  assign new_new_n34461__ = ~new_new_n34458__ & ~new_new_n34460__;
  assign new_new_n34462__ = ~new_new_n34457__ & new_new_n34461__;
  assign new_new_n34463__ = new_new_n34156__ & ~new_new_n34167__;
  assign new_new_n34464__ = ~new_new_n34461__ & ~new_new_n34463__;
  assign new_new_n34465__ = ~new_new_n34462__ & ~new_new_n34464__;
  assign new_new_n34466__ = new_new_n34194__ & ~new_new_n34440__;
  assign new_new_n34467__ = ~new_new_n34441__ & ~new_new_n34466__;
  assign new_new_n34468__ = ~new_new_n34422__ & ~new_new_n34426__;
  assign new_new_n34469__ = new_new_n11378__ & new_new_n32758__;
  assign new_new_n34470__ = ~new_new_n11409__ & ~new_new_n26667__;
  assign new_new_n34471__ = new_new_n10702__ & new_new_n32382__;
  assign new_new_n34472__ = ~new_new_n34470__ & ~new_new_n34471__;
  assign new_new_n34473__ = ~new_new_n34469__ & new_new_n34472__;
  assign new_new_n34474__ = new_new_n10694__ & new_new_n32729__;
  assign new_new_n34475__ = pi08 & ~new_new_n34474__;
  assign new_new_n34476__ = new_new_n12121__ & new_new_n32729__;
  assign new_new_n34477__ = ~new_new_n34475__ & ~new_new_n34476__;
  assign new_new_n34478__ = new_new_n34473__ & ~new_new_n34477__;
  assign new_new_n34479__ = ~pi08 & ~new_new_n34473__;
  assign new_new_n34480__ = ~new_new_n34478__ & ~new_new_n34479__;
  assign new_new_n34481__ = new_new_n34468__ & new_new_n34480__;
  assign new_new_n34482__ = ~new_new_n34468__ & ~new_new_n34480__;
  assign new_new_n34483__ = ~new_new_n34481__ & ~new_new_n34482__;
  assign new_new_n34484__ = new_new_n6985__ & new_new_n26722__;
  assign new_new_n34485__ = new_new_n6991__ & new_new_n26729__;
  assign new_new_n34486__ = ~new_new_n34484__ & ~new_new_n34485__;
  assign new_new_n34487__ = new_new_n6994__ & ~new_new_n27362__;
  assign new_new_n34488__ = pi14 & ~new_new_n34487__;
  assign new_new_n34489__ = new_new_n8388__ & ~new_new_n27242__;
  assign new_new_n34490__ = new_new_n27352__ & new_new_n34489__;
  assign new_new_n34491__ = ~new_new_n34488__ & ~new_new_n34490__;
  assign new_new_n34492__ = new_new_n34486__ & ~new_new_n34491__;
  assign new_new_n34493__ = new_new_n6994__ & new_new_n27353__;
  assign new_new_n34494__ = new_new_n34486__ & ~new_new_n34493__;
  assign new_new_n34495__ = ~pi14 & ~new_new_n34494__;
  assign new_new_n34496__ = new_new_n8820__ & new_new_n27242__;
  assign new_new_n34497__ = new_new_n27352__ & new_new_n34496__;
  assign new_new_n34498__ = ~new_new_n34495__ & ~new_new_n34497__;
  assign new_new_n34499__ = ~new_new_n34492__ & new_new_n34498__;
  assign new_new_n34500__ = new_new_n34344__ & ~new_new_n34407__;
  assign new_new_n34501__ = ~new_new_n34344__ & new_new_n34407__;
  assign new_new_n34502__ = ~new_new_n34500__ & ~new_new_n34501__;
  assign new_new_n34503__ = ~new_new_n34397__ & new_new_n34502__;
  assign new_new_n34504__ = ~new_new_n34398__ & ~new_new_n34503__;
  assign new_new_n34505__ = ~new_new_n34499__ & new_new_n34504__;
  assign new_new_n34506__ = new_new_n34499__ & ~new_new_n34504__;
  assign new_new_n34507__ = ~new_new_n34505__ & ~new_new_n34506__;
  assign new_new_n34508__ = ~new_new_n34343__ & ~new_new_n34407__;
  assign new_new_n34509__ = ~new_new_n34342__ & ~new_new_n34508__;
  assign new_new_n34510__ = new_new_n6634__ & ~new_new_n26741__;
  assign new_new_n34511__ = ~new_new_n6625__ & ~new_new_n26823__;
  assign new_new_n34512__ = new_new_n6629__ & ~new_new_n27221__;
  assign new_new_n34513__ = new_new_n6936__ & new_new_n30393__;
  assign new_new_n34514__ = ~new_new_n34511__ & ~new_new_n34512__;
  assign new_new_n34515__ = ~new_new_n34510__ & new_new_n34514__;
  assign new_new_n34516__ = ~new_new_n34513__ & new_new_n34515__;
  assign new_new_n34517__ = ~pi20 & ~new_new_n34516__;
  assign new_new_n34518__ = pi20 & new_new_n34516__;
  assign new_new_n34519__ = ~new_new_n34517__ & ~new_new_n34518__;
  assign new_new_n34520__ = ~new_new_n34254__ & ~new_new_n34338__;
  assign new_new_n34521__ = ~new_new_n34253__ & ~new_new_n34520__;
  assign new_new_n34522__ = new_new_n34519__ & new_new_n34521__;
  assign new_new_n34523__ = ~new_new_n34519__ & ~new_new_n34521__;
  assign new_new_n34524__ = ~new_new_n34522__ & ~new_new_n34523__;
  assign new_new_n34525__ = new_new_n5213__ & new_new_n26847__;
  assign new_new_n34526__ = new_new_n5191__ & ~new_new_n26888__;
  assign new_new_n34527__ = new_new_n5183__ & ~new_new_n26854__;
  assign new_new_n34528__ = ~new_new_n34526__ & ~new_new_n34527__;
  assign new_new_n34529__ = ~new_new_n34525__ & new_new_n34528__;
  assign new_new_n34530__ = new_new_n5195__ & new_new_n29424__;
  assign new_new_n34531__ = ~pi23 & ~new_new_n34530__;
  assign new_new_n34532__ = new_new_n5974__ & new_new_n29424__;
  assign new_new_n34533__ = ~new_new_n34531__ & ~new_new_n34532__;
  assign new_new_n34534__ = new_new_n34529__ & ~new_new_n34533__;
  assign new_new_n34535__ = pi23 & ~new_new_n34529__;
  assign new_new_n34536__ = ~new_new_n34534__ & ~new_new_n34535__;
  assign new_new_n34537__ = ~new_new_n34267__ & ~new_new_n34333__;
  assign new_new_n34538__ = ~new_new_n34334__ & ~new_new_n34537__;
  assign new_new_n34539__ = ~new_new_n34536__ & new_new_n34538__;
  assign new_new_n34540__ = new_new_n34536__ & ~new_new_n34538__;
  assign new_new_n34541__ = ~new_new_n34539__ & ~new_new_n34540__;
  assign new_new_n34542__ = new_new_n4815__ & new_new_n26928__;
  assign new_new_n34543__ = new_new_n4212__ & ~new_new_n26941__;
  assign new_new_n34544__ = ~new_new_n4818__ & new_new_n27152__;
  assign new_new_n34545__ = new_new_n4813__ & new_new_n27488__;
  assign new_new_n34546__ = ~new_new_n34543__ & ~new_new_n34544__;
  assign new_new_n34547__ = ~new_new_n34542__ & new_new_n34546__;
  assign new_new_n34548__ = ~new_new_n34545__ & new_new_n34547__;
  assign new_new_n34549__ = ~new_new_n333__ & new_new_n26917__;
  assign new_new_n34550__ = new_new_n873__ & ~new_new_n27168__;
  assign new_new_n34551__ = ~new_new_n4900__ & ~new_new_n29366__;
  assign new_new_n34552__ = ~new_new_n34549__ & ~new_new_n34550__;
  assign new_new_n34553__ = ~new_new_n34551__ & new_new_n34552__;
  assign new_new_n34554__ = ~pi26 & ~new_new_n34553__;
  assign new_new_n34555__ = new_new_n4898__ & new_new_n26922__;
  assign new_new_n34556__ = new_new_n801__ & new_new_n26922__;
  assign new_new_n34557__ = pi26 & ~new_new_n34556__;
  assign new_new_n34558__ = ~new_new_n34555__ & ~new_new_n34557__;
  assign new_new_n34559__ = new_new_n34553__ & ~new_new_n34558__;
  assign new_new_n34560__ = ~new_new_n34554__ & ~new_new_n34559__;
  assign new_new_n34561__ = new_new_n161__ & new_new_n26971__;
  assign new_new_n34562__ = new_new_n765__ & ~new_new_n26937__;
  assign new_new_n34563__ = ~new_new_n34561__ & ~new_new_n34562__;
  assign new_new_n34564__ = ~pi31 & ~new_new_n34563__;
  assign new_new_n34565__ = new_new_n71__ & new_new_n26971__;
  assign new_new_n34566__ = new_new_n765__ & new_new_n28005__;
  assign new_new_n34567__ = ~new_new_n34290__ & ~new_new_n34565__;
  assign new_new_n34568__ = ~new_new_n34566__ & new_new_n34567__;
  assign new_new_n34569__ = pi31 & ~new_new_n34568__;
  assign new_new_n34570__ = ~new_new_n34564__ & ~new_new_n34569__;
  assign new_new_n34571__ = ~new_new_n34323__ & ~new_new_n34330__;
  assign new_new_n34572__ = ~new_new_n34322__ & ~new_new_n34571__;
  assign new_new_n34573__ = new_new_n34570__ & new_new_n34572__;
  assign new_new_n34574__ = ~new_new_n34570__ & ~new_new_n34572__;
  assign new_new_n34575__ = ~new_new_n34573__ & ~new_new_n34574__;
  assign new_new_n34576__ = pi02 & ~new_new_n34575__;
  assign new_new_n34577__ = ~pi02 & new_new_n34575__;
  assign new_new_n34578__ = ~new_new_n34576__ & ~new_new_n34577__;
  assign new_new_n34579__ = ~new_new_n34295__ & ~new_new_n34316__;
  assign new_new_n34580__ = ~new_new_n34296__ & ~new_new_n34579__;
  assign new_new_n34581__ = ~new_new_n260__ & ~new_new_n698__;
  assign new_new_n34582__ = new_new_n5567__ & new_new_n34581__;
  assign new_new_n34583__ = new_new_n256__ & new_new_n34582__;
  assign new_new_n34584__ = new_new_n114__ & new_new_n16850__;
  assign new_new_n34585__ = ~new_new_n246__ & new_new_n786__;
  assign new_new_n34586__ = ~new_new_n878__ & ~new_new_n1568__;
  assign new_new_n34587__ = new_new_n34585__ & new_new_n34586__;
  assign new_new_n34588__ = new_new_n307__ & new_new_n1292__;
  assign new_new_n34589__ = new_new_n2913__ & new_new_n4597__;
  assign new_new_n34590__ = new_new_n5366__ & new_new_n16238__;
  assign new_new_n34591__ = ~new_new_n34584__ & new_new_n34590__;
  assign new_new_n34592__ = new_new_n34588__ & new_new_n34589__;
  assign new_new_n34593__ = new_new_n5315__ & new_new_n34587__;
  assign new_new_n34594__ = new_new_n17246__ & new_new_n34593__;
  assign new_new_n34595__ = new_new_n34591__ & new_new_n34592__;
  assign new_new_n34596__ = new_new_n669__ & new_new_n2524__;
  assign new_new_n34597__ = new_new_n34583__ & new_new_n34596__;
  assign new_new_n34598__ = new_new_n34594__ & new_new_n34595__;
  assign new_new_n34599__ = new_new_n34597__ & new_new_n34598__;
  assign new_new_n34600__ = new_new_n2671__ & new_new_n34599__;
  assign new_new_n34601__ = new_new_n19292__ & new_new_n34600__;
  assign new_new_n34602__ = new_new_n34580__ & ~new_new_n34601__;
  assign new_new_n34603__ = ~new_new_n34580__ & new_new_n34601__;
  assign new_new_n34604__ = ~new_new_n34602__ & ~new_new_n34603__;
  assign new_new_n34605__ = new_new_n34578__ & new_new_n34604__;
  assign new_new_n34606__ = ~new_new_n34578__ & ~new_new_n34604__;
  assign new_new_n34607__ = ~new_new_n34605__ & ~new_new_n34606__;
  assign new_new_n34608__ = ~new_new_n34560__ & new_new_n34607__;
  assign new_new_n34609__ = new_new_n34560__ & ~new_new_n34607__;
  assign new_new_n34610__ = ~new_new_n34608__ & ~new_new_n34609__;
  assign new_new_n34611__ = pi29 & ~new_new_n34610__;
  assign new_new_n34612__ = ~pi29 & new_new_n34610__;
  assign new_new_n34613__ = ~new_new_n34611__ & ~new_new_n34612__;
  assign new_new_n34614__ = new_new_n34548__ & new_new_n34613__;
  assign new_new_n34615__ = ~new_new_n34548__ & ~new_new_n34613__;
  assign new_new_n34616__ = ~new_new_n34614__ & ~new_new_n34615__;
  assign new_new_n34617__ = new_new_n34541__ & ~new_new_n34616__;
  assign new_new_n34618__ = ~new_new_n34541__ & new_new_n34616__;
  assign new_new_n34619__ = ~new_new_n34617__ & ~new_new_n34618__;
  assign new_new_n34620__ = ~new_new_n34524__ & new_new_n34619__;
  assign new_new_n34621__ = new_new_n34524__ & ~new_new_n34619__;
  assign new_new_n34622__ = ~new_new_n34620__ & ~new_new_n34621__;
  assign new_new_n34623__ = ~new_new_n34509__ & ~new_new_n34622__;
  assign new_new_n34624__ = new_new_n34509__ & new_new_n34622__;
  assign new_new_n34625__ = ~new_new_n34623__ & ~new_new_n34624__;
  assign new_new_n34626__ = new_new_n7935__ & new_new_n26774__;
  assign new_new_n34627__ = new_new_n6964__ & ~new_new_n26802__;
  assign new_new_n34628__ = new_new_n6968__ & new_new_n26810__;
  assign new_new_n34629__ = ~new_new_n34627__ & ~new_new_n34628__;
  assign new_new_n34630__ = ~new_new_n34626__ & new_new_n34629__;
  assign new_new_n34631__ = new_new_n6958__ & ~new_new_n27373__;
  assign new_new_n34632__ = ~pi17 & ~new_new_n34631__;
  assign new_new_n34633__ = new_new_n8160__ & ~new_new_n27373__;
  assign new_new_n34634__ = ~new_new_n34632__ & ~new_new_n34633__;
  assign new_new_n34635__ = new_new_n34630__ & ~new_new_n34634__;
  assign new_new_n34636__ = pi17 & ~new_new_n34630__;
  assign new_new_n34637__ = ~new_new_n34635__ & ~new_new_n34636__;
  assign new_new_n34638__ = new_new_n34625__ & ~new_new_n34637__;
  assign new_new_n34639__ = ~new_new_n34625__ & new_new_n34637__;
  assign new_new_n34640__ = ~new_new_n34638__ & ~new_new_n34639__;
  assign new_new_n34641__ = new_new_n34507__ & ~new_new_n34640__;
  assign new_new_n34642__ = ~new_new_n34507__ & new_new_n34640__;
  assign new_new_n34643__ = ~new_new_n34641__ & ~new_new_n34642__;
  assign new_new_n34644__ = ~new_new_n34415__ & ~new_new_n34418__;
  assign new_new_n34645__ = ~new_new_n34414__ & ~new_new_n34644__;
  assign new_new_n34646__ = new_new_n34643__ & ~new_new_n34645__;
  assign new_new_n34647__ = ~new_new_n34643__ & new_new_n34645__;
  assign new_new_n34648__ = ~new_new_n34646__ & ~new_new_n34647__;
  assign new_new_n34649__ = new_new_n8858__ & ~new_new_n26674__;
  assign new_new_n34650__ = ~new_new_n8479__ & new_new_n27250__;
  assign new_new_n34651__ = new_new_n8474__ & new_new_n26698__;
  assign new_new_n34652__ = ~new_new_n34650__ & ~new_new_n34651__;
  assign new_new_n34653__ = ~new_new_n34649__ & new_new_n34652__;
  assign new_new_n34654__ = new_new_n8469__ & new_new_n27284__;
  assign new_new_n34655__ = pi11 & ~new_new_n34654__;
  assign new_new_n34656__ = new_new_n11530__ & new_new_n27284__;
  assign new_new_n34657__ = ~new_new_n34655__ & ~new_new_n34656__;
  assign new_new_n34658__ = new_new_n34653__ & ~new_new_n34657__;
  assign new_new_n34659__ = ~pi11 & ~new_new_n34653__;
  assign new_new_n34660__ = ~new_new_n34658__ & ~new_new_n34659__;
  assign new_new_n34661__ = new_new_n34648__ & new_new_n34660__;
  assign new_new_n34662__ = ~new_new_n34648__ & ~new_new_n34660__;
  assign new_new_n34663__ = ~new_new_n34661__ & ~new_new_n34662__;
  assign new_new_n34664__ = new_new_n34483__ & ~new_new_n34663__;
  assign new_new_n34665__ = ~new_new_n34483__ & new_new_n34663__;
  assign new_new_n34666__ = ~new_new_n34664__ & ~new_new_n34665__;
  assign new_new_n34667__ = new_new_n34467__ & new_new_n34666__;
  assign new_new_n34668__ = ~new_new_n34467__ & ~new_new_n34666__;
  assign new_new_n34669__ = ~new_new_n34667__ & ~new_new_n34668__;
  assign new_new_n34670__ = new_new_n11470__ & new_new_n32740__;
  assign new_new_n34671__ = pi05 & ~new_new_n34670__;
  assign new_new_n34672__ = new_new_n12828__ & new_new_n32740__;
  assign new_new_n34673__ = ~new_new_n34671__ & ~new_new_n34672__;
  assign new_new_n34674__ = new_new_n34669__ & new_new_n34673__;
  assign new_new_n34675__ = ~new_new_n34669__ & ~new_new_n34673__;
  assign new_new_n34676__ = ~new_new_n34674__ & ~new_new_n34675__;
  assign new_new_n34677__ = ~new_new_n34458__ & ~new_new_n34459__;
  assign new_new_n34678__ = new_new_n34448__ & ~new_new_n34677__;
  assign new_new_n34679__ = ~new_new_n34457__ & ~new_new_n34678__;
  assign new_new_n34680__ = ~new_new_n34463__ & new_new_n34679__;
  assign new_new_n34681__ = ~new_new_n34465__ & ~new_new_n34676__;
  assign new_new_n34682__ = ~new_new_n34680__ & new_new_n34681__;
  assign new_new_n34683__ = new_new_n34457__ & new_new_n34458__;
  assign new_new_n34684__ = new_new_n34169__ & new_new_n34463__;
  assign new_new_n34685__ = ~new_new_n34445__ & new_new_n34684__;
  assign new_new_n34686__ = ~new_new_n34169__ & ~new_new_n34463__;
  assign new_new_n34687__ = ~new_new_n34457__ & ~new_new_n34686__;
  assign new_new_n34688__ = ~new_new_n34169__ & new_new_n34457__;
  assign new_new_n34689__ = ~new_new_n34445__ & ~new_new_n34688__;
  assign new_new_n34690__ = ~new_new_n34687__ & ~new_new_n34689__;
  assign new_new_n34691__ = new_new_n34184__ & ~new_new_n34690__;
  assign new_new_n34692__ = ~new_new_n34445__ & new_new_n34687__;
  assign new_new_n34693__ = ~new_new_n34184__ & ~new_new_n34684__;
  assign new_new_n34694__ = ~new_new_n34692__ & new_new_n34693__;
  assign new_new_n34695__ = ~new_new_n34691__ & ~new_new_n34694__;
  assign new_new_n34696__ = new_new_n34676__ & ~new_new_n34683__;
  assign new_new_n34697__ = ~new_new_n34685__ & new_new_n34696__;
  assign new_new_n34698__ = ~new_new_n34695__ & new_new_n34697__;
  assign new_new_n34699__ = ~new_new_n34682__ & ~new_new_n34698__;
  assign new_new_n34700__ = new_new_n34456__ & ~new_new_n34699__;
  assign new_new_n34701__ = ~new_new_n34456__ & new_new_n34699__;
  assign po08 = ~new_new_n34700__ & ~new_new_n34701__;
  assign new_new_n34703__ = new_new_n34457__ & ~new_new_n34461__;
  assign new_new_n34704__ = ~new_new_n34462__ & ~new_new_n34676__;
  assign new_new_n34705__ = ~new_new_n34458__ & new_new_n34676__;
  assign new_new_n34706__ = new_new_n34184__ & ~new_new_n34705__;
  assign new_new_n34707__ = ~new_new_n34459__ & ~new_new_n34676__;
  assign new_new_n34708__ = ~new_new_n34706__ & ~new_new_n34707__;
  assign new_new_n34709__ = ~new_new_n34463__ & ~new_new_n34708__;
  assign new_new_n34710__ = ~new_new_n34703__ & ~new_new_n34709__;
  assign new_new_n34711__ = ~new_new_n34704__ & new_new_n34710__;
  assign new_new_n34712__ = new_new_n34700__ & ~new_new_n34711__;
  assign new_new_n34713__ = ~new_new_n34700__ & new_new_n34711__;
  assign new_new_n34714__ = ~new_new_n34712__ & ~new_new_n34713__;
  assign new_new_n34715__ = ~new_new_n34668__ & ~new_new_n34673__;
  assign new_new_n34716__ = ~new_new_n34667__ & ~new_new_n34715__;
  assign new_new_n34717__ = ~new_new_n34481__ & ~new_new_n34663__;
  assign new_new_n34718__ = ~new_new_n34482__ & ~new_new_n34717__;
  assign new_new_n34719__ = ~pi05 & new_new_n34718__;
  assign new_new_n34720__ = pi05 & ~new_new_n34718__;
  assign new_new_n34721__ = ~new_new_n34719__ & ~new_new_n34720__;
  assign new_new_n34722__ = new_new_n10698__ & new_new_n32740__;
  assign new_new_n34723__ = new_new_n10702__ & new_new_n32729__;
  assign new_new_n34724__ = ~new_new_n11409__ & new_new_n32382__;
  assign new_new_n34725__ = ~new_new_n34723__ & ~new_new_n34724__;
  assign new_new_n34726__ = ~new_new_n34722__ & new_new_n34725__;
  assign new_new_n34727__ = new_new_n10694__ & new_new_n33050__;
  assign new_new_n34728__ = ~pi08 & ~new_new_n34727__;
  assign new_new_n34729__ = new_new_n12121__ & new_new_n33050__;
  assign new_new_n34730__ = ~new_new_n34728__ & ~new_new_n34729__;
  assign new_new_n34731__ = new_new_n34726__ & ~new_new_n34730__;
  assign new_new_n34732__ = pi08 & ~new_new_n34726__;
  assign new_new_n34733__ = ~new_new_n34731__ & ~new_new_n34732__;
  assign new_new_n34734__ = new_new_n8858__ & ~new_new_n26667__;
  assign new_new_n34735__ = ~new_new_n8479__ & new_new_n26698__;
  assign new_new_n34736__ = new_new_n8474__ & ~new_new_n26674__;
  assign new_new_n34737__ = new_new_n8470__ & ~new_new_n32340__;
  assign new_new_n34738__ = ~new_new_n34735__ & ~new_new_n34736__;
  assign new_new_n34739__ = ~new_new_n34734__ & new_new_n34738__;
  assign new_new_n34740__ = ~new_new_n34737__ & new_new_n34739__;
  assign new_new_n34741__ = ~new_new_n34624__ & ~new_new_n34637__;
  assign new_new_n34742__ = ~new_new_n34623__ & ~new_new_n34741__;
  assign new_new_n34743__ = new_new_n6991__ & new_new_n26722__;
  assign new_new_n34744__ = new_new_n6985__ & ~new_new_n27242__;
  assign new_new_n34745__ = ~new_new_n34743__ & ~new_new_n34744__;
  assign new_new_n34746__ = new_new_n6994__ & new_new_n27250__;
  assign new_new_n34747__ = ~new_new_n27271__ & new_new_n34746__;
  assign new_new_n34748__ = new_new_n34745__ & ~new_new_n34747__;
  assign new_new_n34749__ = pi14 & ~new_new_n34748__;
  assign new_new_n34750__ = ~pi13 & new_new_n27250__;
  assign new_new_n34751__ = new_new_n6994__ & ~new_new_n27278__;
  assign new_new_n34752__ = pi13 & ~new_new_n27271__;
  assign new_new_n34753__ = ~new_new_n34750__ & ~new_new_n34752__;
  assign new_new_n34754__ = new_new_n34751__ & new_new_n34753__;
  assign new_new_n34755__ = ~pi14 & new_new_n34745__;
  assign new_new_n34756__ = ~new_new_n34751__ & new_new_n34755__;
  assign new_new_n34757__ = ~new_new_n34749__ & ~new_new_n34754__;
  assign new_new_n34758__ = ~new_new_n34756__ & new_new_n34757__;
  assign new_new_n34759__ = ~new_new_n34742__ & new_new_n34758__;
  assign new_new_n34760__ = new_new_n34742__ & ~new_new_n34758__;
  assign new_new_n34761__ = ~new_new_n34759__ & ~new_new_n34760__;
  assign new_new_n34762__ = new_new_n6959__ & new_new_n30644__;
  assign new_new_n34763__ = new_new_n6964__ & new_new_n26810__;
  assign new_new_n34764__ = new_new_n6968__ & new_new_n26774__;
  assign new_new_n34765__ = ~new_new_n34763__ & ~new_new_n34764__;
  assign new_new_n34766__ = ~new_new_n34762__ & new_new_n34765__;
  assign new_new_n34767__ = new_new_n6958__ & new_new_n26729__;
  assign new_new_n34768__ = ~pi17 & ~new_new_n34767__;
  assign new_new_n34769__ = new_new_n7942__ & new_new_n26729__;
  assign new_new_n34770__ = ~new_new_n34768__ & ~new_new_n34769__;
  assign new_new_n34771__ = new_new_n34766__ & ~new_new_n34770__;
  assign new_new_n34772__ = pi17 & ~new_new_n34766__;
  assign new_new_n34773__ = ~new_new_n34771__ & ~new_new_n34772__;
  assign new_new_n34774__ = ~new_new_n34523__ & new_new_n34619__;
  assign new_new_n34775__ = ~new_new_n34522__ & ~new_new_n34774__;
  assign new_new_n34776__ = new_new_n34773__ & new_new_n34775__;
  assign new_new_n34777__ = ~new_new_n34773__ & ~new_new_n34775__;
  assign new_new_n34778__ = ~new_new_n34776__ & ~new_new_n34777__;
  assign new_new_n34779__ = ~new_new_n34539__ & new_new_n34616__;
  assign new_new_n34780__ = ~new_new_n34540__ & ~new_new_n34779__;
  assign new_new_n34781__ = new_new_n5213__ & ~new_new_n26823__;
  assign new_new_n34782__ = new_new_n5191__ & ~new_new_n26854__;
  assign new_new_n34783__ = new_new_n5183__ & new_new_n26847__;
  assign new_new_n34784__ = new_new_n5215__ & ~new_new_n29400__;
  assign new_new_n34785__ = ~new_new_n34782__ & ~new_new_n34783__;
  assign new_new_n34786__ = ~new_new_n34781__ & new_new_n34785__;
  assign new_new_n34787__ = ~new_new_n34784__ & new_new_n34786__;
  assign new_new_n34788__ = pi23 & ~new_new_n34787__;
  assign new_new_n34789__ = ~pi23 & new_new_n34787__;
  assign new_new_n34790__ = ~new_new_n34788__ & ~new_new_n34789__;
  assign new_new_n34791__ = ~new_new_n34609__ & ~new_new_n34616__;
  assign new_new_n34792__ = ~new_new_n34608__ & ~new_new_n34791__;
  assign new_new_n34793__ = ~new_new_n34790__ & new_new_n34792__;
  assign new_new_n34794__ = new_new_n34790__ & ~new_new_n34792__;
  assign new_new_n34795__ = ~new_new_n34793__ & ~new_new_n34794__;
  assign new_new_n34796__ = new_new_n3311__ & ~new_new_n26888__;
  assign new_new_n34797__ = ~new_new_n333__ & ~new_new_n27168__;
  assign new_new_n34798__ = new_new_n873__ & new_new_n26922__;
  assign new_new_n34799__ = ~new_new_n34797__ & ~new_new_n34798__;
  assign new_new_n34800__ = ~new_new_n34796__ & new_new_n34799__;
  assign new_new_n34801__ = pi26 & ~new_new_n34800__;
  assign new_new_n34802__ = new_new_n4898__ & new_new_n27180__;
  assign new_new_n34803__ = new_new_n801__ & new_new_n27180__;
  assign new_new_n34804__ = ~pi26 & ~new_new_n34803__;
  assign new_new_n34805__ = ~new_new_n34802__ & ~new_new_n34804__;
  assign new_new_n34806__ = new_new_n34800__ & ~new_new_n34805__;
  assign new_new_n34807__ = ~new_new_n34801__ & ~new_new_n34806__;
  assign new_new_n34808__ = new_new_n161__ & ~new_new_n26937__;
  assign new_new_n34809__ = new_new_n765__ & new_new_n27152__;
  assign new_new_n34810__ = ~new_new_n34808__ & ~new_new_n34809__;
  assign new_new_n34811__ = ~pi31 & ~new_new_n34810__;
  assign new_new_n34812__ = ~new_new_n71__ & ~new_new_n27480__;
  assign new_new_n34813__ = ~new_new_n161__ & ~new_new_n26937__;
  assign new_new_n34814__ = ~new_new_n34812__ & new_new_n34813__;
  assign new_new_n34815__ = new_new_n161__ & new_new_n27152__;
  assign new_new_n34816__ = new_new_n26937__ & ~new_new_n34815__;
  assign new_new_n34817__ = new_new_n34812__ & new_new_n34816__;
  assign new_new_n34818__ = ~new_new_n34561__ & ~new_new_n34814__;
  assign new_new_n34819__ = ~new_new_n34817__ & new_new_n34818__;
  assign new_new_n34820__ = pi31 & ~new_new_n34819__;
  assign new_new_n34821__ = ~new_new_n34811__ & ~new_new_n34820__;
  assign new_new_n34822__ = ~new_new_n34574__ & new_new_n34607__;
  assign new_new_n34823__ = ~new_new_n34573__ & ~new_new_n34822__;
  assign new_new_n34824__ = new_new_n34821__ & ~new_new_n34823__;
  assign new_new_n34825__ = ~new_new_n34821__ & new_new_n34823__;
  assign new_new_n34826__ = ~new_new_n34824__ & ~new_new_n34825__;
  assign new_new_n34827__ = ~new_new_n34580__ & ~new_new_n34601__;
  assign new_new_n34828__ = ~pi02 & new_new_n34827__;
  assign new_new_n34829__ = new_new_n34580__ & new_new_n34601__;
  assign new_new_n34830__ = pi02 & new_new_n34829__;
  assign new_new_n34831__ = ~new_new_n34828__ & ~new_new_n34830__;
  assign new_new_n34832__ = ~new_new_n250__ & ~new_new_n336__;
  assign new_new_n34833__ = ~new_new_n1372__ & new_new_n34832__;
  assign new_new_n34834__ = ~new_new_n276__ & ~new_new_n961__;
  assign new_new_n34835__ = ~new_new_n2329__ & new_new_n34834__;
  assign new_new_n34836__ = new_new_n748__ & new_new_n34833__;
  assign new_new_n34837__ = ~new_new_n809__ & new_new_n870__;
  assign new_new_n34838__ = new_new_n1665__ & new_new_n2911__;
  assign new_new_n34839__ = new_new_n3202__ & new_new_n34838__;
  assign new_new_n34840__ = new_new_n34836__ & new_new_n34837__;
  assign new_new_n34841__ = new_new_n1805__ & new_new_n34835__;
  assign new_new_n34842__ = new_new_n1826__ & new_new_n4509__;
  assign new_new_n34843__ = new_new_n34841__ & new_new_n34842__;
  assign new_new_n34844__ = new_new_n34839__ & new_new_n34840__;
  assign new_new_n34845__ = new_new_n6247__ & new_new_n34844__;
  assign new_new_n34846__ = new_new_n1305__ & new_new_n34843__;
  assign new_new_n34847__ = new_new_n34845__ & new_new_n34846__;
  assign new_new_n34848__ = new_new_n2864__ & new_new_n34847__;
  assign new_new_n34849__ = new_new_n1446__ & new_new_n34848__;
  assign new_new_n34850__ = new_new_n34831__ & ~new_new_n34849__;
  assign new_new_n34851__ = ~new_new_n34831__ & new_new_n34849__;
  assign new_new_n34852__ = ~new_new_n34850__ & ~new_new_n34851__;
  assign new_new_n34853__ = new_new_n34826__ & new_new_n34852__;
  assign new_new_n34854__ = ~new_new_n34826__ & ~new_new_n34852__;
  assign new_new_n34855__ = ~new_new_n34853__ & ~new_new_n34854__;
  assign new_new_n34856__ = new_new_n34807__ & ~new_new_n34855__;
  assign new_new_n34857__ = ~new_new_n34807__ & new_new_n34855__;
  assign new_new_n34858__ = ~new_new_n34856__ & ~new_new_n34857__;
  assign new_new_n34859__ = new_new_n4815__ & new_new_n26917__;
  assign new_new_n34860__ = ~new_new_n4818__ & ~new_new_n26941__;
  assign new_new_n34861__ = new_new_n4212__ & new_new_n26928__;
  assign new_new_n34862__ = ~new_new_n34860__ & ~new_new_n34861__;
  assign new_new_n34863__ = ~new_new_n34859__ & new_new_n34862__;
  assign new_new_n34864__ = new_new_n4214__ & ~new_new_n27462__;
  assign new_new_n34865__ = ~pi29 & ~new_new_n34864__;
  assign new_new_n34866__ = new_new_n5732__ & ~new_new_n27462__;
  assign new_new_n34867__ = ~new_new_n34865__ & ~new_new_n34866__;
  assign new_new_n34868__ = new_new_n34863__ & ~new_new_n34867__;
  assign new_new_n34869__ = pi29 & ~new_new_n34863__;
  assign new_new_n34870__ = ~new_new_n34868__ & ~new_new_n34869__;
  assign new_new_n34871__ = new_new_n34858__ & ~new_new_n34870__;
  assign new_new_n34872__ = ~new_new_n34858__ & new_new_n34870__;
  assign new_new_n34873__ = ~new_new_n34871__ & ~new_new_n34872__;
  assign new_new_n34874__ = new_new_n34795__ & ~new_new_n34873__;
  assign new_new_n34875__ = ~new_new_n34795__ & new_new_n34873__;
  assign new_new_n34876__ = ~new_new_n34874__ & ~new_new_n34875__;
  assign new_new_n34877__ = ~new_new_n34780__ & new_new_n34876__;
  assign new_new_n34878__ = new_new_n34780__ & ~new_new_n34876__;
  assign new_new_n34879__ = ~new_new_n34877__ & ~new_new_n34878__;
  assign new_new_n34880__ = new_new_n6629__ & ~new_new_n26741__;
  assign new_new_n34881__ = ~new_new_n6625__ & ~new_new_n27221__;
  assign new_new_n34882__ = new_new_n6633__ & new_new_n26802__;
  assign new_new_n34883__ = ~new_new_n6633__ & ~new_new_n30411__;
  assign new_new_n34884__ = new_new_n6631__ & ~new_new_n34882__;
  assign new_new_n34885__ = ~new_new_n34883__ & new_new_n34884__;
  assign new_new_n34886__ = ~new_new_n34880__ & ~new_new_n34881__;
  assign new_new_n34887__ = ~new_new_n34885__ & new_new_n34886__;
  assign new_new_n34888__ = ~pi20 & new_new_n34887__;
  assign new_new_n34889__ = pi20 & ~new_new_n34887__;
  assign new_new_n34890__ = ~new_new_n34888__ & ~new_new_n34889__;
  assign new_new_n34891__ = new_new_n34879__ & new_new_n34890__;
  assign new_new_n34892__ = ~new_new_n34879__ & ~new_new_n34890__;
  assign new_new_n34893__ = ~new_new_n34891__ & ~new_new_n34892__;
  assign new_new_n34894__ = new_new_n34778__ & ~new_new_n34893__;
  assign new_new_n34895__ = ~new_new_n34778__ & new_new_n34893__;
  assign new_new_n34896__ = ~new_new_n34894__ & ~new_new_n34895__;
  assign new_new_n34897__ = new_new_n34761__ & ~new_new_n34896__;
  assign new_new_n34898__ = ~new_new_n34761__ & new_new_n34896__;
  assign new_new_n34899__ = ~new_new_n34897__ & ~new_new_n34898__;
  assign new_new_n34900__ = ~new_new_n34505__ & new_new_n34640__;
  assign new_new_n34901__ = ~new_new_n34506__ & ~new_new_n34900__;
  assign new_new_n34902__ = new_new_n34899__ & ~new_new_n34901__;
  assign new_new_n34903__ = ~new_new_n34899__ & new_new_n34901__;
  assign new_new_n34904__ = ~new_new_n34902__ & ~new_new_n34903__;
  assign new_new_n34905__ = pi11 & ~new_new_n34904__;
  assign new_new_n34906__ = ~pi11 & new_new_n34904__;
  assign new_new_n34907__ = ~new_new_n34905__ & ~new_new_n34906__;
  assign new_new_n34908__ = new_new_n34740__ & new_new_n34907__;
  assign new_new_n34909__ = ~new_new_n34740__ & ~new_new_n34907__;
  assign new_new_n34910__ = ~new_new_n34908__ & ~new_new_n34909__;
  assign new_new_n34911__ = new_new_n34733__ & new_new_n34910__;
  assign new_new_n34912__ = ~new_new_n34733__ & ~new_new_n34910__;
  assign new_new_n34913__ = ~new_new_n34911__ & ~new_new_n34912__;
  assign new_new_n34914__ = ~new_new_n34647__ & ~new_new_n34660__;
  assign new_new_n34915__ = ~new_new_n34646__ & ~new_new_n34914__;
  assign new_new_n34916__ = ~new_new_n34913__ & new_new_n34915__;
  assign new_new_n34917__ = ~new_new_n34912__ & ~new_new_n34915__;
  assign new_new_n34918__ = ~new_new_n34911__ & new_new_n34917__;
  assign new_new_n34919__ = ~new_new_n34916__ & ~new_new_n34918__;
  assign new_new_n34920__ = new_new_n34721__ & ~new_new_n34919__;
  assign new_new_n34921__ = ~new_new_n34721__ & new_new_n34919__;
  assign new_new_n34922__ = ~new_new_n34920__ & ~new_new_n34921__;
  assign new_new_n34923__ = ~new_new_n34716__ & ~new_new_n34922__;
  assign new_new_n34924__ = new_new_n34716__ & new_new_n34922__;
  assign new_new_n34925__ = ~new_new_n34923__ & ~new_new_n34924__;
  assign new_new_n34926__ = new_new_n34714__ & ~new_new_n34925__;
  assign new_new_n34927__ = ~new_new_n34714__ & new_new_n34925__;
  assign po09 = new_new_n34926__ | new_new_n34927__;
  assign new_new_n34929__ = new_new_n34712__ & new_new_n34923__;
  assign new_new_n34930__ = new_new_n34700__ & new_new_n34925__;
  assign new_new_n34931__ = new_new_n34711__ & new_new_n34716__;
  assign new_new_n34932__ = ~new_new_n34930__ & new_new_n34931__;
  assign new_new_n34933__ = ~new_new_n34742__ & ~new_new_n34758__;
  assign new_new_n34934__ = ~new_new_n34898__ & ~new_new_n34933__;
  assign new_new_n34935__ = new_new_n6985__ & new_new_n27250__;
  assign new_new_n34936__ = new_new_n6991__ & ~new_new_n27242__;
  assign new_new_n34937__ = ~new_new_n34935__ & ~new_new_n34936__;
  assign new_new_n34938__ = new_new_n6994__ & new_new_n26698__;
  assign new_new_n34939__ = new_new_n31511__ & new_new_n34938__;
  assign new_new_n34940__ = new_new_n34937__ & ~new_new_n34939__;
  assign new_new_n34941__ = pi14 & ~new_new_n34940__;
  assign new_new_n34942__ = ~pi13 & ~new_new_n34204__;
  assign new_new_n34943__ = pi13 & ~new_new_n31509__;
  assign new_new_n34944__ = new_new_n6994__ & ~new_new_n34942__;
  assign new_new_n34945__ = ~new_new_n34943__ & new_new_n34944__;
  assign new_new_n34946__ = new_new_n6994__ & ~new_new_n31510__;
  assign new_new_n34947__ = ~pi14 & new_new_n34937__;
  assign new_new_n34948__ = ~new_new_n34946__ & new_new_n34947__;
  assign new_new_n34949__ = ~new_new_n34945__ & ~new_new_n34948__;
  assign new_new_n34950__ = ~new_new_n34941__ & new_new_n34949__;
  assign new_new_n34951__ = new_new_n34934__ & ~new_new_n34950__;
  assign new_new_n34952__ = ~new_new_n34934__ & new_new_n34950__;
  assign new_new_n34953__ = ~new_new_n34951__ & ~new_new_n34952__;
  assign new_new_n34954__ = ~new_new_n34776__ & ~new_new_n34893__;
  assign new_new_n34955__ = ~new_new_n34777__ & ~new_new_n34954__;
  assign new_new_n34956__ = new_new_n5213__ & ~new_new_n27221__;
  assign new_new_n34957__ = new_new_n5183__ & ~new_new_n26823__;
  assign new_new_n34958__ = new_new_n5191__ & new_new_n26847__;
  assign new_new_n34959__ = new_new_n5215__ & new_new_n27411__;
  assign new_new_n34960__ = ~new_new_n34957__ & ~new_new_n34958__;
  assign new_new_n34961__ = ~new_new_n34956__ & new_new_n34960__;
  assign new_new_n34962__ = ~new_new_n34959__ & new_new_n34961__;
  assign new_new_n34963__ = pi23 & ~new_new_n34962__;
  assign new_new_n34964__ = ~pi23 & new_new_n34962__;
  assign new_new_n34965__ = ~new_new_n34963__ & ~new_new_n34964__;
  assign new_new_n34966__ = ~new_new_n34793__ & ~new_new_n34873__;
  assign new_new_n34967__ = ~new_new_n34794__ & ~new_new_n34966__;
  assign new_new_n34968__ = new_new_n34965__ & ~new_new_n34967__;
  assign new_new_n34969__ = ~new_new_n34965__ & new_new_n34967__;
  assign new_new_n34970__ = ~new_new_n34968__ & ~new_new_n34969__;
  assign new_new_n34971__ = ~new_new_n4900__ & ~new_new_n27430__;
  assign new_new_n34972__ = ~new_new_n333__ & new_new_n26922__;
  assign new_new_n34973__ = new_new_n873__ & ~new_new_n26888__;
  assign new_new_n34974__ = ~new_new_n34972__ & ~new_new_n34973__;
  assign new_new_n34975__ = ~new_new_n34971__ & new_new_n34974__;
  assign new_new_n34976__ = pi26 & ~new_new_n34975__;
  assign new_new_n34977__ = new_new_n512__ & ~new_new_n26854__;
  assign new_new_n34978__ = new_new_n801__ & ~new_new_n26854__;
  assign new_new_n34979__ = ~pi26 & ~new_new_n34978__;
  assign new_new_n34980__ = ~new_new_n34977__ & ~new_new_n34979__;
  assign new_new_n34981__ = new_new_n34975__ & ~new_new_n34980__;
  assign new_new_n34982__ = ~new_new_n34976__ & ~new_new_n34981__;
  assign new_new_n34983__ = ~new_new_n34857__ & new_new_n34870__;
  assign new_new_n34984__ = ~new_new_n34856__ & ~new_new_n34983__;
  assign new_new_n34985__ = new_new_n4212__ & new_new_n26917__;
  assign new_new_n34986__ = ~new_new_n4818__ & new_new_n26928__;
  assign new_new_n34987__ = new_new_n4815__ & ~new_new_n27168__;
  assign new_new_n34988__ = ~new_new_n34986__ & ~new_new_n34987__;
  assign new_new_n34989__ = ~new_new_n34985__ & new_new_n34988__;
  assign new_new_n34990__ = new_new_n4214__ & ~new_new_n28799__;
  assign new_new_n34991__ = pi29 & ~new_new_n34990__;
  assign new_new_n34992__ = new_new_n4825__ & ~new_new_n28799__;
  assign new_new_n34993__ = ~new_new_n34991__ & ~new_new_n34992__;
  assign new_new_n34994__ = new_new_n34989__ & ~new_new_n34993__;
  assign new_new_n34995__ = ~pi29 & ~new_new_n34989__;
  assign new_new_n34996__ = ~new_new_n34994__ & ~new_new_n34995__;
  assign new_new_n34997__ = ~new_new_n34824__ & ~new_new_n34852__;
  assign new_new_n34998__ = ~new_new_n34825__ & ~new_new_n34997__;
  assign new_new_n34999__ = ~new_new_n34830__ & new_new_n34849__;
  assign new_new_n35000__ = ~new_new_n34828__ & ~new_new_n34849__;
  assign new_new_n35001__ = ~new_new_n34999__ & ~new_new_n35000__;
  assign new_new_n35002__ = ~new_new_n438__ & ~new_new_n603__;
  assign new_new_n35003__ = ~new_new_n843__ & ~new_new_n995__;
  assign new_new_n35004__ = new_new_n35002__ & new_new_n35003__;
  assign new_new_n35005__ = ~new_new_n322__ & new_new_n777__;
  assign new_new_n35006__ = ~new_new_n1217__ & new_new_n1337__;
  assign new_new_n35007__ = new_new_n35005__ & new_new_n35006__;
  assign new_new_n35008__ = new_new_n589__ & new_new_n35004__;
  assign new_new_n35009__ = new_new_n1256__ & new_new_n1849__;
  assign new_new_n35010__ = new_new_n2004__ & new_new_n2322__;
  assign new_new_n35011__ = new_new_n35009__ & new_new_n35010__;
  assign new_new_n35012__ = new_new_n35007__ & new_new_n35008__;
  assign new_new_n35013__ = new_new_n35011__ & new_new_n35012__;
  assign new_new_n35014__ = new_new_n16849__ & new_new_n35013__;
  assign new_new_n35015__ = new_new_n28583__ & new_new_n35014__;
  assign new_new_n35016__ = new_new_n4252__ & new_new_n35015__;
  assign new_new_n35017__ = new_new_n2257__ & new_new_n35016__;
  assign new_new_n35018__ = pi05 & ~new_new_n35017__;
  assign new_new_n35019__ = ~pi05 & new_new_n35017__;
  assign new_new_n35020__ = ~new_new_n35018__ & ~new_new_n35019__;
  assign new_new_n35021__ = ~new_new_n26941__ & new_new_n27152__;
  assign new_new_n35022__ = new_new_n26941__ & new_new_n27128__;
  assign new_new_n35023__ = ~new_new_n27152__ & new_new_n35022__;
  assign new_new_n35024__ = ~new_new_n161__ & ~new_new_n35021__;
  assign new_new_n35025__ = ~new_new_n35023__ & new_new_n35024__;
  assign new_new_n35026__ = ~new_new_n26937__ & ~new_new_n35025__;
  assign new_new_n35027__ = new_new_n26937__ & new_new_n27152__;
  assign new_new_n35028__ = new_new_n26941__ & ~new_new_n35027__;
  assign new_new_n35029__ = ~new_new_n35021__ & ~new_new_n35028__;
  assign new_new_n35030__ = ~new_new_n27128__ & ~new_new_n35029__;
  assign new_new_n35031__ = ~new_new_n161__ & ~new_new_n27476__;
  assign new_new_n35032__ = ~new_new_n35022__ & new_new_n35031__;
  assign new_new_n35033__ = ~new_new_n35030__ & new_new_n35032__;
  assign new_new_n35034__ = new_new_n4147__ & ~new_new_n35026__;
  assign new_new_n35035__ = ~new_new_n35033__ & new_new_n35034__;
  assign new_new_n35036__ = ~new_new_n71__ & new_new_n34815__;
  assign new_new_n35037__ = new_new_n71__ & ~new_new_n27152__;
  assign new_new_n35038__ = pi31 & ~new_new_n35037__;
  assign new_new_n35039__ = ~new_new_n15853__ & ~new_new_n26941__;
  assign new_new_n35040__ = ~new_new_n35036__ & ~new_new_n35039__;
  assign new_new_n35041__ = ~new_new_n35038__ & new_new_n35040__;
  assign new_new_n35042__ = ~new_new_n35035__ & ~new_new_n35041__;
  assign new_new_n35043__ = new_new_n35020__ & ~new_new_n35042__;
  assign new_new_n35044__ = ~new_new_n35020__ & new_new_n35042__;
  assign new_new_n35045__ = ~new_new_n35043__ & ~new_new_n35044__;
  assign new_new_n35046__ = new_new_n35001__ & new_new_n35045__;
  assign new_new_n35047__ = ~new_new_n35001__ & ~new_new_n35045__;
  assign new_new_n35048__ = ~new_new_n35046__ & ~new_new_n35047__;
  assign new_new_n35049__ = ~new_new_n34998__ & ~new_new_n35048__;
  assign new_new_n35050__ = new_new_n34998__ & new_new_n35048__;
  assign new_new_n35051__ = ~new_new_n35049__ & ~new_new_n35050__;
  assign new_new_n35052__ = new_new_n34996__ & new_new_n35051__;
  assign new_new_n35053__ = ~new_new_n34996__ & ~new_new_n35051__;
  assign new_new_n35054__ = ~new_new_n35052__ & ~new_new_n35053__;
  assign new_new_n35055__ = new_new_n34984__ & new_new_n35054__;
  assign new_new_n35056__ = ~new_new_n34984__ & ~new_new_n35054__;
  assign new_new_n35057__ = ~new_new_n35055__ & ~new_new_n35056__;
  assign new_new_n35058__ = new_new_n34982__ & ~new_new_n35057__;
  assign new_new_n35059__ = ~new_new_n34982__ & new_new_n35057__;
  assign new_new_n35060__ = ~new_new_n35058__ & ~new_new_n35059__;
  assign new_new_n35061__ = new_new_n34970__ & ~new_new_n35060__;
  assign new_new_n35062__ = ~new_new_n34970__ & new_new_n35060__;
  assign new_new_n35063__ = ~new_new_n35061__ & ~new_new_n35062__;
  assign new_new_n35064__ = ~new_new_n34877__ & ~new_new_n34890__;
  assign new_new_n35065__ = ~new_new_n34878__ & ~new_new_n35064__;
  assign new_new_n35066__ = ~new_new_n35063__ & ~new_new_n35065__;
  assign new_new_n35067__ = new_new_n35063__ & new_new_n35065__;
  assign new_new_n35068__ = ~new_new_n35066__ & ~new_new_n35067__;
  assign new_new_n35069__ = new_new_n6629__ & ~new_new_n26802__;
  assign new_new_n35070__ = ~new_new_n6625__ & ~new_new_n26741__;
  assign new_new_n35071__ = new_new_n6936__ & new_new_n27395__;
  assign new_new_n35072__ = ~new_new_n35069__ & ~new_new_n35070__;
  assign new_new_n35073__ = ~new_new_n35071__ & new_new_n35072__;
  assign new_new_n35074__ = new_new_n6631__ & new_new_n26810__;
  assign new_new_n35075__ = pi20 & ~new_new_n35074__;
  assign new_new_n35076__ = new_new_n7015__ & new_new_n26810__;
  assign new_new_n35077__ = ~new_new_n35075__ & ~new_new_n35076__;
  assign new_new_n35078__ = new_new_n35073__ & ~new_new_n35077__;
  assign new_new_n35079__ = ~pi20 & ~new_new_n35073__;
  assign new_new_n35080__ = ~new_new_n35078__ & ~new_new_n35079__;
  assign new_new_n35081__ = new_new_n35068__ & ~new_new_n35080__;
  assign new_new_n35082__ = ~new_new_n35068__ & new_new_n35080__;
  assign new_new_n35083__ = ~new_new_n35081__ & ~new_new_n35082__;
  assign new_new_n35084__ = new_new_n7935__ & new_new_n26722__;
  assign new_new_n35085__ = new_new_n6964__ & new_new_n26774__;
  assign new_new_n35086__ = new_new_n6968__ & new_new_n26729__;
  assign new_new_n35087__ = ~new_new_n35085__ & ~new_new_n35086__;
  assign new_new_n35088__ = ~new_new_n35084__ & new_new_n35087__;
  assign new_new_n35089__ = new_new_n6958__ & ~new_new_n27348__;
  assign new_new_n35090__ = ~pi17 & ~new_new_n35089__;
  assign new_new_n35091__ = new_new_n8160__ & ~new_new_n27348__;
  assign new_new_n35092__ = ~new_new_n35090__ & ~new_new_n35091__;
  assign new_new_n35093__ = new_new_n35088__ & ~new_new_n35092__;
  assign new_new_n35094__ = pi17 & ~new_new_n35088__;
  assign new_new_n35095__ = ~new_new_n35093__ & ~new_new_n35094__;
  assign new_new_n35096__ = new_new_n35083__ & new_new_n35095__;
  assign new_new_n35097__ = ~new_new_n35083__ & ~new_new_n35095__;
  assign new_new_n35098__ = ~new_new_n35096__ & ~new_new_n35097__;
  assign new_new_n35099__ = new_new_n34955__ & new_new_n35098__;
  assign new_new_n35100__ = ~new_new_n34955__ & ~new_new_n35098__;
  assign new_new_n35101__ = ~new_new_n35099__ & ~new_new_n35100__;
  assign new_new_n35102__ = ~new_new_n34953__ & ~new_new_n35101__;
  assign new_new_n35103__ = new_new_n34953__ & new_new_n35101__;
  assign new_new_n35104__ = ~new_new_n35102__ & ~new_new_n35103__;
  assign new_new_n35105__ = ~new_new_n34911__ & ~new_new_n34917__;
  assign new_new_n35106__ = ~new_new_n34902__ & ~new_new_n34910__;
  assign new_new_n35107__ = ~new_new_n34903__ & ~new_new_n35106__;
  assign new_new_n35108__ = ~new_new_n35105__ & new_new_n35107__;
  assign new_new_n35109__ = new_new_n35105__ & ~new_new_n35107__;
  assign new_new_n35110__ = ~new_new_n35108__ & ~new_new_n35109__;
  assign new_new_n35111__ = ~new_new_n17566__ & ~new_new_n17567__;
  assign new_new_n35112__ = ~new_new_n32729__ & ~new_new_n35111__;
  assign new_new_n35113__ = ~pi07 & ~new_new_n34178__;
  assign new_new_n35114__ = ~new_new_n9697__ & ~new_new_n10695__;
  assign new_new_n35115__ = ~new_new_n35113__ & new_new_n35114__;
  assign new_new_n35116__ = pi07 & ~new_new_n34178__;
  assign new_new_n35117__ = ~new_new_n9701__ & ~new_new_n10696__;
  assign new_new_n35118__ = ~new_new_n35116__ & new_new_n35117__;
  assign new_new_n35119__ = ~new_new_n34723__ & ~new_new_n35112__;
  assign new_new_n35120__ = ~new_new_n35115__ & new_new_n35119__;
  assign new_new_n35121__ = ~new_new_n35118__ & new_new_n35120__;
  assign new_new_n35122__ = pi08 & ~new_new_n35121__;
  assign new_new_n35123__ = ~pi08 & new_new_n35121__;
  assign new_new_n35124__ = ~new_new_n35122__ & ~new_new_n35123__;
  assign new_new_n35125__ = new_new_n8474__ & ~new_new_n26667__;
  assign new_new_n35126__ = new_new_n8858__ & new_new_n32382__;
  assign new_new_n35127__ = ~new_new_n8479__ & ~new_new_n26674__;
  assign new_new_n35128__ = new_new_n8470__ & ~new_new_n33347__;
  assign new_new_n35129__ = ~new_new_n35126__ & ~new_new_n35127__;
  assign new_new_n35130__ = ~new_new_n35128__ & new_new_n35129__;
  assign new_new_n35131__ = ~new_new_n35125__ & new_new_n35130__;
  assign new_new_n35132__ = ~pi11 & ~new_new_n35131__;
  assign new_new_n35133__ = ~new_new_n8858__ & new_new_n26667__;
  assign new_new_n35134__ = new_new_n8474__ & ~new_new_n35133__;
  assign new_new_n35135__ = pi11 & ~new_new_n35134__;
  assign new_new_n35136__ = new_new_n35130__ & new_new_n35135__;
  assign new_new_n35137__ = ~new_new_n35132__ & ~new_new_n35136__;
  assign new_new_n35138__ = new_new_n35124__ & new_new_n35137__;
  assign new_new_n35139__ = ~new_new_n35124__ & ~new_new_n35137__;
  assign new_new_n35140__ = ~new_new_n35138__ & ~new_new_n35139__;
  assign new_new_n35141__ = new_new_n35110__ & ~new_new_n35140__;
  assign new_new_n35142__ = ~new_new_n35110__ & new_new_n35140__;
  assign new_new_n35143__ = ~new_new_n35141__ & ~new_new_n35142__;
  assign new_new_n35144__ = new_new_n35104__ & new_new_n35143__;
  assign new_new_n35145__ = ~new_new_n35104__ & ~new_new_n35143__;
  assign new_new_n35146__ = ~new_new_n35144__ & ~new_new_n35145__;
  assign new_new_n35147__ = ~new_new_n34719__ & new_new_n34919__;
  assign new_new_n35148__ = ~new_new_n34720__ & ~new_new_n35147__;
  assign new_new_n35149__ = ~new_new_n35146__ & ~new_new_n35148__;
  assign new_new_n35150__ = ~new_new_n34720__ & new_new_n35146__;
  assign new_new_n35151__ = ~new_new_n35147__ & new_new_n35150__;
  assign new_new_n35152__ = ~new_new_n35149__ & ~new_new_n35151__;
  assign new_new_n35153__ = ~new_new_n34700__ & new_new_n34922__;
  assign new_new_n35154__ = po09 & new_new_n35153__;
  assign new_new_n35155__ = ~new_new_n34929__ & new_new_n35152__;
  assign new_new_n35156__ = ~new_new_n34932__ & new_new_n35155__;
  assign new_new_n35157__ = ~new_new_n35154__ & new_new_n35156__;
  assign new_new_n35158__ = ~new_new_n34711__ & ~po09;
  assign new_new_n35159__ = ~new_new_n34923__ & ~new_new_n35158__;
  assign new_new_n35160__ = ~new_new_n34929__ & ~new_new_n35159__;
  assign new_new_n35161__ = ~new_new_n34930__ & ~new_new_n35152__;
  assign new_new_n35162__ = ~new_new_n35160__ & new_new_n35161__;
  assign po10 = ~new_new_n35157__ & ~new_new_n35162__;
  assign new_new_n35164__ = ~new_new_n35105__ & ~new_new_n35124__;
  assign new_new_n35165__ = new_new_n35105__ & new_new_n35124__;
  assign new_new_n35166__ = ~new_new_n35104__ & ~new_new_n35107__;
  assign new_new_n35167__ = new_new_n35104__ & new_new_n35107__;
  assign new_new_n35168__ = ~new_new_n35166__ & ~new_new_n35167__;
  assign new_new_n35169__ = ~new_new_n35137__ & new_new_n35168__;
  assign new_new_n35170__ = new_new_n35137__ & ~new_new_n35168__;
  assign new_new_n35171__ = ~new_new_n35169__ & ~new_new_n35170__;
  assign new_new_n35172__ = ~new_new_n35165__ & new_new_n35171__;
  assign new_new_n35173__ = ~new_new_n35164__ & ~new_new_n35172__;
  assign new_new_n35174__ = ~new_new_n35137__ & ~new_new_n35167__;
  assign new_new_n35175__ = ~new_new_n35166__ & ~new_new_n35174__;
  assign new_new_n35176__ = new_new_n19825__ & new_new_n26698__;
  assign new_new_n35177__ = new_new_n19829__ & new_new_n27250__;
  assign new_new_n35178__ = ~new_new_n6994__ & ~new_new_n35177__;
  assign new_new_n35179__ = ~new_new_n35176__ & new_new_n35178__;
  assign new_new_n35180__ = new_new_n6994__ & new_new_n26674__;
  assign new_new_n35181__ = ~new_new_n27284__ & new_new_n35180__;
  assign new_new_n35182__ = ~new_new_n35179__ & ~new_new_n35181__;
  assign new_new_n35183__ = ~pi14 & ~new_new_n35182__;
  assign new_new_n35184__ = new_new_n6994__ & ~new_new_n27284__;
  assign new_new_n35185__ = pi14 & ~new_new_n35179__;
  assign new_new_n35186__ = ~new_new_n35180__ & new_new_n35185__;
  assign new_new_n35187__ = ~new_new_n35184__ & new_new_n35186__;
  assign new_new_n35188__ = new_new_n26674__ & new_new_n27284__;
  assign new_new_n35189__ = ~pi13 & ~new_new_n35188__;
  assign new_new_n35190__ = pi13 & ~new_new_n27288__;
  assign new_new_n35191__ = new_new_n6994__ & ~new_new_n35189__;
  assign new_new_n35192__ = ~new_new_n35190__ & new_new_n35191__;
  assign new_new_n35193__ = ~new_new_n35183__ & ~new_new_n35187__;
  assign new_new_n35194__ = ~new_new_n35192__ & new_new_n35193__;
  assign new_new_n35195__ = new_new_n6968__ & new_new_n26722__;
  assign new_new_n35196__ = new_new_n6964__ & new_new_n26729__;
  assign new_new_n35197__ = ~new_new_n35195__ & ~new_new_n35196__;
  assign new_new_n35198__ = new_new_n6958__ & ~new_new_n27362__;
  assign new_new_n35199__ = pi17 & ~new_new_n35198__;
  assign new_new_n35200__ = ~pi16 & new_new_n27242__;
  assign new_new_n35201__ = pi16 & ~new_new_n27242__;
  assign new_new_n35202__ = new_new_n6958__ & ~new_new_n35200__;
  assign new_new_n35203__ = ~new_new_n35201__ & new_new_n35202__;
  assign new_new_n35204__ = new_new_n27352__ & new_new_n35203__;
  assign new_new_n35205__ = ~new_new_n35199__ & ~new_new_n35204__;
  assign new_new_n35206__ = new_new_n35197__ & ~new_new_n35205__;
  assign new_new_n35207__ = new_new_n6958__ & new_new_n27353__;
  assign new_new_n35208__ = new_new_n35197__ & ~new_new_n35207__;
  assign new_new_n35209__ = ~pi17 & ~new_new_n35208__;
  assign new_new_n35210__ = ~new_new_n35206__ & ~new_new_n35209__;
  assign new_new_n35211__ = ~new_new_n35067__ & ~new_new_n35081__;
  assign new_new_n35212__ = new_new_n6634__ & new_new_n26774__;
  assign new_new_n35213__ = new_new_n6629__ & new_new_n26810__;
  assign new_new_n35214__ = ~new_new_n6625__ & ~new_new_n26802__;
  assign new_new_n35215__ = new_new_n6936__ & ~new_new_n27373__;
  assign new_new_n35216__ = ~new_new_n35213__ & ~new_new_n35214__;
  assign new_new_n35217__ = ~new_new_n35212__ & new_new_n35216__;
  assign new_new_n35218__ = ~new_new_n35215__ & new_new_n35217__;
  assign new_new_n35219__ = ~new_new_n34968__ & new_new_n35060__;
  assign new_new_n35220__ = ~new_new_n34969__ & ~new_new_n35219__;
  assign new_new_n35221__ = new_new_n5213__ & ~new_new_n26741__;
  assign new_new_n35222__ = new_new_n5191__ & ~new_new_n26823__;
  assign new_new_n35223__ = new_new_n5183__ & ~new_new_n27221__;
  assign new_new_n35224__ = new_new_n5215__ & new_new_n30393__;
  assign new_new_n35225__ = ~new_new_n35222__ & ~new_new_n35223__;
  assign new_new_n35226__ = ~new_new_n35221__ & new_new_n35225__;
  assign new_new_n35227__ = ~new_new_n35224__ & new_new_n35226__;
  assign new_new_n35228__ = pi23 & ~new_new_n35227__;
  assign new_new_n35229__ = ~pi23 & new_new_n35227__;
  assign new_new_n35230__ = ~new_new_n35228__ & ~new_new_n35229__;
  assign new_new_n35231__ = new_new_n180__ & new_new_n766__;
  assign new_new_n35232__ = ~new_new_n602__ & ~new_new_n1080__;
  assign new_new_n35233__ = ~new_new_n35231__ & new_new_n35232__;
  assign new_new_n35234__ = ~new_new_n1105__ & new_new_n2994__;
  assign new_new_n35235__ = new_new_n3026__ & new_new_n18536__;
  assign new_new_n35236__ = new_new_n35234__ & new_new_n35235__;
  assign new_new_n35237__ = new_new_n347__ & new_new_n35233__;
  assign new_new_n35238__ = ~new_new_n1539__ & new_new_n3560__;
  assign new_new_n35239__ = new_new_n35237__ & new_new_n35238__;
  assign new_new_n35240__ = new_new_n1175__ & new_new_n35236__;
  assign new_new_n35241__ = new_new_n7092__ & new_new_n7604__;
  assign new_new_n35242__ = new_new_n35240__ & new_new_n35241__;
  assign new_new_n35243__ = new_new_n35239__ & new_new_n35242__;
  assign new_new_n35244__ = ~new_new_n106__ & ~new_new_n249__;
  assign new_new_n35245__ = ~new_new_n472__ & new_new_n35244__;
  assign new_new_n35246__ = ~new_new_n166__ & ~new_new_n258__;
  assign new_new_n35247__ = ~new_new_n732__ & new_new_n948__;
  assign new_new_n35248__ = new_new_n2711__ & new_new_n35247__;
  assign new_new_n35249__ = new_new_n35245__ & new_new_n35246__;
  assign new_new_n35250__ = ~new_new_n809__ & new_new_n2379__;
  assign new_new_n35251__ = new_new_n2470__ & new_new_n3012__;
  assign new_new_n35252__ = new_new_n4236__ & new_new_n5282__;
  assign new_new_n35253__ = new_new_n35251__ & new_new_n35252__;
  assign new_new_n35254__ = new_new_n35249__ & new_new_n35250__;
  assign new_new_n35255__ = new_new_n7650__ & new_new_n35248__;
  assign new_new_n35256__ = new_new_n35254__ & new_new_n35255__;
  assign new_new_n35257__ = new_new_n1504__ & new_new_n35253__;
  assign new_new_n35258__ = new_new_n35256__ & new_new_n35257__;
  assign new_new_n35259__ = new_new_n2075__ & new_new_n35258__;
  assign new_new_n35260__ = new_new_n35243__ & new_new_n35259__;
  assign new_new_n35261__ = new_new_n1249__ & new_new_n35260__;
  assign new_new_n35262__ = ~new_new_n6811__ & ~new_new_n35017__;
  assign new_new_n35263__ = ~new_new_n6810__ & ~new_new_n35262__;
  assign new_new_n35264__ = new_new_n71__ & new_new_n26941__;
  assign new_new_n35265__ = new_new_n27441__ & ~new_new_n27481__;
  assign new_new_n35266__ = ~new_new_n161__ & ~new_new_n27159__;
  assign new_new_n35267__ = ~new_new_n35265__ & new_new_n35266__;
  assign new_new_n35268__ = ~new_new_n27152__ & ~new_new_n35267__;
  assign new_new_n35269__ = ~new_new_n26928__ & new_new_n28980__;
  assign new_new_n35270__ = new_new_n26928__ & ~new_new_n28980__;
  assign new_new_n35271__ = ~new_new_n161__ & ~new_new_n27483__;
  assign new_new_n35272__ = ~new_new_n35269__ & ~new_new_n35270__;
  assign new_new_n35273__ = new_new_n35271__ & new_new_n35272__;
  assign new_new_n35274__ = ~new_new_n35268__ & ~new_new_n35273__;
  assign new_new_n35275__ = ~new_new_n71__ & ~new_new_n35274__;
  assign new_new_n35276__ = pi31 & ~new_new_n35264__;
  assign new_new_n35277__ = ~new_new_n35275__ & new_new_n35276__;
  assign new_new_n35278__ = new_new_n161__ & new_new_n26941__;
  assign new_new_n35279__ = ~new_new_n161__ & ~new_new_n26928__;
  assign new_new_n35280__ = new_new_n4876__ & ~new_new_n35278__;
  assign new_new_n35281__ = ~new_new_n35279__ & new_new_n35280__;
  assign new_new_n35282__ = ~new_new_n35277__ & ~new_new_n35281__;
  assign new_new_n35283__ = ~new_new_n35263__ & new_new_n35282__;
  assign new_new_n35284__ = new_new_n35263__ & ~new_new_n35282__;
  assign new_new_n35285__ = ~new_new_n35283__ & ~new_new_n35284__;
  assign new_new_n35286__ = new_new_n35261__ & new_new_n35285__;
  assign new_new_n35287__ = ~new_new_n35261__ & ~new_new_n35285__;
  assign new_new_n35288__ = ~new_new_n35286__ & ~new_new_n35287__;
  assign new_new_n35289__ = pi02 & ~new_new_n35020__;
  assign new_new_n35290__ = new_new_n34827__ & ~new_new_n34849__;
  assign new_new_n35291__ = new_new_n35042__ & new_new_n35290__;
  assign new_new_n35292__ = ~new_new_n35289__ & ~new_new_n35291__;
  assign new_new_n35293__ = new_new_n34829__ & new_new_n34849__;
  assign new_new_n35294__ = ~new_new_n35042__ & new_new_n35293__;
  assign new_new_n35295__ = ~new_new_n35292__ & ~new_new_n35294__;
  assign new_new_n35296__ = ~new_new_n34830__ & new_new_n35042__;
  assign new_new_n35297__ = new_new_n34849__ & ~new_new_n35296__;
  assign new_new_n35298__ = ~new_new_n34828__ & ~new_new_n35042__;
  assign new_new_n35299__ = new_new_n35020__ & ~new_new_n35298__;
  assign new_new_n35300__ = ~new_new_n35297__ & new_new_n35299__;
  assign new_new_n35301__ = ~new_new_n35295__ & ~new_new_n35300__;
  assign new_new_n35302__ = ~new_new_n4818__ & new_new_n26917__;
  assign new_new_n35303__ = new_new_n4212__ & ~new_new_n27168__;
  assign new_new_n35304__ = new_new_n4815__ & new_new_n26922__;
  assign new_new_n35305__ = ~new_new_n35302__ & ~new_new_n35303__;
  assign new_new_n35306__ = ~new_new_n35304__ & new_new_n35305__;
  assign new_new_n35307__ = new_new_n4214__ & ~new_new_n29366__;
  assign new_new_n35308__ = pi29 & ~new_new_n35307__;
  assign new_new_n35309__ = new_new_n4825__ & ~new_new_n29366__;
  assign new_new_n35310__ = ~new_new_n35308__ & ~new_new_n35309__;
  assign new_new_n35311__ = new_new_n35306__ & ~new_new_n35310__;
  assign new_new_n35312__ = ~pi29 & ~new_new_n35306__;
  assign new_new_n35313__ = ~new_new_n35311__ & ~new_new_n35312__;
  assign new_new_n35314__ = ~new_new_n35301__ & ~new_new_n35313__;
  assign new_new_n35315__ = new_new_n35301__ & new_new_n35313__;
  assign new_new_n35316__ = ~new_new_n35314__ & ~new_new_n35315__;
  assign new_new_n35317__ = new_new_n35288__ & new_new_n35316__;
  assign new_new_n35318__ = ~new_new_n35288__ & ~new_new_n35316__;
  assign new_new_n35319__ = ~new_new_n35317__ & ~new_new_n35318__;
  assign new_new_n35320__ = ~new_new_n34996__ & ~new_new_n35050__;
  assign new_new_n35321__ = ~new_new_n35049__ & ~new_new_n35320__;
  assign new_new_n35322__ = ~new_new_n35319__ & ~new_new_n35321__;
  assign new_new_n35323__ = new_new_n35319__ & new_new_n35321__;
  assign new_new_n35324__ = ~new_new_n35322__ & ~new_new_n35323__;
  assign new_new_n35325__ = new_new_n3311__ & new_new_n26847__;
  assign new_new_n35326__ = new_new_n873__ & ~new_new_n26854__;
  assign new_new_n35327__ = ~new_new_n333__ & ~new_new_n26888__;
  assign new_new_n35328__ = ~new_new_n4900__ & new_new_n29424__;
  assign new_new_n35329__ = ~new_new_n35326__ & ~new_new_n35327__;
  assign new_new_n35330__ = ~new_new_n35325__ & new_new_n35329__;
  assign new_new_n35331__ = ~new_new_n35328__ & new_new_n35330__;
  assign new_new_n35332__ = pi26 & ~new_new_n35331__;
  assign new_new_n35333__ = ~pi26 & new_new_n35331__;
  assign new_new_n35334__ = ~new_new_n35332__ & ~new_new_n35333__;
  assign new_new_n35335__ = new_new_n35324__ & new_new_n35334__;
  assign new_new_n35336__ = ~new_new_n35324__ & ~new_new_n35334__;
  assign new_new_n35337__ = ~new_new_n35335__ & ~new_new_n35336__;
  assign new_new_n35338__ = ~new_new_n35230__ & ~new_new_n35337__;
  assign new_new_n35339__ = new_new_n35230__ & new_new_n35337__;
  assign new_new_n35340__ = ~new_new_n35338__ & ~new_new_n35339__;
  assign new_new_n35341__ = new_new_n34982__ & ~new_new_n35055__;
  assign new_new_n35342__ = ~new_new_n35056__ & ~new_new_n35341__;
  assign new_new_n35343__ = new_new_n35340__ & ~new_new_n35342__;
  assign new_new_n35344__ = ~new_new_n35340__ & new_new_n35342__;
  assign new_new_n35345__ = ~new_new_n35343__ & ~new_new_n35344__;
  assign new_new_n35346__ = new_new_n35220__ & new_new_n35345__;
  assign new_new_n35347__ = ~new_new_n35220__ & ~new_new_n35345__;
  assign new_new_n35348__ = ~new_new_n35346__ & ~new_new_n35347__;
  assign new_new_n35349__ = pi20 & ~new_new_n35348__;
  assign new_new_n35350__ = ~pi20 & new_new_n35348__;
  assign new_new_n35351__ = ~new_new_n35349__ & ~new_new_n35350__;
  assign new_new_n35352__ = new_new_n35218__ & new_new_n35351__;
  assign new_new_n35353__ = ~new_new_n35218__ & ~new_new_n35351__;
  assign new_new_n35354__ = ~new_new_n35352__ & ~new_new_n35353__;
  assign new_new_n35355__ = new_new_n35211__ & ~new_new_n35354__;
  assign new_new_n35356__ = ~new_new_n35211__ & new_new_n35354__;
  assign new_new_n35357__ = ~new_new_n35355__ & ~new_new_n35356__;
  assign new_new_n35358__ = new_new_n35210__ & ~new_new_n35357__;
  assign new_new_n35359__ = ~new_new_n35210__ & new_new_n35357__;
  assign new_new_n35360__ = ~new_new_n35358__ & ~new_new_n35359__;
  assign new_new_n35361__ = new_new_n35194__ & new_new_n35360__;
  assign new_new_n35362__ = ~new_new_n35194__ & ~new_new_n35360__;
  assign new_new_n35363__ = ~new_new_n35361__ & ~new_new_n35362__;
  assign new_new_n35364__ = ~new_new_n34955__ & ~new_new_n35096__;
  assign new_new_n35365__ = ~new_new_n35097__ & ~new_new_n35364__;
  assign new_new_n35366__ = ~new_new_n35363__ & new_new_n35365__;
  assign new_new_n35367__ = new_new_n35363__ & ~new_new_n35365__;
  assign new_new_n35368__ = ~new_new_n35366__ & ~new_new_n35367__;
  assign new_new_n35369__ = ~new_new_n34934__ & ~new_new_n34950__;
  assign new_new_n35370__ = new_new_n34934__ & new_new_n34950__;
  assign new_new_n35371__ = ~new_new_n35101__ & ~new_new_n35370__;
  assign new_new_n35372__ = ~new_new_n35369__ & ~new_new_n35371__;
  assign new_new_n35373__ = new_new_n35368__ & ~new_new_n35372__;
  assign new_new_n35374__ = ~new_new_n35368__ & new_new_n35372__;
  assign new_new_n35375__ = ~new_new_n35373__ & ~new_new_n35374__;
  assign new_new_n35376__ = new_new_n8474__ & new_new_n32382__;
  assign new_new_n35377__ = ~new_new_n8479__ & ~new_new_n26667__;
  assign new_new_n35378__ = new_new_n8858__ & new_new_n32729__;
  assign new_new_n35379__ = ~new_new_n35376__ & ~new_new_n35377__;
  assign new_new_n35380__ = ~new_new_n35378__ & new_new_n35379__;
  assign new_new_n35381__ = new_new_n8469__ & new_new_n32758__;
  assign new_new_n35382__ = pi11 & ~new_new_n35381__;
  assign new_new_n35383__ = new_new_n11530__ & new_new_n32758__;
  assign new_new_n35384__ = ~new_new_n35382__ & ~new_new_n35383__;
  assign new_new_n35385__ = new_new_n35380__ & ~new_new_n35384__;
  assign new_new_n35386__ = ~pi11 & ~new_new_n35380__;
  assign new_new_n35387__ = ~new_new_n35385__ & ~new_new_n35386__;
  assign new_new_n35388__ = ~new_new_n35375__ & new_new_n35387__;
  assign new_new_n35389__ = new_new_n35375__ & ~new_new_n35387__;
  assign new_new_n35390__ = ~new_new_n35388__ & ~new_new_n35389__;
  assign new_new_n35391__ = ~new_new_n35175__ & new_new_n35390__;
  assign new_new_n35392__ = new_new_n35175__ & ~new_new_n35390__;
  assign new_new_n35393__ = ~new_new_n35391__ & ~new_new_n35392__;
  assign new_new_n35394__ = ~new_new_n11409__ & new_new_n32740__;
  assign new_new_n35395__ = ~pi08 & new_new_n35394__;
  assign new_new_n35396__ = pi08 & ~new_new_n35394__;
  assign new_new_n35397__ = ~new_new_n35395__ & ~new_new_n35396__;
  assign new_new_n35398__ = new_new_n35393__ & new_new_n35397__;
  assign new_new_n35399__ = ~new_new_n35393__ & ~new_new_n35397__;
  assign new_new_n35400__ = ~new_new_n35398__ & ~new_new_n35399__;
  assign new_new_n35401__ = new_new_n35173__ & new_new_n35400__;
  assign new_new_n35402__ = ~new_new_n35173__ & ~new_new_n35400__;
  assign new_new_n35403__ = ~new_new_n35401__ & ~new_new_n35402__;
  assign new_new_n35404__ = ~new_new_n34719__ & ~new_new_n35146__;
  assign new_new_n35405__ = new_new_n34919__ & ~new_new_n35150__;
  assign new_new_n35406__ = ~new_new_n35404__ & ~new_new_n35405__;
  assign new_new_n35407__ = ~new_new_n34931__ & ~new_new_n35406__;
  assign new_new_n35408__ = ~new_new_n34716__ & ~new_new_n35151__;
  assign new_new_n35409__ = ~new_new_n34711__ & new_new_n35408__;
  assign new_new_n35410__ = ~new_new_n35149__ & ~new_new_n35409__;
  assign new_new_n35411__ = ~new_new_n35407__ & new_new_n35410__;
  assign new_new_n35412__ = ~new_new_n34711__ & ~new_new_n34922__;
  assign new_new_n35413__ = new_new_n35152__ & ~new_new_n35412__;
  assign new_new_n35414__ = new_new_n34700__ & new_new_n35413__;
  assign new_new_n35415__ = new_new_n34923__ & ~new_new_n35152__;
  assign new_new_n35416__ = ~new_new_n34711__ & new_new_n35415__;
  assign new_new_n35417__ = ~new_new_n35414__ & ~new_new_n35416__;
  assign new_new_n35418__ = ~po09 & ~new_new_n35417__;
  assign new_new_n35419__ = new_new_n35411__ & ~new_new_n35418__;
  assign new_new_n35420__ = ~new_new_n35411__ & new_new_n35418__;
  assign new_new_n35421__ = ~new_new_n35419__ & ~new_new_n35420__;
  assign new_new_n35422__ = new_new_n35403__ & ~new_new_n35421__;
  assign new_new_n35423__ = ~new_new_n35403__ & new_new_n35421__;
  assign po11 = new_new_n35422__ | new_new_n35423__;
  assign new_new_n35425__ = new_new_n8470__ & new_new_n33050__;
  assign new_new_n35426__ = new_new_n8858__ & new_new_n32740__;
  assign new_new_n35427__ = new_new_n8474__ & new_new_n32729__;
  assign new_new_n35428__ = ~new_new_n8479__ & new_new_n32382__;
  assign new_new_n35429__ = ~new_new_n35427__ & ~new_new_n35428__;
  assign new_new_n35430__ = ~new_new_n35426__ & new_new_n35429__;
  assign new_new_n35431__ = ~new_new_n35425__ & new_new_n35430__;
  assign new_new_n35432__ = pi11 & ~new_new_n35431__;
  assign new_new_n35433__ = ~pi11 & new_new_n35431__;
  assign new_new_n35434__ = ~new_new_n35432__ & ~new_new_n35433__;
  assign new_new_n35435__ = ~new_new_n35361__ & ~new_new_n35365__;
  assign new_new_n35436__ = ~new_new_n35362__ & ~new_new_n35435__;
  assign new_new_n35437__ = new_new_n6991__ & new_new_n26698__;
  assign new_new_n35438__ = new_new_n6985__ & ~new_new_n26674__;
  assign new_new_n35439__ = ~new_new_n35437__ & ~new_new_n35438__;
  assign new_new_n35440__ = ~new_new_n26667__ & ~new_new_n32340__;
  assign new_new_n35441__ = new_new_n6994__ & new_new_n35440__;
  assign new_new_n35442__ = new_new_n35439__ & ~new_new_n35441__;
  assign new_new_n35443__ = pi14 & ~new_new_n35442__;
  assign new_new_n35444__ = ~pi13 & ~new_new_n32338__;
  assign new_new_n35445__ = pi13 & ~new_new_n32341__;
  assign new_new_n35446__ = new_new_n6994__ & ~new_new_n35444__;
  assign new_new_n35447__ = ~new_new_n35445__ & new_new_n35446__;
  assign new_new_n35448__ = new_new_n26667__ & new_new_n32337__;
  assign new_new_n35449__ = new_new_n6994__ & ~new_new_n35448__;
  assign new_new_n35450__ = ~pi14 & new_new_n35439__;
  assign new_new_n35451__ = ~new_new_n35449__ & new_new_n35450__;
  assign new_new_n35452__ = ~new_new_n35447__ & ~new_new_n35451__;
  assign new_new_n35453__ = ~new_new_n35443__ & new_new_n35452__;
  assign new_new_n35454__ = new_new_n35210__ & ~new_new_n35356__;
  assign new_new_n35455__ = ~new_new_n35355__ & ~new_new_n35454__;
  assign new_new_n35456__ = ~new_new_n35453__ & ~new_new_n35455__;
  assign new_new_n35457__ = new_new_n35453__ & new_new_n35455__;
  assign new_new_n35458__ = ~new_new_n35456__ & ~new_new_n35457__;
  assign new_new_n35459__ = ~new_new_n35346__ & new_new_n35354__;
  assign new_new_n35460__ = ~new_new_n35347__ & ~new_new_n35459__;
  assign new_new_n35461__ = new_new_n6629__ & new_new_n26774__;
  assign new_new_n35462__ = ~new_new_n6625__ & new_new_n26810__;
  assign new_new_n35463__ = new_new_n6633__ & ~new_new_n26729__;
  assign new_new_n35464__ = ~new_new_n6633__ & ~new_new_n30644__;
  assign new_new_n35465__ = new_new_n6631__ & ~new_new_n35463__;
  assign new_new_n35466__ = ~new_new_n35464__ & new_new_n35465__;
  assign new_new_n35467__ = ~new_new_n35462__ & ~new_new_n35466__;
  assign new_new_n35468__ = ~new_new_n35461__ & new_new_n35467__;
  assign new_new_n35469__ = ~pi20 & ~new_new_n35468__;
  assign new_new_n35470__ = new_new_n6625__ & ~new_new_n26774__;
  assign new_new_n35471__ = new_new_n6629__ & ~new_new_n35470__;
  assign new_new_n35472__ = pi20 & ~new_new_n35471__;
  assign new_new_n35473__ = new_new_n35467__ & new_new_n35472__;
  assign new_new_n35474__ = ~new_new_n35469__ & ~new_new_n35473__;
  assign new_new_n35475__ = ~new_new_n35338__ & ~new_new_n35342__;
  assign new_new_n35476__ = ~new_new_n35339__ & ~new_new_n35475__;
  assign new_new_n35477__ = ~new_new_n35474__ & ~new_new_n35476__;
  assign new_new_n35478__ = new_new_n35474__ & new_new_n35476__;
  assign new_new_n35479__ = ~new_new_n35477__ & ~new_new_n35478__;
  assign new_new_n35480__ = ~new_new_n4900__ & ~new_new_n29400__;
  assign new_new_n35481__ = ~new_new_n333__ & ~new_new_n26854__;
  assign new_new_n35482__ = new_new_n873__ & new_new_n26847__;
  assign new_new_n35483__ = ~new_new_n35481__ & ~new_new_n35482__;
  assign new_new_n35484__ = ~new_new_n35480__ & new_new_n35483__;
  assign new_new_n35485__ = pi26 & ~new_new_n35484__;
  assign new_new_n35486__ = new_new_n512__ & ~new_new_n26823__;
  assign new_new_n35487__ = new_new_n801__ & ~new_new_n26823__;
  assign new_new_n35488__ = ~pi26 & ~new_new_n35487__;
  assign new_new_n35489__ = ~new_new_n35486__ & ~new_new_n35488__;
  assign new_new_n35490__ = new_new_n35484__ & ~new_new_n35489__;
  assign new_new_n35491__ = ~new_new_n35485__ & ~new_new_n35490__;
  assign new_new_n35492__ = new_new_n161__ & new_new_n26928__;
  assign new_new_n35493__ = new_new_n765__ & new_new_n26917__;
  assign new_new_n35494__ = ~new_new_n35492__ & ~new_new_n35493__;
  assign new_new_n35495__ = ~pi31 & ~new_new_n35494__;
  assign new_new_n35496__ = new_new_n765__ & new_new_n27462__;
  assign new_new_n35497__ = new_new_n71__ & ~new_new_n26928__;
  assign new_new_n35498__ = pi31 & ~new_new_n35278__;
  assign new_new_n35499__ = ~new_new_n35497__ & new_new_n35498__;
  assign new_new_n35500__ = ~new_new_n35496__ & new_new_n35499__;
  assign new_new_n35501__ = ~new_new_n35495__ & ~new_new_n35500__;
  assign new_new_n35502__ = ~new_new_n35288__ & ~new_new_n35315__;
  assign new_new_n35503__ = ~new_new_n35314__ & ~new_new_n35502__;
  assign new_new_n35504__ = new_new_n35501__ & new_new_n35503__;
  assign new_new_n35505__ = ~new_new_n35501__ & ~new_new_n35503__;
  assign new_new_n35506__ = ~new_new_n35504__ & ~new_new_n35505__;
  assign new_new_n35507__ = new_new_n590__ & ~new_new_n765__;
  assign new_new_n35508__ = ~new_new_n723__ & ~new_new_n990__;
  assign new_new_n35509__ = ~new_new_n189__ & new_new_n35508__;
  assign new_new_n35510__ = new_new_n2166__ & new_new_n3775__;
  assign new_new_n35511__ = ~new_new_n35507__ & new_new_n35510__;
  assign new_new_n35512__ = ~new_new_n115__ & new_new_n35509__;
  assign new_new_n35513__ = new_new_n1710__ & new_new_n2909__;
  assign new_new_n35514__ = new_new_n35512__ & new_new_n35513__;
  assign new_new_n35515__ = new_new_n1149__ & new_new_n35511__;
  assign new_new_n35516__ = new_new_n5412__ & new_new_n35515__;
  assign new_new_n35517__ = new_new_n2926__ & new_new_n35514__;
  assign new_new_n35518__ = new_new_n28573__ & new_new_n35517__;
  assign new_new_n35519__ = new_new_n35516__ & new_new_n35518__;
  assign new_new_n35520__ = ~new_new_n600__ & ~new_new_n843__;
  assign new_new_n35521__ = ~new_new_n346__ & new_new_n35520__;
  assign new_new_n35522__ = ~new_new_n959__ & ~new_new_n961__;
  assign new_new_n35523__ = new_new_n35521__ & new_new_n35522__;
  assign new_new_n35524__ = new_new_n1472__ & new_new_n1637__;
  assign new_new_n35525__ = new_new_n35523__ & new_new_n35524__;
  assign new_new_n35526__ = ~new_new_n249__ & ~new_new_n585__;
  assign new_new_n35527__ = ~new_new_n634__ & ~new_new_n768__;
  assign new_new_n35528__ = ~new_new_n845__ & ~new_new_n947__;
  assign new_new_n35529__ = new_new_n35527__ & new_new_n35528__;
  assign new_new_n35530__ = ~new_new_n143__ & new_new_n35526__;
  assign new_new_n35531__ = ~new_new_n894__ & new_new_n17525__;
  assign new_new_n35532__ = new_new_n35530__ & new_new_n35531__;
  assign new_new_n35533__ = new_new_n16128__ & new_new_n35529__;
  assign new_new_n35534__ = new_new_n35532__ & new_new_n35533__;
  assign new_new_n35535__ = new_new_n3275__ & new_new_n35534__;
  assign new_new_n35536__ = new_new_n4259__ & new_new_n35525__;
  assign new_new_n35537__ = new_new_n35535__ & new_new_n35536__;
  assign new_new_n35538__ = new_new_n4628__ & new_new_n35537__;
  assign new_new_n35539__ = new_new_n35519__ & new_new_n35538__;
  assign new_new_n35540__ = new_new_n16875__ & new_new_n35539__;
  assign new_new_n35541__ = ~new_new_n35282__ & ~new_new_n35540__;
  assign new_new_n35542__ = new_new_n35282__ & new_new_n35540__;
  assign new_new_n35543__ = ~new_new_n35541__ & ~new_new_n35542__;
  assign new_new_n35544__ = ~new_new_n35284__ & ~new_new_n35286__;
  assign new_new_n35545__ = new_new_n35543__ & ~new_new_n35544__;
  assign new_new_n35546__ = ~new_new_n35543__ & new_new_n35544__;
  assign new_new_n35547__ = ~new_new_n35545__ & ~new_new_n35546__;
  assign new_new_n35548__ = new_new_n35506__ & new_new_n35547__;
  assign new_new_n35549__ = ~new_new_n35506__ & ~new_new_n35547__;
  assign new_new_n35550__ = ~new_new_n35548__ & ~new_new_n35549__;
  assign new_new_n35551__ = ~new_new_n35491__ & ~new_new_n35550__;
  assign new_new_n35552__ = new_new_n35491__ & new_new_n35550__;
  assign new_new_n35553__ = ~new_new_n35551__ & ~new_new_n35552__;
  assign new_new_n35554__ = new_new_n4815__ & ~new_new_n26888__;
  assign new_new_n35555__ = new_new_n4212__ & new_new_n26922__;
  assign new_new_n35556__ = ~new_new_n4818__ & ~new_new_n27168__;
  assign new_new_n35557__ = new_new_n4813__ & new_new_n27180__;
  assign new_new_n35558__ = ~new_new_n35555__ & ~new_new_n35556__;
  assign new_new_n35559__ = ~new_new_n35554__ & new_new_n35558__;
  assign new_new_n35560__ = ~new_new_n35557__ & new_new_n35559__;
  assign new_new_n35561__ = pi29 & ~new_new_n35560__;
  assign new_new_n35562__ = ~pi29 & new_new_n35560__;
  assign new_new_n35563__ = ~new_new_n35561__ & ~new_new_n35562__;
  assign new_new_n35564__ = new_new_n35553__ & new_new_n35563__;
  assign new_new_n35565__ = ~new_new_n35553__ & ~new_new_n35563__;
  assign new_new_n35566__ = ~new_new_n35564__ & ~new_new_n35565__;
  assign new_new_n35567__ = new_new_n5191__ & ~new_new_n27221__;
  assign new_new_n35568__ = new_new_n5183__ & ~new_new_n26741__;
  assign new_new_n35569__ = ~new_new_n35567__ & ~new_new_n35568__;
  assign new_new_n35570__ = new_new_n5195__ & ~new_new_n27391__;
  assign new_new_n35571__ = pi23 & ~new_new_n35570__;
  assign new_new_n35572__ = ~pi22 & ~new_new_n30410__;
  assign new_new_n35573__ = pi22 & ~new_new_n30692__;
  assign new_new_n35574__ = new_new_n5195__ & ~new_new_n35572__;
  assign new_new_n35575__ = ~new_new_n35573__ & new_new_n35574__;
  assign new_new_n35576__ = ~new_new_n35571__ & ~new_new_n35575__;
  assign new_new_n35577__ = new_new_n35569__ & ~new_new_n35576__;
  assign new_new_n35578__ = new_new_n5195__ & ~new_new_n26802__;
  assign new_new_n35579__ = new_new_n30411__ & new_new_n35578__;
  assign new_new_n35580__ = new_new_n35569__ & ~new_new_n35579__;
  assign new_new_n35581__ = ~pi23 & ~new_new_n35580__;
  assign new_new_n35582__ = ~new_new_n35577__ & ~new_new_n35581__;
  assign new_new_n35583__ = ~new_new_n35323__ & new_new_n35334__;
  assign new_new_n35584__ = ~new_new_n35322__ & ~new_new_n35583__;
  assign new_new_n35585__ = ~new_new_n35582__ & ~new_new_n35584__;
  assign new_new_n35586__ = new_new_n35582__ & new_new_n35584__;
  assign new_new_n35587__ = ~new_new_n35566__ & ~new_new_n35585__;
  assign new_new_n35588__ = ~new_new_n35586__ & ~new_new_n35587__;
  assign new_new_n35589__ = ~new_new_n35585__ & new_new_n35588__;
  assign new_new_n35590__ = new_new_n35566__ & ~new_new_n35589__;
  assign new_new_n35591__ = ~new_new_n35586__ & new_new_n35587__;
  assign new_new_n35592__ = ~new_new_n35590__ & ~new_new_n35591__;
  assign new_new_n35593__ = ~new_new_n35479__ & new_new_n35592__;
  assign new_new_n35594__ = new_new_n35479__ & ~new_new_n35592__;
  assign new_new_n35595__ = ~new_new_n35593__ & ~new_new_n35594__;
  assign new_new_n35596__ = ~new_new_n35460__ & ~new_new_n35595__;
  assign new_new_n35597__ = new_new_n35460__ & new_new_n35595__;
  assign new_new_n35598__ = ~new_new_n35596__ & ~new_new_n35597__;
  assign new_new_n35599__ = new_new_n6964__ & new_new_n26722__;
  assign new_new_n35600__ = new_new_n6968__ & ~new_new_n27242__;
  assign new_new_n35601__ = new_new_n7935__ & new_new_n27250__;
  assign new_new_n35602__ = ~new_new_n35599__ & ~new_new_n35600__;
  assign new_new_n35603__ = ~new_new_n35601__ & new_new_n35602__;
  assign new_new_n35604__ = new_new_n6958__ & ~new_new_n27271__;
  assign new_new_n35605__ = pi17 & ~new_new_n35604__;
  assign new_new_n35606__ = new_new_n7942__ & ~new_new_n27271__;
  assign new_new_n35607__ = ~new_new_n35605__ & ~new_new_n35606__;
  assign new_new_n35608__ = new_new_n35603__ & ~new_new_n35607__;
  assign new_new_n35609__ = ~pi17 & ~new_new_n35603__;
  assign new_new_n35610__ = ~new_new_n35608__ & ~new_new_n35609__;
  assign new_new_n35611__ = new_new_n35598__ & ~new_new_n35610__;
  assign new_new_n35612__ = ~new_new_n35598__ & new_new_n35610__;
  assign new_new_n35613__ = ~new_new_n35611__ & ~new_new_n35612__;
  assign new_new_n35614__ = new_new_n35458__ & new_new_n35613__;
  assign new_new_n35615__ = ~new_new_n35458__ & ~new_new_n35613__;
  assign new_new_n35616__ = ~new_new_n35614__ & ~new_new_n35615__;
  assign new_new_n35617__ = new_new_n35436__ & new_new_n35616__;
  assign new_new_n35618__ = ~new_new_n35436__ & ~new_new_n35616__;
  assign new_new_n35619__ = ~new_new_n35617__ & ~new_new_n35618__;
  assign new_new_n35620__ = new_new_n35434__ & ~new_new_n35619__;
  assign new_new_n35621__ = ~new_new_n35434__ & new_new_n35619__;
  assign new_new_n35622__ = ~new_new_n35620__ & ~new_new_n35621__;
  assign new_new_n35623__ = pi08 & ~new_new_n35622__;
  assign new_new_n35624__ = ~pi08 & new_new_n35622__;
  assign new_new_n35625__ = ~new_new_n35623__ & ~new_new_n35624__;
  assign new_new_n35626__ = ~new_new_n35374__ & new_new_n35387__;
  assign new_new_n35627__ = ~new_new_n35373__ & ~new_new_n35626__;
  assign new_new_n35628__ = new_new_n35625__ & ~new_new_n35627__;
  assign new_new_n35629__ = ~new_new_n35625__ & new_new_n35627__;
  assign new_new_n35630__ = ~new_new_n35628__ & ~new_new_n35629__;
  assign new_new_n35631__ = pi08 & ~new_new_n35392__;
  assign new_new_n35632__ = new_new_n35630__ & new_new_n35631__;
  assign new_new_n35633__ = ~pi08 & ~new_new_n35391__;
  assign new_new_n35634__ = ~new_new_n35630__ & new_new_n35633__;
  assign new_new_n35635__ = ~new_new_n35632__ & ~new_new_n35634__;
  assign new_new_n35636__ = ~new_new_n35394__ & ~new_new_n35635__;
  assign new_new_n35637__ = ~new_new_n35391__ & ~new_new_n35395__;
  assign new_new_n35638__ = ~new_new_n35392__ & ~new_new_n35637__;
  assign new_new_n35639__ = new_new_n35630__ & new_new_n35638__;
  assign new_new_n35640__ = pi08 & new_new_n35394__;
  assign new_new_n35641__ = ~new_new_n35392__ & ~new_new_n35640__;
  assign new_new_n35642__ = ~new_new_n35391__ & ~new_new_n35641__;
  assign new_new_n35643__ = ~new_new_n35630__ & new_new_n35642__;
  assign new_new_n35644__ = ~new_new_n35639__ & ~new_new_n35643__;
  assign new_new_n35645__ = ~new_new_n35636__ & new_new_n35644__;
  assign new_new_n35646__ = ~new_new_n35402__ & ~new_new_n35411__;
  assign new_new_n35647__ = ~po11 & new_new_n35646__;
  assign new_new_n35648__ = ~new_new_n35402__ & ~new_new_n35418__;
  assign new_new_n35649__ = new_new_n35402__ & new_new_n35420__;
  assign new_new_n35650__ = ~new_new_n35401__ & ~new_new_n35648__;
  assign new_new_n35651__ = ~new_new_n35649__ & new_new_n35650__;
  assign new_new_n35652__ = ~new_new_n35647__ & ~new_new_n35651__;
  assign new_new_n35653__ = new_new_n35645__ & ~new_new_n35652__;
  assign new_new_n35654__ = new_new_n35173__ & new_new_n35411__;
  assign new_new_n35655__ = po11 & new_new_n35654__;
  assign new_new_n35656__ = ~new_new_n35401__ & ~new_new_n35411__;
  assign new_new_n35657__ = ~new_new_n35402__ & ~new_new_n35656__;
  assign new_new_n35658__ = ~new_new_n35418__ & new_new_n35657__;
  assign new_new_n35659__ = ~new_new_n35649__ & ~new_new_n35658__;
  assign new_new_n35660__ = ~new_new_n35655__ & new_new_n35659__;
  assign new_new_n35661__ = ~new_new_n35645__ & ~new_new_n35660__;
  assign po12 = new_new_n35653__ | new_new_n35661__;
  assign new_new_n35663__ = ~new_new_n35173__ & ~new_new_n35411__;
  assign new_new_n35664__ = ~new_new_n35645__ & ~new_new_n35663__;
  assign new_new_n35665__ = new_new_n35418__ & new_new_n35664__;
  assign new_new_n35666__ = new_new_n35402__ & new_new_n35645__;
  assign new_new_n35667__ = ~new_new_n35411__ & new_new_n35666__;
  assign new_new_n35668__ = ~new_new_n35665__ & ~new_new_n35667__;
  assign new_new_n35669__ = ~po11 & ~new_new_n35668__;
  assign new_new_n35670__ = new_new_n6991__ & ~new_new_n26674__;
  assign new_new_n35671__ = new_new_n6985__ & ~new_new_n26667__;
  assign new_new_n35672__ = ~new_new_n35670__ & ~new_new_n35671__;
  assign new_new_n35673__ = new_new_n6994__ & new_new_n32382__;
  assign new_new_n35674__ = ~new_new_n33347__ & new_new_n35673__;
  assign new_new_n35675__ = new_new_n35672__ & ~new_new_n35674__;
  assign new_new_n35676__ = pi14 & ~new_new_n35675__;
  assign new_new_n35677__ = ~pi13 & new_new_n32382__;
  assign new_new_n35678__ = pi13 & ~new_new_n33347__;
  assign new_new_n35679__ = ~new_new_n32382__ & new_new_n33346__;
  assign new_new_n35680__ = new_new_n6994__ & ~new_new_n35679__;
  assign new_new_n35681__ = ~new_new_n35677__ & ~new_new_n35678__;
  assign new_new_n35682__ = new_new_n35680__ & new_new_n35681__;
  assign new_new_n35683__ = ~pi14 & new_new_n35672__;
  assign new_new_n35684__ = ~new_new_n35680__ & new_new_n35683__;
  assign new_new_n35685__ = ~new_new_n35676__ & ~new_new_n35684__;
  assign new_new_n35686__ = ~new_new_n35682__ & new_new_n35685__;
  assign new_new_n35687__ = ~new_new_n35457__ & ~new_new_n35613__;
  assign new_new_n35688__ = ~new_new_n35456__ & ~new_new_n35687__;
  assign new_new_n35689__ = ~new_new_n35686__ & ~new_new_n35688__;
  assign new_new_n35690__ = new_new_n35686__ & new_new_n35688__;
  assign new_new_n35691__ = ~new_new_n35689__ & ~new_new_n35690__;
  assign new_new_n35692__ = new_new_n6968__ & new_new_n27250__;
  assign new_new_n35693__ = new_new_n6964__ & ~new_new_n27242__;
  assign new_new_n35694__ = ~new_new_n35692__ & ~new_new_n35693__;
  assign new_new_n35695__ = new_new_n6958__ & new_new_n26698__;
  assign new_new_n35696__ = new_new_n31511__ & new_new_n35695__;
  assign new_new_n35697__ = new_new_n35694__ & ~new_new_n35696__;
  assign new_new_n35698__ = pi17 & ~new_new_n35697__;
  assign new_new_n35699__ = new_new_n6958__ & ~new_new_n31510__;
  assign new_new_n35700__ = ~pi17 & ~new_new_n35699__;
  assign new_new_n35701__ = ~pi16 & ~new_new_n34204__;
  assign new_new_n35702__ = pi16 & ~new_new_n31509__;
  assign new_new_n35703__ = new_new_n6958__ & ~new_new_n35701__;
  assign new_new_n35704__ = ~new_new_n35702__ & new_new_n35703__;
  assign new_new_n35705__ = ~new_new_n35700__ & ~new_new_n35704__;
  assign new_new_n35706__ = new_new_n35694__ & ~new_new_n35705__;
  assign new_new_n35707__ = ~new_new_n35698__ & ~new_new_n35706__;
  assign new_new_n35708__ = ~new_new_n35597__ & new_new_n35610__;
  assign new_new_n35709__ = ~new_new_n35596__ & ~new_new_n35708__;
  assign new_new_n35710__ = ~new_new_n35478__ & ~new_new_n35592__;
  assign new_new_n35711__ = ~new_new_n35477__ & ~new_new_n35710__;
  assign new_new_n35712__ = new_new_n6629__ & new_new_n26729__;
  assign new_new_n35713__ = ~new_new_n6625__ & new_new_n26774__;
  assign new_new_n35714__ = new_new_n6634__ & new_new_n26722__;
  assign new_new_n35715__ = ~new_new_n35712__ & ~new_new_n35713__;
  assign new_new_n35716__ = ~new_new_n35714__ & new_new_n35715__;
  assign new_new_n35717__ = new_new_n6631__ & ~new_new_n27348__;
  assign new_new_n35718__ = ~pi20 & ~new_new_n35717__;
  assign new_new_n35719__ = new_new_n7015__ & ~new_new_n27348__;
  assign new_new_n35720__ = ~new_new_n35718__ & ~new_new_n35719__;
  assign new_new_n35721__ = new_new_n35716__ & ~new_new_n35720__;
  assign new_new_n35722__ = pi20 & ~new_new_n35716__;
  assign new_new_n35723__ = ~new_new_n35721__ & ~new_new_n35722__;
  assign new_new_n35724__ = ~new_new_n35711__ & new_new_n35723__;
  assign new_new_n35725__ = new_new_n35711__ & ~new_new_n35723__;
  assign new_new_n35726__ = ~new_new_n35724__ & ~new_new_n35725__;
  assign new_new_n35727__ = new_new_n5183__ & ~new_new_n26802__;
  assign new_new_n35728__ = new_new_n5191__ & ~new_new_n26741__;
  assign new_new_n35729__ = new_new_n5213__ & new_new_n26810__;
  assign new_new_n35730__ = ~new_new_n35727__ & ~new_new_n35728__;
  assign new_new_n35731__ = ~new_new_n35729__ & new_new_n35730__;
  assign new_new_n35732__ = new_new_n5195__ & new_new_n27395__;
  assign new_new_n35733__ = new_new_n3311__ & ~new_new_n27221__;
  assign new_new_n35734__ = ~new_new_n333__ & new_new_n26847__;
  assign new_new_n35735__ = new_new_n873__ & ~new_new_n26823__;
  assign new_new_n35736__ = ~new_new_n35734__ & ~new_new_n35735__;
  assign new_new_n35737__ = ~new_new_n35733__ & new_new_n35736__;
  assign new_new_n35738__ = ~pi26 & ~new_new_n35737__;
  assign new_new_n35739__ = new_new_n512__ & new_new_n27411__;
  assign new_new_n35740__ = new_new_n801__ & new_new_n27411__;
  assign new_new_n35741__ = pi26 & ~new_new_n35740__;
  assign new_new_n35742__ = ~new_new_n35739__ & ~new_new_n35741__;
  assign new_new_n35743__ = new_new_n35737__ & ~new_new_n35742__;
  assign new_new_n35744__ = ~new_new_n35738__ & ~new_new_n35743__;
  assign new_new_n35745__ = ~new_new_n35551__ & new_new_n35563__;
  assign new_new_n35746__ = ~new_new_n35552__ & ~new_new_n35745__;
  assign new_new_n35747__ = new_new_n35744__ & new_new_n35746__;
  assign new_new_n35748__ = ~new_new_n35744__ & ~new_new_n35746__;
  assign new_new_n35749__ = ~new_new_n35747__ & ~new_new_n35748__;
  assign new_new_n35750__ = new_new_n4813__ & ~new_new_n27430__;
  assign new_new_n35751__ = ~new_new_n4818__ & new_new_n26922__;
  assign new_new_n35752__ = new_new_n4212__ & ~new_new_n26888__;
  assign new_new_n35753__ = ~new_new_n35751__ & ~new_new_n35752__;
  assign new_new_n35754__ = ~new_new_n35750__ & new_new_n35753__;
  assign new_new_n35755__ = new_new_n4214__ & ~new_new_n26854__;
  assign new_new_n35756__ = pi29 & ~new_new_n35755__;
  assign new_new_n35757__ = new_new_n5732__ & ~new_new_n26854__;
  assign new_new_n35758__ = ~new_new_n35756__ & ~new_new_n35757__;
  assign new_new_n35759__ = new_new_n35754__ & ~new_new_n35758__;
  assign new_new_n35760__ = ~pi29 & ~new_new_n35754__;
  assign new_new_n35761__ = ~new_new_n35759__ & ~new_new_n35760__;
  assign new_new_n35762__ = ~new_new_n35504__ & new_new_n35547__;
  assign new_new_n35763__ = ~new_new_n35505__ & ~new_new_n35762__;
  assign new_new_n35764__ = ~new_new_n35761__ & ~new_new_n35763__;
  assign new_new_n35765__ = new_new_n35761__ & new_new_n35763__;
  assign new_new_n35766__ = ~new_new_n35764__ & ~new_new_n35765__;
  assign new_new_n35767__ = new_new_n161__ & new_new_n26917__;
  assign new_new_n35768__ = new_new_n765__ & ~new_new_n27168__;
  assign new_new_n35769__ = ~new_new_n35767__ & ~new_new_n35768__;
  assign new_new_n35770__ = ~pi31 & ~new_new_n35769__;
  assign new_new_n35771__ = new_new_n71__ & new_new_n26917__;
  assign new_new_n35772__ = new_new_n765__ & ~new_new_n28799__;
  assign new_new_n35773__ = ~new_new_n35492__ & ~new_new_n35771__;
  assign new_new_n35774__ = ~new_new_n35772__ & new_new_n35773__;
  assign new_new_n35775__ = pi31 & ~new_new_n35774__;
  assign new_new_n35776__ = ~new_new_n35770__ & ~new_new_n35775__;
  assign new_new_n35777__ = new_new_n35261__ & ~new_new_n35542__;
  assign new_new_n35778__ = new_new_n35263__ & ~new_new_n35777__;
  assign new_new_n35779__ = ~new_new_n35261__ & ~new_new_n35541__;
  assign new_new_n35780__ = ~new_new_n35778__ & ~new_new_n35779__;
  assign new_new_n35781__ = new_new_n35776__ & ~new_new_n35780__;
  assign new_new_n35782__ = ~new_new_n35776__ & new_new_n35780__;
  assign new_new_n35783__ = ~new_new_n35781__ & ~new_new_n35782__;
  assign new_new_n35784__ = ~new_new_n509__ & ~new_new_n785__;
  assign new_new_n35785__ = new_new_n1154__ & new_new_n35784__;
  assign new_new_n35786__ = new_new_n1156__ & new_new_n2158__;
  assign new_new_n35787__ = new_new_n35785__ & new_new_n35786__;
  assign new_new_n35788__ = new_new_n744__ & new_new_n1223__;
  assign new_new_n35789__ = new_new_n1707__ & new_new_n2992__;
  assign new_new_n35790__ = new_new_n3076__ & new_new_n18162__;
  assign new_new_n35791__ = new_new_n35789__ & new_new_n35790__;
  assign new_new_n35792__ = new_new_n35787__ & new_new_n35788__;
  assign new_new_n35793__ = new_new_n116__ & new_new_n932__;
  assign new_new_n35794__ = new_new_n35792__ & new_new_n35793__;
  assign new_new_n35795__ = new_new_n2091__ & new_new_n35791__;
  assign new_new_n35796__ = new_new_n16296__ & new_new_n35795__;
  assign new_new_n35797__ = new_new_n35794__ & new_new_n35796__;
  assign new_new_n35798__ = new_new_n1030__ & new_new_n2618__;
  assign new_new_n35799__ = new_new_n35797__ & new_new_n35798__;
  assign new_new_n35800__ = new_new_n2987__ & new_new_n35799__;
  assign new_new_n35801__ = ~new_new_n35261__ & ~new_new_n35800__;
  assign new_new_n35802__ = new_new_n35261__ & new_new_n35800__;
  assign new_new_n35803__ = ~pi08 & ~new_new_n35802__;
  assign new_new_n35804__ = ~new_new_n35801__ & ~new_new_n35803__;
  assign new_new_n35805__ = ~new_new_n35801__ & ~new_new_n35804__;
  assign new_new_n35806__ = ~new_new_n35802__ & new_new_n35804__;
  assign new_new_n35807__ = pi08 & ~new_new_n35806__;
  assign new_new_n35808__ = ~new_new_n35805__ & ~new_new_n35807__;
  assign new_new_n35809__ = new_new_n35783__ & ~new_new_n35808__;
  assign new_new_n35810__ = ~new_new_n35783__ & new_new_n35808__;
  assign new_new_n35811__ = ~new_new_n35809__ & ~new_new_n35810__;
  assign new_new_n35812__ = new_new_n35766__ & new_new_n35811__;
  assign new_new_n35813__ = ~new_new_n35766__ & ~new_new_n35811__;
  assign new_new_n35814__ = ~new_new_n35812__ & ~new_new_n35813__;
  assign new_new_n35815__ = new_new_n35749__ & ~new_new_n35814__;
  assign new_new_n35816__ = ~new_new_n35749__ & new_new_n35814__;
  assign new_new_n35817__ = ~new_new_n35815__ & ~new_new_n35816__;
  assign new_new_n35818__ = pi23 & new_new_n35817__;
  assign new_new_n35819__ = ~pi23 & ~new_new_n35817__;
  assign new_new_n35820__ = ~new_new_n35818__ & ~new_new_n35819__;
  assign new_new_n35821__ = ~new_new_n35732__ & ~new_new_n35820__;
  assign new_new_n35822__ = pi22 & new_new_n35817__;
  assign new_new_n35823__ = ~pi22 & ~new_new_n35817__;
  assign new_new_n35824__ = ~new_new_n35822__ & ~new_new_n35823__;
  assign new_new_n35825__ = new_new_n35732__ & ~new_new_n35824__;
  assign new_new_n35826__ = ~new_new_n35821__ & ~new_new_n35825__;
  assign new_new_n35827__ = new_new_n35731__ & ~new_new_n35826__;
  assign new_new_n35828__ = ~new_new_n35731__ & new_new_n35820__;
  assign new_new_n35829__ = ~new_new_n35827__ & ~new_new_n35828__;
  assign new_new_n35830__ = new_new_n35588__ & ~new_new_n35829__;
  assign new_new_n35831__ = ~new_new_n35588__ & new_new_n35829__;
  assign new_new_n35832__ = ~new_new_n35830__ & ~new_new_n35831__;
  assign new_new_n35833__ = new_new_n35726__ & ~new_new_n35832__;
  assign new_new_n35834__ = ~new_new_n35726__ & new_new_n35832__;
  assign new_new_n35835__ = ~new_new_n35833__ & ~new_new_n35834__;
  assign new_new_n35836__ = ~new_new_n35709__ & ~new_new_n35835__;
  assign new_new_n35837__ = new_new_n35709__ & new_new_n35835__;
  assign new_new_n35838__ = ~new_new_n35836__ & ~new_new_n35837__;
  assign new_new_n35839__ = new_new_n35707__ & ~new_new_n35838__;
  assign new_new_n35840__ = ~new_new_n35707__ & new_new_n35838__;
  assign new_new_n35841__ = ~new_new_n35839__ & ~new_new_n35840__;
  assign new_new_n35842__ = new_new_n35691__ & ~new_new_n35841__;
  assign new_new_n35843__ = ~new_new_n35691__ & new_new_n35841__;
  assign new_new_n35844__ = ~new_new_n35842__ & ~new_new_n35843__;
  assign new_new_n35845__ = new_new_n35434__ & ~new_new_n35618__;
  assign new_new_n35846__ = ~new_new_n35617__ & ~new_new_n35845__;
  assign new_new_n35847__ = ~new_new_n35844__ & new_new_n35846__;
  assign new_new_n35848__ = new_new_n35844__ & ~new_new_n35846__;
  assign new_new_n35849__ = ~new_new_n35847__ & ~new_new_n35848__;
  assign new_new_n35850__ = ~new_new_n8479__ & new_new_n32729__;
  assign new_new_n35851__ = new_new_n8474__ & new_new_n32740__;
  assign new_new_n35852__ = ~new_new_n35850__ & ~new_new_n35851__;
  assign new_new_n35853__ = new_new_n8469__ & ~new_new_n34178__;
  assign new_new_n35854__ = pi11 & ~new_new_n35853__;
  assign new_new_n35855__ = new_new_n11530__ & ~new_new_n34178__;
  assign new_new_n35856__ = ~new_new_n35854__ & ~new_new_n35855__;
  assign new_new_n35857__ = new_new_n35852__ & ~new_new_n35856__;
  assign new_new_n35858__ = ~pi11 & ~new_new_n35852__;
  assign new_new_n35859__ = ~new_new_n35857__ & ~new_new_n35858__;
  assign new_new_n35860__ = ~new_new_n35624__ & new_new_n35627__;
  assign new_new_n35861__ = ~new_new_n35623__ & ~new_new_n35860__;
  assign new_new_n35862__ = ~new_new_n35859__ & new_new_n35861__;
  assign new_new_n35863__ = new_new_n35859__ & ~new_new_n35861__;
  assign new_new_n35864__ = ~new_new_n35862__ & ~new_new_n35863__;
  assign new_new_n35865__ = new_new_n35849__ & ~new_new_n35864__;
  assign new_new_n35866__ = ~new_new_n35849__ & new_new_n35864__;
  assign new_new_n35867__ = ~new_new_n35865__ & ~new_new_n35866__;
  assign new_new_n35868__ = new_new_n35630__ & new_new_n35645__;
  assign new_new_n35869__ = ~new_new_n35645__ & new_new_n35657__;
  assign new_new_n35870__ = ~new_new_n35868__ & ~new_new_n35869__;
  assign new_new_n35871__ = new_new_n35867__ & new_new_n35870__;
  assign new_new_n35872__ = ~new_new_n35867__ & ~new_new_n35870__;
  assign new_new_n35873__ = ~new_new_n35871__ & ~new_new_n35872__;
  assign new_new_n35874__ = new_new_n35669__ & ~new_new_n35873__;
  assign new_new_n35875__ = ~new_new_n35669__ & new_new_n35873__;
  assign po13 = new_new_n35874__ | new_new_n35875__;
  assign new_new_n35877__ = new_new_n35846__ & ~new_new_n35870__;
  assign new_new_n35878__ = new_new_n35844__ & ~new_new_n35861__;
  assign new_new_n35879__ = ~new_new_n35844__ & new_new_n35861__;
  assign new_new_n35880__ = ~new_new_n35859__ & ~new_new_n35879__;
  assign new_new_n35881__ = ~new_new_n35878__ & ~new_new_n35880__;
  assign new_new_n35882__ = ~new_new_n35877__ & ~new_new_n35881__;
  assign new_new_n35883__ = ~new_new_n35846__ & new_new_n35870__;
  assign new_new_n35884__ = new_new_n35881__ & ~new_new_n35883__;
  assign new_new_n35885__ = ~new_new_n35882__ & ~new_new_n35884__;
  assign new_new_n35886__ = ~new_new_n8479__ & new_new_n32740__;
  assign new_new_n35887__ = ~pi11 & ~new_new_n35886__;
  assign new_new_n35888__ = pi11 & new_new_n35886__;
  assign new_new_n35889__ = ~new_new_n35887__ & ~new_new_n35888__;
  assign new_new_n35890__ = ~new_new_n35689__ & ~new_new_n35841__;
  assign new_new_n35891__ = ~new_new_n35690__ & ~new_new_n35890__;
  assign new_new_n35892__ = ~new_new_n35707__ & ~new_new_n35837__;
  assign new_new_n35893__ = ~new_new_n35836__ & ~new_new_n35892__;
  assign new_new_n35894__ = new_new_n6991__ & ~new_new_n26667__;
  assign new_new_n35895__ = new_new_n6985__ & new_new_n32382__;
  assign new_new_n35896__ = ~new_new_n35894__ & ~new_new_n35895__;
  assign new_new_n35897__ = new_new_n6994__ & new_new_n32729__;
  assign new_new_n35898__ = new_new_n32758__ & new_new_n35897__;
  assign new_new_n35899__ = new_new_n35896__ & ~new_new_n35898__;
  assign new_new_n35900__ = pi14 & ~new_new_n35899__;
  assign new_new_n35901__ = new_new_n6994__ & ~new_new_n33614__;
  assign new_new_n35902__ = ~pi14 & new_new_n35896__;
  assign new_new_n35903__ = ~new_new_n35901__ & new_new_n35902__;
  assign new_new_n35904__ = ~pi13 & ~new_new_n33617__;
  assign new_new_n35905__ = pi13 & ~new_new_n33619__;
  assign new_new_n35906__ = new_new_n6994__ & ~new_new_n35904__;
  assign new_new_n35907__ = ~new_new_n35905__ & new_new_n35906__;
  assign new_new_n35908__ = ~new_new_n35900__ & ~new_new_n35903__;
  assign new_new_n35909__ = ~new_new_n35907__ & new_new_n35908__;
  assign new_new_n35910__ = new_new_n6968__ & new_new_n26698__;
  assign new_new_n35911__ = new_new_n6964__ & new_new_n27250__;
  assign new_new_n35912__ = new_new_n7935__ & ~new_new_n26674__;
  assign new_new_n35913__ = ~new_new_n35910__ & ~new_new_n35911__;
  assign new_new_n35914__ = ~new_new_n35912__ & new_new_n35913__;
  assign new_new_n35915__ = new_new_n6958__ & new_new_n27284__;
  assign new_new_n35916__ = pi17 & ~new_new_n35915__;
  assign new_new_n35917__ = new_new_n7942__ & new_new_n27284__;
  assign new_new_n35918__ = ~new_new_n35916__ & ~new_new_n35917__;
  assign new_new_n35919__ = new_new_n35914__ & ~new_new_n35918__;
  assign new_new_n35920__ = ~pi17 & ~new_new_n35914__;
  assign new_new_n35921__ = ~new_new_n35919__ & ~new_new_n35920__;
  assign new_new_n35922__ = new_new_n6629__ & new_new_n26722__;
  assign new_new_n35923__ = ~new_new_n6625__ & new_new_n26729__;
  assign new_new_n35924__ = ~new_new_n35922__ & ~new_new_n35923__;
  assign new_new_n35925__ = new_new_n6631__ & ~new_new_n27362__;
  assign new_new_n35926__ = pi20 & ~new_new_n35925__;
  assign new_new_n35927__ = ~pi19 & new_new_n27242__;
  assign new_new_n35928__ = pi19 & ~new_new_n27242__;
  assign new_new_n35929__ = new_new_n6631__ & ~new_new_n35927__;
  assign new_new_n35930__ = ~new_new_n35928__ & new_new_n35929__;
  assign new_new_n35931__ = new_new_n27352__ & new_new_n35930__;
  assign new_new_n35932__ = ~new_new_n35926__ & ~new_new_n35931__;
  assign new_new_n35933__ = new_new_n35924__ & ~new_new_n35932__;
  assign new_new_n35934__ = new_new_n6631__ & new_new_n27353__;
  assign new_new_n35935__ = new_new_n35924__ & ~new_new_n35934__;
  assign new_new_n35936__ = ~pi20 & ~new_new_n35935__;
  assign new_new_n35937__ = ~new_new_n35933__ & ~new_new_n35936__;
  assign new_new_n35938__ = ~new_new_n35588__ & ~new_new_n35817__;
  assign new_new_n35939__ = new_new_n35588__ & new_new_n35817__;
  assign new_new_n35940__ = new_new_n5215__ & new_new_n27395__;
  assign new_new_n35941__ = new_new_n35731__ & ~new_new_n35940__;
  assign new_new_n35942__ = pi23 & ~new_new_n35941__;
  assign new_new_n35943__ = ~pi23 & new_new_n35941__;
  assign new_new_n35944__ = ~new_new_n35942__ & ~new_new_n35943__;
  assign new_new_n35945__ = ~new_new_n35939__ & ~new_new_n35944__;
  assign new_new_n35946__ = ~new_new_n35938__ & ~new_new_n35945__;
  assign new_new_n35947__ = new_new_n35937__ & ~new_new_n35946__;
  assign new_new_n35948__ = ~new_new_n35937__ & new_new_n35946__;
  assign new_new_n35949__ = ~new_new_n35947__ & ~new_new_n35948__;
  assign new_new_n35950__ = new_new_n873__ & ~new_new_n27221__;
  assign new_new_n35951__ = ~new_new_n333__ & ~new_new_n26823__;
  assign new_new_n35952__ = new_new_n3311__ & ~new_new_n26741__;
  assign new_new_n35953__ = ~new_new_n35950__ & ~new_new_n35951__;
  assign new_new_n35954__ = ~new_new_n35952__ & new_new_n35953__;
  assign new_new_n35955__ = ~pi26 & ~new_new_n35954__;
  assign new_new_n35956__ = new_new_n512__ & new_new_n30393__;
  assign new_new_n35957__ = new_new_n801__ & new_new_n30393__;
  assign new_new_n35958__ = pi26 & ~new_new_n35957__;
  assign new_new_n35959__ = ~new_new_n35956__ & ~new_new_n35958__;
  assign new_new_n35960__ = new_new_n35954__ & ~new_new_n35959__;
  assign new_new_n35961__ = ~new_new_n35955__ & ~new_new_n35960__;
  assign new_new_n35962__ = new_new_n4815__ & new_new_n26847__;
  assign new_new_n35963__ = ~new_new_n4818__ & ~new_new_n26888__;
  assign new_new_n35964__ = new_new_n4212__ & ~new_new_n26854__;
  assign new_new_n35965__ = ~new_new_n35963__ & ~new_new_n35964__;
  assign new_new_n35966__ = ~new_new_n35962__ & new_new_n35965__;
  assign new_new_n35967__ = new_new_n4214__ & new_new_n29424__;
  assign new_new_n35968__ = pi29 & ~new_new_n35967__;
  assign new_new_n35969__ = new_new_n4825__ & new_new_n29424__;
  assign new_new_n35970__ = ~new_new_n35968__ & ~new_new_n35969__;
  assign new_new_n35971__ = new_new_n35966__ & ~new_new_n35970__;
  assign new_new_n35972__ = ~pi29 & ~new_new_n35966__;
  assign new_new_n35973__ = ~new_new_n35971__ & ~new_new_n35972__;
  assign new_new_n35974__ = ~new_new_n35782__ & ~new_new_n35808__;
  assign new_new_n35975__ = ~new_new_n35781__ & ~new_new_n35974__;
  assign new_new_n35976__ = ~new_new_n35973__ & new_new_n35975__;
  assign new_new_n35977__ = new_new_n35973__ & ~new_new_n35975__;
  assign new_new_n35978__ = ~new_new_n35976__ & ~new_new_n35977__;
  assign new_new_n35979__ = ~new_new_n351__ & ~new_new_n482__;
  assign new_new_n35980__ = ~new_new_n933__ & ~new_new_n937__;
  assign new_new_n35981__ = ~new_new_n1031__ & new_new_n35980__;
  assign new_new_n35982__ = new_new_n1559__ & new_new_n35979__;
  assign new_new_n35983__ = new_new_n3077__ & new_new_n35982__;
  assign new_new_n35984__ = new_new_n1806__ & new_new_n35981__;
  assign new_new_n35985__ = new_new_n3989__ & new_new_n6322__;
  assign new_new_n35986__ = new_new_n35984__ & new_new_n35985__;
  assign new_new_n35987__ = new_new_n2989__ & new_new_n35983__;
  assign new_new_n35988__ = new_new_n3025__ & new_new_n35987__;
  assign new_new_n35989__ = new_new_n5589__ & new_new_n35986__;
  assign new_new_n35990__ = new_new_n17428__ & new_new_n35989__;
  assign new_new_n35991__ = new_new_n35988__ & new_new_n35990__;
  assign new_new_n35992__ = new_new_n798__ & new_new_n35991__;
  assign new_new_n35993__ = new_new_n2375__ & new_new_n35992__;
  assign new_new_n35994__ = new_new_n71__ & ~new_new_n27168__;
  assign new_new_n35995__ = new_new_n765__ & ~new_new_n29366__;
  assign new_new_n35996__ = ~new_new_n35767__ & ~new_new_n35994__;
  assign new_new_n35997__ = ~new_new_n35995__ & new_new_n35996__;
  assign new_new_n35998__ = pi31 & ~new_new_n35997__;
  assign new_new_n35999__ = new_new_n161__ & new_new_n27168__;
  assign new_new_n36000__ = ~new_new_n161__ & ~new_new_n26922__;
  assign new_new_n36001__ = new_new_n4876__ & ~new_new_n35999__;
  assign new_new_n36002__ = ~new_new_n36000__ & new_new_n36001__;
  assign new_new_n36003__ = ~new_new_n35998__ & ~new_new_n36002__;
  assign new_new_n36004__ = ~new_new_n35993__ & new_new_n36003__;
  assign new_new_n36005__ = new_new_n35993__ & ~new_new_n36003__;
  assign new_new_n36006__ = ~new_new_n36004__ & ~new_new_n36005__;
  assign new_new_n36007__ = ~new_new_n35804__ & ~new_new_n36006__;
  assign new_new_n36008__ = new_new_n35804__ & new_new_n36006__;
  assign new_new_n36009__ = ~new_new_n36007__ & ~new_new_n36008__;
  assign new_new_n36010__ = new_new_n35978__ & new_new_n36009__;
  assign new_new_n36011__ = ~new_new_n35978__ & ~new_new_n36009__;
  assign new_new_n36012__ = ~new_new_n36010__ & ~new_new_n36011__;
  assign new_new_n36013__ = ~new_new_n35961__ & ~new_new_n36012__;
  assign new_new_n36014__ = new_new_n35961__ & new_new_n36012__;
  assign new_new_n36015__ = ~new_new_n36013__ & ~new_new_n36014__;
  assign new_new_n36016__ = ~new_new_n35765__ & ~new_new_n35811__;
  assign new_new_n36017__ = ~new_new_n35764__ & ~new_new_n36016__;
  assign new_new_n36018__ = new_new_n36015__ & ~new_new_n36017__;
  assign new_new_n36019__ = ~new_new_n36015__ & new_new_n36017__;
  assign new_new_n36020__ = ~new_new_n36018__ & ~new_new_n36019__;
  assign new_new_n36021__ = new_new_n5183__ & new_new_n26810__;
  assign new_new_n36022__ = new_new_n5191__ & ~new_new_n26802__;
  assign new_new_n36023__ = ~new_new_n36021__ & ~new_new_n36022__;
  assign new_new_n36024__ = new_new_n5195__ & new_new_n33688__;
  assign new_new_n36025__ = new_new_n36023__ & ~new_new_n36024__;
  assign new_new_n36026__ = ~pi23 & ~new_new_n36025__;
  assign new_new_n36027__ = new_new_n5195__ & ~new_new_n33698__;
  assign new_new_n36028__ = pi23 & ~new_new_n36027__;
  assign new_new_n36029__ = ~pi22 & ~new_new_n33692__;
  assign new_new_n36030__ = pi22 & ~new_new_n33694__;
  assign new_new_n36031__ = new_new_n5195__ & ~new_new_n36029__;
  assign new_new_n36032__ = ~new_new_n36030__ & new_new_n36031__;
  assign new_new_n36033__ = ~new_new_n36028__ & ~new_new_n36032__;
  assign new_new_n36034__ = new_new_n36023__ & ~new_new_n36033__;
  assign new_new_n36035__ = ~new_new_n36026__ & ~new_new_n36034__;
  assign new_new_n36036__ = ~new_new_n35747__ & ~new_new_n35814__;
  assign new_new_n36037__ = ~new_new_n35748__ & ~new_new_n36036__;
  assign new_new_n36038__ = ~new_new_n36035__ & ~new_new_n36037__;
  assign new_new_n36039__ = new_new_n36035__ & new_new_n36037__;
  assign new_new_n36040__ = ~new_new_n36038__ & ~new_new_n36039__;
  assign new_new_n36041__ = ~new_new_n36020__ & new_new_n36040__;
  assign new_new_n36042__ = new_new_n36020__ & ~new_new_n36040__;
  assign new_new_n36043__ = ~new_new_n36041__ & ~new_new_n36042__;
  assign new_new_n36044__ = new_new_n35949__ & ~new_new_n36043__;
  assign new_new_n36045__ = ~new_new_n35949__ & new_new_n36043__;
  assign new_new_n36046__ = ~new_new_n36044__ & ~new_new_n36045__;
  assign new_new_n36047__ = ~new_new_n35921__ & new_new_n36046__;
  assign new_new_n36048__ = new_new_n35921__ & ~new_new_n36046__;
  assign new_new_n36049__ = ~new_new_n36047__ & ~new_new_n36048__;
  assign new_new_n36050__ = ~new_new_n35724__ & new_new_n35832__;
  assign new_new_n36051__ = ~new_new_n35725__ & ~new_new_n36050__;
  assign new_new_n36052__ = new_new_n36049__ & new_new_n36051__;
  assign new_new_n36053__ = ~new_new_n36049__ & ~new_new_n36051__;
  assign new_new_n36054__ = ~new_new_n36052__ & ~new_new_n36053__;
  assign new_new_n36055__ = new_new_n35909__ & new_new_n36054__;
  assign new_new_n36056__ = ~new_new_n35909__ & ~new_new_n36054__;
  assign new_new_n36057__ = ~new_new_n36055__ & ~new_new_n36056__;
  assign new_new_n36058__ = new_new_n35893__ & ~new_new_n36057__;
  assign new_new_n36059__ = ~new_new_n35893__ & new_new_n36057__;
  assign new_new_n36060__ = ~new_new_n36058__ & ~new_new_n36059__;
  assign new_new_n36061__ = ~new_new_n35891__ & ~new_new_n36060__;
  assign new_new_n36062__ = new_new_n35891__ & new_new_n36060__;
  assign new_new_n36063__ = ~new_new_n36061__ & ~new_new_n36062__;
  assign new_new_n36064__ = new_new_n35889__ & new_new_n36063__;
  assign new_new_n36065__ = ~new_new_n35889__ & ~new_new_n36063__;
  assign new_new_n36066__ = ~new_new_n36064__ & ~new_new_n36065__;
  assign new_new_n36067__ = ~new_new_n35878__ & ~new_new_n35879__;
  assign new_new_n36068__ = new_new_n35864__ & ~new_new_n36067__;
  assign new_new_n36069__ = ~new_new_n35877__ & ~new_new_n36068__;
  assign new_new_n36070__ = ~new_new_n35883__ & new_new_n36069__;
  assign new_new_n36071__ = ~new_new_n35885__ & ~new_new_n36066__;
  assign new_new_n36072__ = ~new_new_n36070__ & new_new_n36071__;
  assign new_new_n36073__ = new_new_n35878__ & new_new_n35883__;
  assign new_new_n36074__ = ~new_new_n35844__ & ~new_new_n35883__;
  assign new_new_n36075__ = ~new_new_n35877__ & ~new_new_n36074__;
  assign new_new_n36076__ = ~new_new_n35861__ & new_new_n36075__;
  assign new_new_n36077__ = new_new_n35848__ & new_new_n35870__;
  assign new_new_n36078__ = ~new_new_n36076__ & ~new_new_n36077__;
  assign new_new_n36079__ = ~new_new_n35859__ & ~new_new_n36078__;
  assign new_new_n36080__ = new_new_n35861__ & ~new_new_n36075__;
  assign new_new_n36081__ = new_new_n35847__ & ~new_new_n35870__;
  assign new_new_n36082__ = ~new_new_n36080__ & ~new_new_n36081__;
  assign new_new_n36083__ = new_new_n35859__ & ~new_new_n36082__;
  assign new_new_n36084__ = new_new_n35877__ & new_new_n35879__;
  assign new_new_n36085__ = new_new_n36066__ & ~new_new_n36073__;
  assign new_new_n36086__ = ~new_new_n36084__ & new_new_n36085__;
  assign new_new_n36087__ = ~new_new_n36079__ & new_new_n36086__;
  assign new_new_n36088__ = ~new_new_n36083__ & new_new_n36087__;
  assign new_new_n36089__ = ~new_new_n36072__ & ~new_new_n36088__;
  assign new_new_n36090__ = new_new_n35669__ & new_new_n35873__;
  assign new_new_n36091__ = new_new_n36089__ & new_new_n36090__;
  assign new_new_n36092__ = ~new_new_n36089__ & ~new_new_n36090__;
  assign po14 = ~new_new_n36091__ & ~new_new_n36092__;
  assign new_new_n36094__ = ~new_new_n35893__ & ~new_new_n36055__;
  assign new_new_n36095__ = ~new_new_n36056__ & ~new_new_n36094__;
  assign new_new_n36096__ = pi14 & new_new_n32740__;
  assign new_new_n36097__ = ~pi13 & ~new_new_n32740__;
  assign new_new_n36098__ = new_new_n33050__ & new_new_n36097__;
  assign new_new_n36099__ = ~new_new_n36096__ & ~new_new_n36098__;
  assign new_new_n36100__ = new_new_n6994__ & ~new_new_n36099__;
  assign new_new_n36101__ = new_new_n18717__ & new_new_n33050__;
  assign new_new_n36102__ = new_new_n6991__ & new_new_n32382__;
  assign new_new_n36103__ = new_new_n6985__ & new_new_n32729__;
  assign new_new_n36104__ = ~new_new_n36102__ & ~new_new_n36103__;
  assign new_new_n36105__ = ~pi14 & ~new_new_n36104__;
  assign new_new_n36106__ = pi14 & new_new_n36104__;
  assign new_new_n36107__ = ~new_new_n36105__ & ~new_new_n36106__;
  assign new_new_n36108__ = ~new_new_n36101__ & new_new_n36107__;
  assign new_new_n36109__ = ~new_new_n36100__ & ~new_new_n36108__;
  assign new_new_n36110__ = ~new_new_n36047__ & ~new_new_n36051__;
  assign new_new_n36111__ = ~new_new_n36048__ & ~new_new_n36110__;
  assign new_new_n36112__ = ~new_new_n36109__ & ~new_new_n36111__;
  assign new_new_n36113__ = new_new_n36109__ & new_new_n36111__;
  assign new_new_n36114__ = ~new_new_n36112__ & ~new_new_n36113__;
  assign new_new_n36115__ = ~new_new_n36020__ & ~new_new_n36038__;
  assign new_new_n36116__ = ~new_new_n36039__ & ~new_new_n36115__;
  assign new_new_n36117__ = new_new_n5213__ & new_new_n26729__;
  assign new_new_n36118__ = new_new_n5191__ & new_new_n26810__;
  assign new_new_n36119__ = new_new_n5183__ & new_new_n26774__;
  assign new_new_n36120__ = ~new_new_n36117__ & ~new_new_n36118__;
  assign new_new_n36121__ = ~new_new_n36119__ & new_new_n36120__;
  assign new_new_n36122__ = new_new_n5195__ & new_new_n30644__;
  assign new_new_n36123__ = pi23 & ~new_new_n36122__;
  assign new_new_n36124__ = new_new_n7878__ & new_new_n30644__;
  assign new_new_n36125__ = ~new_new_n36123__ & ~new_new_n36124__;
  assign new_new_n36126__ = new_new_n36121__ & ~new_new_n36125__;
  assign new_new_n36127__ = ~pi23 & ~new_new_n36121__;
  assign new_new_n36128__ = ~new_new_n36126__ & ~new_new_n36127__;
  assign new_new_n36129__ = ~new_new_n36014__ & ~new_new_n36017__;
  assign new_new_n36130__ = ~new_new_n36013__ & ~new_new_n36129__;
  assign new_new_n36131__ = ~new_new_n36128__ & ~new_new_n36130__;
  assign new_new_n36132__ = new_new_n36128__ & new_new_n36130__;
  assign new_new_n36133__ = ~new_new_n36131__ & ~new_new_n36132__;
  assign new_new_n36134__ = ~new_new_n333__ & ~new_new_n27221__;
  assign new_new_n36135__ = new_new_n873__ & ~new_new_n26741__;
  assign new_new_n36136__ = ~new_new_n36134__ & ~new_new_n36135__;
  assign new_new_n36137__ = ~new_new_n110__ & ~new_new_n26802__;
  assign new_new_n36138__ = new_new_n30411__ & new_new_n36137__;
  assign new_new_n36139__ = new_new_n36136__ & ~new_new_n36138__;
  assign new_new_n36140__ = ~pi26 & ~new_new_n36139__;
  assign new_new_n36141__ = new_new_n801__ & ~new_new_n27391__;
  assign new_new_n36142__ = pi26 & ~new_new_n36141__;
  assign new_new_n36143__ = ~pi25 & ~new_new_n30410__;
  assign new_new_n36144__ = pi25 & ~new_new_n30692__;
  assign new_new_n36145__ = ~new_new_n110__ & ~new_new_n36143__;
  assign new_new_n36146__ = ~new_new_n36144__ & new_new_n36145__;
  assign new_new_n36147__ = ~new_new_n36142__ & ~new_new_n36146__;
  assign new_new_n36148__ = new_new_n36136__ & ~new_new_n36147__;
  assign new_new_n36149__ = ~new_new_n36140__ & ~new_new_n36148__;
  assign new_new_n36150__ = new_new_n4813__ & ~new_new_n29400__;
  assign new_new_n36151__ = ~new_new_n4818__ & ~new_new_n26854__;
  assign new_new_n36152__ = new_new_n4212__ & new_new_n26847__;
  assign new_new_n36153__ = new_new_n4815__ & ~new_new_n26823__;
  assign new_new_n36154__ = ~new_new_n36151__ & ~new_new_n36152__;
  assign new_new_n36155__ = ~new_new_n36153__ & new_new_n36154__;
  assign new_new_n36156__ = ~new_new_n36150__ & new_new_n36155__;
  assign new_new_n36157__ = new_new_n765__ & ~new_new_n27180__;
  assign new_new_n36158__ = ~new_new_n35999__ & ~new_new_n36157__;
  assign new_new_n36159__ = pi31 & ~new_new_n36158__;
  assign new_new_n36160__ = new_new_n161__ & new_new_n26922__;
  assign new_new_n36161__ = ~new_new_n71__ & new_new_n36160__;
  assign new_new_n36162__ = new_new_n71__ & ~new_new_n26922__;
  assign new_new_n36163__ = pi31 & ~new_new_n36162__;
  assign new_new_n36164__ = ~new_new_n15853__ & ~new_new_n26888__;
  assign new_new_n36165__ = ~new_new_n36161__ & ~new_new_n36163__;
  assign new_new_n36166__ = ~new_new_n36164__ & new_new_n36165__;
  assign new_new_n36167__ = ~new_new_n36159__ & ~new_new_n36166__;
  assign new_new_n36168__ = ~new_new_n232__ & ~new_new_n238__;
  assign new_new_n36169__ = ~new_new_n488__ & ~new_new_n588__;
  assign new_new_n36170__ = ~new_new_n919__ & new_new_n1106__;
  assign new_new_n36171__ = new_new_n1424__ & new_new_n1711__;
  assign new_new_n36172__ = new_new_n1859__ & new_new_n2383__;
  assign new_new_n36173__ = new_new_n36171__ & new_new_n36172__;
  assign new_new_n36174__ = new_new_n36169__ & new_new_n36170__;
  assign new_new_n36175__ = ~new_new_n254__ & new_new_n36168__;
  assign new_new_n36176__ = ~new_new_n630__ & new_new_n1145__;
  assign new_new_n36177__ = new_new_n1599__ & new_new_n2549__;
  assign new_new_n36178__ = new_new_n36176__ & new_new_n36177__;
  assign new_new_n36179__ = new_new_n36174__ & new_new_n36175__;
  assign new_new_n36180__ = new_new_n709__ & new_new_n36173__;
  assign new_new_n36181__ = new_new_n2641__ & new_new_n36180__;
  assign new_new_n36182__ = new_new_n36178__ & new_new_n36179__;
  assign new_new_n36183__ = new_new_n36181__ & new_new_n36182__;
  assign new_new_n36184__ = new_new_n16789__ & new_new_n18522__;
  assign new_new_n36185__ = new_new_n36183__ & new_new_n36184__;
  assign new_new_n36186__ = new_new_n6181__ & new_new_n36185__;
  assign new_new_n36187__ = new_new_n35243__ & new_new_n36186__;
  assign new_new_n36188__ = ~new_new_n35993__ & ~new_new_n36187__;
  assign new_new_n36189__ = new_new_n35993__ & new_new_n36187__;
  assign new_new_n36190__ = ~new_new_n36188__ & ~new_new_n36189__;
  assign new_new_n36191__ = ~new_new_n35804__ & ~new_new_n36004__;
  assign new_new_n36192__ = ~new_new_n36005__ & ~new_new_n36191__;
  assign new_new_n36193__ = ~new_new_n36190__ & new_new_n36192__;
  assign new_new_n36194__ = new_new_n36190__ & ~new_new_n36192__;
  assign new_new_n36195__ = ~new_new_n36193__ & ~new_new_n36194__;
  assign new_new_n36196__ = ~new_new_n36167__ & new_new_n36195__;
  assign new_new_n36197__ = new_new_n36167__ & ~new_new_n36195__;
  assign new_new_n36198__ = ~new_new_n36196__ & ~new_new_n36197__;
  assign new_new_n36199__ = pi29 & ~new_new_n36198__;
  assign new_new_n36200__ = ~pi29 & new_new_n36198__;
  assign new_new_n36201__ = ~new_new_n36199__ & ~new_new_n36200__;
  assign new_new_n36202__ = new_new_n36156__ & new_new_n36201__;
  assign new_new_n36203__ = ~new_new_n36156__ & ~new_new_n36201__;
  assign new_new_n36204__ = ~new_new_n36202__ & ~new_new_n36203__;
  assign new_new_n36205__ = ~new_new_n36149__ & new_new_n36204__;
  assign new_new_n36206__ = new_new_n36149__ & ~new_new_n36204__;
  assign new_new_n36207__ = ~new_new_n36205__ & ~new_new_n36206__;
  assign new_new_n36208__ = ~new_new_n35976__ & new_new_n36009__;
  assign new_new_n36209__ = ~new_new_n35977__ & ~new_new_n36208__;
  assign new_new_n36210__ = new_new_n36207__ & new_new_n36209__;
  assign new_new_n36211__ = ~new_new_n36207__ & ~new_new_n36209__;
  assign new_new_n36212__ = ~new_new_n36210__ & ~new_new_n36211__;
  assign new_new_n36213__ = new_new_n36133__ & ~new_new_n36212__;
  assign new_new_n36214__ = ~new_new_n36133__ & new_new_n36212__;
  assign new_new_n36215__ = ~new_new_n36213__ & ~new_new_n36214__;
  assign new_new_n36216__ = ~new_new_n36116__ & new_new_n36215__;
  assign new_new_n36217__ = new_new_n36116__ & ~new_new_n36215__;
  assign new_new_n36218__ = ~new_new_n36216__ & ~new_new_n36217__;
  assign new_new_n36219__ = new_new_n6634__ & new_new_n27250__;
  assign new_new_n36220__ = ~new_new_n6625__ & new_new_n26722__;
  assign new_new_n36221__ = new_new_n6629__ & ~new_new_n27242__;
  assign new_new_n36222__ = new_new_n6936__ & ~new_new_n27271__;
  assign new_new_n36223__ = ~new_new_n36220__ & ~new_new_n36221__;
  assign new_new_n36224__ = ~new_new_n36219__ & new_new_n36223__;
  assign new_new_n36225__ = ~new_new_n36222__ & new_new_n36224__;
  assign new_new_n36226__ = ~pi20 & ~new_new_n36225__;
  assign new_new_n36227__ = pi20 & new_new_n36225__;
  assign new_new_n36228__ = ~new_new_n36226__ & ~new_new_n36227__;
  assign new_new_n36229__ = new_new_n36218__ & new_new_n36228__;
  assign new_new_n36230__ = ~new_new_n36218__ & ~new_new_n36228__;
  assign new_new_n36231__ = ~new_new_n36229__ & ~new_new_n36230__;
  assign new_new_n36232__ = new_new_n6959__ & ~new_new_n32340__;
  assign new_new_n36233__ = new_new_n6964__ & new_new_n26698__;
  assign new_new_n36234__ = new_new_n6968__ & ~new_new_n26674__;
  assign new_new_n36235__ = ~new_new_n36233__ & ~new_new_n36234__;
  assign new_new_n36236__ = ~new_new_n36232__ & new_new_n36235__;
  assign new_new_n36237__ = new_new_n6958__ & ~new_new_n26667__;
  assign new_new_n36238__ = pi17 & ~new_new_n36237__;
  assign new_new_n36239__ = new_new_n8160__ & ~new_new_n26667__;
  assign new_new_n36240__ = ~new_new_n36238__ & ~new_new_n36239__;
  assign new_new_n36241__ = new_new_n36236__ & ~new_new_n36240__;
  assign new_new_n36242__ = ~pi17 & ~new_new_n36236__;
  assign new_new_n36243__ = ~new_new_n36241__ & ~new_new_n36242__;
  assign new_new_n36244__ = ~new_new_n35948__ & new_new_n36043__;
  assign new_new_n36245__ = ~new_new_n35947__ & ~new_new_n36244__;
  assign new_new_n36246__ = ~new_new_n36243__ & new_new_n36245__;
  assign new_new_n36247__ = new_new_n36243__ & ~new_new_n36245__;
  assign new_new_n36248__ = ~new_new_n36231__ & ~new_new_n36247__;
  assign new_new_n36249__ = ~new_new_n36246__ & new_new_n36248__;
  assign new_new_n36250__ = ~new_new_n36231__ & ~new_new_n36249__;
  assign new_new_n36251__ = ~new_new_n36246__ & ~new_new_n36248__;
  assign new_new_n36252__ = ~new_new_n36247__ & new_new_n36251__;
  assign new_new_n36253__ = ~new_new_n36250__ & ~new_new_n36252__;
  assign new_new_n36254__ = new_new_n36114__ & ~new_new_n36253__;
  assign new_new_n36255__ = ~new_new_n36114__ & new_new_n36253__;
  assign new_new_n36256__ = ~new_new_n36254__ & ~new_new_n36255__;
  assign new_new_n36257__ = ~new_new_n36095__ & ~new_new_n36256__;
  assign new_new_n36258__ = new_new_n36095__ & new_new_n36256__;
  assign new_new_n36259__ = ~new_new_n36257__ & ~new_new_n36258__;
  assign new_new_n36260__ = new_new_n35889__ & ~new_new_n36062__;
  assign new_new_n36261__ = ~new_new_n36061__ & ~new_new_n36260__;
  assign new_new_n36262__ = new_new_n35877__ & new_new_n35881__;
  assign new_new_n36263__ = ~new_new_n35882__ & ~new_new_n36066__;
  assign new_new_n36264__ = ~new_new_n35859__ & new_new_n35878__;
  assign new_new_n36265__ = ~new_new_n36066__ & ~new_new_n36264__;
  assign new_new_n36266__ = new_new_n35859__ & new_new_n35879__;
  assign new_new_n36267__ = ~new_new_n36265__ & ~new_new_n36266__;
  assign new_new_n36268__ = ~new_new_n35883__ & ~new_new_n36267__;
  assign new_new_n36269__ = ~new_new_n36262__ & ~new_new_n36268__;
  assign new_new_n36270__ = ~new_new_n36263__ & new_new_n36269__;
  assign new_new_n36271__ = ~new_new_n36261__ & new_new_n36270__;
  assign new_new_n36272__ = ~pi11 & new_new_n36271__;
  assign new_new_n36273__ = new_new_n36261__ & ~new_new_n36270__;
  assign new_new_n36274__ = ~new_new_n36271__ & ~new_new_n36273__;
  assign new_new_n36275__ = pi11 & ~new_new_n36274__;
  assign new_new_n36276__ = ~pi11 & new_new_n36274__;
  assign new_new_n36277__ = ~new_new_n36275__ & ~new_new_n36276__;
  assign new_new_n36278__ = new_new_n36091__ & new_new_n36277__;
  assign new_new_n36279__ = ~new_new_n36091__ & ~new_new_n36277__;
  assign new_new_n36280__ = ~new_new_n36278__ & ~new_new_n36279__;
  assign new_new_n36281__ = ~new_new_n36272__ & ~new_new_n36280__;
  assign new_new_n36282__ = new_new_n36259__ & new_new_n36281__;
  assign new_new_n36283__ = ~new_new_n36259__ & ~new_new_n36281__;
  assign po15 = ~new_new_n36282__ & ~new_new_n36283__;
  assign new_new_n36285__ = ~new_new_n36256__ & new_new_n36261__;
  assign new_new_n36286__ = ~new_new_n36095__ & ~new_new_n36270__;
  assign new_new_n36287__ = new_new_n36285__ & new_new_n36286__;
  assign new_new_n36288__ = ~new_new_n36113__ & new_new_n36253__;
  assign new_new_n36289__ = ~new_new_n36112__ & ~new_new_n36288__;
  assign new_new_n36290__ = ~new_new_n6989__ & ~new_new_n34178__;
  assign new_new_n36291__ = pi14 & ~new_new_n36290__;
  assign new_new_n36292__ = ~pi14 & ~new_new_n6984__;
  assign new_new_n36293__ = ~new_new_n23485__ & new_new_n36292__;
  assign new_new_n36294__ = ~new_new_n34178__ & new_new_n36293__;
  assign new_new_n36295__ = ~new_new_n36291__ & ~new_new_n36294__;
  assign new_new_n36296__ = ~new_new_n32729__ & ~new_new_n36295__;
  assign new_new_n36297__ = ~pi14 & ~new_new_n34177__;
  assign new_new_n36298__ = ~pi13 & ~new_new_n34178__;
  assign new_new_n36299__ = ~new_new_n6981__ & ~new_new_n36297__;
  assign new_new_n36300__ = ~new_new_n36298__ & new_new_n36299__;
  assign new_new_n36301__ = ~new_new_n6984__ & ~new_new_n6988__;
  assign new_new_n36302__ = new_new_n32729__ & new_new_n36301__;
  assign new_new_n36303__ = ~new_new_n36300__ & ~new_new_n36302__;
  assign new_new_n36304__ = ~new_new_n36296__ & new_new_n36303__;
  assign new_new_n36305__ = new_new_n6959__ & ~new_new_n33347__;
  assign new_new_n36306__ = new_new_n6964__ & ~new_new_n26674__;
  assign new_new_n36307__ = new_new_n6968__ & ~new_new_n26667__;
  assign new_new_n36308__ = new_new_n7935__ & new_new_n32382__;
  assign new_new_n36309__ = ~new_new_n36306__ & ~new_new_n36307__;
  assign new_new_n36310__ = ~new_new_n36308__ & new_new_n36309__;
  assign new_new_n36311__ = ~new_new_n36305__ & new_new_n36310__;
  assign new_new_n36312__ = ~pi17 & ~new_new_n36311__;
  assign new_new_n36313__ = pi17 & new_new_n36311__;
  assign new_new_n36314__ = ~new_new_n36312__ & ~new_new_n36313__;
  assign new_new_n36315__ = new_new_n6634__ & new_new_n26698__;
  assign new_new_n36316__ = new_new_n6629__ & new_new_n27250__;
  assign new_new_n36317__ = ~new_new_n6625__ & ~new_new_n27242__;
  assign new_new_n36318__ = new_new_n6936__ & new_new_n31511__;
  assign new_new_n36319__ = ~new_new_n36316__ & ~new_new_n36317__;
  assign new_new_n36320__ = ~new_new_n36315__ & new_new_n36319__;
  assign new_new_n36321__ = ~new_new_n36318__ & new_new_n36320__;
  assign new_new_n36322__ = pi20 & ~new_new_n36321__;
  assign new_new_n36323__ = ~pi20 & new_new_n36321__;
  assign new_new_n36324__ = ~new_new_n36322__ & ~new_new_n36323__;
  assign new_new_n36325__ = ~new_new_n36216__ & ~new_new_n36228__;
  assign new_new_n36326__ = ~new_new_n36217__ & ~new_new_n36325__;
  assign new_new_n36327__ = ~new_new_n36324__ & new_new_n36326__;
  assign new_new_n36328__ = new_new_n36324__ & ~new_new_n36326__;
  assign new_new_n36329__ = ~new_new_n36327__ & ~new_new_n36328__;
  assign new_new_n36330__ = ~new_new_n36205__ & ~new_new_n36209__;
  assign new_new_n36331__ = ~new_new_n36206__ & ~new_new_n36330__;
  assign new_new_n36332__ = new_new_n4815__ & ~new_new_n27221__;
  assign new_new_n36333__ = new_new_n4212__ & ~new_new_n26823__;
  assign new_new_n36334__ = ~new_new_n4818__ & new_new_n26847__;
  assign new_new_n36335__ = new_new_n4813__ & new_new_n27411__;
  assign new_new_n36336__ = ~new_new_n36333__ & ~new_new_n36334__;
  assign new_new_n36337__ = ~new_new_n36332__ & new_new_n36336__;
  assign new_new_n36338__ = ~new_new_n36335__ & new_new_n36337__;
  assign new_new_n36339__ = pi29 & ~new_new_n36338__;
  assign new_new_n36340__ = ~pi29 & new_new_n36338__;
  assign new_new_n36341__ = ~new_new_n36339__ & ~new_new_n36340__;
  assign new_new_n36342__ = new_new_n35804__ & new_new_n36187__;
  assign new_new_n36343__ = new_new_n36003__ & new_new_n36342__;
  assign new_new_n36344__ = new_new_n35993__ & ~new_new_n36343__;
  assign new_new_n36345__ = ~new_new_n35804__ & ~new_new_n36187__;
  assign new_new_n36346__ = ~new_new_n36003__ & new_new_n36345__;
  assign new_new_n36347__ = ~new_new_n35993__ & ~new_new_n36346__;
  assign new_new_n36348__ = ~new_new_n36344__ & ~new_new_n36347__;
  assign new_new_n36349__ = new_new_n161__ & ~new_new_n26888__;
  assign new_new_n36350__ = new_new_n765__ & ~new_new_n26854__;
  assign new_new_n36351__ = ~new_new_n36349__ & ~new_new_n36350__;
  assign new_new_n36352__ = ~pi31 & ~new_new_n36351__;
  assign new_new_n36353__ = new_new_n71__ & ~new_new_n26888__;
  assign new_new_n36354__ = new_new_n765__ & ~new_new_n27430__;
  assign new_new_n36355__ = ~new_new_n36160__ & ~new_new_n36353__;
  assign new_new_n36356__ = ~new_new_n36354__ & new_new_n36355__;
  assign new_new_n36357__ = pi31 & ~new_new_n36356__;
  assign new_new_n36358__ = ~new_new_n36352__ & ~new_new_n36357__;
  assign new_new_n36359__ = ~new_new_n235__ & ~new_new_n302__;
  assign new_new_n36360__ = ~new_new_n511__ & ~new_new_n634__;
  assign new_new_n36361__ = ~new_new_n1031__ & new_new_n36360__;
  assign new_new_n36362__ = ~new_new_n143__ & new_new_n36359__;
  assign new_new_n36363__ = ~new_new_n277__ & ~new_new_n300__;
  assign new_new_n36364__ = new_new_n3010__ & new_new_n36363__;
  assign new_new_n36365__ = new_new_n36361__ & new_new_n36362__;
  assign new_new_n36366__ = new_new_n589__ & new_new_n989__;
  assign new_new_n36367__ = new_new_n1153__ & new_new_n1523__;
  assign new_new_n36368__ = new_new_n6122__ & new_new_n36367__;
  assign new_new_n36369__ = new_new_n36365__ & new_new_n36366__;
  assign new_new_n36370__ = new_new_n36364__ & new_new_n36369__;
  assign new_new_n36371__ = new_new_n2871__ & new_new_n36368__;
  assign new_new_n36372__ = new_new_n6105__ & new_new_n36371__;
  assign new_new_n36373__ = new_new_n2047__ & new_new_n36370__;
  assign new_new_n36374__ = new_new_n36372__ & new_new_n36373__;
  assign new_new_n36375__ = new_new_n1128__ & new_new_n36374__;
  assign new_new_n36376__ = new_new_n2115__ & new_new_n36375__;
  assign new_new_n36377__ = ~pi11 & ~new_new_n36376__;
  assign new_new_n36378__ = pi11 & new_new_n36376__;
  assign new_new_n36379__ = ~new_new_n36377__ & ~new_new_n36378__;
  assign new_new_n36380__ = new_new_n36358__ & ~new_new_n36379__;
  assign new_new_n36381__ = ~new_new_n36358__ & new_new_n36379__;
  assign new_new_n36382__ = ~new_new_n36380__ & ~new_new_n36381__;
  assign new_new_n36383__ = new_new_n36348__ & new_new_n36382__;
  assign new_new_n36384__ = ~new_new_n36348__ & ~new_new_n36382__;
  assign new_new_n36385__ = ~new_new_n36383__ & ~new_new_n36384__;
  assign new_new_n36386__ = ~new_new_n36197__ & new_new_n36204__;
  assign new_new_n36387__ = ~new_new_n36196__ & ~new_new_n36386__;
  assign new_new_n36388__ = ~new_new_n36385__ & new_new_n36387__;
  assign new_new_n36389__ = new_new_n36385__ & ~new_new_n36387__;
  assign new_new_n36390__ = ~new_new_n36388__ & ~new_new_n36389__;
  assign new_new_n36391__ = new_new_n36341__ & ~new_new_n36390__;
  assign new_new_n36392__ = ~new_new_n36341__ & new_new_n36390__;
  assign new_new_n36393__ = ~new_new_n36391__ & ~new_new_n36392__;
  assign new_new_n36394__ = ~new_new_n36331__ & new_new_n36393__;
  assign new_new_n36395__ = new_new_n36331__ & ~new_new_n36393__;
  assign new_new_n36396__ = ~new_new_n36394__ & ~new_new_n36395__;
  assign new_new_n36397__ = new_new_n3311__ & new_new_n26810__;
  assign new_new_n36398__ = new_new_n873__ & ~new_new_n26802__;
  assign new_new_n36399__ = ~new_new_n4900__ & new_new_n27395__;
  assign new_new_n36400__ = ~new_new_n36397__ & ~new_new_n36398__;
  assign new_new_n36401__ = ~new_new_n36399__ & new_new_n36400__;
  assign new_new_n36402__ = new_new_n303__ & ~new_new_n26741__;
  assign new_new_n36403__ = pi26 & ~new_new_n36402__;
  assign new_new_n36404__ = new_new_n145__ & ~new_new_n26741__;
  assign new_new_n36405__ = ~pi26 & ~new_new_n36404__;
  assign new_new_n36406__ = pi23 & ~new_new_n36405__;
  assign new_new_n36407__ = ~new_new_n36403__ & ~new_new_n36406__;
  assign new_new_n36408__ = new_new_n36401__ & ~new_new_n36407__;
  assign new_new_n36409__ = ~pi26 & ~new_new_n36401__;
  assign new_new_n36410__ = ~new_new_n36408__ & ~new_new_n36409__;
  assign new_new_n36411__ = new_new_n36396__ & ~new_new_n36410__;
  assign new_new_n36412__ = ~new_new_n36396__ & new_new_n36410__;
  assign new_new_n36413__ = ~new_new_n36411__ & ~new_new_n36412__;
  assign new_new_n36414__ = new_new_n5213__ & new_new_n26722__;
  assign new_new_n36415__ = new_new_n5191__ & new_new_n26774__;
  assign new_new_n36416__ = new_new_n5183__ & new_new_n26729__;
  assign new_new_n36417__ = ~new_new_n36415__ & ~new_new_n36416__;
  assign new_new_n36418__ = ~new_new_n36414__ & new_new_n36417__;
  assign new_new_n36419__ = new_new_n5195__ & ~new_new_n27348__;
  assign new_new_n36420__ = ~pi23 & ~new_new_n36419__;
  assign new_new_n36421__ = new_new_n5974__ & ~new_new_n27348__;
  assign new_new_n36422__ = ~new_new_n36420__ & ~new_new_n36421__;
  assign new_new_n36423__ = new_new_n36418__ & ~new_new_n36422__;
  assign new_new_n36424__ = pi23 & ~new_new_n36418__;
  assign new_new_n36425__ = ~new_new_n36423__ & ~new_new_n36424__;
  assign new_new_n36426__ = ~new_new_n36132__ & new_new_n36212__;
  assign new_new_n36427__ = ~new_new_n36131__ & ~new_new_n36426__;
  assign new_new_n36428__ = ~new_new_n36425__ & new_new_n36427__;
  assign new_new_n36429__ = new_new_n36425__ & ~new_new_n36427__;
  assign new_new_n36430__ = ~new_new_n36428__ & ~new_new_n36429__;
  assign new_new_n36431__ = ~new_new_n36413__ & ~new_new_n36430__;
  assign new_new_n36432__ = new_new_n36413__ & new_new_n36430__;
  assign new_new_n36433__ = ~new_new_n36431__ & ~new_new_n36432__;
  assign new_new_n36434__ = ~new_new_n36329__ & new_new_n36433__;
  assign new_new_n36435__ = new_new_n36329__ & ~new_new_n36433__;
  assign new_new_n36436__ = ~new_new_n36434__ & ~new_new_n36435__;
  assign new_new_n36437__ = new_new_n36251__ & new_new_n36436__;
  assign new_new_n36438__ = ~new_new_n36251__ & ~new_new_n36436__;
  assign new_new_n36439__ = ~new_new_n36437__ & ~new_new_n36438__;
  assign new_new_n36440__ = new_new_n36314__ & ~new_new_n36439__;
  assign new_new_n36441__ = ~new_new_n36314__ & new_new_n36439__;
  assign new_new_n36442__ = ~new_new_n36440__ & ~new_new_n36441__;
  assign new_new_n36443__ = ~new_new_n36304__ & new_new_n36442__;
  assign new_new_n36444__ = new_new_n36304__ & ~new_new_n36442__;
  assign new_new_n36445__ = ~new_new_n36443__ & ~new_new_n36444__;
  assign new_new_n36446__ = new_new_n36289__ & new_new_n36445__;
  assign new_new_n36447__ = ~new_new_n36289__ & ~new_new_n36445__;
  assign new_new_n36448__ = ~new_new_n36446__ & ~new_new_n36447__;
  assign new_new_n36449__ = new_new_n36256__ & new_new_n36271__;
  assign new_new_n36450__ = ~new_new_n36256__ & ~new_new_n36271__;
  assign new_new_n36451__ = ~new_new_n36273__ & ~new_new_n36450__;
  assign new_new_n36452__ = new_new_n36095__ & new_new_n36451__;
  assign new_new_n36453__ = pi11 & ~new_new_n36449__;
  assign new_new_n36454__ = ~new_new_n36452__ & new_new_n36453__;
  assign new_new_n36455__ = ~new_new_n36256__ & new_new_n36273__;
  assign new_new_n36456__ = ~new_new_n36095__ & ~new_new_n36451__;
  assign new_new_n36457__ = ~pi11 & ~new_new_n36455__;
  assign new_new_n36458__ = ~new_new_n36456__ & new_new_n36457__;
  assign new_new_n36459__ = ~new_new_n36454__ & ~new_new_n36458__;
  assign new_new_n36460__ = new_new_n36095__ & new_new_n36270__;
  assign new_new_n36461__ = new_new_n36256__ & ~new_new_n36261__;
  assign new_new_n36462__ = new_new_n36460__ & new_new_n36461__;
  assign new_new_n36463__ = ~new_new_n36287__ & ~new_new_n36448__;
  assign new_new_n36464__ = ~new_new_n36462__ & new_new_n36463__;
  assign new_new_n36465__ = ~new_new_n36459__ & new_new_n36464__;
  assign new_new_n36466__ = ~pi11 & ~new_new_n36258__;
  assign new_new_n36467__ = ~new_new_n36257__ & ~new_new_n36466__;
  assign new_new_n36468__ = new_new_n36273__ & new_new_n36467__;
  assign new_new_n36469__ = pi11 & ~new_new_n36095__;
  assign new_new_n36470__ = ~pi11 & new_new_n36095__;
  assign new_new_n36471__ = ~new_new_n36469__ & ~new_new_n36470__;
  assign new_new_n36472__ = ~new_new_n36259__ & new_new_n36471__;
  assign new_new_n36473__ = new_new_n36274__ & ~new_new_n36472__;
  assign new_new_n36474__ = new_new_n36271__ & ~new_new_n36467__;
  assign new_new_n36475__ = new_new_n36448__ & ~new_new_n36468__;
  assign new_new_n36476__ = ~new_new_n36474__ & new_new_n36475__;
  assign new_new_n36477__ = ~new_new_n36473__ & new_new_n36476__;
  assign new_new_n36478__ = ~new_new_n36465__ & ~new_new_n36477__;
  assign new_new_n36479__ = pi11 & ~new_new_n36271__;
  assign new_new_n36480__ = new_new_n36273__ & ~new_new_n36479__;
  assign new_new_n36481__ = ~new_new_n36273__ & new_new_n36479__;
  assign new_new_n36482__ = ~new_new_n36480__ & ~new_new_n36481__;
  assign new_new_n36483__ = new_new_n36259__ & new_new_n36482__;
  assign new_new_n36484__ = ~new_new_n36259__ & ~new_new_n36482__;
  assign new_new_n36485__ = ~new_new_n36483__ & ~new_new_n36484__;
  assign new_new_n36486__ = new_new_n36091__ & new_new_n36485__;
  assign new_new_n36487__ = ~new_new_n36478__ & new_new_n36486__;
  assign new_new_n36488__ = new_new_n36478__ & ~new_new_n36486__;
  assign po16 = ~new_new_n36487__ & ~new_new_n36488__;
  assign new_new_n36490__ = pi11 & ~new_new_n36285__;
  assign new_new_n36491__ = ~new_new_n36461__ & ~new_new_n36490__;
  assign new_new_n36492__ = ~new_new_n36448__ & new_new_n36491__;
  assign new_new_n36493__ = new_new_n36460__ & ~new_new_n36492__;
  assign new_new_n36494__ = ~new_new_n36285__ & new_new_n36448__;
  assign new_new_n36495__ = ~new_new_n36448__ & ~new_new_n36461__;
  assign new_new_n36496__ = pi11 & ~new_new_n36495__;
  assign new_new_n36497__ = ~new_new_n36494__ & ~new_new_n36496__;
  assign new_new_n36498__ = ~new_new_n36286__ & ~new_new_n36497__;
  assign new_new_n36499__ = new_new_n36448__ & ~new_new_n36491__;
  assign new_new_n36500__ = ~new_new_n36493__ & ~new_new_n36499__;
  assign new_new_n36501__ = ~new_new_n36498__ & new_new_n36500__;
  assign new_new_n36502__ = ~new_new_n36487__ & new_new_n36501__;
  assign new_new_n36503__ = ~new_new_n36327__ & new_new_n36433__;
  assign new_new_n36504__ = ~new_new_n36328__ & ~new_new_n36503__;
  assign new_new_n36505__ = new_new_n5183__ & new_new_n26722__;
  assign new_new_n36506__ = new_new_n5191__ & new_new_n26729__;
  assign new_new_n36507__ = ~new_new_n36505__ & ~new_new_n36506__;
  assign new_new_n36508__ = new_new_n5195__ & new_new_n27353__;
  assign new_new_n36509__ = new_new_n36507__ & ~new_new_n36508__;
  assign new_new_n36510__ = pi23 & ~new_new_n36509__;
  assign new_new_n36511__ = new_new_n5195__ & ~new_new_n27362__;
  assign new_new_n36512__ = ~pi23 & ~new_new_n36511__;
  assign new_new_n36513__ = pi22 & ~new_new_n27242__;
  assign new_new_n36514__ = ~pi22 & new_new_n27242__;
  assign new_new_n36515__ = ~new_new_n36513__ & ~new_new_n36514__;
  assign new_new_n36516__ = new_new_n5195__ & ~new_new_n36515__;
  assign new_new_n36517__ = new_new_n27352__ & new_new_n36516__;
  assign new_new_n36518__ = ~new_new_n36512__ & ~new_new_n36517__;
  assign new_new_n36519__ = new_new_n36507__ & ~new_new_n36518__;
  assign new_new_n36520__ = ~new_new_n36510__ & ~new_new_n36519__;
  assign new_new_n36521__ = new_new_n3311__ & new_new_n26774__;
  assign new_new_n36522__ = ~new_new_n333__ & ~new_new_n26802__;
  assign new_new_n36523__ = new_new_n873__ & new_new_n26810__;
  assign new_new_n36524__ = ~new_new_n36522__ & ~new_new_n36523__;
  assign new_new_n36525__ = ~new_new_n36521__ & new_new_n36524__;
  assign new_new_n36526__ = ~pi26 & ~new_new_n36525__;
  assign new_new_n36527__ = new_new_n512__ & ~new_new_n27373__;
  assign new_new_n36528__ = new_new_n801__ & ~new_new_n27373__;
  assign new_new_n36529__ = pi26 & ~new_new_n36528__;
  assign new_new_n36530__ = ~new_new_n36527__ & ~new_new_n36529__;
  assign new_new_n36531__ = new_new_n36525__ & ~new_new_n36530__;
  assign new_new_n36532__ = ~new_new_n36526__ & ~new_new_n36531__;
  assign new_new_n36533__ = new_new_n36341__ & ~new_new_n36389__;
  assign new_new_n36534__ = ~new_new_n36388__ & ~new_new_n36533__;
  assign new_new_n36535__ = new_new_n36532__ & new_new_n36534__;
  assign new_new_n36536__ = ~new_new_n36532__ & ~new_new_n36534__;
  assign new_new_n36537__ = ~new_new_n36535__ & ~new_new_n36536__;
  assign new_new_n36538__ = ~new_new_n36395__ & ~new_new_n36411__;
  assign new_new_n36539__ = ~new_new_n35993__ & ~new_new_n36378__;
  assign new_new_n36540__ = ~new_new_n36377__ & new_new_n36539__;
  assign new_new_n36541__ = ~new_new_n36343__ & ~new_new_n36540__;
  assign new_new_n36542__ = ~new_new_n36347__ & new_new_n36541__;
  assign new_new_n36543__ = new_new_n36358__ & ~new_new_n36542__;
  assign new_new_n36544__ = ~new_new_n36346__ & new_new_n36540__;
  assign new_new_n36545__ = ~new_new_n36343__ & ~new_new_n36358__;
  assign new_new_n36546__ = new_new_n35993__ & ~new_new_n36379__;
  assign new_new_n36547__ = ~new_new_n36545__ & new_new_n36546__;
  assign new_new_n36548__ = ~new_new_n36543__ & ~new_new_n36544__;
  assign new_new_n36549__ = ~new_new_n36547__ & new_new_n36548__;
  assign new_new_n36550__ = new_new_n4212__ & ~new_new_n27221__;
  assign new_new_n36551__ = ~new_new_n4818__ & ~new_new_n26823__;
  assign new_new_n36552__ = new_new_n4815__ & ~new_new_n26741__;
  assign new_new_n36553__ = ~new_new_n36550__ & ~new_new_n36551__;
  assign new_new_n36554__ = ~new_new_n36552__ & new_new_n36553__;
  assign new_new_n36555__ = new_new_n4214__ & new_new_n30393__;
  assign new_new_n36556__ = pi29 & ~new_new_n36555__;
  assign new_new_n36557__ = new_new_n4825__ & new_new_n30393__;
  assign new_new_n36558__ = ~new_new_n36556__ & ~new_new_n36557__;
  assign new_new_n36559__ = new_new_n36554__ & ~new_new_n36558__;
  assign new_new_n36560__ = ~pi29 & ~new_new_n36554__;
  assign new_new_n36561__ = ~new_new_n36559__ & ~new_new_n36560__;
  assign new_new_n36562__ = new_new_n71__ & ~new_new_n26854__;
  assign new_new_n36563__ = new_new_n765__ & new_new_n29424__;
  assign new_new_n36564__ = ~new_new_n36349__ & ~new_new_n36562__;
  assign new_new_n36565__ = ~new_new_n36563__ & new_new_n36564__;
  assign new_new_n36566__ = pi31 & ~new_new_n36565__;
  assign new_new_n36567__ = new_new_n161__ & new_new_n26854__;
  assign new_new_n36568__ = ~new_new_n161__ & ~new_new_n26847__;
  assign new_new_n36569__ = new_new_n4876__ & ~new_new_n36567__;
  assign new_new_n36570__ = ~new_new_n36568__ & new_new_n36569__;
  assign new_new_n36571__ = ~new_new_n36566__ & ~new_new_n36570__;
  assign new_new_n36572__ = ~new_new_n36561__ & ~new_new_n36571__;
  assign new_new_n36573__ = new_new_n36561__ & new_new_n36571__;
  assign new_new_n36574__ = ~new_new_n36572__ & ~new_new_n36573__;
  assign new_new_n36575__ = ~new_new_n36377__ & ~new_new_n36539__;
  assign new_new_n36576__ = ~new_new_n96__ & ~new_new_n127__;
  assign new_new_n36577__ = ~new_new_n309__ & new_new_n36576__;
  assign new_new_n36578__ = ~new_new_n952__ & ~new_new_n1130__;
  assign new_new_n36579__ = new_new_n6123__ & new_new_n36578__;
  assign new_new_n36580__ = ~new_new_n373__ & new_new_n36577__;
  assign new_new_n36581__ = ~new_new_n519__ & new_new_n1905__;
  assign new_new_n36582__ = new_new_n2643__ & new_new_n3793__;
  assign new_new_n36583__ = new_new_n36581__ & new_new_n36582__;
  assign new_new_n36584__ = new_new_n36579__ & new_new_n36580__;
  assign new_new_n36585__ = new_new_n4601__ & new_new_n36584__;
  assign new_new_n36586__ = new_new_n16489__ & new_new_n36583__;
  assign new_new_n36587__ = new_new_n36585__ & new_new_n36586__;
  assign new_new_n36588__ = new_new_n33421__ & new_new_n34004__;
  assign new_new_n36589__ = new_new_n36587__ & new_new_n36588__;
  assign new_new_n36590__ = new_new_n16202__ & new_new_n36589__;
  assign new_new_n36591__ = new_new_n18535__ & new_new_n36590__;
  assign new_new_n36592__ = new_new_n36575__ & ~new_new_n36591__;
  assign new_new_n36593__ = ~new_new_n36575__ & new_new_n36591__;
  assign new_new_n36594__ = ~new_new_n36592__ & ~new_new_n36593__;
  assign new_new_n36595__ = new_new_n36574__ & ~new_new_n36594__;
  assign new_new_n36596__ = ~new_new_n36574__ & new_new_n36594__;
  assign new_new_n36597__ = ~new_new_n36595__ & ~new_new_n36596__;
  assign new_new_n36598__ = new_new_n36549__ & new_new_n36597__;
  assign new_new_n36599__ = ~new_new_n36549__ & ~new_new_n36597__;
  assign new_new_n36600__ = ~new_new_n36598__ & ~new_new_n36599__;
  assign new_new_n36601__ = new_new_n36538__ & ~new_new_n36600__;
  assign new_new_n36602__ = ~new_new_n36538__ & new_new_n36600__;
  assign new_new_n36603__ = ~new_new_n36601__ & ~new_new_n36602__;
  assign new_new_n36604__ = new_new_n36537__ & new_new_n36603__;
  assign new_new_n36605__ = ~new_new_n36537__ & ~new_new_n36603__;
  assign new_new_n36606__ = ~new_new_n36604__ & ~new_new_n36605__;
  assign new_new_n36607__ = new_new_n36520__ & new_new_n36606__;
  assign new_new_n36608__ = ~new_new_n36520__ & ~new_new_n36606__;
  assign new_new_n36609__ = ~new_new_n36607__ & ~new_new_n36608__;
  assign new_new_n36610__ = new_new_n7935__ & new_new_n32729__;
  assign new_new_n36611__ = new_new_n6964__ & ~new_new_n26667__;
  assign new_new_n36612__ = new_new_n6968__ & new_new_n32382__;
  assign new_new_n36613__ = ~new_new_n36610__ & ~new_new_n36611__;
  assign new_new_n36614__ = ~new_new_n36612__ & new_new_n36613__;
  assign new_new_n36615__ = new_new_n6958__ & new_new_n32758__;
  assign new_new_n36616__ = pi17 & ~new_new_n36615__;
  assign new_new_n36617__ = new_new_n7942__ & new_new_n32758__;
  assign new_new_n36618__ = ~new_new_n36616__ & ~new_new_n36617__;
  assign new_new_n36619__ = new_new_n36614__ & ~new_new_n36618__;
  assign new_new_n36620__ = ~pi17 & ~new_new_n36614__;
  assign new_new_n36621__ = ~new_new_n36619__ & ~new_new_n36620__;
  assign new_new_n36622__ = ~new_new_n36609__ & new_new_n36621__;
  assign new_new_n36623__ = new_new_n36609__ & ~new_new_n36621__;
  assign new_new_n36624__ = ~new_new_n36622__ & ~new_new_n36623__;
  assign new_new_n36625__ = new_new_n6936__ & new_new_n27284__;
  assign new_new_n36626__ = new_new_n6629__ & new_new_n26698__;
  assign new_new_n36627__ = ~new_new_n6625__ & new_new_n27250__;
  assign new_new_n36628__ = new_new_n6634__ & ~new_new_n26674__;
  assign new_new_n36629__ = ~new_new_n36626__ & ~new_new_n36627__;
  assign new_new_n36630__ = ~new_new_n36628__ & new_new_n36629__;
  assign new_new_n36631__ = ~new_new_n36625__ & new_new_n36630__;
  assign new_new_n36632__ = pi20 & ~new_new_n36631__;
  assign new_new_n36633__ = ~pi20 & new_new_n36631__;
  assign new_new_n36634__ = ~new_new_n36632__ & ~new_new_n36633__;
  assign new_new_n36635__ = ~new_new_n36413__ & ~new_new_n36429__;
  assign new_new_n36636__ = ~new_new_n36428__ & ~new_new_n36635__;
  assign new_new_n36637__ = ~new_new_n36634__ & ~new_new_n36636__;
  assign new_new_n36638__ = new_new_n36634__ & new_new_n36636__;
  assign new_new_n36639__ = ~new_new_n36637__ & ~new_new_n36638__;
  assign new_new_n36640__ = new_new_n36624__ & ~new_new_n36639__;
  assign new_new_n36641__ = ~new_new_n36624__ & new_new_n36639__;
  assign new_new_n36642__ = ~new_new_n36640__ & ~new_new_n36641__;
  assign new_new_n36643__ = new_new_n36504__ & new_new_n36642__;
  assign new_new_n36644__ = ~new_new_n36504__ & ~new_new_n36642__;
  assign new_new_n36645__ = ~new_new_n36643__ & ~new_new_n36644__;
  assign new_new_n36646__ = ~new_new_n36314__ & ~new_new_n36437__;
  assign new_new_n36647__ = ~new_new_n36438__ & ~new_new_n36646__;
  assign new_new_n36648__ = ~new_new_n36645__ & ~new_new_n36647__;
  assign new_new_n36649__ = new_new_n36645__ & new_new_n36647__;
  assign new_new_n36650__ = ~new_new_n36648__ & ~new_new_n36649__;
  assign new_new_n36651__ = new_new_n6991__ & new_new_n32740__;
  assign new_new_n36652__ = ~pi14 & ~new_new_n36651__;
  assign new_new_n36653__ = new_new_n6991__ & new_new_n36096__;
  assign new_new_n36654__ = ~new_new_n36652__ & ~new_new_n36653__;
  assign new_new_n36655__ = ~new_new_n36650__ & new_new_n36654__;
  assign new_new_n36656__ = new_new_n36650__ & ~new_new_n36654__;
  assign new_new_n36657__ = ~new_new_n36655__ & ~new_new_n36656__;
  assign new_new_n36658__ = new_new_n36502__ & ~new_new_n36657__;
  assign new_new_n36659__ = new_new_n36444__ & new_new_n36658__;
  assign new_new_n36660__ = new_new_n36487__ & ~new_new_n36501__;
  assign new_new_n36661__ = ~new_new_n36502__ & ~new_new_n36660__;
  assign new_new_n36662__ = new_new_n36657__ & new_new_n36661__;
  assign new_new_n36663__ = ~new_new_n36658__ & ~new_new_n36662__;
  assign new_new_n36664__ = ~new_new_n36289__ & ~new_new_n36663__;
  assign new_new_n36665__ = ~new_new_n36657__ & new_new_n36660__;
  assign new_new_n36666__ = ~new_new_n36664__ & ~new_new_n36665__;
  assign new_new_n36667__ = ~new_new_n36443__ & ~new_new_n36666__;
  assign new_new_n36668__ = ~new_new_n36289__ & ~new_new_n36443__;
  assign new_new_n36669__ = ~new_new_n36444__ & ~new_new_n36668__;
  assign new_new_n36670__ = new_new_n36502__ & new_new_n36669__;
  assign new_new_n36671__ = new_new_n36289__ & ~new_new_n36304__;
  assign new_new_n36672__ = new_new_n36660__ & new_new_n36671__;
  assign new_new_n36673__ = ~new_new_n36670__ & ~new_new_n36672__;
  assign new_new_n36674__ = new_new_n36657__ & ~new_new_n36673__;
  assign new_new_n36675__ = ~new_new_n36657__ & ~new_new_n36669__;
  assign new_new_n36676__ = ~new_new_n36444__ & new_new_n36657__;
  assign new_new_n36677__ = ~new_new_n36675__ & ~new_new_n36676__;
  assign new_new_n36678__ = new_new_n36661__ & new_new_n36677__;
  assign new_new_n36679__ = ~new_new_n36659__ & ~new_new_n36678__;
  assign new_new_n36680__ = ~new_new_n36674__ & new_new_n36679__;
  assign po17 = new_new_n36667__ | ~new_new_n36680__;
  assign new_new_n36682__ = ~new_new_n36501__ & ~new_new_n36657__;
  assign new_new_n36683__ = new_new_n36671__ & new_new_n36682__;
  assign new_new_n36684__ = ~new_new_n36444__ & ~new_new_n36657__;
  assign new_new_n36685__ = new_new_n36657__ & ~new_new_n36669__;
  assign new_new_n36686__ = ~new_new_n36684__ & ~new_new_n36685__;
  assign new_new_n36687__ = new_new_n36501__ & new_new_n36686__;
  assign new_new_n36688__ = new_new_n36501__ & new_new_n36657__;
  assign new_new_n36689__ = new_new_n36289__ & ~new_new_n36657__;
  assign new_new_n36690__ = ~new_new_n36443__ & ~new_new_n36689__;
  assign new_new_n36691__ = ~new_new_n36682__ & new_new_n36690__;
  assign new_new_n36692__ = ~new_new_n36688__ & new_new_n36691__;
  assign new_new_n36693__ = ~new_new_n36683__ & ~new_new_n36687__;
  assign new_new_n36694__ = ~new_new_n36692__ & new_new_n36693__;
  assign new_new_n36695__ = new_new_n36487__ & ~new_new_n36694__;
  assign new_new_n36696__ = new_new_n7935__ & ~new_new_n32382__;
  assign new_new_n36697__ = pi17 & new_new_n36696__;
  assign new_new_n36698__ = new_new_n6959__ & new_new_n33050__;
  assign new_new_n36699__ = new_new_n6964__ & new_new_n32382__;
  assign new_new_n36700__ = ~new_new_n36698__ & ~new_new_n36699__;
  assign new_new_n36701__ = pi17 & new_new_n36700__;
  assign new_new_n36702__ = ~new_new_n36696__ & ~new_new_n36701__;
  assign new_new_n36703__ = ~new_new_n32729__ & ~new_new_n36697__;
  assign new_new_n36704__ = ~new_new_n36702__ & new_new_n36703__;
  assign new_new_n36705__ = new_new_n6968__ & new_new_n32729__;
  assign new_new_n36706__ = new_new_n36700__ & ~new_new_n36705__;
  assign new_new_n36707__ = ~pi17 & ~new_new_n36706__;
  assign new_new_n36708__ = ~new_new_n6968__ & new_new_n32729__;
  assign new_new_n36709__ = new_new_n36701__ & new_new_n36708__;
  assign new_new_n36710__ = ~new_new_n36707__ & ~new_new_n36709__;
  assign new_new_n36711__ = ~new_new_n36704__ & new_new_n36710__;
  assign new_new_n36712__ = new_new_n36538__ & new_new_n36606__;
  assign new_new_n36713__ = ~new_new_n36608__ & ~new_new_n36712__;
  assign new_new_n36714__ = new_new_n6629__ & ~new_new_n26674__;
  assign new_new_n36715__ = ~new_new_n6625__ & new_new_n26698__;
  assign new_new_n36716__ = new_new_n6936__ & ~new_new_n32340__;
  assign new_new_n36717__ = ~new_new_n36714__ & ~new_new_n36715__;
  assign new_new_n36718__ = ~new_new_n36716__ & new_new_n36717__;
  assign new_new_n36719__ = new_new_n6631__ & ~new_new_n26667__;
  assign new_new_n36720__ = ~pi20 & ~new_new_n36719__;
  assign new_new_n36721__ = new_new_n6640__ & ~new_new_n26667__;
  assign new_new_n36722__ = ~new_new_n36720__ & ~new_new_n36721__;
  assign new_new_n36723__ = new_new_n36718__ & ~new_new_n36722__;
  assign new_new_n36724__ = pi20 & ~new_new_n36718__;
  assign new_new_n36725__ = ~new_new_n36723__ & ~new_new_n36724__;
  assign new_new_n36726__ = new_new_n5191__ & new_new_n26722__;
  assign new_new_n36727__ = new_new_n5183__ & ~new_new_n27242__;
  assign new_new_n36728__ = new_new_n5215__ & ~new_new_n27271__;
  assign new_new_n36729__ = ~new_new_n36726__ & ~new_new_n36727__;
  assign new_new_n36730__ = ~new_new_n36728__ & new_new_n36729__;
  assign new_new_n36731__ = new_new_n5195__ & new_new_n27250__;
  assign new_new_n36732__ = pi23 & ~new_new_n36731__;
  assign new_new_n36733__ = new_new_n5974__ & new_new_n27250__;
  assign new_new_n36734__ = ~new_new_n36732__ & ~new_new_n36733__;
  assign new_new_n36735__ = new_new_n36730__ & ~new_new_n36734__;
  assign new_new_n36736__ = ~pi23 & ~new_new_n36730__;
  assign new_new_n36737__ = ~new_new_n36735__ & ~new_new_n36736__;
  assign new_new_n36738__ = ~new_new_n36536__ & new_new_n36600__;
  assign new_new_n36739__ = ~new_new_n36535__ & ~new_new_n36738__;
  assign new_new_n36740__ = new_new_n36737__ & ~new_new_n36739__;
  assign new_new_n36741__ = ~new_new_n36737__ & new_new_n36739__;
  assign new_new_n36742__ = ~new_new_n36740__ & ~new_new_n36741__;
  assign new_new_n36743__ = new_new_n873__ & new_new_n26774__;
  assign new_new_n36744__ = ~new_new_n333__ & new_new_n26810__;
  assign new_new_n36745__ = new_new_n3311__ & new_new_n26729__;
  assign new_new_n36746__ = ~new_new_n36743__ & ~new_new_n36744__;
  assign new_new_n36747__ = ~new_new_n36745__ & new_new_n36746__;
  assign new_new_n36748__ = ~pi26 & ~new_new_n36747__;
  assign new_new_n36749__ = new_new_n512__ & new_new_n30644__;
  assign new_new_n36750__ = new_new_n801__ & new_new_n30644__;
  assign new_new_n36751__ = pi26 & ~new_new_n36750__;
  assign new_new_n36752__ = ~new_new_n36749__ & ~new_new_n36751__;
  assign new_new_n36753__ = new_new_n36747__ & ~new_new_n36752__;
  assign new_new_n36754__ = ~new_new_n36748__ & ~new_new_n36753__;
  assign new_new_n36755__ = new_new_n36549__ & ~new_new_n36575__;
  assign new_new_n36756__ = ~new_new_n36549__ & new_new_n36575__;
  assign new_new_n36757__ = ~new_new_n36755__ & ~new_new_n36756__;
  assign new_new_n36758__ = ~new_new_n36594__ & ~new_new_n36757__;
  assign new_new_n36759__ = new_new_n36574__ & ~new_new_n36758__;
  assign new_new_n36760__ = ~new_new_n36549__ & ~new_new_n36593__;
  assign new_new_n36761__ = ~new_new_n36592__ & ~new_new_n36760__;
  assign new_new_n36762__ = ~new_new_n36573__ & new_new_n36761__;
  assign new_new_n36763__ = ~new_new_n36572__ & ~new_new_n36761__;
  assign new_new_n36764__ = ~new_new_n36762__ & ~new_new_n36763__;
  assign new_new_n36765__ = ~new_new_n36759__ & ~new_new_n36764__;
  assign new_new_n36766__ = new_new_n765__ & new_new_n29400__;
  assign new_new_n36767__ = ~new_new_n36567__ & ~new_new_n36766__;
  assign new_new_n36768__ = pi31 & ~new_new_n36767__;
  assign new_new_n36769__ = new_new_n161__ & new_new_n26847__;
  assign new_new_n36770__ = ~new_new_n71__ & new_new_n36769__;
  assign new_new_n36771__ = new_new_n71__ & ~new_new_n26847__;
  assign new_new_n36772__ = pi31 & ~new_new_n36771__;
  assign new_new_n36773__ = ~new_new_n15853__ & ~new_new_n26823__;
  assign new_new_n36774__ = ~new_new_n36770__ & ~new_new_n36772__;
  assign new_new_n36775__ = ~new_new_n36773__ & new_new_n36774__;
  assign new_new_n36776__ = ~new_new_n36768__ & ~new_new_n36775__;
  assign new_new_n36777__ = ~new_new_n375__ & ~new_new_n715__;
  assign new_new_n36778__ = ~new_new_n749__ & ~new_new_n933__;
  assign new_new_n36779__ = ~new_new_n1080__ & new_new_n36778__;
  assign new_new_n36780__ = ~new_new_n1167__ & new_new_n36777__;
  assign new_new_n36781__ = new_new_n36779__ & new_new_n36780__;
  assign new_new_n36782__ = ~new_new_n218__ & new_new_n1917__;
  assign new_new_n36783__ = new_new_n1947__ & new_new_n4458__;
  assign new_new_n36784__ = new_new_n36782__ & new_new_n36783__;
  assign new_new_n36785__ = new_new_n347__ & new_new_n36781__;
  assign new_new_n36786__ = new_new_n2867__ & new_new_n36785__;
  assign new_new_n36787__ = new_new_n36784__ & new_new_n36786__;
  assign new_new_n36788__ = new_new_n3647__ & new_new_n3803__;
  assign new_new_n36789__ = new_new_n3988__ & new_new_n6255__;
  assign new_new_n36790__ = new_new_n36788__ & new_new_n36789__;
  assign new_new_n36791__ = new_new_n36787__ & new_new_n36790__;
  assign new_new_n36792__ = new_new_n3090__ & new_new_n4436__;
  assign new_new_n36793__ = new_new_n36791__ & new_new_n36792__;
  assign new_new_n36794__ = ~new_new_n36776__ & new_new_n36793__;
  assign new_new_n36795__ = new_new_n36776__ & ~new_new_n36793__;
  assign new_new_n36796__ = ~new_new_n36794__ & ~new_new_n36795__;
  assign new_new_n36797__ = ~new_new_n36591__ & ~new_new_n36796__;
  assign new_new_n36798__ = ~new_new_n3090__ & new_new_n36776__;
  assign new_new_n36799__ = new_new_n36796__ & ~new_new_n36798__;
  assign new_new_n36800__ = new_new_n36591__ & new_new_n36799__;
  assign new_new_n36801__ = ~new_new_n36797__ & ~new_new_n36800__;
  assign new_new_n36802__ = ~new_new_n36765__ & ~new_new_n36801__;
  assign new_new_n36803__ = new_new_n36573__ & new_new_n36756__;
  assign new_new_n36804__ = ~new_new_n36549__ & new_new_n36573__;
  assign new_new_n36805__ = new_new_n36549__ & ~new_new_n36573__;
  assign new_new_n36806__ = ~new_new_n36572__ & new_new_n36575__;
  assign new_new_n36807__ = ~new_new_n36805__ & new_new_n36806__;
  assign new_new_n36808__ = ~new_new_n36804__ & ~new_new_n36807__;
  assign new_new_n36809__ = ~new_new_n36591__ & ~new_new_n36808__;
  assign new_new_n36810__ = new_new_n36572__ & new_new_n36755__;
  assign new_new_n36811__ = new_new_n36572__ & ~new_new_n36756__;
  assign new_new_n36812__ = ~new_new_n36573__ & new_new_n36755__;
  assign new_new_n36813__ = ~new_new_n36811__ & ~new_new_n36812__;
  assign new_new_n36814__ = new_new_n36591__ & ~new_new_n36813__;
  assign new_new_n36815__ = ~new_new_n36803__ & ~new_new_n36810__;
  assign new_new_n36816__ = ~new_new_n36814__ & new_new_n36815__;
  assign new_new_n36817__ = ~new_new_n36809__ & new_new_n36816__;
  assign new_new_n36818__ = new_new_n36801__ & ~new_new_n36817__;
  assign new_new_n36819__ = ~new_new_n36802__ & ~new_new_n36818__;
  assign new_new_n36820__ = new_new_n36754__ & new_new_n36819__;
  assign new_new_n36821__ = ~new_new_n36754__ & ~new_new_n36819__;
  assign new_new_n36822__ = ~new_new_n36820__ & ~new_new_n36821__;
  assign new_new_n36823__ = new_new_n4815__ & ~new_new_n26802__;
  assign new_new_n36824__ = ~new_new_n4818__ & ~new_new_n27221__;
  assign new_new_n36825__ = new_new_n4212__ & ~new_new_n26741__;
  assign new_new_n36826__ = ~new_new_n36824__ & ~new_new_n36825__;
  assign new_new_n36827__ = ~new_new_n36823__ & new_new_n36826__;
  assign new_new_n36828__ = new_new_n4214__ & new_new_n30411__;
  assign new_new_n36829__ = pi29 & ~new_new_n36828__;
  assign new_new_n36830__ = new_new_n4825__ & new_new_n30411__;
  assign new_new_n36831__ = ~new_new_n36829__ & ~new_new_n36830__;
  assign new_new_n36832__ = new_new_n36827__ & ~new_new_n36831__;
  assign new_new_n36833__ = ~pi29 & ~new_new_n36827__;
  assign new_new_n36834__ = ~new_new_n36832__ & ~new_new_n36833__;
  assign new_new_n36835__ = new_new_n36822__ & ~new_new_n36834__;
  assign new_new_n36836__ = ~new_new_n36822__ & new_new_n36834__;
  assign new_new_n36837__ = ~new_new_n36835__ & ~new_new_n36836__;
  assign new_new_n36838__ = new_new_n36742__ & new_new_n36837__;
  assign new_new_n36839__ = ~new_new_n36742__ & ~new_new_n36837__;
  assign new_new_n36840__ = ~new_new_n36838__ & ~new_new_n36839__;
  assign new_new_n36841__ = new_new_n36725__ & new_new_n36840__;
  assign new_new_n36842__ = ~new_new_n36725__ & ~new_new_n36840__;
  assign new_new_n36843__ = ~new_new_n36841__ & ~new_new_n36842__;
  assign new_new_n36844__ = ~new_new_n36713__ & ~new_new_n36843__;
  assign new_new_n36845__ = new_new_n36713__ & new_new_n36843__;
  assign new_new_n36846__ = ~new_new_n36844__ & ~new_new_n36845__;
  assign new_new_n36847__ = new_new_n36711__ & ~new_new_n36846__;
  assign new_new_n36848__ = ~new_new_n36711__ & new_new_n36846__;
  assign new_new_n36849__ = ~new_new_n36847__ & ~new_new_n36848__;
  assign new_new_n36850__ = ~new_new_n36609__ & ~new_new_n36637__;
  assign new_new_n36851__ = ~new_new_n36638__ & ~new_new_n36850__;
  assign new_new_n36852__ = ~new_new_n36849__ & new_new_n36851__;
  assign new_new_n36853__ = new_new_n36849__ & ~new_new_n36851__;
  assign new_new_n36854__ = ~new_new_n36852__ & ~new_new_n36853__;
  assign new_new_n36855__ = ~new_new_n36504__ & ~new_new_n36621__;
  assign new_new_n36856__ = new_new_n36504__ & new_new_n36621__;
  assign new_new_n36857__ = ~new_new_n36609__ & ~new_new_n36639__;
  assign new_new_n36858__ = new_new_n36609__ & new_new_n36639__;
  assign new_new_n36859__ = ~new_new_n36857__ & ~new_new_n36858__;
  assign new_new_n36860__ = ~new_new_n36856__ & ~new_new_n36859__;
  assign new_new_n36861__ = ~new_new_n36855__ & ~new_new_n36860__;
  assign new_new_n36862__ = ~new_new_n36854__ & new_new_n36861__;
  assign new_new_n36863__ = new_new_n36854__ & ~new_new_n36861__;
  assign new_new_n36864__ = ~new_new_n36862__ & ~new_new_n36863__;
  assign new_new_n36865__ = pi14 & new_new_n36864__;
  assign new_new_n36866__ = ~pi14 & ~new_new_n36864__;
  assign new_new_n36867__ = ~new_new_n36865__ & ~new_new_n36866__;
  assign new_new_n36868__ = new_new_n36669__ & ~new_new_n36688__;
  assign new_new_n36869__ = ~new_new_n36682__ & ~new_new_n36868__;
  assign new_new_n36870__ = ~new_new_n36867__ & new_new_n36869__;
  assign new_new_n36871__ = new_new_n36867__ & ~new_new_n36869__;
  assign new_new_n36872__ = ~new_new_n36870__ & ~new_new_n36871__;
  assign new_new_n36873__ = ~new_new_n36648__ & ~new_new_n36654__;
  assign new_new_n36874__ = ~new_new_n36649__ & ~new_new_n36873__;
  assign new_new_n36875__ = ~new_new_n36872__ & ~new_new_n36874__;
  assign new_new_n36876__ = new_new_n36872__ & new_new_n36874__;
  assign new_new_n36877__ = ~new_new_n36875__ & ~new_new_n36876__;
  assign new_new_n36878__ = new_new_n36695__ & new_new_n36877__;
  assign new_new_n36879__ = ~new_new_n36695__ & ~new_new_n36877__;
  assign po18 = ~new_new_n36878__ & ~new_new_n36879__;
  assign new_new_n36881__ = new_new_n36867__ & new_new_n36874__;
  assign new_new_n36882__ = ~new_new_n36869__ & new_new_n36881__;
  assign new_new_n36883__ = ~po18 & new_new_n36882__;
  assign new_new_n36884__ = ~new_new_n36874__ & new_new_n36877__;
  assign new_new_n36885__ = ~new_new_n36870__ & ~new_new_n36884__;
  assign new_new_n36886__ = ~new_new_n36878__ & ~new_new_n36885__;
  assign new_new_n36887__ = ~new_new_n36883__ & ~new_new_n36886__;
  assign new_new_n36888__ = ~new_new_n36848__ & new_new_n36851__;
  assign new_new_n36889__ = ~new_new_n36847__ & ~new_new_n36888__;
  assign new_new_n36890__ = new_new_n6936__ & ~new_new_n33347__;
  assign new_new_n36891__ = new_new_n6629__ & ~new_new_n26667__;
  assign new_new_n36892__ = ~new_new_n6625__ & ~new_new_n26674__;
  assign new_new_n36893__ = new_new_n6634__ & new_new_n32382__;
  assign new_new_n36894__ = ~new_new_n36891__ & ~new_new_n36892__;
  assign new_new_n36895__ = ~new_new_n36893__ & new_new_n36894__;
  assign new_new_n36896__ = ~new_new_n36890__ & new_new_n36895__;
  assign new_new_n36897__ = ~pi20 & ~new_new_n36896__;
  assign new_new_n36898__ = pi20 & new_new_n36896__;
  assign new_new_n36899__ = ~new_new_n36897__ & ~new_new_n36898__;
  assign new_new_n36900__ = ~new_new_n36841__ & ~new_new_n36845__;
  assign new_new_n36901__ = ~new_new_n36899__ & ~new_new_n36900__;
  assign new_new_n36902__ = new_new_n36899__ & new_new_n36900__;
  assign new_new_n36903__ = ~new_new_n36901__ & ~new_new_n36902__;
  assign new_new_n36904__ = new_new_n5183__ & new_new_n27250__;
  assign new_new_n36905__ = new_new_n5191__ & ~new_new_n27242__;
  assign new_new_n36906__ = ~new_new_n36904__ & ~new_new_n36905__;
  assign new_new_n36907__ = new_new_n5195__ & new_new_n26698__;
  assign new_new_n36908__ = new_new_n31511__ & new_new_n36907__;
  assign new_new_n36909__ = new_new_n36906__ & ~new_new_n36908__;
  assign new_new_n36910__ = pi23 & ~new_new_n36909__;
  assign new_new_n36911__ = new_new_n5195__ & ~new_new_n31510__;
  assign new_new_n36912__ = ~pi23 & ~new_new_n36911__;
  assign new_new_n36913__ = ~pi22 & ~new_new_n34204__;
  assign new_new_n36914__ = pi22 & ~new_new_n31509__;
  assign new_new_n36915__ = new_new_n5195__ & ~new_new_n36913__;
  assign new_new_n36916__ = ~new_new_n36914__ & new_new_n36915__;
  assign new_new_n36917__ = ~new_new_n36912__ & ~new_new_n36916__;
  assign new_new_n36918__ = new_new_n36906__ & ~new_new_n36917__;
  assign new_new_n36919__ = ~new_new_n36910__ & ~new_new_n36918__;
  assign new_new_n36920__ = ~new_new_n36741__ & ~new_new_n36837__;
  assign new_new_n36921__ = ~new_new_n36740__ & ~new_new_n36920__;
  assign new_new_n36922__ = ~new_new_n36919__ & ~new_new_n36921__;
  assign new_new_n36923__ = new_new_n36919__ & new_new_n36921__;
  assign new_new_n36924__ = ~new_new_n36922__ & ~new_new_n36923__;
  assign new_new_n36925__ = new_new_n3311__ & new_new_n26722__;
  assign new_new_n36926__ = ~new_new_n333__ & new_new_n26774__;
  assign new_new_n36927__ = new_new_n873__ & new_new_n26729__;
  assign new_new_n36928__ = ~new_new_n36926__ & ~new_new_n36927__;
  assign new_new_n36929__ = ~new_new_n36925__ & new_new_n36928__;
  assign new_new_n36930__ = pi26 & ~new_new_n36929__;
  assign new_new_n36931__ = new_new_n4898__ & ~new_new_n27348__;
  assign new_new_n36932__ = new_new_n801__ & ~new_new_n27348__;
  assign new_new_n36933__ = ~pi26 & ~new_new_n36932__;
  assign new_new_n36934__ = ~new_new_n36931__ & ~new_new_n36933__;
  assign new_new_n36935__ = new_new_n36929__ & ~new_new_n36934__;
  assign new_new_n36936__ = ~new_new_n36930__ & ~new_new_n36935__;
  assign new_new_n36937__ = new_new_n4815__ & new_new_n26810__;
  assign new_new_n36938__ = new_new_n4212__ & ~new_new_n26802__;
  assign new_new_n36939__ = new_new_n4813__ & new_new_n27395__;
  assign new_new_n36940__ = ~new_new_n36937__ & ~new_new_n36938__;
  assign new_new_n36941__ = ~new_new_n36939__ & new_new_n36940__;
  assign new_new_n36942__ = new_new_n67__ & ~new_new_n26741__;
  assign new_new_n36943__ = pi29 & ~new_new_n36942__;
  assign new_new_n36944__ = new_new_n65__ & ~new_new_n26741__;
  assign new_new_n36945__ = ~pi29 & ~new_new_n36944__;
  assign new_new_n36946__ = pi26 & ~new_new_n36945__;
  assign new_new_n36947__ = ~new_new_n36943__ & ~new_new_n36946__;
  assign new_new_n36948__ = new_new_n36941__ & ~new_new_n36947__;
  assign new_new_n36949__ = ~pi29 & ~new_new_n36941__;
  assign new_new_n36950__ = ~new_new_n36948__ & ~new_new_n36949__;
  assign new_new_n36951__ = ~new_new_n36762__ & ~new_new_n36801__;
  assign new_new_n36952__ = new_new_n36573__ & ~new_new_n36761__;
  assign new_new_n36953__ = ~new_new_n36755__ & ~new_new_n36801__;
  assign new_new_n36954__ = ~new_new_n36591__ & new_new_n36756__;
  assign new_new_n36955__ = ~new_new_n36797__ & ~new_new_n36954__;
  assign new_new_n36956__ = ~new_new_n36953__ & new_new_n36955__;
  assign new_new_n36957__ = ~new_new_n36572__ & ~new_new_n36956__;
  assign new_new_n36958__ = ~new_new_n36951__ & ~new_new_n36952__;
  assign new_new_n36959__ = ~new_new_n36957__ & new_new_n36958__;
  assign new_new_n36960__ = ~new_new_n36950__ & new_new_n36959__;
  assign new_new_n36961__ = new_new_n36950__ & ~new_new_n36959__;
  assign new_new_n36962__ = ~new_new_n36960__ & ~new_new_n36961__;
  assign new_new_n36963__ = ~pi14 & ~new_new_n36776__;
  assign new_new_n36964__ = pi14 & ~new_new_n36794__;
  assign new_new_n36965__ = new_new_n36591__ & ~new_new_n36963__;
  assign new_new_n36966__ = ~new_new_n36964__ & new_new_n36965__;
  assign new_new_n36967__ = ~pi14 & new_new_n36799__;
  assign new_new_n36968__ = pi14 & new_new_n36795__;
  assign new_new_n36969__ = ~new_new_n36963__ & ~new_new_n36968__;
  assign new_new_n36970__ = ~new_new_n36591__ & ~new_new_n36969__;
  assign new_new_n36971__ = new_new_n161__ & ~new_new_n26823__;
  assign new_new_n36972__ = new_new_n765__ & ~new_new_n27221__;
  assign new_new_n36973__ = ~new_new_n36971__ & ~new_new_n36972__;
  assign new_new_n36974__ = ~pi31 & ~new_new_n36973__;
  assign new_new_n36975__ = new_new_n71__ & ~new_new_n26823__;
  assign new_new_n36976__ = new_new_n765__ & new_new_n27411__;
  assign new_new_n36977__ = ~new_new_n36769__ & ~new_new_n36975__;
  assign new_new_n36978__ = ~new_new_n36976__ & new_new_n36977__;
  assign new_new_n36979__ = pi31 & ~new_new_n36978__;
  assign new_new_n36980__ = ~new_new_n36974__ & ~new_new_n36979__;
  assign new_new_n36981__ = ~new_new_n322__ & ~new_new_n785__;
  assign new_new_n36982__ = ~new_new_n329__ & new_new_n934__;
  assign new_new_n36983__ = new_new_n1740__ & new_new_n36982__;
  assign new_new_n36984__ = ~new_new_n676__ & new_new_n36981__;
  assign new_new_n36985__ = new_new_n4233__ & new_new_n36984__;
  assign new_new_n36986__ = new_new_n1001__ & new_new_n36983__;
  assign new_new_n36987__ = new_new_n3132__ & new_new_n36986__;
  assign new_new_n36988__ = new_new_n1644__ & new_new_n36985__;
  assign new_new_n36989__ = new_new_n36987__ & new_new_n36988__;
  assign new_new_n36990__ = new_new_n7613__ & new_new_n17601__;
  assign new_new_n36991__ = new_new_n36989__ & new_new_n36990__;
  assign new_new_n36992__ = new_new_n17274__ & new_new_n36991__;
  assign new_new_n36993__ = new_new_n3512__ & new_new_n36992__;
  assign new_new_n36994__ = ~new_new_n36980__ & new_new_n36993__;
  assign new_new_n36995__ = new_new_n36980__ & ~new_new_n36993__;
  assign new_new_n36996__ = ~new_new_n36994__ & ~new_new_n36995__;
  assign new_new_n36997__ = ~new_new_n36966__ & new_new_n36996__;
  assign new_new_n36998__ = ~new_new_n36967__ & new_new_n36997__;
  assign new_new_n36999__ = ~new_new_n36970__ & new_new_n36998__;
  assign new_new_n37000__ = new_new_n36591__ & ~new_new_n36794__;
  assign new_new_n37001__ = ~new_new_n36591__ & ~new_new_n36795__;
  assign new_new_n37002__ = ~new_new_n36798__ & new_new_n37001__;
  assign new_new_n37003__ = ~new_new_n37000__ & ~new_new_n37002__;
  assign new_new_n37004__ = pi14 & ~new_new_n37003__;
  assign new_new_n37005__ = ~pi14 & ~new_new_n37000__;
  assign new_new_n37006__ = ~new_new_n37001__ & new_new_n37005__;
  assign new_new_n37007__ = ~new_new_n36996__ & ~new_new_n37006__;
  assign new_new_n37008__ = ~new_new_n37004__ & new_new_n37007__;
  assign new_new_n37009__ = ~new_new_n36999__ & ~new_new_n37008__;
  assign new_new_n37010__ = ~new_new_n36962__ & new_new_n37009__;
  assign new_new_n37011__ = new_new_n36962__ & ~new_new_n37009__;
  assign new_new_n37012__ = ~new_new_n37010__ & ~new_new_n37011__;
  assign new_new_n37013__ = ~new_new_n36936__ & ~new_new_n37012__;
  assign new_new_n37014__ = new_new_n36936__ & new_new_n37012__;
  assign new_new_n37015__ = ~new_new_n37013__ & ~new_new_n37014__;
  assign new_new_n37016__ = ~new_new_n36820__ & ~new_new_n36834__;
  assign new_new_n37017__ = ~new_new_n36821__ & ~new_new_n37016__;
  assign new_new_n37018__ = new_new_n37015__ & ~new_new_n37017__;
  assign new_new_n37019__ = ~new_new_n37015__ & new_new_n37017__;
  assign new_new_n37020__ = ~new_new_n37018__ & ~new_new_n37019__;
  assign new_new_n37021__ = new_new_n36924__ & ~new_new_n37020__;
  assign new_new_n37022__ = ~new_new_n36924__ & new_new_n37020__;
  assign new_new_n37023__ = ~new_new_n37021__ & ~new_new_n37022__;
  assign new_new_n37024__ = new_new_n36903__ & new_new_n37023__;
  assign new_new_n37025__ = ~new_new_n36903__ & ~new_new_n37023__;
  assign new_new_n37026__ = ~new_new_n37024__ & ~new_new_n37025__;
  assign new_new_n37027__ = ~new_new_n36889__ & new_new_n37026__;
  assign new_new_n37028__ = new_new_n36889__ & ~new_new_n37026__;
  assign new_new_n37029__ = ~new_new_n37027__ & ~new_new_n37028__;
  assign new_new_n37030__ = new_new_n6964__ & new_new_n32729__;
  assign new_new_n37031__ = new_new_n6968__ & new_new_n32740__;
  assign new_new_n37032__ = ~new_new_n37030__ & ~new_new_n37031__;
  assign new_new_n37033__ = new_new_n6958__ & ~new_new_n34178__;
  assign new_new_n37034__ = pi17 & ~new_new_n37033__;
  assign new_new_n37035__ = new_new_n7942__ & ~new_new_n34178__;
  assign new_new_n37036__ = ~new_new_n37034__ & ~new_new_n37035__;
  assign new_new_n37037__ = new_new_n37032__ & ~new_new_n37036__;
  assign new_new_n37038__ = ~pi17 & ~new_new_n37032__;
  assign new_new_n37039__ = ~new_new_n37037__ & ~new_new_n37038__;
  assign new_new_n37040__ = new_new_n37029__ & new_new_n37039__;
  assign new_new_n37041__ = ~new_new_n37029__ & ~new_new_n37039__;
  assign new_new_n37042__ = ~new_new_n37040__ & ~new_new_n37041__;
  assign new_new_n37043__ = ~pi14 & ~new_new_n36863__;
  assign new_new_n37044__ = ~new_new_n36862__ & ~new_new_n37043__;
  assign new_new_n37045__ = new_new_n37042__ & new_new_n37044__;
  assign new_new_n37046__ = ~new_new_n37042__ & ~new_new_n37044__;
  assign new_new_n37047__ = ~new_new_n37045__ & ~new_new_n37046__;
  assign new_new_n37048__ = ~new_new_n36887__ & ~new_new_n37047__;
  assign new_new_n37049__ = new_new_n36870__ & ~new_new_n36874__;
  assign new_new_n37050__ = ~new_new_n36882__ & ~new_new_n37049__;
  assign new_new_n37051__ = new_new_n36695__ & ~new_new_n37050__;
  assign new_new_n37052__ = ~new_new_n36869__ & ~new_new_n36877__;
  assign new_new_n37053__ = ~new_new_n36695__ & ~new_new_n36881__;
  assign new_new_n37054__ = ~new_new_n37052__ & new_new_n37053__;
  assign new_new_n37055__ = new_new_n37047__ & ~new_new_n37051__;
  assign new_new_n37056__ = ~new_new_n37054__ & new_new_n37055__;
  assign po19 = new_new_n37048__ | new_new_n37056__;
  assign new_new_n37058__ = new_new_n36861__ & ~new_new_n36874__;
  assign new_new_n37059__ = ~new_new_n36861__ & new_new_n36874__;
  assign new_new_n37060__ = ~pi14 & ~new_new_n37059__;
  assign new_new_n37061__ = new_new_n36854__ & ~new_new_n36869__;
  assign new_new_n37062__ = new_new_n37042__ & ~new_new_n37061__;
  assign new_new_n37063__ = ~new_new_n37058__ & ~new_new_n37060__;
  assign new_new_n37064__ = ~new_new_n37062__ & new_new_n37063__;
  assign new_new_n37065__ = ~new_new_n36854__ & new_new_n36869__;
  assign new_new_n37066__ = ~new_new_n37042__ & ~new_new_n37058__;
  assign new_new_n37067__ = new_new_n37042__ & ~new_new_n37059__;
  assign new_new_n37068__ = pi14 & ~new_new_n37067__;
  assign new_new_n37069__ = ~new_new_n37066__ & ~new_new_n37068__;
  assign new_new_n37070__ = ~new_new_n37065__ & ~new_new_n37069__;
  assign new_new_n37071__ = ~new_new_n37042__ & new_new_n37061__;
  assign new_new_n37072__ = ~new_new_n37070__ & ~new_new_n37071__;
  assign new_new_n37073__ = ~new_new_n37064__ & new_new_n37072__;
  assign new_new_n37074__ = ~new_new_n36902__ & ~new_new_n37023__;
  assign new_new_n37075__ = ~new_new_n36901__ & ~new_new_n37074__;
  assign new_new_n37076__ = new_new_n6629__ & new_new_n32382__;
  assign new_new_n37077__ = ~new_new_n6625__ & ~new_new_n26667__;
  assign new_new_n37078__ = new_new_n6634__ & new_new_n32729__;
  assign new_new_n37079__ = ~new_new_n37076__ & ~new_new_n37077__;
  assign new_new_n37080__ = ~new_new_n37078__ & new_new_n37079__;
  assign new_new_n37081__ = new_new_n6631__ & new_new_n32758__;
  assign new_new_n37082__ = ~pi20 & ~new_new_n37081__;
  assign new_new_n37083__ = new_new_n7015__ & new_new_n32758__;
  assign new_new_n37084__ = ~new_new_n37082__ & ~new_new_n37083__;
  assign new_new_n37085__ = new_new_n37080__ & ~new_new_n37084__;
  assign new_new_n37086__ = pi20 & ~new_new_n37080__;
  assign new_new_n37087__ = ~new_new_n37085__ & ~new_new_n37086__;
  assign new_new_n37088__ = new_new_n5213__ & ~new_new_n26674__;
  assign new_new_n37089__ = new_new_n5183__ & new_new_n26698__;
  assign new_new_n37090__ = new_new_n5215__ & new_new_n27284__;
  assign new_new_n37091__ = ~new_new_n37088__ & ~new_new_n37089__;
  assign new_new_n37092__ = ~new_new_n37090__ & new_new_n37091__;
  assign new_new_n37093__ = new_new_n5185__ & new_new_n27250__;
  assign new_new_n37094__ = pi23 & ~new_new_n37093__;
  assign new_new_n37095__ = new_new_n5188__ & new_new_n27250__;
  assign new_new_n37096__ = ~pi23 & ~new_new_n37095__;
  assign new_new_n37097__ = pi20 & ~new_new_n37096__;
  assign new_new_n37098__ = ~new_new_n37094__ & ~new_new_n37097__;
  assign new_new_n37099__ = new_new_n37092__ & ~new_new_n37098__;
  assign new_new_n37100__ = ~pi23 & ~new_new_n37092__;
  assign new_new_n37101__ = ~new_new_n37099__ & ~new_new_n37100__;
  assign new_new_n37102__ = ~new_new_n333__ & new_new_n26729__;
  assign new_new_n37103__ = new_new_n873__ & new_new_n26722__;
  assign new_new_n37104__ = ~new_new_n37102__ & ~new_new_n37103__;
  assign new_new_n37105__ = new_new_n801__ & new_new_n27353__;
  assign new_new_n37106__ = new_new_n37104__ & ~new_new_n37105__;
  assign new_new_n37107__ = pi26 & ~new_new_n37106__;
  assign new_new_n37108__ = pi25 & new_new_n27242__;
  assign new_new_n37109__ = ~pi25 & ~new_new_n27242__;
  assign new_new_n37110__ = ~new_new_n110__ & ~new_new_n37108__;
  assign new_new_n37111__ = ~new_new_n37109__ & new_new_n37110__;
  assign new_new_n37112__ = new_new_n27352__ & new_new_n37111__;
  assign new_new_n37113__ = new_new_n801__ & ~new_new_n27362__;
  assign new_new_n37114__ = ~pi26 & ~new_new_n37113__;
  assign new_new_n37115__ = ~new_new_n37112__ & ~new_new_n37114__;
  assign new_new_n37116__ = new_new_n37104__ & ~new_new_n37115__;
  assign new_new_n37117__ = ~new_new_n37107__ & ~new_new_n37116__;
  assign new_new_n37118__ = ~new_new_n130__ & ~new_new_n438__;
  assign new_new_n37119__ = new_new_n1085__ & new_new_n37118__;
  assign new_new_n37120__ = new_new_n2332__ & new_new_n3430__;
  assign new_new_n37121__ = new_new_n4253__ & new_new_n7155__;
  assign new_new_n37122__ = new_new_n37120__ & new_new_n37121__;
  assign new_new_n37123__ = new_new_n960__ & new_new_n37119__;
  assign new_new_n37124__ = ~new_new_n1105__ & new_new_n1943__;
  assign new_new_n37125__ = new_new_n2453__ & new_new_n37124__;
  assign new_new_n37126__ = new_new_n37122__ & new_new_n37123__;
  assign new_new_n37127__ = new_new_n3099__ & new_new_n3649__;
  assign new_new_n37128__ = new_new_n37126__ & new_new_n37127__;
  assign new_new_n37129__ = new_new_n6817__ & new_new_n37125__;
  assign new_new_n37130__ = new_new_n37128__ & new_new_n37129__;
  assign new_new_n37131__ = new_new_n17544__ & new_new_n37130__;
  assign new_new_n37132__ = new_new_n6121__ & new_new_n37131__;
  assign new_new_n37133__ = new_new_n2987__ & new_new_n37132__;
  assign new_new_n37134__ = ~pi14 & ~new_new_n36993__;
  assign new_new_n37135__ = pi14 & new_new_n36993__;
  assign new_new_n37136__ = ~new_new_n36591__ & ~new_new_n37135__;
  assign new_new_n37137__ = ~new_new_n37134__ & ~new_new_n37136__;
  assign new_new_n37138__ = new_new_n37133__ & new_new_n37137__;
  assign new_new_n37139__ = ~new_new_n37133__ & ~new_new_n37137__;
  assign new_new_n37140__ = ~new_new_n37138__ & ~new_new_n37139__;
  assign new_new_n37141__ = new_new_n5021__ & ~new_new_n26741__;
  assign new_new_n37142__ = new_new_n765__ & new_new_n30393__;
  assign new_new_n37143__ = ~new_new_n36971__ & ~new_new_n37142__;
  assign new_new_n37144__ = pi31 & ~new_new_n37143__;
  assign new_new_n37145__ = new_new_n5053__ & ~new_new_n27221__;
  assign new_new_n37146__ = ~new_new_n37141__ & ~new_new_n37145__;
  assign new_new_n37147__ = ~new_new_n37144__ & new_new_n37146__;
  assign new_new_n37148__ = ~new_new_n37140__ & new_new_n37147__;
  assign new_new_n37149__ = new_new_n37140__ & ~new_new_n37147__;
  assign new_new_n37150__ = ~new_new_n37148__ & ~new_new_n37149__;
  assign new_new_n37151__ = new_new_n4813__ & ~new_new_n27373__;
  assign new_new_n37152__ = ~new_new_n4818__ & ~new_new_n26802__;
  assign new_new_n37153__ = new_new_n4212__ & new_new_n26810__;
  assign new_new_n37154__ = ~new_new_n37152__ & ~new_new_n37153__;
  assign new_new_n37155__ = ~new_new_n37151__ & new_new_n37154__;
  assign new_new_n37156__ = new_new_n4214__ & new_new_n26774__;
  assign new_new_n37157__ = ~pi29 & ~new_new_n37156__;
  assign new_new_n37158__ = new_new_n4825__ & new_new_n26774__;
  assign new_new_n37159__ = ~new_new_n37157__ & ~new_new_n37158__;
  assign new_new_n37160__ = new_new_n37155__ & ~new_new_n37159__;
  assign new_new_n37161__ = pi29 & ~new_new_n37155__;
  assign new_new_n37162__ = ~new_new_n37160__ & ~new_new_n37161__;
  assign new_new_n37163__ = new_new_n36795__ & ~new_new_n36980__;
  assign new_new_n37164__ = new_new_n36794__ & new_new_n36980__;
  assign new_new_n37165__ = ~new_new_n36794__ & ~new_new_n36980__;
  assign new_new_n37166__ = ~new_new_n37134__ & ~new_new_n37135__;
  assign new_new_n37167__ = ~new_new_n37165__ & ~new_new_n37166__;
  assign new_new_n37168__ = new_new_n36591__ & ~new_new_n37164__;
  assign new_new_n37169__ = ~new_new_n37167__ & new_new_n37168__;
  assign new_new_n37170__ = ~new_new_n36795__ & new_new_n36980__;
  assign new_new_n37171__ = ~new_new_n36591__ & ~new_new_n37166__;
  assign new_new_n37172__ = ~new_new_n37170__ & new_new_n37171__;
  assign new_new_n37173__ = ~new_new_n37163__ & ~new_new_n37172__;
  assign new_new_n37174__ = ~new_new_n37169__ & new_new_n37173__;
  assign new_new_n37175__ = ~new_new_n37162__ & new_new_n37174__;
  assign new_new_n37176__ = new_new_n37162__ & ~new_new_n37174__;
  assign new_new_n37177__ = ~new_new_n37175__ & ~new_new_n37176__;
  assign new_new_n37178__ = new_new_n37150__ & new_new_n37177__;
  assign new_new_n37179__ = ~new_new_n37150__ & ~new_new_n37177__;
  assign new_new_n37180__ = ~new_new_n37178__ & ~new_new_n37179__;
  assign new_new_n37181__ = new_new_n37117__ & ~new_new_n37180__;
  assign new_new_n37182__ = ~new_new_n37117__ & new_new_n37180__;
  assign new_new_n37183__ = ~new_new_n37181__ & ~new_new_n37182__;
  assign new_new_n37184__ = ~new_new_n36960__ & new_new_n37009__;
  assign new_new_n37185__ = ~new_new_n36961__ & ~new_new_n37184__;
  assign new_new_n37186__ = new_new_n37183__ & ~new_new_n37185__;
  assign new_new_n37187__ = ~new_new_n37183__ & new_new_n37185__;
  assign new_new_n37188__ = ~new_new_n37186__ & ~new_new_n37187__;
  assign new_new_n37189__ = ~new_new_n37101__ & ~new_new_n37188__;
  assign new_new_n37190__ = new_new_n37101__ & new_new_n37188__;
  assign new_new_n37191__ = ~new_new_n37189__ & ~new_new_n37190__;
  assign new_new_n37192__ = ~new_new_n37013__ & ~new_new_n37017__;
  assign new_new_n37193__ = ~new_new_n37014__ & ~new_new_n37192__;
  assign new_new_n37194__ = new_new_n37191__ & ~new_new_n37193__;
  assign new_new_n37195__ = ~new_new_n37191__ & new_new_n37193__;
  assign new_new_n37196__ = ~new_new_n37194__ & ~new_new_n37195__;
  assign new_new_n37197__ = new_new_n37087__ & new_new_n37196__;
  assign new_new_n37198__ = ~new_new_n37087__ & ~new_new_n37196__;
  assign new_new_n37199__ = ~new_new_n37197__ & ~new_new_n37198__;
  assign new_new_n37200__ = ~new_new_n36923__ & ~new_new_n37020__;
  assign new_new_n37201__ = ~new_new_n36922__ & ~new_new_n37200__;
  assign new_new_n37202__ = new_new_n37199__ & ~new_new_n37201__;
  assign new_new_n37203__ = ~new_new_n37199__ & new_new_n37201__;
  assign new_new_n37204__ = ~new_new_n37202__ & ~new_new_n37203__;
  assign new_new_n37205__ = ~new_new_n37075__ & ~new_new_n37204__;
  assign new_new_n37206__ = new_new_n37075__ & new_new_n37204__;
  assign new_new_n37207__ = ~new_new_n37205__ & ~new_new_n37206__;
  assign new_new_n37208__ = new_new_n6962__ & new_new_n32740__;
  assign new_new_n37209__ = new_new_n6961__ & new_new_n32740__;
  assign new_new_n37210__ = pi17 & ~new_new_n37209__;
  assign new_new_n37211__ = ~new_new_n37208__ & ~new_new_n37210__;
  assign new_new_n37212__ = new_new_n37207__ & ~new_new_n37211__;
  assign new_new_n37213__ = ~new_new_n37207__ & new_new_n37211__;
  assign new_new_n37214__ = ~new_new_n37212__ & ~new_new_n37213__;
  assign new_new_n37215__ = ~new_new_n37027__ & ~new_new_n37039__;
  assign new_new_n37216__ = ~new_new_n37028__ & ~new_new_n37215__;
  assign new_new_n37217__ = new_new_n37214__ & new_new_n37216__;
  assign new_new_n37218__ = ~new_new_n37214__ & ~new_new_n37216__;
  assign new_new_n37219__ = ~new_new_n37217__ & ~new_new_n37218__;
  assign new_new_n37220__ = new_new_n37073__ & ~new_new_n37219__;
  assign new_new_n37221__ = ~new_new_n37073__ & new_new_n37219__;
  assign new_new_n37222__ = ~new_new_n37220__ & ~new_new_n37221__;
  assign new_new_n37223__ = ~new_new_n36881__ & new_new_n37047__;
  assign new_new_n37224__ = new_new_n36881__ & ~new_new_n37047__;
  assign new_new_n37225__ = ~new_new_n37223__ & ~new_new_n37224__;
  assign new_new_n37226__ = new_new_n36878__ & new_new_n37225__;
  assign new_new_n37227__ = ~new_new_n37222__ & new_new_n37226__;
  assign new_new_n37228__ = ~new_new_n36882__ & new_new_n37047__;
  assign new_new_n37229__ = ~new_new_n36870__ & new_new_n36874__;
  assign new_new_n37230__ = ~new_new_n36875__ & ~new_new_n37229__;
  assign new_new_n37231__ = ~new_new_n37047__ & ~new_new_n37230__;
  assign new_new_n37232__ = new_new_n36695__ & ~new_new_n37228__;
  assign new_new_n37233__ = ~new_new_n37231__ & new_new_n37232__;
  assign new_new_n37234__ = new_new_n37222__ & ~new_new_n37233__;
  assign po20 = ~new_new_n37227__ & ~new_new_n37234__;
  assign new_new_n37236__ = ~new_new_n37206__ & ~new_new_n37211__;
  assign new_new_n37237__ = ~new_new_n37205__ & ~new_new_n37236__;
  assign new_new_n37238__ = ~new_new_n37214__ & new_new_n37216__;
  assign new_new_n37239__ = ~new_new_n37220__ & ~new_new_n37238__;
  assign new_new_n37240__ = new_new_n37237__ & ~new_new_n37239__;
  assign new_new_n37241__ = ~new_new_n37237__ & new_new_n37239__;
  assign new_new_n37242__ = ~new_new_n37240__ & ~new_new_n37241__;
  assign new_new_n37243__ = ~new_new_n37222__ & new_new_n37233__;
  assign new_new_n37244__ = ~new_new_n37197__ & ~new_new_n37201__;
  assign new_new_n37245__ = ~new_new_n37198__ & ~new_new_n37244__;
  assign new_new_n37246__ = new_new_n6634__ & new_new_n32740__;
  assign new_new_n37247__ = new_new_n6629__ & new_new_n32729__;
  assign new_new_n37248__ = ~new_new_n6625__ & new_new_n32382__;
  assign new_new_n37249__ = ~new_new_n37247__ & ~new_new_n37248__;
  assign new_new_n37250__ = ~new_new_n37246__ & new_new_n37249__;
  assign new_new_n37251__ = new_new_n6631__ & new_new_n33050__;
  assign new_new_n37252__ = ~pi20 & ~new_new_n37251__;
  assign new_new_n37253__ = new_new_n7015__ & new_new_n33050__;
  assign new_new_n37254__ = ~new_new_n37252__ & ~new_new_n37253__;
  assign new_new_n37255__ = new_new_n37250__ & ~new_new_n37254__;
  assign new_new_n37256__ = pi20 & ~new_new_n37250__;
  assign new_new_n37257__ = ~new_new_n37255__ & ~new_new_n37256__;
  assign new_new_n37258__ = ~new_new_n37190__ & ~new_new_n37193__;
  assign new_new_n37259__ = ~new_new_n37189__ & ~new_new_n37258__;
  assign new_new_n37260__ = ~new_new_n37257__ & new_new_n37259__;
  assign new_new_n37261__ = new_new_n37257__ & ~new_new_n37259__;
  assign new_new_n37262__ = ~new_new_n37260__ & ~new_new_n37261__;
  assign new_new_n37263__ = ~new_new_n333__ & new_new_n26722__;
  assign new_new_n37264__ = new_new_n873__ & ~new_new_n27242__;
  assign new_new_n37265__ = new_new_n3311__ & new_new_n27250__;
  assign new_new_n37266__ = ~new_new_n37263__ & ~new_new_n37264__;
  assign new_new_n37267__ = ~new_new_n37265__ & new_new_n37266__;
  assign new_new_n37268__ = pi26 & ~new_new_n37267__;
  assign new_new_n37269__ = new_new_n4898__ & ~new_new_n27271__;
  assign new_new_n37270__ = new_new_n801__ & ~new_new_n27271__;
  assign new_new_n37271__ = ~pi26 & ~new_new_n37270__;
  assign new_new_n37272__ = ~new_new_n37269__ & ~new_new_n37271__;
  assign new_new_n37273__ = new_new_n37267__ & ~new_new_n37272__;
  assign new_new_n37274__ = ~new_new_n37268__ & ~new_new_n37273__;
  assign new_new_n37275__ = ~new_new_n37150__ & ~new_new_n37175__;
  assign new_new_n37276__ = ~new_new_n37176__ & ~new_new_n37275__;
  assign new_new_n37277__ = ~new_new_n37274__ & new_new_n37276__;
  assign new_new_n37278__ = new_new_n37274__ & ~new_new_n37276__;
  assign new_new_n37279__ = ~new_new_n37277__ & ~new_new_n37278__;
  assign new_new_n37280__ = ~new_new_n4818__ & new_new_n26810__;
  assign new_new_n37281__ = new_new_n4212__ & new_new_n26774__;
  assign new_new_n37282__ = ~new_new_n37280__ & ~new_new_n37281__;
  assign new_new_n37283__ = new_new_n4214__ & new_new_n26729__;
  assign new_new_n37284__ = new_new_n30644__ & new_new_n37283__;
  assign new_new_n37285__ = new_new_n37282__ & ~new_new_n37284__;
  assign new_new_n37286__ = pi29 & ~new_new_n37285__;
  assign new_new_n37287__ = new_new_n4214__ & ~new_new_n33918__;
  assign new_new_n37288__ = ~pi29 & ~new_new_n37287__;
  assign new_new_n37289__ = pi28 & ~new_new_n33922__;
  assign new_new_n37290__ = ~pi28 & ~new_new_n33924__;
  assign new_new_n37291__ = new_new_n4214__ & ~new_new_n37289__;
  assign new_new_n37292__ = ~new_new_n37290__ & new_new_n37291__;
  assign new_new_n37293__ = ~new_new_n37288__ & ~new_new_n37292__;
  assign new_new_n37294__ = new_new_n37282__ & ~new_new_n37293__;
  assign new_new_n37295__ = ~new_new_n37286__ & ~new_new_n37294__;
  assign new_new_n37296__ = new_new_n71__ & new_new_n26741__;
  assign new_new_n37297__ = new_new_n161__ & ~new_new_n26741__;
  assign new_new_n37298__ = ~new_new_n161__ & ~new_new_n26802__;
  assign new_new_n37299__ = ~new_new_n37297__ & ~new_new_n37298__;
  assign new_new_n37300__ = new_new_n4876__ & ~new_new_n37299__;
  assign new_new_n37301__ = new_new_n161__ & ~new_new_n27221__;
  assign new_new_n37302__ = ~new_new_n161__ & new_new_n30411__;
  assign new_new_n37303__ = ~new_new_n71__ & ~new_new_n37301__;
  assign new_new_n37304__ = ~new_new_n37302__ & new_new_n37303__;
  assign new_new_n37305__ = pi31 & ~new_new_n37304__;
  assign new_new_n37306__ = ~new_new_n37300__ & ~new_new_n37305__;
  assign new_new_n37307__ = ~new_new_n37296__ & ~new_new_n37306__;
  assign new_new_n37308__ = new_new_n37138__ & new_new_n37147__;
  assign new_new_n37309__ = new_new_n37139__ & ~new_new_n37147__;
  assign new_new_n37310__ = ~new_new_n37308__ & ~new_new_n37309__;
  assign new_new_n37311__ = ~new_new_n952__ & new_new_n1218__;
  assign new_new_n37312__ = ~new_new_n1506__ & new_new_n1944__;
  assign new_new_n37313__ = new_new_n3168__ & new_new_n4727__;
  assign new_new_n37314__ = new_new_n37312__ & new_new_n37313__;
  assign new_new_n37315__ = new_new_n2098__ & new_new_n37311__;
  assign new_new_n37316__ = new_new_n2586__ & new_new_n3262__;
  assign new_new_n37317__ = new_new_n3280__ & new_new_n3318__;
  assign new_new_n37318__ = new_new_n37316__ & new_new_n37317__;
  assign new_new_n37319__ = new_new_n37314__ & new_new_n37315__;
  assign new_new_n37320__ = new_new_n37318__ & new_new_n37319__;
  assign new_new_n37321__ = new_new_n343__ & new_new_n3095__;
  assign new_new_n37322__ = new_new_n37320__ & new_new_n37321__;
  assign new_new_n37323__ = new_new_n3903__ & new_new_n37322__;
  assign new_new_n37324__ = new_new_n1874__ & new_new_n37323__;
  assign new_new_n37325__ = new_new_n6228__ & new_new_n37324__;
  assign new_new_n37326__ = ~new_new_n37310__ & new_new_n37325__;
  assign new_new_n37327__ = new_new_n37310__ & ~new_new_n37325__;
  assign new_new_n37328__ = ~new_new_n37326__ & ~new_new_n37327__;
  assign new_new_n37329__ = ~new_new_n37307__ & new_new_n37328__;
  assign new_new_n37330__ = new_new_n37307__ & ~new_new_n37328__;
  assign new_new_n37331__ = ~new_new_n37329__ & ~new_new_n37330__;
  assign new_new_n37332__ = new_new_n37295__ & ~new_new_n37331__;
  assign new_new_n37333__ = ~new_new_n37295__ & new_new_n37331__;
  assign new_new_n37334__ = ~new_new_n37332__ & ~new_new_n37333__;
  assign new_new_n37335__ = new_new_n37279__ & ~new_new_n37334__;
  assign new_new_n37336__ = ~new_new_n37279__ & new_new_n37334__;
  assign new_new_n37337__ = ~new_new_n37335__ & ~new_new_n37336__;
  assign new_new_n37338__ = ~new_new_n37182__ & new_new_n37185__;
  assign new_new_n37339__ = ~new_new_n37181__ & ~new_new_n37338__;
  assign new_new_n37340__ = new_new_n37337__ & ~new_new_n37339__;
  assign new_new_n37341__ = ~new_new_n37337__ & new_new_n37339__;
  assign new_new_n37342__ = new_new_n5191__ & new_new_n26698__;
  assign new_new_n37343__ = new_new_n5183__ & ~new_new_n26674__;
  assign new_new_n37344__ = ~new_new_n37342__ & ~new_new_n37343__;
  assign new_new_n37345__ = new_new_n5195__ & new_new_n35440__;
  assign new_new_n37346__ = new_new_n37344__ & ~new_new_n37345__;
  assign new_new_n37347__ = ~pi23 & ~new_new_n37346__;
  assign new_new_n37348__ = new_new_n5195__ & ~new_new_n35448__;
  assign new_new_n37349__ = pi23 & ~new_new_n37348__;
  assign new_new_n37350__ = pi22 & ~new_new_n32338__;
  assign new_new_n37351__ = ~pi22 & ~new_new_n32341__;
  assign new_new_n37352__ = new_new_n5195__ & ~new_new_n37350__;
  assign new_new_n37353__ = ~new_new_n37351__ & new_new_n37352__;
  assign new_new_n37354__ = ~new_new_n37349__ & ~new_new_n37353__;
  assign new_new_n37355__ = new_new_n37344__ & ~new_new_n37354__;
  assign new_new_n37356__ = ~new_new_n37347__ & ~new_new_n37355__;
  assign new_new_n37357__ = ~new_new_n37340__ & new_new_n37356__;
  assign new_new_n37358__ = ~new_new_n37341__ & ~new_new_n37357__;
  assign new_new_n37359__ = ~new_new_n37340__ & new_new_n37358__;
  assign new_new_n37360__ = ~new_new_n37341__ & new_new_n37357__;
  assign new_new_n37361__ = new_new_n37356__ & ~new_new_n37360__;
  assign new_new_n37362__ = ~new_new_n37359__ & ~new_new_n37361__;
  assign new_new_n37363__ = new_new_n37262__ & ~new_new_n37362__;
  assign new_new_n37364__ = ~new_new_n37262__ & new_new_n37362__;
  assign new_new_n37365__ = ~new_new_n37363__ & ~new_new_n37364__;
  assign new_new_n37366__ = ~new_new_n37245__ & new_new_n37365__;
  assign new_new_n37367__ = new_new_n37245__ & ~new_new_n37365__;
  assign new_new_n37368__ = ~new_new_n37366__ & ~new_new_n37367__;
  assign new_new_n37369__ = ~pi17 & ~new_new_n37368__;
  assign new_new_n37370__ = pi17 & new_new_n37368__;
  assign new_new_n37371__ = ~new_new_n37369__ & ~new_new_n37370__;
  assign new_new_n37372__ = new_new_n37243__ & new_new_n37371__;
  assign new_new_n37373__ = ~new_new_n37243__ & ~new_new_n37371__;
  assign new_new_n37374__ = ~new_new_n37372__ & ~new_new_n37373__;
  assign new_new_n37375__ = new_new_n37242__ & new_new_n37374__;
  assign new_new_n37376__ = ~new_new_n37242__ & ~new_new_n37374__;
  assign po21 = ~new_new_n37375__ & ~new_new_n37376__;
  assign new_new_n37378__ = pi17 & ~new_new_n37366__;
  assign new_new_n37379__ = ~new_new_n37367__ & ~new_new_n37378__;
  assign new_new_n37380__ = ~new_new_n9921__ & ~new_new_n32729__;
  assign new_new_n37381__ = pi19 & ~new_new_n34178__;
  assign new_new_n37382__ = ~new_new_n6619__ & ~new_new_n6632__;
  assign new_new_n37383__ = ~new_new_n37381__ & new_new_n37382__;
  assign new_new_n37384__ = ~pi19 & ~new_new_n34178__;
  assign new_new_n37385__ = ~new_new_n6620__ & ~new_new_n6622__;
  assign new_new_n37386__ = ~new_new_n37384__ & new_new_n37385__;
  assign new_new_n37387__ = ~new_new_n37247__ & ~new_new_n37380__;
  assign new_new_n37388__ = ~new_new_n37383__ & new_new_n37387__;
  assign new_new_n37389__ = ~new_new_n37386__ & new_new_n37388__;
  assign new_new_n37390__ = ~pi20 & new_new_n37389__;
  assign new_new_n37391__ = pi20 & ~new_new_n37389__;
  assign new_new_n37392__ = ~new_new_n37390__ & ~new_new_n37391__;
  assign new_new_n37393__ = ~new_new_n37260__ & new_new_n37362__;
  assign new_new_n37394__ = ~new_new_n37261__ & ~new_new_n37393__;
  assign new_new_n37395__ = new_new_n5215__ & ~new_new_n33347__;
  assign new_new_n37396__ = new_new_n5191__ & ~new_new_n26674__;
  assign new_new_n37397__ = new_new_n5183__ & ~new_new_n26667__;
  assign new_new_n37398__ = new_new_n5213__ & new_new_n32382__;
  assign new_new_n37399__ = ~new_new_n37396__ & ~new_new_n37397__;
  assign new_new_n37400__ = ~new_new_n37398__ & new_new_n37399__;
  assign new_new_n37401__ = ~new_new_n37395__ & new_new_n37400__;
  assign new_new_n37402__ = ~new_new_n333__ & ~new_new_n27242__;
  assign new_new_n37403__ = new_new_n873__ & new_new_n27250__;
  assign new_new_n37404__ = ~new_new_n37402__ & ~new_new_n37403__;
  assign new_new_n37405__ = ~new_new_n110__ & new_new_n26698__;
  assign new_new_n37406__ = new_new_n31511__ & new_new_n37405__;
  assign new_new_n37407__ = new_new_n37404__ & ~new_new_n37406__;
  assign new_new_n37408__ = pi26 & ~new_new_n37407__;
  assign new_new_n37409__ = new_new_n801__ & ~new_new_n31510__;
  assign new_new_n37410__ = ~pi26 & ~new_new_n37409__;
  assign new_new_n37411__ = ~pi25 & ~new_new_n34204__;
  assign new_new_n37412__ = pi25 & ~new_new_n31509__;
  assign new_new_n37413__ = ~new_new_n110__ & ~new_new_n37411__;
  assign new_new_n37414__ = ~new_new_n37412__ & new_new_n37413__;
  assign new_new_n37415__ = ~new_new_n37410__ & ~new_new_n37414__;
  assign new_new_n37416__ = new_new_n37404__ & ~new_new_n37415__;
  assign new_new_n37417__ = ~new_new_n37408__ & ~new_new_n37416__;
  assign new_new_n37418__ = ~new_new_n37278__ & new_new_n37334__;
  assign new_new_n37419__ = ~new_new_n37277__ & ~new_new_n37418__;
  assign new_new_n37420__ = ~new_new_n37417__ & ~new_new_n37419__;
  assign new_new_n37421__ = new_new_n37417__ & new_new_n37419__;
  assign new_new_n37422__ = ~new_new_n37420__ & ~new_new_n37421__;
  assign new_new_n37423__ = new_new_n4815__ & new_new_n26722__;
  assign new_new_n37424__ = ~new_new_n4818__ & new_new_n26774__;
  assign new_new_n37425__ = new_new_n4212__ & new_new_n26729__;
  assign new_new_n37426__ = ~new_new_n37424__ & ~new_new_n37425__;
  assign new_new_n37427__ = ~new_new_n37423__ & new_new_n37426__;
  assign new_new_n37428__ = new_new_n4214__ & ~new_new_n27348__;
  assign new_new_n37429__ = ~pi29 & ~new_new_n37428__;
  assign new_new_n37430__ = new_new_n5732__ & ~new_new_n27348__;
  assign new_new_n37431__ = ~new_new_n37429__ & ~new_new_n37430__;
  assign new_new_n37432__ = new_new_n37427__ & ~new_new_n37431__;
  assign new_new_n37433__ = pi29 & ~new_new_n37427__;
  assign new_new_n37434__ = ~new_new_n37432__ & ~new_new_n37433__;
  assign new_new_n37435__ = ~new_new_n37309__ & ~new_new_n37325__;
  assign new_new_n37436__ = ~new_new_n37308__ & ~new_new_n37435__;
  assign new_new_n37437__ = new_new_n5021__ & new_new_n26810__;
  assign new_new_n37438__ = new_new_n765__ & new_new_n27395__;
  assign new_new_n37439__ = ~new_new_n37297__ & ~new_new_n37438__;
  assign new_new_n37440__ = pi31 & ~new_new_n37439__;
  assign new_new_n37441__ = new_new_n5053__ & ~new_new_n26802__;
  assign new_new_n37442__ = ~new_new_n37437__ & ~new_new_n37441__;
  assign new_new_n37443__ = ~new_new_n37440__ & new_new_n37442__;
  assign new_new_n37444__ = ~new_new_n37436__ & new_new_n37443__;
  assign new_new_n37445__ = new_new_n37436__ & ~new_new_n37443__;
  assign new_new_n37446__ = ~new_new_n37444__ & ~new_new_n37445__;
  assign new_new_n37447__ = ~new_new_n308__ & ~new_new_n947__;
  assign new_new_n37448__ = ~new_new_n1007__ & new_new_n37447__;
  assign new_new_n37449__ = ~new_new_n317__ & ~new_new_n380__;
  assign new_new_n37450__ = new_new_n966__ & new_new_n1663__;
  assign new_new_n37451__ = new_new_n5430__ & new_new_n37450__;
  assign new_new_n37452__ = new_new_n37448__ & new_new_n37449__;
  assign new_new_n37453__ = new_new_n1294__ & new_new_n1993__;
  assign new_new_n37454__ = new_new_n2290__ & new_new_n37453__;
  assign new_new_n37455__ = new_new_n37451__ & new_new_n37452__;
  assign new_new_n37456__ = new_new_n347__ & ~new_new_n1539__;
  assign new_new_n37457__ = new_new_n37455__ & new_new_n37456__;
  assign new_new_n37458__ = new_new_n1717__ & new_new_n37454__;
  assign new_new_n37459__ = new_new_n16152__ & new_new_n37458__;
  assign new_new_n37460__ = new_new_n37457__ & new_new_n37459__;
  assign new_new_n37461__ = new_new_n1237__ & new_new_n37460__;
  assign new_new_n37462__ = new_new_n4978__ & new_new_n5584__;
  assign new_new_n37463__ = new_new_n37461__ & new_new_n37462__;
  assign new_new_n37464__ = new_new_n37325__ & new_new_n37463__;
  assign new_new_n37465__ = ~new_new_n37325__ & ~new_new_n37463__;
  assign new_new_n37466__ = ~pi17 & ~new_new_n37464__;
  assign new_new_n37467__ = ~new_new_n37465__ & ~new_new_n37466__;
  assign new_new_n37468__ = ~new_new_n37464__ & new_new_n37467__;
  assign new_new_n37469__ = pi17 & ~new_new_n37468__;
  assign new_new_n37470__ = ~new_new_n37465__ & new_new_n37466__;
  assign new_new_n37471__ = ~new_new_n37469__ & ~new_new_n37470__;
  assign new_new_n37472__ = new_new_n37446__ & ~new_new_n37471__;
  assign new_new_n37473__ = ~new_new_n37446__ & new_new_n37471__;
  assign new_new_n37474__ = ~new_new_n37472__ & ~new_new_n37473__;
  assign new_new_n37475__ = ~new_new_n37434__ & new_new_n37474__;
  assign new_new_n37476__ = new_new_n37434__ & ~new_new_n37474__;
  assign new_new_n37477__ = ~new_new_n37475__ & ~new_new_n37476__;
  assign new_new_n37478__ = new_new_n37295__ & ~new_new_n37329__;
  assign new_new_n37479__ = ~new_new_n37330__ & ~new_new_n37478__;
  assign new_new_n37480__ = new_new_n37477__ & new_new_n37479__;
  assign new_new_n37481__ = ~new_new_n37477__ & ~new_new_n37479__;
  assign new_new_n37482__ = ~new_new_n37480__ & ~new_new_n37481__;
  assign new_new_n37483__ = new_new_n37422__ & ~new_new_n37482__;
  assign new_new_n37484__ = ~new_new_n37422__ & new_new_n37482__;
  assign new_new_n37485__ = ~new_new_n37483__ & ~new_new_n37484__;
  assign new_new_n37486__ = new_new_n37358__ & new_new_n37485__;
  assign new_new_n37487__ = ~new_new_n37358__ & ~new_new_n37485__;
  assign new_new_n37488__ = ~new_new_n37486__ & ~new_new_n37487__;
  assign new_new_n37489__ = pi23 & ~new_new_n37488__;
  assign new_new_n37490__ = ~pi23 & new_new_n37488__;
  assign new_new_n37491__ = ~new_new_n37489__ & ~new_new_n37490__;
  assign new_new_n37492__ = new_new_n37401__ & new_new_n37491__;
  assign new_new_n37493__ = ~new_new_n37401__ & ~new_new_n37491__;
  assign new_new_n37494__ = ~new_new_n37492__ & ~new_new_n37493__;
  assign new_new_n37495__ = new_new_n37394__ & ~new_new_n37494__;
  assign new_new_n37496__ = ~new_new_n37394__ & new_new_n37494__;
  assign new_new_n37497__ = ~new_new_n37495__ & ~new_new_n37496__;
  assign new_new_n37498__ = new_new_n37392__ & new_new_n37497__;
  assign new_new_n37499__ = ~new_new_n37392__ & ~new_new_n37497__;
  assign new_new_n37500__ = ~new_new_n37498__ & ~new_new_n37499__;
  assign new_new_n37501__ = ~new_new_n37379__ & ~new_new_n37500__;
  assign new_new_n37502__ = ~new_new_n37367__ & new_new_n37500__;
  assign new_new_n37503__ = ~new_new_n37378__ & new_new_n37502__;
  assign new_new_n37504__ = ~new_new_n37501__ & ~new_new_n37503__;
  assign new_new_n37505__ = new_new_n37240__ & ~new_new_n37372__;
  assign new_new_n37506__ = ~new_new_n37241__ & new_new_n37373__;
  assign new_new_n37507__ = new_new_n37241__ & new_new_n37372__;
  assign new_new_n37508__ = ~new_new_n37505__ & ~new_new_n37506__;
  assign new_new_n37509__ = ~new_new_n37507__ & new_new_n37508__;
  assign new_new_n37510__ = new_new_n37504__ & ~new_new_n37509__;
  assign new_new_n37511__ = ~new_new_n37239__ & po21;
  assign new_new_n37512__ = new_new_n37243__ & ~new_new_n37511__;
  assign new_new_n37513__ = ~new_new_n37237__ & new_new_n37371__;
  assign new_new_n37514__ = new_new_n37239__ & ~po21;
  assign new_new_n37515__ = ~new_new_n37513__ & ~new_new_n37514__;
  assign new_new_n37516__ = ~new_new_n37512__ & new_new_n37515__;
  assign new_new_n37517__ = ~new_new_n37504__ & ~new_new_n37507__;
  assign new_new_n37518__ = ~new_new_n37516__ & new_new_n37517__;
  assign po22 = new_new_n37510__ | new_new_n37518__;
  assign new_new_n37520__ = ~new_new_n37392__ & ~new_new_n37495__;
  assign new_new_n37521__ = ~new_new_n37496__ & ~new_new_n37520__;
  assign new_new_n37522__ = ~new_new_n6625__ & new_new_n32740__;
  assign new_new_n37523__ = pi20 & ~new_new_n37522__;
  assign new_new_n37524__ = ~pi20 & new_new_n37522__;
  assign new_new_n37525__ = ~new_new_n37523__ & ~new_new_n37524__;
  assign new_new_n37526__ = ~new_new_n37486__ & new_new_n37494__;
  assign new_new_n37527__ = ~new_new_n37487__ & ~new_new_n37526__;
  assign new_new_n37528__ = new_new_n5191__ & ~new_new_n26667__;
  assign new_new_n37529__ = new_new_n5183__ & new_new_n32382__;
  assign new_new_n37530__ = ~new_new_n37528__ & ~new_new_n37529__;
  assign new_new_n37531__ = new_new_n5195__ & new_new_n32729__;
  assign new_new_n37532__ = new_new_n32758__ & new_new_n37531__;
  assign new_new_n37533__ = new_new_n37530__ & ~new_new_n37532__;
  assign new_new_n37534__ = pi23 & ~new_new_n37533__;
  assign new_new_n37535__ = new_new_n5195__ & ~new_new_n33614__;
  assign new_new_n37536__ = ~pi23 & ~new_new_n37535__;
  assign new_new_n37537__ = ~pi22 & ~new_new_n33617__;
  assign new_new_n37538__ = pi22 & ~new_new_n33619__;
  assign new_new_n37539__ = new_new_n5195__ & ~new_new_n37537__;
  assign new_new_n37540__ = ~new_new_n37538__ & new_new_n37539__;
  assign new_new_n37541__ = ~new_new_n37536__ & ~new_new_n37540__;
  assign new_new_n37542__ = new_new_n37530__ & ~new_new_n37541__;
  assign new_new_n37543__ = ~new_new_n37534__ & ~new_new_n37542__;
  assign new_new_n37544__ = new_new_n873__ & new_new_n26698__;
  assign new_new_n37545__ = ~new_new_n333__ & new_new_n27250__;
  assign new_new_n37546__ = new_new_n3311__ & ~new_new_n26674__;
  assign new_new_n37547__ = ~new_new_n37544__ & ~new_new_n37545__;
  assign new_new_n37548__ = ~new_new_n37546__ & new_new_n37547__;
  assign new_new_n37549__ = ~pi26 & ~new_new_n37548__;
  assign new_new_n37550__ = new_new_n512__ & new_new_n27284__;
  assign new_new_n37551__ = new_new_n801__ & new_new_n27284__;
  assign new_new_n37552__ = pi26 & ~new_new_n37551__;
  assign new_new_n37553__ = ~new_new_n37550__ & ~new_new_n37552__;
  assign new_new_n37554__ = new_new_n37548__ & ~new_new_n37553__;
  assign new_new_n37555__ = ~new_new_n37549__ & ~new_new_n37554__;
  assign new_new_n37556__ = ~new_new_n4818__ & new_new_n26729__;
  assign new_new_n37557__ = new_new_n4212__ & new_new_n26722__;
  assign new_new_n37558__ = ~new_new_n37556__ & ~new_new_n37557__;
  assign new_new_n37559__ = new_new_n4214__ & ~new_new_n27362__;
  assign new_new_n37560__ = pi29 & ~new_new_n37559__;
  assign new_new_n37561__ = ~pi28 & new_new_n27242__;
  assign new_new_n37562__ = pi28 & ~new_new_n27242__;
  assign new_new_n37563__ = new_new_n4214__ & ~new_new_n37561__;
  assign new_new_n37564__ = ~new_new_n37562__ & new_new_n37563__;
  assign new_new_n37565__ = new_new_n27352__ & new_new_n37564__;
  assign new_new_n37566__ = ~new_new_n37560__ & ~new_new_n37565__;
  assign new_new_n37567__ = new_new_n37558__ & ~new_new_n37566__;
  assign new_new_n37568__ = new_new_n4214__ & new_new_n27353__;
  assign new_new_n37569__ = new_new_n37558__ & ~new_new_n37568__;
  assign new_new_n37570__ = ~pi29 & ~new_new_n37569__;
  assign new_new_n37571__ = ~new_new_n37567__ & ~new_new_n37570__;
  assign new_new_n37572__ = new_new_n37555__ & ~new_new_n37571__;
  assign new_new_n37573__ = ~new_new_n37555__ & new_new_n37571__;
  assign new_new_n37574__ = ~new_new_n37572__ & ~new_new_n37573__;
  assign new_new_n37575__ = ~new_new_n92__ & ~new_new_n717__;
  assign new_new_n37576__ = ~new_new_n1031__ & new_new_n37575__;
  assign new_new_n37577__ = ~new_new_n322__ & ~new_new_n334__;
  assign new_new_n37578__ = new_new_n1154__ & new_new_n1213__;
  assign new_new_n37579__ = new_new_n2589__ & new_new_n37578__;
  assign new_new_n37580__ = new_new_n37576__ & new_new_n37577__;
  assign new_new_n37581__ = new_new_n3101__ & new_new_n3368__;
  assign new_new_n37582__ = new_new_n5566__ & new_new_n37581__;
  assign new_new_n37583__ = new_new_n37579__ & new_new_n37580__;
  assign new_new_n37584__ = new_new_n37582__ & new_new_n37583__;
  assign new_new_n37585__ = new_new_n16266__ & new_new_n37584__;
  assign new_new_n37586__ = new_new_n1104__ & new_new_n3137__;
  assign new_new_n37587__ = new_new_n37585__ & new_new_n37586__;
  assign new_new_n37588__ = new_new_n7743__ & new_new_n37587__;
  assign new_new_n37589__ = new_new_n35519__ & new_new_n37588__;
  assign new_new_n37590__ = new_new_n37467__ & ~new_new_n37589__;
  assign new_new_n37591__ = ~new_new_n37467__ & new_new_n37589__;
  assign new_new_n37592__ = ~new_new_n37590__ & ~new_new_n37591__;
  assign new_new_n37593__ = new_new_n161__ & new_new_n26810__;
  assign new_new_n37594__ = new_new_n765__ & new_new_n26774__;
  assign new_new_n37595__ = ~new_new_n37593__ & ~new_new_n37594__;
  assign new_new_n37596__ = ~pi31 & ~new_new_n37595__;
  assign new_new_n37597__ = ~new_new_n71__ & new_new_n31581__;
  assign new_new_n37598__ = new_new_n26810__ & new_new_n37597__;
  assign new_new_n37599__ = ~new_new_n26810__ & ~new_new_n37597__;
  assign new_new_n37600__ = ~new_new_n37598__ & ~new_new_n37599__;
  assign new_new_n37601__ = ~new_new_n161__ & ~new_new_n37600__;
  assign new_new_n37602__ = new_new_n161__ & new_new_n26802__;
  assign new_new_n37603__ = pi31 & ~new_new_n37602__;
  assign new_new_n37604__ = ~new_new_n37601__ & new_new_n37603__;
  assign new_new_n37605__ = ~new_new_n37596__ & ~new_new_n37604__;
  assign new_new_n37606__ = ~new_new_n37445__ & ~new_new_n37471__;
  assign new_new_n37607__ = ~new_new_n37444__ & ~new_new_n37606__;
  assign new_new_n37608__ = new_new_n37605__ & ~new_new_n37607__;
  assign new_new_n37609__ = ~new_new_n37605__ & new_new_n37607__;
  assign new_new_n37610__ = ~new_new_n37608__ & ~new_new_n37609__;
  assign new_new_n37611__ = new_new_n37592__ & new_new_n37610__;
  assign new_new_n37612__ = ~new_new_n37592__ & ~new_new_n37610__;
  assign new_new_n37613__ = ~new_new_n37611__ & ~new_new_n37612__;
  assign new_new_n37614__ = ~new_new_n37475__ & ~new_new_n37479__;
  assign new_new_n37615__ = ~new_new_n37476__ & ~new_new_n37614__;
  assign new_new_n37616__ = new_new_n37613__ & ~new_new_n37615__;
  assign new_new_n37617__ = ~new_new_n37613__ & new_new_n37615__;
  assign new_new_n37618__ = ~new_new_n37616__ & ~new_new_n37617__;
  assign new_new_n37619__ = new_new_n37574__ & new_new_n37618__;
  assign new_new_n37620__ = ~new_new_n37574__ & ~new_new_n37618__;
  assign new_new_n37621__ = ~new_new_n37619__ & ~new_new_n37620__;
  assign new_new_n37622__ = new_new_n37543__ & ~new_new_n37621__;
  assign new_new_n37623__ = ~new_new_n37543__ & new_new_n37621__;
  assign new_new_n37624__ = ~new_new_n37622__ & ~new_new_n37623__;
  assign new_new_n37625__ = ~new_new_n37420__ & ~new_new_n37482__;
  assign new_new_n37626__ = ~new_new_n37421__ & ~new_new_n37625__;
  assign new_new_n37627__ = new_new_n37624__ & ~new_new_n37626__;
  assign new_new_n37628__ = ~new_new_n37624__ & new_new_n37626__;
  assign new_new_n37629__ = ~new_new_n37627__ & ~new_new_n37628__;
  assign new_new_n37630__ = new_new_n37527__ & new_new_n37629__;
  assign new_new_n37631__ = ~new_new_n37527__ & ~new_new_n37629__;
  assign new_new_n37632__ = ~new_new_n37630__ & ~new_new_n37631__;
  assign new_new_n37633__ = new_new_n32382__ & new_new_n37522__;
  assign new_new_n37634__ = new_new_n37632__ & ~new_new_n37633__;
  assign new_new_n37635__ = new_new_n37525__ & ~new_new_n37634__;
  assign new_new_n37636__ = ~new_new_n37525__ & new_new_n37632__;
  assign new_new_n37637__ = ~new_new_n37635__ & ~new_new_n37636__;
  assign new_new_n37638__ = new_new_n37521__ & ~new_new_n37637__;
  assign new_new_n37639__ = ~new_new_n37521__ & new_new_n37637__;
  assign new_new_n37640__ = ~new_new_n37638__ & ~new_new_n37639__;
  assign new_new_n37641__ = new_new_n37239__ & new_new_n37371__;
  assign new_new_n37642__ = new_new_n37243__ & new_new_n37504__;
  assign new_new_n37643__ = ~new_new_n37641__ & new_new_n37642__;
  assign new_new_n37644__ = ~new_new_n37504__ & new_new_n37513__;
  assign new_new_n37645__ = new_new_n37239__ & new_new_n37644__;
  assign new_new_n37646__ = ~new_new_n37643__ & ~new_new_n37645__;
  assign new_new_n37647__ = ~po21 & ~new_new_n37646__;
  assign new_new_n37648__ = new_new_n37240__ & ~new_new_n37501__;
  assign new_new_n37649__ = pi17 & ~new_new_n37502__;
  assign new_new_n37650__ = ~new_new_n37366__ & ~new_new_n37500__;
  assign new_new_n37651__ = ~new_new_n37649__ & ~new_new_n37650__;
  assign new_new_n37652__ = ~new_new_n37241__ & new_new_n37651__;
  assign new_new_n37653__ = ~new_new_n37503__ & ~new_new_n37648__;
  assign new_new_n37654__ = ~new_new_n37652__ & new_new_n37653__;
  assign new_new_n37655__ = new_new_n37647__ & new_new_n37654__;
  assign new_new_n37656__ = ~new_new_n37647__ & ~new_new_n37654__;
  assign new_new_n37657__ = ~new_new_n37655__ & ~new_new_n37656__;
  assign new_new_n37658__ = new_new_n37640__ & new_new_n37657__;
  assign new_new_n37659__ = ~new_new_n37640__ & ~new_new_n37657__;
  assign po23 = ~new_new_n37658__ & ~new_new_n37659__;
  assign new_new_n37661__ = new_new_n37639__ & ~new_new_n37647__;
  assign new_new_n37662__ = ~new_new_n37638__ & new_new_n37657__;
  assign new_new_n37663__ = ~new_new_n37639__ & new_new_n37655__;
  assign new_new_n37664__ = new_new_n37525__ & ~new_new_n37630__;
  assign new_new_n37665__ = ~new_new_n37631__ & ~new_new_n37664__;
  assign new_new_n37666__ = new_new_n5213__ & new_new_n32740__;
  assign new_new_n37667__ = new_new_n5183__ & new_new_n32729__;
  assign new_new_n37668__ = new_new_n5191__ & new_new_n32382__;
  assign new_new_n37669__ = ~new_new_n37667__ & ~new_new_n37668__;
  assign new_new_n37670__ = ~new_new_n37666__ & new_new_n37669__;
  assign new_new_n37671__ = new_new_n5195__ & new_new_n33050__;
  assign new_new_n37672__ = ~pi23 & ~new_new_n37671__;
  assign new_new_n37673__ = new_new_n5974__ & new_new_n33050__;
  assign new_new_n37674__ = ~new_new_n37672__ & ~new_new_n37673__;
  assign new_new_n37675__ = new_new_n37670__ & ~new_new_n37674__;
  assign new_new_n37676__ = pi23 & ~new_new_n37670__;
  assign new_new_n37677__ = ~new_new_n37675__ & ~new_new_n37676__;
  assign new_new_n37678__ = ~new_new_n37555__ & ~new_new_n37615__;
  assign new_new_n37679__ = new_new_n37555__ & new_new_n37615__;
  assign new_new_n37680__ = new_new_n37571__ & ~new_new_n37613__;
  assign new_new_n37681__ = ~new_new_n37571__ & new_new_n37613__;
  assign new_new_n37682__ = ~new_new_n37680__ & ~new_new_n37681__;
  assign new_new_n37683__ = ~new_new_n37679__ & new_new_n37682__;
  assign new_new_n37684__ = ~new_new_n37678__ & ~new_new_n37683__;
  assign new_new_n37685__ = new_new_n37677__ & ~new_new_n37684__;
  assign new_new_n37686__ = ~new_new_n37677__ & new_new_n37684__;
  assign new_new_n37687__ = ~new_new_n37685__ & ~new_new_n37686__;
  assign new_new_n37688__ = ~new_new_n37622__ & new_new_n37626__;
  assign new_new_n37689__ = ~new_new_n37623__ & ~new_new_n37688__;
  assign new_new_n37690__ = new_new_n37687__ & ~new_new_n37689__;
  assign new_new_n37691__ = ~new_new_n37687__ & new_new_n37689__;
  assign new_new_n37692__ = ~new_new_n37690__ & ~new_new_n37691__;
  assign new_new_n37693__ = ~new_new_n37571__ & new_new_n37607__;
  assign new_new_n37694__ = ~new_new_n37591__ & new_new_n37605__;
  assign new_new_n37695__ = ~new_new_n37590__ & ~new_new_n37694__;
  assign new_new_n37696__ = new_new_n37693__ & ~new_new_n37695__;
  assign new_new_n37697__ = new_new_n37590__ & new_new_n37605__;
  assign new_new_n37698__ = new_new_n37571__ & ~new_new_n37607__;
  assign new_new_n37699__ = new_new_n37591__ & ~new_new_n37605__;
  assign new_new_n37700__ = ~new_new_n37697__ & ~new_new_n37699__;
  assign new_new_n37701__ = ~new_new_n37693__ & new_new_n37700__;
  assign new_new_n37702__ = ~new_new_n37698__ & new_new_n37701__;
  assign new_new_n37703__ = new_new_n37695__ & new_new_n37698__;
  assign new_new_n37704__ = ~new_new_n160__ & ~new_new_n253__;
  assign new_new_n37705__ = ~new_new_n785__ & ~new_new_n1031__;
  assign new_new_n37706__ = new_new_n37704__ & new_new_n37705__;
  assign new_new_n37707__ = ~new_new_n591__ & ~new_new_n673__;
  assign new_new_n37708__ = new_new_n1702__ & new_new_n19504__;
  assign new_new_n37709__ = new_new_n37707__ & new_new_n37708__;
  assign new_new_n37710__ = new_new_n836__ & new_new_n37706__;
  assign new_new_n37711__ = new_new_n16471__ & new_new_n37710__;
  assign new_new_n37712__ = new_new_n2705__ & new_new_n37709__;
  assign new_new_n37713__ = new_new_n37711__ & new_new_n37712__;
  assign new_new_n37714__ = new_new_n18159__ & new_new_n34583__;
  assign new_new_n37715__ = new_new_n37713__ & new_new_n37714__;
  assign new_new_n37716__ = new_new_n4955__ & new_new_n5310__;
  assign new_new_n37717__ = new_new_n37715__ & new_new_n37716__;
  assign new_new_n37718__ = new_new_n7415__ & new_new_n37717__;
  assign new_new_n37719__ = new_new_n1249__ & new_new_n37718__;
  assign new_new_n37720__ = new_new_n71__ & new_new_n26774__;
  assign new_new_n37721__ = ~new_new_n37593__ & ~new_new_n37720__;
  assign new_new_n37722__ = pi31 & ~new_new_n37721__;
  assign new_new_n37723__ = new_new_n161__ & ~new_new_n26774__;
  assign new_new_n37724__ = ~new_new_n161__ & ~new_new_n26729__;
  assign new_new_n37725__ = new_new_n4876__ & ~new_new_n37723__;
  assign new_new_n37726__ = ~new_new_n37724__ & new_new_n37725__;
  assign new_new_n37727__ = ~new_new_n161__ & new_new_n4147__;
  assign new_new_n37728__ = new_new_n30644__ & new_new_n37727__;
  assign new_new_n37729__ = ~new_new_n37722__ & ~new_new_n37726__;
  assign new_new_n37730__ = ~new_new_n37728__ & new_new_n37729__;
  assign new_new_n37731__ = ~new_new_n37719__ & ~new_new_n37730__;
  assign new_new_n37732__ = new_new_n37719__ & new_new_n37730__;
  assign new_new_n37733__ = ~new_new_n37731__ & ~new_new_n37732__;
  assign new_new_n37734__ = new_new_n37589__ & ~new_new_n37733__;
  assign new_new_n37735__ = ~new_new_n37589__ & new_new_n37733__;
  assign new_new_n37736__ = ~new_new_n37734__ & ~new_new_n37735__;
  assign new_new_n37737__ = ~new_new_n37696__ & new_new_n37736__;
  assign new_new_n37738__ = ~new_new_n37703__ & new_new_n37737__;
  assign new_new_n37739__ = ~new_new_n37702__ & new_new_n37738__;
  assign new_new_n37740__ = new_new_n37571__ & new_new_n37608__;
  assign new_new_n37741__ = new_new_n37467__ & new_new_n37740__;
  assign new_new_n37742__ = ~new_new_n37571__ & ~new_new_n37608__;
  assign new_new_n37743__ = ~new_new_n37609__ & ~new_new_n37742__;
  assign new_new_n37744__ = new_new_n37467__ & new_new_n37743__;
  assign new_new_n37745__ = ~new_new_n37740__ & ~new_new_n37744__;
  assign new_new_n37746__ = ~new_new_n37589__ & ~new_new_n37745__;
  assign new_new_n37747__ = ~new_new_n37571__ & new_new_n37609__;
  assign new_new_n37748__ = new_new_n37467__ & ~new_new_n37747__;
  assign new_new_n37749__ = new_new_n37589__ & ~new_new_n37743__;
  assign new_new_n37750__ = ~new_new_n37748__ & new_new_n37749__;
  assign new_new_n37751__ = ~new_new_n37467__ & ~new_new_n37571__;
  assign new_new_n37752__ = new_new_n37609__ & new_new_n37751__;
  assign new_new_n37753__ = ~new_new_n37736__ & ~new_new_n37741__;
  assign new_new_n37754__ = ~new_new_n37752__ & new_new_n37753__;
  assign new_new_n37755__ = ~new_new_n37750__ & new_new_n37754__;
  assign new_new_n37756__ = ~new_new_n37746__ & new_new_n37755__;
  assign new_new_n37757__ = ~new_new_n37739__ & ~new_new_n37756__;
  assign new_new_n37758__ = ~pi20 & ~new_new_n37757__;
  assign new_new_n37759__ = pi20 & new_new_n37757__;
  assign new_new_n37760__ = ~new_new_n37758__ & ~new_new_n37759__;
  assign new_new_n37761__ = ~new_new_n4818__ & new_new_n26722__;
  assign new_new_n37762__ = new_new_n4212__ & ~new_new_n27242__;
  assign new_new_n37763__ = new_new_n4813__ & ~new_new_n27271__;
  assign new_new_n37764__ = ~new_new_n37761__ & ~new_new_n37762__;
  assign new_new_n37765__ = ~new_new_n37763__ & new_new_n37764__;
  assign new_new_n37766__ = new_new_n4214__ & new_new_n27250__;
  assign new_new_n37767__ = ~new_new_n4900__ & ~new_new_n32340__;
  assign new_new_n37768__ = ~new_new_n333__ & new_new_n26698__;
  assign new_new_n37769__ = new_new_n873__ & ~new_new_n26674__;
  assign new_new_n37770__ = ~new_new_n37768__ & ~new_new_n37769__;
  assign new_new_n37771__ = ~new_new_n37767__ & new_new_n37770__;
  assign new_new_n37772__ = pi26 & ~new_new_n37771__;
  assign new_new_n37773__ = new_new_n512__ & ~new_new_n26667__;
  assign new_new_n37774__ = new_new_n801__ & ~new_new_n26667__;
  assign new_new_n37775__ = ~pi26 & ~new_new_n37774__;
  assign new_new_n37776__ = ~new_new_n37773__ & ~new_new_n37775__;
  assign new_new_n37777__ = new_new_n37771__ & ~new_new_n37776__;
  assign new_new_n37778__ = ~new_new_n37772__ & ~new_new_n37777__;
  assign new_new_n37779__ = ~pi28 & ~new_new_n37778__;
  assign new_new_n37780__ = pi28 & new_new_n37778__;
  assign new_new_n37781__ = ~new_new_n37779__ & ~new_new_n37780__;
  assign new_new_n37782__ = new_new_n37766__ & ~new_new_n37781__;
  assign new_new_n37783__ = pi29 & ~new_new_n37778__;
  assign new_new_n37784__ = ~pi29 & new_new_n37778__;
  assign new_new_n37785__ = ~new_new_n37783__ & ~new_new_n37784__;
  assign new_new_n37786__ = ~new_new_n37766__ & ~new_new_n37785__;
  assign new_new_n37787__ = ~new_new_n37782__ & ~new_new_n37786__;
  assign new_new_n37788__ = new_new_n37765__ & ~new_new_n37787__;
  assign new_new_n37789__ = ~new_new_n37765__ & new_new_n37785__;
  assign new_new_n37790__ = ~new_new_n37788__ & ~new_new_n37789__;
  assign new_new_n37791__ = new_new_n37760__ & ~new_new_n37790__;
  assign new_new_n37792__ = ~new_new_n37760__ & new_new_n37790__;
  assign new_new_n37793__ = ~new_new_n37791__ & ~new_new_n37792__;
  assign new_new_n37794__ = new_new_n37692__ & new_new_n37793__;
  assign new_new_n37795__ = ~new_new_n37692__ & ~new_new_n37793__;
  assign new_new_n37796__ = ~new_new_n37794__ & ~new_new_n37795__;
  assign new_new_n37797__ = new_new_n37665__ & ~new_new_n37796__;
  assign new_new_n37798__ = ~new_new_n37665__ & new_new_n37796__;
  assign new_new_n37799__ = ~new_new_n37797__ & ~new_new_n37798__;
  assign new_new_n37800__ = ~new_new_n37661__ & ~new_new_n37799__;
  assign new_new_n37801__ = ~new_new_n37663__ & new_new_n37800__;
  assign new_new_n37802__ = ~new_new_n37662__ & new_new_n37801__;
  assign new_new_n37803__ = ~new_new_n37637__ & new_new_n37656__;
  assign new_new_n37804__ = new_new_n37637__ & ~new_new_n37656__;
  assign new_new_n37805__ = new_new_n37521__ & ~new_new_n37655__;
  assign new_new_n37806__ = ~new_new_n37804__ & new_new_n37805__;
  assign new_new_n37807__ = new_new_n37639__ & new_new_n37655__;
  assign new_new_n37808__ = new_new_n37799__ & ~new_new_n37803__;
  assign new_new_n37809__ = ~new_new_n37807__ & new_new_n37808__;
  assign new_new_n37810__ = ~new_new_n37806__ & new_new_n37809__;
  assign po24 = ~new_new_n37802__ & ~new_new_n37810__;
  assign new_new_n37812__ = new_new_n37637__ & new_new_n37654__;
  assign new_new_n37813__ = ~new_new_n37665__ & ~new_new_n37812__;
  assign new_new_n37814__ = ~new_new_n37637__ & ~new_new_n37654__;
  assign new_new_n37815__ = ~new_new_n37812__ & ~new_new_n37814__;
  assign new_new_n37816__ = new_new_n37521__ & ~new_new_n37815__;
  assign new_new_n37817__ = ~new_new_n37521__ & ~new_new_n37814__;
  assign new_new_n37818__ = new_new_n37665__ & new_new_n37817__;
  assign new_new_n37819__ = new_new_n37796__ & ~new_new_n37813__;
  assign new_new_n37820__ = ~new_new_n37816__ & new_new_n37819__;
  assign new_new_n37821__ = ~new_new_n37818__ & new_new_n37820__;
  assign new_new_n37822__ = ~new_new_n37665__ & new_new_n37817__;
  assign new_new_n37823__ = new_new_n37665__ & ~new_new_n37812__;
  assign new_new_n37824__ = ~new_new_n37796__ & ~new_new_n37823__;
  assign new_new_n37825__ = ~new_new_n37816__ & new_new_n37824__;
  assign new_new_n37826__ = ~new_new_n37822__ & new_new_n37825__;
  assign new_new_n37827__ = ~new_new_n37821__ & ~new_new_n37826__;
  assign new_new_n37828__ = new_new_n37647__ & ~new_new_n37827__;
  assign new_new_n37829__ = ~new_new_n37797__ & ~new_new_n37812__;
  assign new_new_n37830__ = ~new_new_n37817__ & new_new_n37829__;
  assign new_new_n37831__ = ~new_new_n37798__ & ~new_new_n37830__;
  assign new_new_n37832__ = new_new_n37828__ & new_new_n37831__;
  assign new_new_n37833__ = ~new_new_n37828__ & ~new_new_n37831__;
  assign new_new_n37834__ = ~new_new_n37832__ & ~new_new_n37833__;
  assign new_new_n37835__ = pi22 & new_new_n34178__;
  assign new_new_n37836__ = ~new_new_n5210__ & ~new_new_n37835__;
  assign new_new_n37837__ = ~new_new_n5181__ & ~new_new_n37836__;
  assign new_new_n37838__ = ~new_new_n5186__ & ~new_new_n5189__;
  assign new_new_n37839__ = ~new_new_n32729__ & ~new_new_n37838__;
  assign new_new_n37840__ = ~pi22 & new_new_n34178__;
  assign new_new_n37841__ = ~new_new_n5211__ & ~new_new_n37840__;
  assign new_new_n37842__ = ~new_new_n5179__ & ~new_new_n37841__;
  assign new_new_n37843__ = ~new_new_n37667__ & ~new_new_n37839__;
  assign new_new_n37844__ = ~new_new_n37837__ & new_new_n37843__;
  assign new_new_n37845__ = ~new_new_n37842__ & new_new_n37844__;
  assign new_new_n37846__ = ~pi23 & ~new_new_n37845__;
  assign new_new_n37847__ = pi23 & new_new_n37845__;
  assign new_new_n37848__ = ~new_new_n37846__ & ~new_new_n37847__;
  assign new_new_n37849__ = ~new_new_n37757__ & new_new_n37790__;
  assign new_new_n37850__ = new_new_n37757__ & ~new_new_n37790__;
  assign new_new_n37851__ = ~new_new_n37849__ & ~new_new_n37850__;
  assign new_new_n37852__ = ~new_new_n37686__ & new_new_n37851__;
  assign new_new_n37853__ = ~new_new_n37685__ & ~new_new_n37852__;
  assign new_new_n37854__ = ~new_new_n4900__ & ~new_new_n33347__;
  assign new_new_n37855__ = ~new_new_n333__ & ~new_new_n26674__;
  assign new_new_n37856__ = new_new_n873__ & ~new_new_n26667__;
  assign new_new_n37857__ = ~new_new_n37855__ & ~new_new_n37856__;
  assign new_new_n37858__ = ~new_new_n37854__ & new_new_n37857__;
  assign new_new_n37859__ = ~pi26 & ~new_new_n37858__;
  assign new_new_n37860__ = new_new_n4898__ & new_new_n32382__;
  assign new_new_n37861__ = new_new_n801__ & new_new_n32382__;
  assign new_new_n37862__ = pi26 & ~new_new_n37861__;
  assign new_new_n37863__ = ~new_new_n37860__ & ~new_new_n37862__;
  assign new_new_n37864__ = new_new_n37858__ & ~new_new_n37863__;
  assign new_new_n37865__ = ~new_new_n37859__ & ~new_new_n37864__;
  assign new_new_n37866__ = ~new_new_n37757__ & ~new_new_n37778__;
  assign new_new_n37867__ = new_new_n37757__ & new_new_n37778__;
  assign new_new_n37868__ = new_new_n4815__ & new_new_n27250__;
  assign new_new_n37869__ = new_new_n37765__ & ~new_new_n37868__;
  assign new_new_n37870__ = pi29 & ~new_new_n37869__;
  assign new_new_n37871__ = ~pi29 & new_new_n37869__;
  assign new_new_n37872__ = ~new_new_n37870__ & ~new_new_n37871__;
  assign new_new_n37873__ = ~new_new_n37867__ & ~new_new_n37872__;
  assign new_new_n37874__ = ~new_new_n37866__ & ~new_new_n37873__;
  assign new_new_n37875__ = new_new_n37865__ & ~new_new_n37874__;
  assign new_new_n37876__ = ~new_new_n37865__ & new_new_n37874__;
  assign new_new_n37877__ = ~new_new_n37875__ & ~new_new_n37876__;
  assign new_new_n37878__ = new_new_n4813__ & new_new_n31511__;
  assign new_new_n37879__ = ~new_new_n4818__ & ~new_new_n27242__;
  assign new_new_n37880__ = new_new_n4212__ & new_new_n27250__;
  assign new_new_n37881__ = ~new_new_n37879__ & ~new_new_n37880__;
  assign new_new_n37882__ = ~new_new_n37878__ & new_new_n37881__;
  assign new_new_n37883__ = new_new_n4214__ & new_new_n26698__;
  assign new_new_n37884__ = ~pi29 & ~new_new_n37883__;
  assign new_new_n37885__ = new_new_n4825__ & new_new_n26698__;
  assign new_new_n37886__ = ~new_new_n37884__ & ~new_new_n37885__;
  assign new_new_n37887__ = new_new_n37882__ & ~new_new_n37886__;
  assign new_new_n37888__ = pi29 & ~new_new_n37882__;
  assign new_new_n37889__ = ~new_new_n37887__ & ~new_new_n37888__;
  assign new_new_n37890__ = ~new_new_n37736__ & new_new_n37751__;
  assign new_new_n37891__ = new_new_n37467__ & new_new_n37571__;
  assign new_new_n37892__ = ~new_new_n37609__ & new_new_n37733__;
  assign new_new_n37893__ = new_new_n37589__ & ~new_new_n37892__;
  assign new_new_n37894__ = ~new_new_n37608__ & new_new_n37735__;
  assign new_new_n37895__ = ~new_new_n37893__ & ~new_new_n37894__;
  assign new_new_n37896__ = ~new_new_n37891__ & ~new_new_n37895__;
  assign new_new_n37897__ = ~new_new_n37589__ & ~new_new_n37609__;
  assign new_new_n37898__ = new_new_n37736__ & ~new_new_n37751__;
  assign new_new_n37899__ = ~new_new_n37608__ & ~new_new_n37897__;
  assign new_new_n37900__ = ~new_new_n37898__ & new_new_n37899__;
  assign new_new_n37901__ = ~new_new_n37890__ & ~new_new_n37896__;
  assign new_new_n37902__ = ~new_new_n37900__ & new_new_n37901__;
  assign new_new_n37903__ = ~new_new_n37889__ & new_new_n37902__;
  assign new_new_n37904__ = new_new_n37889__ & ~new_new_n37902__;
  assign new_new_n37905__ = ~new_new_n37903__ & ~new_new_n37904__;
  assign new_new_n37906__ = ~new_new_n96__ & ~new_new_n240__;
  assign new_new_n37907__ = ~new_new_n315__ & new_new_n37906__;
  assign new_new_n37908__ = ~new_new_n306__ & new_new_n672__;
  assign new_new_n37909__ = new_new_n1077__ & ~new_new_n1167__;
  assign new_new_n37910__ = ~new_new_n1265__ & new_new_n3689__;
  assign new_new_n37911__ = new_new_n37909__ & new_new_n37910__;
  assign new_new_n37912__ = new_new_n37907__ & new_new_n37908__;
  assign new_new_n37913__ = new_new_n1331__ & new_new_n4413__;
  assign new_new_n37914__ = new_new_n17501__ & new_new_n37913__;
  assign new_new_n37915__ = new_new_n37911__ & new_new_n37912__;
  assign new_new_n37916__ = new_new_n2480__ & new_new_n37915__;
  assign new_new_n37917__ = new_new_n3095__ & new_new_n37914__;
  assign new_new_n37918__ = new_new_n37916__ & new_new_n37917__;
  assign new_new_n37919__ = new_new_n18161__ & new_new_n19323__;
  assign new_new_n37920__ = new_new_n37918__ & new_new_n37919__;
  assign new_new_n37921__ = new_new_n1596__ & new_new_n37920__;
  assign new_new_n37922__ = new_new_n5410__ & new_new_n37921__;
  assign new_new_n37923__ = ~pi20 & ~new_new_n37922__;
  assign new_new_n37924__ = pi20 & new_new_n37922__;
  assign new_new_n37925__ = ~new_new_n37923__ & ~new_new_n37924__;
  assign new_new_n37926__ = new_new_n5021__ & new_new_n26722__;
  assign new_new_n37927__ = new_new_n765__ & new_new_n27348__;
  assign new_new_n37928__ = ~new_new_n37723__ & ~new_new_n37927__;
  assign new_new_n37929__ = new_new_n4147__ & new_new_n37928__;
  assign new_new_n37930__ = pi31 & ~new_new_n37928__;
  assign new_new_n37931__ = ~new_new_n5052__ & new_new_n26729__;
  assign new_new_n37932__ = ~new_new_n37930__ & new_new_n37931__;
  assign new_new_n37933__ = ~new_new_n37926__ & ~new_new_n37929__;
  assign new_new_n37934__ = ~new_new_n37932__ & new_new_n37933__;
  assign new_new_n37935__ = new_new_n37925__ & new_new_n37934__;
  assign new_new_n37936__ = ~new_new_n37925__ & ~new_new_n37934__;
  assign new_new_n37937__ = ~new_new_n37935__ & ~new_new_n37936__;
  assign new_new_n37938__ = new_new_n37589__ & ~new_new_n37732__;
  assign new_new_n37939__ = ~new_new_n37589__ & ~new_new_n37731__;
  assign new_new_n37940__ = ~new_new_n37938__ & ~new_new_n37939__;
  assign new_new_n37941__ = new_new_n37937__ & ~new_new_n37940__;
  assign new_new_n37942__ = ~new_new_n37937__ & new_new_n37940__;
  assign new_new_n37943__ = ~new_new_n37941__ & ~new_new_n37942__;
  assign new_new_n37944__ = new_new_n37905__ & ~new_new_n37943__;
  assign new_new_n37945__ = ~new_new_n37905__ & new_new_n37943__;
  assign new_new_n37946__ = ~new_new_n37944__ & ~new_new_n37945__;
  assign new_new_n37947__ = new_new_n37877__ & new_new_n37946__;
  assign new_new_n37948__ = ~new_new_n37877__ & ~new_new_n37946__;
  assign new_new_n37949__ = ~new_new_n37947__ & ~new_new_n37948__;
  assign new_new_n37950__ = new_new_n37853__ & ~new_new_n37949__;
  assign new_new_n37951__ = ~new_new_n37853__ & new_new_n37949__;
  assign new_new_n37952__ = ~new_new_n37950__ & ~new_new_n37951__;
  assign new_new_n37953__ = ~new_new_n37848__ & ~new_new_n37952__;
  assign new_new_n37954__ = new_new_n37848__ & new_new_n37952__;
  assign new_new_n37955__ = ~new_new_n37953__ & ~new_new_n37954__;
  assign new_new_n37956__ = pi20 & new_new_n37689__;
  assign new_new_n37957__ = ~pi20 & ~new_new_n37689__;
  assign new_new_n37958__ = new_new_n37687__ & new_new_n37851__;
  assign new_new_n37959__ = ~new_new_n37687__ & ~new_new_n37851__;
  assign new_new_n37960__ = ~new_new_n37957__ & ~new_new_n37958__;
  assign new_new_n37961__ = ~new_new_n37959__ & new_new_n37960__;
  assign new_new_n37962__ = ~new_new_n37956__ & ~new_new_n37961__;
  assign new_new_n37963__ = ~new_new_n37955__ & new_new_n37962__;
  assign new_new_n37964__ = new_new_n37955__ & ~new_new_n37962__;
  assign new_new_n37965__ = ~new_new_n37963__ & ~new_new_n37964__;
  assign new_new_n37966__ = ~new_new_n37834__ & ~new_new_n37965__;
  assign new_new_n37967__ = new_new_n37834__ & new_new_n37965__;
  assign po25 = ~new_new_n37966__ & ~new_new_n37967__;
  assign new_new_n37969__ = new_new_n37834__ & ~new_new_n37963__;
  assign new_new_n37970__ = new_new_n37832__ & ~new_new_n37964__;
  assign new_new_n37971__ = ~new_new_n37828__ & new_new_n37964__;
  assign new_new_n37972__ = ~new_new_n37970__ & ~new_new_n37971__;
  assign new_new_n37973__ = ~new_new_n37969__ & new_new_n37972__;
  assign new_new_n37974__ = ~new_new_n37848__ & ~new_new_n37951__;
  assign new_new_n37975__ = ~new_new_n37950__ & ~new_new_n37974__;
  assign new_new_n37976__ = new_new_n3311__ & new_new_n32729__;
  assign new_new_n37977__ = ~new_new_n333__ & ~new_new_n26667__;
  assign new_new_n37978__ = new_new_n873__ & new_new_n32382__;
  assign new_new_n37979__ = ~new_new_n37976__ & ~new_new_n37977__;
  assign new_new_n37980__ = ~new_new_n37978__ & new_new_n37979__;
  assign new_new_n37981__ = ~pi26 & ~new_new_n37980__;
  assign new_new_n37982__ = new_new_n512__ & new_new_n32758__;
  assign new_new_n37983__ = new_new_n801__ & new_new_n32758__;
  assign new_new_n37984__ = pi26 & ~new_new_n37983__;
  assign new_new_n37985__ = ~new_new_n37982__ & ~new_new_n37984__;
  assign new_new_n37986__ = new_new_n37980__ & ~new_new_n37985__;
  assign new_new_n37987__ = ~new_new_n37981__ & ~new_new_n37986__;
  assign new_new_n37988__ = new_new_n4212__ & new_new_n26698__;
  assign new_new_n37989__ = ~new_new_n4818__ & new_new_n27250__;
  assign new_new_n37990__ = new_new_n4815__ & ~new_new_n26674__;
  assign new_new_n37991__ = ~new_new_n37988__ & ~new_new_n37989__;
  assign new_new_n37992__ = ~new_new_n37990__ & new_new_n37991__;
  assign new_new_n37993__ = new_new_n4214__ & new_new_n27284__;
  assign new_new_n37994__ = pi29 & ~new_new_n37993__;
  assign new_new_n37995__ = new_new_n4825__ & new_new_n27284__;
  assign new_new_n37996__ = ~new_new_n37994__ & ~new_new_n37995__;
  assign new_new_n37997__ = new_new_n37992__ & ~new_new_n37996__;
  assign new_new_n37998__ = ~pi29 & ~new_new_n37992__;
  assign new_new_n37999__ = ~new_new_n37997__ & ~new_new_n37998__;
  assign new_new_n38000__ = new_new_n37732__ & new_new_n37934__;
  assign new_new_n38001__ = ~new_new_n37732__ & ~new_new_n37934__;
  assign new_new_n38002__ = new_new_n37589__ & ~new_new_n37925__;
  assign new_new_n38003__ = ~new_new_n38001__ & new_new_n38002__;
  assign new_new_n38004__ = new_new_n37731__ & ~new_new_n37935__;
  assign new_new_n38005__ = ~new_new_n37589__ & ~new_new_n37936__;
  assign new_new_n38006__ = ~new_new_n38004__ & new_new_n38005__;
  assign new_new_n38007__ = ~new_new_n38000__ & ~new_new_n38003__;
  assign new_new_n38008__ = ~new_new_n38006__ & new_new_n38007__;
  assign new_new_n38009__ = new_new_n37999__ & ~new_new_n38008__;
  assign new_new_n38010__ = ~new_new_n37999__ & new_new_n38008__;
  assign new_new_n38011__ = ~new_new_n38009__ & ~new_new_n38010__;
  assign new_new_n38012__ = ~new_new_n37589__ & ~new_new_n37924__;
  assign new_new_n38013__ = ~new_new_n37923__ & ~new_new_n38012__;
  assign new_new_n38014__ = ~new_new_n26729__ & ~new_new_n27348__;
  assign new_new_n38015__ = ~new_new_n15853__ & ~new_new_n27350__;
  assign new_new_n38016__ = ~new_new_n38014__ & new_new_n38015__;
  assign new_new_n38017__ = ~new_new_n27334__ & ~new_new_n38016__;
  assign new_new_n38018__ = new_new_n27242__ & ~new_new_n38017__;
  assign new_new_n38019__ = new_new_n26729__ & ~new_new_n27242__;
  assign new_new_n38020__ = new_new_n27348__ & new_new_n38019__;
  assign new_new_n38021__ = ~new_new_n71__ & ~new_new_n38020__;
  assign new_new_n38022__ = ~new_new_n161__ & ~new_new_n26722__;
  assign new_new_n38023__ = ~new_new_n38021__ & new_new_n38022__;
  assign new_new_n38024__ = ~new_new_n27242__ & new_new_n27349__;
  assign new_new_n38025__ = ~new_new_n161__ & ~new_new_n38024__;
  assign new_new_n38026__ = ~new_new_n71__ & ~new_new_n26729__;
  assign new_new_n38027__ = ~new_new_n38025__ & new_new_n38026__;
  assign new_new_n38028__ = pi31 & ~new_new_n38023__;
  assign new_new_n38029__ = ~new_new_n38027__ & new_new_n38028__;
  assign new_new_n38030__ = ~new_new_n38018__ & new_new_n38029__;
  assign new_new_n38031__ = new_new_n161__ & new_new_n26722__;
  assign new_new_n38032__ = new_new_n765__ & ~new_new_n27242__;
  assign new_new_n38033__ = ~new_new_n38031__ & ~new_new_n38032__;
  assign new_new_n38034__ = ~pi31 & ~new_new_n38033__;
  assign new_new_n38035__ = ~new_new_n38030__ & ~new_new_n38034__;
  assign new_new_n38036__ = ~new_new_n247__ & ~new_new_n253__;
  assign new_new_n38037__ = ~new_new_n473__ & new_new_n38036__;
  assign new_new_n38038__ = ~new_new_n192__ & ~new_new_n198__;
  assign new_new_n38039__ = ~new_new_n1073__ & new_new_n4000__;
  assign new_new_n38040__ = new_new_n17421__ & new_new_n38039__;
  assign new_new_n38041__ = new_new_n38037__ & new_new_n38038__;
  assign new_new_n38042__ = new_new_n38040__ & new_new_n38041__;
  assign new_new_n38043__ = new_new_n1076__ & new_new_n4341__;
  assign new_new_n38044__ = new_new_n38042__ & new_new_n38043__;
  assign new_new_n38045__ = new_new_n2201__ & new_new_n38044__;
  assign new_new_n38046__ = new_new_n19280__ & new_new_n38045__;
  assign new_new_n38047__ = new_new_n2354__ & new_new_n4240__;
  assign new_new_n38048__ = new_new_n16294__ & new_new_n38047__;
  assign new_new_n38049__ = new_new_n4978__ & new_new_n38046__;
  assign new_new_n38050__ = new_new_n38048__ & new_new_n38049__;
  assign new_new_n38051__ = new_new_n38035__ & ~new_new_n38050__;
  assign new_new_n38052__ = ~new_new_n38035__ & new_new_n38050__;
  assign new_new_n38053__ = ~new_new_n38051__ & ~new_new_n38052__;
  assign new_new_n38054__ = new_new_n38013__ & new_new_n38053__;
  assign new_new_n38055__ = ~new_new_n38013__ & ~new_new_n38053__;
  assign new_new_n38056__ = ~new_new_n38054__ & ~new_new_n38055__;
  assign new_new_n38057__ = new_new_n38011__ & new_new_n38056__;
  assign new_new_n38058__ = ~new_new_n38011__ & ~new_new_n38056__;
  assign new_new_n38059__ = ~new_new_n38057__ & ~new_new_n38058__;
  assign new_new_n38060__ = ~new_new_n37987__ & ~new_new_n38059__;
  assign new_new_n38061__ = new_new_n37987__ & new_new_n38059__;
  assign new_new_n38062__ = ~new_new_n38060__ & ~new_new_n38061__;
  assign new_new_n38063__ = ~new_new_n37904__ & new_new_n37943__;
  assign new_new_n38064__ = ~new_new_n37903__ & ~new_new_n38063__;
  assign new_new_n38065__ = new_new_n38062__ & ~new_new_n38064__;
  assign new_new_n38066__ = ~new_new_n38062__ & new_new_n38064__;
  assign new_new_n38067__ = ~new_new_n38065__ & ~new_new_n38066__;
  assign new_new_n38068__ = ~new_new_n37876__ & ~new_new_n37946__;
  assign new_new_n38069__ = ~new_new_n37875__ & ~new_new_n38068__;
  assign new_new_n38070__ = ~new_new_n38067__ & new_new_n38069__;
  assign new_new_n38071__ = new_new_n38067__ & ~new_new_n38069__;
  assign new_new_n38072__ = ~new_new_n38070__ & ~new_new_n38071__;
  assign new_new_n38073__ = new_new_n5191__ & new_new_n32740__;
  assign new_new_n38074__ = ~pi23 & new_new_n38073__;
  assign new_new_n38075__ = pi23 & ~new_new_n38073__;
  assign new_new_n38076__ = ~new_new_n38074__ & ~new_new_n38075__;
  assign new_new_n38077__ = new_new_n38072__ & new_new_n38076__;
  assign new_new_n38078__ = ~new_new_n38072__ & ~new_new_n38076__;
  assign new_new_n38079__ = ~new_new_n38077__ & ~new_new_n38078__;
  assign new_new_n38080__ = new_new_n37975__ & new_new_n38079__;
  assign new_new_n38081__ = ~new_new_n37975__ & ~new_new_n38079__;
  assign new_new_n38082__ = ~new_new_n38080__ & ~new_new_n38081__;
  assign new_new_n38083__ = ~new_new_n37973__ & new_new_n38082__;
  assign new_new_n38084__ = ~new_new_n37833__ & ~new_new_n37964__;
  assign new_new_n38085__ = ~new_new_n37832__ & new_new_n37955__;
  assign new_new_n38086__ = ~new_new_n38084__ & ~new_new_n38085__;
  assign new_new_n38087__ = ~new_new_n37833__ & new_new_n37955__;
  assign new_new_n38088__ = ~new_new_n37832__ & new_new_n37962__;
  assign new_new_n38089__ = ~new_new_n38087__ & new_new_n38088__;
  assign new_new_n38090__ = ~new_new_n38086__ & ~new_new_n38089__;
  assign new_new_n38091__ = ~new_new_n38082__ & ~new_new_n38090__;
  assign po26 = new_new_n38083__ | new_new_n38091__;
  assign new_new_n38093__ = new_new_n37831__ & ~new_new_n37963__;
  assign new_new_n38094__ = ~new_new_n37964__ & ~new_new_n38093__;
  assign new_new_n38095__ = new_new_n37975__ & ~new_new_n38094__;
  assign new_new_n38096__ = ~new_new_n38060__ & ~new_new_n38064__;
  assign new_new_n38097__ = ~new_new_n38061__ & ~new_new_n38096__;
  assign new_new_n38098__ = pi23 & new_new_n38097__;
  assign new_new_n38099__ = ~pi23 & ~new_new_n38097__;
  assign new_new_n38100__ = ~new_new_n38098__ & ~new_new_n38099__;
  assign new_new_n38101__ = new_new_n4813__ & ~new_new_n32340__;
  assign new_new_n38102__ = ~new_new_n4818__ & new_new_n26698__;
  assign new_new_n38103__ = new_new_n4212__ & ~new_new_n26674__;
  assign new_new_n38104__ = ~new_new_n38102__ & ~new_new_n38103__;
  assign new_new_n38105__ = ~new_new_n38101__ & new_new_n38104__;
  assign new_new_n38106__ = new_new_n4214__ & ~new_new_n26667__;
  assign new_new_n38107__ = pi29 & ~new_new_n38106__;
  assign new_new_n38108__ = new_new_n5732__ & ~new_new_n26667__;
  assign new_new_n38109__ = ~new_new_n38107__ & ~new_new_n38108__;
  assign new_new_n38110__ = new_new_n38105__ & ~new_new_n38109__;
  assign new_new_n38111__ = ~pi29 & ~new_new_n38105__;
  assign new_new_n38112__ = ~new_new_n38110__ & ~new_new_n38111__;
  assign new_new_n38113__ = new_new_n3311__ & ~new_new_n32382__;
  assign new_new_n38114__ = ~pi26 & new_new_n38113__;
  assign new_new_n38115__ = ~new_new_n4900__ & new_new_n33050__;
  assign new_new_n38116__ = ~new_new_n333__ & new_new_n32382__;
  assign new_new_n38117__ = ~new_new_n38115__ & ~new_new_n38116__;
  assign new_new_n38118__ = ~pi26 & new_new_n38117__;
  assign new_new_n38119__ = ~new_new_n38113__ & ~new_new_n38118__;
  assign new_new_n38120__ = ~new_new_n32729__ & ~new_new_n38114__;
  assign new_new_n38121__ = ~new_new_n38119__ & new_new_n38120__;
  assign new_new_n38122__ = new_new_n873__ & new_new_n32729__;
  assign new_new_n38123__ = new_new_n38117__ & ~new_new_n38122__;
  assign new_new_n38124__ = pi26 & ~new_new_n38123__;
  assign new_new_n38125__ = ~new_new_n9023__ & new_new_n32729__;
  assign new_new_n38126__ = new_new_n38118__ & new_new_n38125__;
  assign new_new_n38127__ = ~new_new_n38124__ & ~new_new_n38126__;
  assign new_new_n38128__ = ~new_new_n38121__ & new_new_n38127__;
  assign new_new_n38129__ = new_new_n161__ & ~new_new_n27242__;
  assign new_new_n38130__ = ~new_new_n15853__ & new_new_n27250__;
  assign new_new_n38131__ = ~new_new_n38129__ & ~new_new_n38130__;
  assign new_new_n38132__ = ~pi31 & ~new_new_n38131__;
  assign new_new_n38133__ = new_new_n71__ & ~new_new_n27242__;
  assign new_new_n38134__ = new_new_n765__ & ~new_new_n27271__;
  assign new_new_n38135__ = ~new_new_n38031__ & ~new_new_n38133__;
  assign new_new_n38136__ = ~new_new_n38134__ & new_new_n38135__;
  assign new_new_n38137__ = pi31 & ~new_new_n38136__;
  assign new_new_n38138__ = ~new_new_n38132__ & ~new_new_n38137__;
  assign new_new_n38139__ = ~new_new_n38009__ & ~new_new_n38056__;
  assign new_new_n38140__ = ~new_new_n38010__ & ~new_new_n38139__;
  assign new_new_n38141__ = ~new_new_n38138__ & ~new_new_n38140__;
  assign new_new_n38142__ = new_new_n38138__ & new_new_n38140__;
  assign new_new_n38143__ = ~new_new_n38141__ & ~new_new_n38142__;
  assign new_new_n38144__ = new_new_n38013__ & new_new_n38050__;
  assign new_new_n38145__ = new_new_n38035__ & new_new_n38144__;
  assign new_new_n38146__ = ~new_new_n38013__ & ~new_new_n38050__;
  assign new_new_n38147__ = ~new_new_n38035__ & new_new_n38146__;
  assign new_new_n38148__ = ~new_new_n38145__ & ~new_new_n38147__;
  assign new_new_n38149__ = new_new_n169__ & ~new_new_n598__;
  assign new_new_n38150__ = new_new_n114__ & ~new_new_n310__;
  assign new_new_n38151__ = new_new_n100__ & ~new_new_n1700__;
  assign new_new_n38152__ = ~new_new_n209__ & ~new_new_n384__;
  assign new_new_n38153__ = ~new_new_n472__ & new_new_n38152__;
  assign new_new_n38154__ = ~new_new_n276__ & ~new_new_n993__;
  assign new_new_n38155__ = new_new_n4062__ & ~new_new_n38149__;
  assign new_new_n38156__ = ~new_new_n38151__ & new_new_n38155__;
  assign new_new_n38157__ = new_new_n38153__ & new_new_n38154__;
  assign new_new_n38158__ = new_new_n1145__ & new_new_n2653__;
  assign new_new_n38159__ = new_new_n3059__ & new_new_n3484__;
  assign new_new_n38160__ = ~new_new_n38150__ & new_new_n38159__;
  assign new_new_n38161__ = new_new_n38157__ & new_new_n38158__;
  assign new_new_n38162__ = new_new_n256__ & new_new_n38156__;
  assign new_new_n38163__ = new_new_n38161__ & new_new_n38162__;
  assign new_new_n38164__ = new_new_n35525__ & new_new_n38160__;
  assign new_new_n38165__ = new_new_n38163__ & new_new_n38164__;
  assign new_new_n38166__ = new_new_n15949__ & new_new_n38165__;
  assign new_new_n38167__ = new_new_n28572__ & new_new_n38166__;
  assign new_new_n38168__ = new_new_n4107__ & new_new_n38167__;
  assign new_new_n38169__ = new_new_n38148__ & ~new_new_n38168__;
  assign new_new_n38170__ = ~new_new_n38148__ & new_new_n38168__;
  assign new_new_n38171__ = ~new_new_n38169__ & ~new_new_n38170__;
  assign new_new_n38172__ = new_new_n38143__ & new_new_n38171__;
  assign new_new_n38173__ = ~new_new_n38143__ & ~new_new_n38171__;
  assign new_new_n38174__ = ~new_new_n38172__ & ~new_new_n38173__;
  assign new_new_n38175__ = ~new_new_n38128__ & new_new_n38174__;
  assign new_new_n38176__ = new_new_n38128__ & ~new_new_n38174__;
  assign new_new_n38177__ = ~new_new_n38112__ & ~new_new_n38175__;
  assign new_new_n38178__ = ~new_new_n38176__ & ~new_new_n38177__;
  assign new_new_n38179__ = ~new_new_n38175__ & new_new_n38178__;
  assign new_new_n38180__ = new_new_n38112__ & ~new_new_n38179__;
  assign new_new_n38181__ = ~new_new_n38176__ & new_new_n38177__;
  assign new_new_n38182__ = ~new_new_n38180__ & ~new_new_n38181__;
  assign new_new_n38183__ = new_new_n38100__ & ~new_new_n38182__;
  assign new_new_n38184__ = ~new_new_n38100__ & new_new_n38182__;
  assign new_new_n38185__ = ~new_new_n38183__ & ~new_new_n38184__;
  assign new_new_n38186__ = ~pi23 & ~new_new_n38070__;
  assign new_new_n38187__ = new_new_n38185__ & new_new_n38186__;
  assign new_new_n38188__ = ~new_new_n38071__ & ~new_new_n38185__;
  assign new_new_n38189__ = pi23 & new_new_n38188__;
  assign new_new_n38190__ = ~new_new_n38187__ & ~new_new_n38189__;
  assign new_new_n38191__ = ~new_new_n38073__ & ~new_new_n38190__;
  assign new_new_n38192__ = pi23 & new_new_n38073__;
  assign new_new_n38193__ = ~new_new_n38070__ & new_new_n38192__;
  assign new_new_n38194__ = ~new_new_n38071__ & ~new_new_n38193__;
  assign new_new_n38195__ = new_new_n38185__ & ~new_new_n38194__;
  assign new_new_n38196__ = ~new_new_n38070__ & ~new_new_n38074__;
  assign new_new_n38197__ = new_new_n38188__ & ~new_new_n38196__;
  assign new_new_n38198__ = ~new_new_n38195__ & ~new_new_n38197__;
  assign new_new_n38199__ = ~new_new_n38191__ & new_new_n38198__;
  assign new_new_n38200__ = new_new_n38095__ & new_new_n38199__;
  assign new_new_n38201__ = ~new_new_n38095__ & ~new_new_n38199__;
  assign new_new_n38202__ = new_new_n38082__ & ~new_new_n38094__;
  assign new_new_n38203__ = ~new_new_n38082__ & new_new_n38094__;
  assign new_new_n38204__ = ~new_new_n38202__ & ~new_new_n38203__;
  assign new_new_n38205__ = ~new_new_n38200__ & ~new_new_n38201__;
  assign new_new_n38206__ = ~new_new_n38204__ & new_new_n38205__;
  assign new_new_n38207__ = ~po26 & new_new_n38206__;
  assign new_new_n38208__ = ~new_new_n37975__ & new_new_n38094__;
  assign new_new_n38209__ = ~new_new_n38079__ & ~new_new_n38208__;
  assign new_new_n38210__ = ~new_new_n38079__ & ~po26;
  assign new_new_n38211__ = ~new_new_n38095__ & new_new_n38199__;
  assign new_new_n38212__ = ~new_new_n38210__ & ~new_new_n38211__;
  assign new_new_n38213__ = ~new_new_n38209__ & ~new_new_n38212__;
  assign new_new_n38214__ = new_new_n38079__ & ~new_new_n38095__;
  assign new_new_n38215__ = po26 & new_new_n38214__;
  assign new_new_n38216__ = ~new_new_n38199__ & ~new_new_n38208__;
  assign new_new_n38217__ = ~new_new_n38215__ & new_new_n38216__;
  assign new_new_n38218__ = ~new_new_n38213__ & ~new_new_n38217__;
  assign new_new_n38219__ = ~new_new_n38207__ & ~new_new_n38218__;
  assign new_new_n38220__ = new_new_n38200__ & new_new_n38210__;
  assign po27 = new_new_n38219__ | new_new_n38220__;
  assign new_new_n38222__ = new_new_n4212__ & ~new_new_n26667__;
  assign new_new_n38223__ = ~new_new_n4818__ & ~new_new_n26674__;
  assign new_new_n38224__ = new_new_n4815__ & new_new_n32382__;
  assign new_new_n38225__ = ~new_new_n38222__ & ~new_new_n38223__;
  assign new_new_n38226__ = ~new_new_n38224__ & new_new_n38225__;
  assign new_new_n38227__ = new_new_n4214__ & ~new_new_n33347__;
  assign new_new_n38228__ = ~pi29 & ~new_new_n38227__;
  assign new_new_n38229__ = new_new_n5732__ & ~new_new_n33347__;
  assign new_new_n38230__ = ~new_new_n38228__ & ~new_new_n38229__;
  assign new_new_n38231__ = new_new_n38226__ & ~new_new_n38230__;
  assign new_new_n38232__ = pi29 & ~new_new_n38226__;
  assign new_new_n38233__ = ~new_new_n38231__ & ~new_new_n38232__;
  assign new_new_n38234__ = ~new_new_n38142__ & ~new_new_n38171__;
  assign new_new_n38235__ = ~new_new_n38141__ & ~new_new_n38234__;
  assign new_new_n38236__ = ~new_new_n38233__ & new_new_n38235__;
  assign new_new_n38237__ = new_new_n38233__ & ~new_new_n38235__;
  assign new_new_n38238__ = ~new_new_n38236__ & ~new_new_n38237__;
  assign new_new_n38239__ = ~new_new_n164__ & ~new_new_n718__;
  assign new_new_n38240__ = ~new_new_n251__ & ~new_new_n670__;
  assign new_new_n38241__ = ~new_new_n724__ & ~new_new_n826__;
  assign new_new_n38242__ = new_new_n38240__ & new_new_n38241__;
  assign new_new_n38243__ = ~new_new_n993__ & new_new_n38239__;
  assign new_new_n38244__ = new_new_n1709__ & ~new_new_n1921__;
  assign new_new_n38245__ = new_new_n38243__ & new_new_n38244__;
  assign new_new_n38246__ = ~new_new_n809__ & new_new_n38242__;
  assign new_new_n38247__ = new_new_n941__ & new_new_n2771__;
  assign new_new_n38248__ = new_new_n16793__ & new_new_n38247__;
  assign new_new_n38249__ = new_new_n38245__ & new_new_n38246__;
  assign new_new_n38250__ = new_new_n5593__ & new_new_n38249__;
  assign new_new_n38251__ = new_new_n38248__ & new_new_n38250__;
  assign new_new_n38252__ = new_new_n565__ & new_new_n38251__;
  assign new_new_n38253__ = new_new_n3835__ & new_new_n38252__;
  assign new_new_n38254__ = new_new_n38168__ & new_new_n38253__;
  assign new_new_n38255__ = ~new_new_n38168__ & ~new_new_n38253__;
  assign new_new_n38256__ = ~new_new_n38254__ & ~new_new_n38255__;
  assign new_new_n38257__ = ~pi23 & ~new_new_n38256__;
  assign new_new_n38258__ = pi23 & new_new_n38256__;
  assign new_new_n38259__ = ~new_new_n38257__ & ~new_new_n38258__;
  assign new_new_n38260__ = new_new_n161__ & new_new_n27250__;
  assign new_new_n38261__ = new_new_n765__ & new_new_n26698__;
  assign new_new_n38262__ = ~new_new_n38260__ & ~new_new_n38261__;
  assign new_new_n38263__ = ~pi31 & ~new_new_n38262__;
  assign new_new_n38264__ = new_new_n161__ & new_new_n27242__;
  assign new_new_n38265__ = ~new_new_n71__ & ~new_new_n32299__;
  assign new_new_n38266__ = ~new_new_n161__ & ~new_new_n27250__;
  assign new_new_n38267__ = ~new_new_n38265__ & new_new_n38266__;
  assign new_new_n38268__ = ~new_new_n32299__ & new_new_n38130__;
  assign new_new_n38269__ = pi31 & ~new_new_n38264__;
  assign new_new_n38270__ = ~new_new_n38268__ & new_new_n38269__;
  assign new_new_n38271__ = ~new_new_n38267__ & new_new_n38270__;
  assign new_new_n38272__ = ~new_new_n38263__ & ~new_new_n38271__;
  assign new_new_n38273__ = ~new_new_n38147__ & ~new_new_n38168__;
  assign new_new_n38274__ = ~new_new_n38145__ & ~new_new_n38273__;
  assign new_new_n38275__ = ~new_new_n38272__ & new_new_n38274__;
  assign new_new_n38276__ = new_new_n38272__ & ~new_new_n38274__;
  assign new_new_n38277__ = ~new_new_n38275__ & ~new_new_n38276__;
  assign new_new_n38278__ = new_new_n38259__ & new_new_n38277__;
  assign new_new_n38279__ = ~new_new_n38259__ & ~new_new_n38277__;
  assign new_new_n38280__ = ~new_new_n38278__ & ~new_new_n38279__;
  assign new_new_n38281__ = new_new_n38238__ & new_new_n38280__;
  assign new_new_n38282__ = ~new_new_n38238__ & ~new_new_n38280__;
  assign new_new_n38283__ = ~new_new_n38281__ & ~new_new_n38282__;
  assign new_new_n38284__ = ~new_new_n38098__ & ~new_new_n38182__;
  assign new_new_n38285__ = ~new_new_n38099__ & ~new_new_n38284__;
  assign new_new_n38286__ = new_new_n38185__ & ~new_new_n38199__;
  assign new_new_n38287__ = ~new_new_n38209__ & new_new_n38211__;
  assign new_new_n38288__ = ~new_new_n38286__ & ~new_new_n38287__;
  assign new_new_n38289__ = ~new_new_n349__ & ~new_new_n34178__;
  assign new_new_n38290__ = pi26 & ~new_new_n38289__;
  assign new_new_n38291__ = pi25 & new_new_n99__;
  assign new_new_n38292__ = ~pi26 & ~new_new_n389__;
  assign new_new_n38293__ = ~new_new_n38291__ & new_new_n38292__;
  assign new_new_n38294__ = ~new_new_n34178__ & new_new_n38293__;
  assign new_new_n38295__ = ~new_new_n38290__ & ~new_new_n38294__;
  assign new_new_n38296__ = ~new_new_n32729__ & ~new_new_n38295__;
  assign new_new_n38297__ = ~pi25 & ~new_new_n34178__;
  assign new_new_n38298__ = ~pi26 & ~new_new_n34177__;
  assign new_new_n38299__ = ~new_new_n104__ & ~new_new_n38298__;
  assign new_new_n38300__ = ~new_new_n38297__ & new_new_n38299__;
  assign new_new_n38301__ = ~new_new_n430__ & ~new_new_n4780__;
  assign new_new_n38302__ = new_new_n32729__ & new_new_n38301__;
  assign new_new_n38303__ = ~new_new_n38300__ & ~new_new_n38302__;
  assign new_new_n38304__ = ~new_new_n38296__ & new_new_n38303__;
  assign new_new_n38305__ = new_new_n38178__ & ~new_new_n38304__;
  assign new_new_n38306__ = ~new_new_n38178__ & new_new_n38304__;
  assign new_new_n38307__ = ~new_new_n38305__ & ~new_new_n38306__;
  assign new_new_n38308__ = new_new_n38288__ & ~new_new_n38307__;
  assign new_new_n38309__ = ~new_new_n38288__ & new_new_n38307__;
  assign new_new_n38310__ = ~new_new_n38308__ & ~new_new_n38309__;
  assign new_new_n38311__ = new_new_n38207__ & new_new_n38310__;
  assign new_new_n38312__ = ~new_new_n38207__ & ~new_new_n38310__;
  assign new_new_n38313__ = ~new_new_n38311__ & ~new_new_n38312__;
  assign new_new_n38314__ = new_new_n38285__ & ~new_new_n38313__;
  assign new_new_n38315__ = ~new_new_n38285__ & new_new_n38313__;
  assign new_new_n38316__ = ~new_new_n38314__ & ~new_new_n38315__;
  assign new_new_n38317__ = new_new_n38283__ & new_new_n38316__;
  assign new_new_n38318__ = ~new_new_n38283__ & ~new_new_n38316__;
  assign po28 = ~new_new_n38317__ & ~new_new_n38318__;
  assign new_new_n38320__ = new_new_n4813__ & new_new_n32758__;
  assign new_new_n38321__ = ~new_new_n4818__ & ~new_new_n26667__;
  assign new_new_n38322__ = new_new_n4212__ & new_new_n32382__;
  assign new_new_n38323__ = ~new_new_n38321__ & ~new_new_n38322__;
  assign new_new_n38324__ = ~new_new_n38320__ & new_new_n38323__;
  assign new_new_n38325__ = new_new_n4214__ & new_new_n32729__;
  assign new_new_n38326__ = ~pi29 & ~new_new_n38325__;
  assign new_new_n38327__ = new_new_n4825__ & new_new_n32729__;
  assign new_new_n38328__ = ~new_new_n38326__ & ~new_new_n38327__;
  assign new_new_n38329__ = new_new_n38324__ & ~new_new_n38328__;
  assign new_new_n38330__ = pi29 & ~new_new_n38324__;
  assign new_new_n38331__ = ~new_new_n38329__ & ~new_new_n38330__;
  assign new_new_n38332__ = ~new_new_n38259__ & ~new_new_n38276__;
  assign new_new_n38333__ = ~new_new_n38275__ & ~new_new_n38332__;
  assign new_new_n38334__ = new_new_n38331__ & ~new_new_n38333__;
  assign new_new_n38335__ = ~new_new_n38331__ & new_new_n38333__;
  assign new_new_n38336__ = ~new_new_n38334__ & ~new_new_n38335__;
  assign new_new_n38337__ = new_new_n26674__ & new_new_n32298__;
  assign new_new_n38338__ = ~new_new_n161__ & ~new_new_n27287__;
  assign new_new_n38339__ = ~new_new_n38337__ & new_new_n38338__;
  assign new_new_n38340__ = new_new_n27250__ & ~new_new_n38339__;
  assign new_new_n38341__ = new_new_n27250__ & ~new_new_n27275__;
  assign new_new_n38342__ = ~new_new_n26674__ & new_new_n32297__;
  assign new_new_n38343__ = new_new_n26674__ & ~new_new_n32297__;
  assign new_new_n38344__ = ~new_new_n161__ & ~new_new_n38341__;
  assign new_new_n38345__ = ~new_new_n38342__ & ~new_new_n38343__;
  assign new_new_n38346__ = new_new_n38344__ & new_new_n38345__;
  assign new_new_n38347__ = new_new_n4147__ & ~new_new_n38340__;
  assign new_new_n38348__ = ~new_new_n38346__ & new_new_n38347__;
  assign new_new_n38349__ = new_new_n161__ & new_new_n26698__;
  assign new_new_n38350__ = ~new_new_n71__ & new_new_n38349__;
  assign new_new_n38351__ = new_new_n71__ & ~new_new_n26698__;
  assign new_new_n38352__ = pi31 & ~new_new_n38351__;
  assign new_new_n38353__ = ~new_new_n15853__ & ~new_new_n26674__;
  assign new_new_n38354__ = ~new_new_n38350__ & ~new_new_n38352__;
  assign new_new_n38355__ = ~new_new_n38353__ & new_new_n38354__;
  assign new_new_n38356__ = ~new_new_n38348__ & ~new_new_n38355__;
  assign new_new_n38357__ = ~pi23 & ~new_new_n38254__;
  assign new_new_n38358__ = ~new_new_n38255__ & ~new_new_n38357__;
  assign new_new_n38359__ = ~new_new_n168__ & ~new_new_n240__;
  assign new_new_n38360__ = ~new_new_n996__ & new_new_n38359__;
  assign new_new_n38361__ = ~new_new_n192__ & new_new_n1218__;
  assign new_new_n38362__ = new_new_n2640__ & new_new_n38361__;
  assign new_new_n38363__ = new_new_n227__ & new_new_n38360__;
  assign new_new_n38364__ = new_new_n281__ & new_new_n330__;
  assign new_new_n38365__ = new_new_n1097__ & new_new_n1611__;
  assign new_new_n38366__ = new_new_n2453__ & new_new_n4073__;
  assign new_new_n38367__ = new_new_n38365__ & new_new_n38366__;
  assign new_new_n38368__ = new_new_n38363__ & new_new_n38364__;
  assign new_new_n38369__ = new_new_n554__ & new_new_n38362__;
  assign new_new_n38370__ = new_new_n4573__ & new_new_n5432__;
  assign new_new_n38371__ = new_new_n15933__ & new_new_n38370__;
  assign new_new_n38372__ = new_new_n38368__ & new_new_n38369__;
  assign new_new_n38373__ = new_new_n38367__ & new_new_n38372__;
  assign new_new_n38374__ = new_new_n667__ & new_new_n38371__;
  assign new_new_n38375__ = new_new_n38373__ & new_new_n38374__;
  assign new_new_n38376__ = new_new_n19142__ & new_new_n38375__;
  assign new_new_n38377__ = new_new_n38358__ & ~new_new_n38376__;
  assign new_new_n38378__ = ~new_new_n38358__ & new_new_n38376__;
  assign new_new_n38379__ = ~new_new_n38377__ & ~new_new_n38378__;
  assign new_new_n38380__ = ~new_new_n38356__ & ~new_new_n38379__;
  assign new_new_n38381__ = new_new_n38356__ & new_new_n38379__;
  assign new_new_n38382__ = ~new_new_n38380__ & ~new_new_n38381__;
  assign new_new_n38383__ = new_new_n38336__ & ~new_new_n38382__;
  assign new_new_n38384__ = ~new_new_n38336__ & new_new_n38382__;
  assign new_new_n38385__ = ~new_new_n38383__ & ~new_new_n38384__;
  assign new_new_n38386__ = ~new_new_n38236__ & ~new_new_n38280__;
  assign new_new_n38387__ = ~new_new_n38237__ & ~new_new_n38386__;
  assign new_new_n38388__ = ~new_new_n38385__ & ~new_new_n38387__;
  assign new_new_n38389__ = new_new_n38385__ & new_new_n38387__;
  assign new_new_n38390__ = ~new_new_n38388__ & ~new_new_n38389__;
  assign new_new_n38391__ = ~new_new_n333__ & new_new_n32740__;
  assign new_new_n38392__ = ~pi26 & ~new_new_n38391__;
  assign new_new_n38393__ = pi26 & new_new_n38391__;
  assign new_new_n38394__ = ~new_new_n38392__ & ~new_new_n38393__;
  assign new_new_n38395__ = new_new_n38390__ & ~new_new_n38394__;
  assign new_new_n38396__ = ~new_new_n38390__ & new_new_n38394__;
  assign new_new_n38397__ = ~new_new_n38395__ & ~new_new_n38396__;
  assign new_new_n38398__ = ~new_new_n38178__ & ~new_new_n38283__;
  assign new_new_n38399__ = new_new_n38178__ & new_new_n38283__;
  assign new_new_n38400__ = ~new_new_n38398__ & ~new_new_n38399__;
  assign new_new_n38401__ = new_new_n38307__ & ~new_new_n38400__;
  assign new_new_n38402__ = new_new_n38285__ & new_new_n38288__;
  assign new_new_n38403__ = ~new_new_n38285__ & ~new_new_n38288__;
  assign new_new_n38404__ = ~new_new_n38401__ & ~new_new_n38402__;
  assign new_new_n38405__ = ~new_new_n38403__ & new_new_n38404__;
  assign new_new_n38406__ = ~new_new_n38304__ & ~new_new_n38399__;
  assign new_new_n38407__ = ~new_new_n38398__ & ~new_new_n38406__;
  assign new_new_n38408__ = new_new_n38403__ & ~new_new_n38407__;
  assign new_new_n38409__ = new_new_n38402__ & new_new_n38407__;
  assign new_new_n38410__ = ~new_new_n38408__ & ~new_new_n38409__;
  assign new_new_n38411__ = ~new_new_n38405__ & new_new_n38410__;
  assign new_new_n38412__ = ~new_new_n38397__ & ~new_new_n38411__;
  assign new_new_n38413__ = new_new_n38283__ & ~new_new_n38288__;
  assign new_new_n38414__ = ~new_new_n38283__ & new_new_n38288__;
  assign new_new_n38415__ = ~new_new_n38285__ & ~new_new_n38414__;
  assign new_new_n38416__ = ~new_new_n38413__ & ~new_new_n38415__;
  assign new_new_n38417__ = ~new_new_n38178__ & new_new_n38416__;
  assign new_new_n38418__ = new_new_n38285__ & new_new_n38414__;
  assign new_new_n38419__ = ~new_new_n38417__ & ~new_new_n38418__;
  assign new_new_n38420__ = ~new_new_n38304__ & ~new_new_n38419__;
  assign new_new_n38421__ = ~new_new_n38178__ & new_new_n38285__;
  assign new_new_n38422__ = new_new_n38414__ & new_new_n38421__;
  assign new_new_n38423__ = ~new_new_n38285__ & new_new_n38413__;
  assign new_new_n38424__ = new_new_n38178__ & new_new_n38423__;
  assign new_new_n38425__ = ~new_new_n38178__ & ~new_new_n38423__;
  assign new_new_n38426__ = new_new_n38304__ & ~new_new_n38416__;
  assign new_new_n38427__ = ~new_new_n38425__ & new_new_n38426__;
  assign new_new_n38428__ = ~new_new_n38422__ & ~new_new_n38424__;
  assign new_new_n38429__ = ~new_new_n38427__ & new_new_n38428__;
  assign new_new_n38430__ = ~new_new_n38420__ & new_new_n38429__;
  assign new_new_n38431__ = new_new_n38397__ & ~new_new_n38430__;
  assign new_new_n38432__ = ~new_new_n38412__ & ~new_new_n38431__;
  assign new_new_n38433__ = new_new_n38207__ & ~po28;
  assign new_new_n38434__ = new_new_n38432__ & new_new_n38433__;
  assign new_new_n38435__ = ~new_new_n38432__ & ~new_new_n38433__;
  assign po29 = ~new_new_n38434__ & ~new_new_n38435__;
  assign new_new_n38437__ = new_new_n38178__ & ~new_new_n38285__;
  assign new_new_n38438__ = new_new_n38397__ & ~new_new_n38421__;
  assign new_new_n38439__ = ~new_new_n38304__ & ~new_new_n38438__;
  assign new_new_n38440__ = ~new_new_n38414__ & ~new_new_n38439__;
  assign new_new_n38441__ = new_new_n38437__ & new_new_n38440__;
  assign new_new_n38442__ = ~new_new_n38413__ & ~new_new_n38440__;
  assign new_new_n38443__ = new_new_n38397__ & ~new_new_n38442__;
  assign new_new_n38444__ = ~new_new_n38304__ & ~new_new_n38437__;
  assign new_new_n38445__ = ~new_new_n38397__ & ~new_new_n38413__;
  assign new_new_n38446__ = ~new_new_n38421__ & ~new_new_n38444__;
  assign new_new_n38447__ = ~new_new_n38445__ & new_new_n38446__;
  assign new_new_n38448__ = ~new_new_n38441__ & ~new_new_n38447__;
  assign new_new_n38449__ = ~new_new_n38443__ & new_new_n38448__;
  assign new_new_n38450__ = ~new_new_n164__ & ~new_new_n541__;
  assign new_new_n38451__ = new_new_n177__ & new_new_n38450__;
  assign new_new_n38452__ = new_new_n421__ & new_new_n38451__;
  assign new_new_n38453__ = ~new_new_n805__ & new_new_n15933__;
  assign new_new_n38454__ = new_new_n38452__ & new_new_n38453__;
  assign new_new_n38455__ = new_new_n2753__ & new_new_n38454__;
  assign new_new_n38456__ = new_new_n3859__ & new_new_n38455__;
  assign new_new_n38457__ = new_new_n38376__ & ~new_new_n38456__;
  assign new_new_n38458__ = ~new_new_n38376__ & new_new_n38456__;
  assign new_new_n38459__ = ~new_new_n38457__ & ~new_new_n38458__;
  assign new_new_n38460__ = ~new_new_n38356__ & ~new_new_n38378__;
  assign new_new_n38461__ = ~new_new_n38377__ & ~new_new_n38460__;
  assign new_new_n38462__ = new_new_n38459__ & new_new_n38461__;
  assign new_new_n38463__ = ~new_new_n38459__ & ~new_new_n38461__;
  assign new_new_n38464__ = ~new_new_n38462__ & ~new_new_n38463__;
  assign new_new_n38465__ = pi26 & new_new_n38464__;
  assign new_new_n38466__ = ~pi26 & ~new_new_n38464__;
  assign new_new_n38467__ = ~new_new_n38465__ & ~new_new_n38466__;
  assign new_new_n38468__ = new_new_n4813__ & new_new_n33050__;
  assign new_new_n38469__ = new_new_n4815__ & new_new_n32740__;
  assign new_new_n38470__ = new_new_n4212__ & new_new_n32729__;
  assign new_new_n38471__ = ~new_new_n38469__ & ~new_new_n38470__;
  assign new_new_n38472__ = ~new_new_n38468__ & new_new_n38471__;
  assign new_new_n38473__ = new_new_n67__ & new_new_n32382__;
  assign new_new_n38474__ = pi29 & ~new_new_n38473__;
  assign new_new_n38475__ = new_new_n65__ & new_new_n32382__;
  assign new_new_n38476__ = ~pi29 & ~new_new_n38475__;
  assign new_new_n38477__ = pi26 & ~new_new_n38476__;
  assign new_new_n38478__ = ~new_new_n38474__ & ~new_new_n38477__;
  assign new_new_n38479__ = new_new_n38472__ & ~new_new_n38478__;
  assign new_new_n38480__ = ~pi29 & ~new_new_n38472__;
  assign new_new_n38481__ = ~new_new_n38479__ & ~new_new_n38480__;
  assign new_new_n38482__ = new_new_n5053__ & ~new_new_n26674__;
  assign new_new_n38483__ = ~new_new_n161__ & ~new_new_n32340__;
  assign new_new_n38484__ = ~new_new_n38349__ & ~new_new_n38483__;
  assign new_new_n38485__ = pi31 & ~new_new_n38484__;
  assign new_new_n38486__ = new_new_n5052__ & ~new_new_n26667__;
  assign new_new_n38487__ = ~new_new_n38485__ & ~new_new_n38486__;
  assign new_new_n38488__ = ~new_new_n71__ & ~new_new_n38487__;
  assign new_new_n38489__ = ~new_new_n38482__ & ~new_new_n38488__;
  assign new_new_n38490__ = ~new_new_n38335__ & new_new_n38382__;
  assign new_new_n38491__ = ~new_new_n38334__ & ~new_new_n38490__;
  assign new_new_n38492__ = new_new_n38489__ & new_new_n38491__;
  assign new_new_n38493__ = ~new_new_n38489__ & ~new_new_n38491__;
  assign new_new_n38494__ = ~new_new_n38492__ & ~new_new_n38493__;
  assign new_new_n38495__ = new_new_n38481__ & ~new_new_n38494__;
  assign new_new_n38496__ = ~new_new_n38481__ & new_new_n38494__;
  assign new_new_n38497__ = ~new_new_n38495__ & ~new_new_n38496__;
  assign new_new_n38498__ = new_new_n38467__ & new_new_n38497__;
  assign new_new_n38499__ = ~new_new_n38467__ & ~new_new_n38497__;
  assign new_new_n38500__ = ~new_new_n38498__ & ~new_new_n38499__;
  assign new_new_n38501__ = ~new_new_n38434__ & new_new_n38500__;
  assign new_new_n38502__ = new_new_n38434__ & ~new_new_n38500__;
  assign new_new_n38503__ = ~new_new_n38501__ & ~new_new_n38502__;
  assign new_new_n38504__ = ~new_new_n38389__ & new_new_n38394__;
  assign new_new_n38505__ = ~new_new_n38388__ & ~new_new_n38504__;
  assign new_new_n38506__ = new_new_n38503__ & ~new_new_n38505__;
  assign new_new_n38507__ = ~new_new_n38503__ & new_new_n38505__;
  assign new_new_n38508__ = ~new_new_n38506__ & ~new_new_n38507__;
  assign new_new_n38509__ = new_new_n38449__ & ~new_new_n38508__;
  assign new_new_n38510__ = ~new_new_n38449__ & new_new_n38508__;
  assign po30 = ~new_new_n38509__ & ~new_new_n38510__;
  assign new_new_n38512__ = new_new_n38434__ & ~new_new_n38449__;
  assign new_new_n38513__ = ~new_new_n38501__ & ~new_new_n38512__;
  assign new_new_n38514__ = new_new_n38500__ & ~new_new_n38505__;
  assign new_new_n38515__ = new_new_n38449__ & ~new_new_n38514__;
  assign new_new_n38516__ = new_new_n38513__ & ~new_new_n38515__;
  assign new_new_n38517__ = ~new_new_n38449__ & ~new_new_n38500__;
  assign new_new_n38518__ = ~new_new_n38434__ & new_new_n38505__;
  assign new_new_n38519__ = ~new_new_n38517__ & ~new_new_n38518__;
  assign new_new_n38520__ = po30 & ~new_new_n38519__;
  assign new_new_n38521__ = ~new_new_n38516__ & ~new_new_n38520__;
  assign new_new_n38522__ = ~new_new_n38465__ & new_new_n38481__;
  assign new_new_n38523__ = ~new_new_n38466__ & ~new_new_n38522__;
  assign new_new_n38524__ = new_new_n38492__ & new_new_n38523__;
  assign new_new_n38525__ = new_new_n38464__ & ~new_new_n38481__;
  assign new_new_n38526__ = ~new_new_n38464__ & new_new_n38481__;
  assign new_new_n38527__ = ~new_new_n38525__ & ~new_new_n38526__;
  assign new_new_n38528__ = ~new_new_n38467__ & ~new_new_n38527__;
  assign new_new_n38529__ = new_new_n38494__ & ~new_new_n38528__;
  assign new_new_n38530__ = new_new_n38493__ & ~new_new_n38523__;
  assign new_new_n38531__ = ~pi29 & new_new_n462__;
  assign new_new_n38532__ = ~pi26 & new_new_n38531__;
  assign new_new_n38533__ = pi26 & ~new_new_n38531__;
  assign new_new_n38534__ = ~new_new_n38376__ & new_new_n38533__;
  assign new_new_n38535__ = new_new_n38376__ & ~new_new_n38533__;
  assign new_new_n38536__ = new_new_n3765__ & ~new_new_n38532__;
  assign new_new_n38537__ = ~new_new_n38534__ & new_new_n38536__;
  assign new_new_n38538__ = ~new_new_n38535__ & new_new_n38537__;
  assign new_new_n38539__ = new_new_n264__ & new_new_n38376__;
  assign new_new_n38540__ = pi29 & ~new_new_n38376__;
  assign new_new_n38541__ = pi26 & ~new_new_n3765__;
  assign new_new_n38542__ = new_new_n38540__ & new_new_n38541__;
  assign new_new_n38543__ = ~new_new_n38539__ & ~new_new_n38542__;
  assign new_new_n38544__ = new_new_n462__ & ~new_new_n38543__;
  assign new_new_n38545__ = ~pi26 & ~new_new_n3765__;
  assign new_new_n38546__ = ~new_new_n38540__ & new_new_n38545__;
  assign new_new_n38547__ = ~new_new_n38538__ & ~new_new_n38546__;
  assign new_new_n38548__ = ~new_new_n38544__ & new_new_n38547__;
  assign new_new_n38549__ = ~new_new_n76__ & ~new_new_n38548__;
  assign new_new_n38550__ = new_new_n5053__ & ~new_new_n26667__;
  assign new_new_n38551__ = new_new_n5059__ & ~new_new_n26674__;
  assign new_new_n38552__ = pi31 & new_new_n33347__;
  assign new_new_n38553__ = ~pi31 & ~new_new_n32382__;
  assign new_new_n38554__ = new_new_n765__ & ~new_new_n38553__;
  assign new_new_n38555__ = ~new_new_n38552__ & new_new_n38554__;
  assign new_new_n38556__ = ~new_new_n38550__ & ~new_new_n38551__;
  assign new_new_n38557__ = ~new_new_n38555__ & new_new_n38556__;
  assign new_new_n38558__ = ~new_new_n38549__ & ~new_new_n38557__;
  assign new_new_n38559__ = new_new_n38549__ & new_new_n38557__;
  assign new_new_n38560__ = ~new_new_n38558__ & ~new_new_n38559__;
  assign new_new_n38561__ = new_new_n4813__ & ~new_new_n34178__;
  assign new_new_n38562__ = new_new_n4818__ & ~new_new_n38561__;
  assign new_new_n38563__ = ~new_new_n4813__ & ~new_new_n32729__;
  assign new_new_n38564__ = ~new_new_n38562__ & ~new_new_n38563__;
  assign new_new_n38565__ = new_new_n38560__ & ~new_new_n38564__;
  assign new_new_n38566__ = ~new_new_n32729__ & ~new_new_n38561__;
  assign new_new_n38567__ = ~new_new_n38562__ & ~new_new_n38566__;
  assign new_new_n38568__ = ~new_new_n38560__ & new_new_n38567__;
  assign new_new_n38569__ = ~new_new_n38565__ & ~new_new_n38568__;
  assign new_new_n38570__ = ~new_new_n38457__ & ~new_new_n38461__;
  assign new_new_n38571__ = ~new_new_n38458__ & ~new_new_n38570__;
  assign new_new_n38572__ = new_new_n38569__ & ~new_new_n38571__;
  assign new_new_n38573__ = ~new_new_n38569__ & new_new_n38571__;
  assign new_new_n38574__ = ~new_new_n38572__ & ~new_new_n38573__;
  assign new_new_n38575__ = ~new_new_n38524__ & ~new_new_n38530__;
  assign new_new_n38576__ = new_new_n38574__ & new_new_n38575__;
  assign new_new_n38577__ = ~new_new_n38529__ & new_new_n38576__;
  assign new_new_n38578__ = new_new_n38481__ & new_new_n38492__;
  assign new_new_n38579__ = ~new_new_n38464__ & new_new_n38578__;
  assign new_new_n38580__ = ~new_new_n38481__ & ~new_new_n38492__;
  assign new_new_n38581__ = ~new_new_n38464__ & ~new_new_n38493__;
  assign new_new_n38582__ = ~new_new_n38580__ & new_new_n38581__;
  assign new_new_n38583__ = ~new_new_n38578__ & ~new_new_n38582__;
  assign new_new_n38584__ = ~pi26 & ~new_new_n38583__;
  assign new_new_n38585__ = new_new_n38493__ & new_new_n38525__;
  assign new_new_n38586__ = new_new_n38493__ & ~new_new_n38526__;
  assign new_new_n38587__ = new_new_n38464__ & new_new_n38580__;
  assign new_new_n38588__ = ~new_new_n38586__ & ~new_new_n38587__;
  assign new_new_n38589__ = pi26 & ~new_new_n38588__;
  assign new_new_n38590__ = ~new_new_n38574__ & ~new_new_n38585__;
  assign new_new_n38591__ = ~new_new_n38579__ & new_new_n38590__;
  assign new_new_n38592__ = ~new_new_n38584__ & new_new_n38591__;
  assign new_new_n38593__ = ~new_new_n38589__ & new_new_n38592__;
  assign new_new_n38594__ = ~new_new_n38577__ & ~new_new_n38593__;
  assign new_new_n38595__ = ~new_new_n38521__ & new_new_n38594__;
  assign new_new_n38596__ = ~new_new_n38505__ & ~new_new_n38513__;
  assign new_new_n38597__ = ~new_new_n38434__ & new_new_n38509__;
  assign new_new_n38598__ = new_new_n38449__ & new_new_n38514__;
  assign new_new_n38599__ = ~new_new_n38517__ & ~new_new_n38598__;
  assign new_new_n38600__ = new_new_n38434__ & new_new_n38599__;
  assign new_new_n38601__ = ~new_new_n38596__ & ~new_new_n38600__;
  assign new_new_n38602__ = ~new_new_n38597__ & new_new_n38601__;
  assign new_new_n38603__ = ~new_new_n38594__ & ~new_new_n38602__;
  assign po31 = new_new_n38595__ | new_new_n38603__;
endmodule


