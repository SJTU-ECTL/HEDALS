// Benchmark "square" written by ABC on Wed Jul 13 18:49:40 2022

module square ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47,
    pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45,
    pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57,
    pi58, pi59, pi60, pi61, pi62, pi63;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127;
  wire new_new_n195__, new_new_n196__, new_new_n197__, new_new_n199__,
    new_new_n200__, new_new_n201__, new_new_n202__, new_new_n203__,
    new_new_n204__, new_new_n206__, new_new_n207__, new_new_n208__,
    new_new_n209__, new_new_n210__, new_new_n211__, new_new_n212__,
    new_new_n214__, new_new_n215__, new_new_n216__, new_new_n217__,
    new_new_n218__, new_new_n219__, new_new_n220__, new_new_n221__,
    new_new_n222__, new_new_n223__, new_new_n224__, new_new_n225__,
    new_new_n226__, new_new_n227__, new_new_n228__, new_new_n229__,
    new_new_n230__, new_new_n231__, new_new_n232__, new_new_n233__,
    new_new_n234__, new_new_n235__, new_new_n236__, new_new_n237__,
    new_new_n238__, new_new_n239__, new_new_n241__, new_new_n242__,
    new_new_n243__, new_new_n244__, new_new_n245__, new_new_n246__,
    new_new_n247__, new_new_n248__, new_new_n249__, new_new_n250__,
    new_new_n251__, new_new_n252__, new_new_n253__, new_new_n254__,
    new_new_n255__, new_new_n256__, new_new_n257__, new_new_n258__,
    new_new_n259__, new_new_n260__, new_new_n261__, new_new_n262__,
    new_new_n263__, new_new_n264__, new_new_n265__, new_new_n266__,
    new_new_n267__, new_new_n269__, new_new_n270__, new_new_n271__,
    new_new_n272__, new_new_n273__, new_new_n274__, new_new_n275__,
    new_new_n276__, new_new_n277__, new_new_n278__, new_new_n279__,
    new_new_n280__, new_new_n281__, new_new_n282__, new_new_n283__,
    new_new_n284__, new_new_n285__, new_new_n286__, new_new_n287__,
    new_new_n288__, new_new_n289__, new_new_n290__, new_new_n291__,
    new_new_n292__, new_new_n293__, new_new_n294__, new_new_n295__,
    new_new_n296__, new_new_n297__, new_new_n298__, new_new_n299__,
    new_new_n300__, new_new_n301__, new_new_n302__, new_new_n303__,
    new_new_n304__, new_new_n305__, new_new_n306__, new_new_n307__,
    new_new_n308__, new_new_n309__, new_new_n310__, new_new_n311__,
    new_new_n312__, new_new_n314__, new_new_n315__, new_new_n316__,
    new_new_n317__, new_new_n318__, new_new_n319__, new_new_n320__,
    new_new_n321__, new_new_n322__, new_new_n323__, new_new_n324__,
    new_new_n325__, new_new_n326__, new_new_n327__, new_new_n328__,
    new_new_n329__, new_new_n330__, new_new_n331__, new_new_n332__,
    new_new_n333__, new_new_n334__, new_new_n335__, new_new_n336__,
    new_new_n337__, new_new_n338__, new_new_n339__, new_new_n340__,
    new_new_n341__, new_new_n342__, new_new_n343__, new_new_n344__,
    new_new_n345__, new_new_n346__, new_new_n347__, new_new_n348__,
    new_new_n349__, new_new_n350__, new_new_n351__, new_new_n352__,
    new_new_n353__, new_new_n355__, new_new_n356__, new_new_n357__,
    new_new_n358__, new_new_n359__, new_new_n360__, new_new_n361__,
    new_new_n362__, new_new_n363__, new_new_n364__, new_new_n365__,
    new_new_n366__, new_new_n367__, new_new_n368__, new_new_n369__,
    new_new_n370__, new_new_n371__, new_new_n372__, new_new_n373__,
    new_new_n374__, new_new_n375__, new_new_n376__, new_new_n377__,
    new_new_n378__, new_new_n379__, new_new_n380__, new_new_n381__,
    new_new_n382__, new_new_n383__, new_new_n384__, new_new_n385__,
    new_new_n386__, new_new_n387__, new_new_n388__, new_new_n389__,
    new_new_n390__, new_new_n391__, new_new_n392__, new_new_n393__,
    new_new_n394__, new_new_n395__, new_new_n396__, new_new_n397__,
    new_new_n398__, new_new_n399__, new_new_n400__, new_new_n401__,
    new_new_n402__, new_new_n403__, new_new_n404__, new_new_n405__,
    new_new_n406__, new_new_n407__, new_new_n408__, new_new_n409__,
    new_new_n410__, new_new_n411__, new_new_n412__, new_new_n413__,
    new_new_n414__, new_new_n415__, new_new_n416__, new_new_n418__,
    new_new_n419__, new_new_n420__, new_new_n421__, new_new_n422__,
    new_new_n423__, new_new_n424__, new_new_n425__, new_new_n426__,
    new_new_n427__, new_new_n428__, new_new_n429__, new_new_n430__,
    new_new_n431__, new_new_n432__, new_new_n433__, new_new_n434__,
    new_new_n435__, new_new_n436__, new_new_n437__, new_new_n438__,
    new_new_n439__, new_new_n440__, new_new_n441__, new_new_n442__,
    new_new_n443__, new_new_n444__, new_new_n445__, new_new_n446__,
    new_new_n447__, new_new_n448__, new_new_n449__, new_new_n450__,
    new_new_n451__, new_new_n452__, new_new_n453__, new_new_n454__,
    new_new_n455__, new_new_n456__, new_new_n457__, new_new_n458__,
    new_new_n459__, new_new_n460__, new_new_n461__, new_new_n462__,
    new_new_n463__, new_new_n464__, new_new_n465__, new_new_n466__,
    new_new_n467__, new_new_n468__, new_new_n469__, new_new_n470__,
    new_new_n471__, new_new_n473__, new_new_n474__, new_new_n475__,
    new_new_n476__, new_new_n477__, new_new_n478__, new_new_n479__,
    new_new_n480__, new_new_n481__, new_new_n482__, new_new_n483__,
    new_new_n484__, new_new_n485__, new_new_n486__, new_new_n487__,
    new_new_n488__, new_new_n489__, new_new_n490__, new_new_n491__,
    new_new_n492__, new_new_n493__, new_new_n494__, new_new_n495__,
    new_new_n496__, new_new_n497__, new_new_n498__, new_new_n499__,
    new_new_n500__, new_new_n501__, new_new_n502__, new_new_n503__,
    new_new_n504__, new_new_n505__, new_new_n506__, new_new_n507__,
    new_new_n508__, new_new_n509__, new_new_n510__, new_new_n511__,
    new_new_n512__, new_new_n513__, new_new_n514__, new_new_n515__,
    new_new_n516__, new_new_n517__, new_new_n518__, new_new_n519__,
    new_new_n520__, new_new_n521__, new_new_n522__, new_new_n523__,
    new_new_n524__, new_new_n525__, new_new_n526__, new_new_n527__,
    new_new_n528__, new_new_n529__, new_new_n530__, new_new_n531__,
    new_new_n532__, new_new_n533__, new_new_n534__, new_new_n535__,
    new_new_n536__, new_new_n537__, new_new_n538__, new_new_n539__,
    new_new_n540__, new_new_n541__, new_new_n542__, new_new_n543__,
    new_new_n544__, new_new_n545__, new_new_n547__, new_new_n548__,
    new_new_n549__, new_new_n550__, new_new_n551__, new_new_n552__,
    new_new_n553__, new_new_n554__, new_new_n555__, new_new_n556__,
    new_new_n557__, new_new_n558__, new_new_n559__, new_new_n560__,
    new_new_n561__, new_new_n562__, new_new_n563__, new_new_n564__,
    new_new_n565__, new_new_n566__, new_new_n567__, new_new_n568__,
    new_new_n569__, new_new_n570__, new_new_n571__, new_new_n572__,
    new_new_n573__, new_new_n574__, new_new_n575__, new_new_n576__,
    new_new_n577__, new_new_n578__, new_new_n579__, new_new_n580__,
    new_new_n581__, new_new_n582__, new_new_n583__, new_new_n584__,
    new_new_n585__, new_new_n586__, new_new_n587__, new_new_n588__,
    new_new_n589__, new_new_n590__, new_new_n591__, new_new_n592__,
    new_new_n593__, new_new_n594__, new_new_n595__, new_new_n596__,
    new_new_n597__, new_new_n598__, new_new_n599__, new_new_n600__,
    new_new_n601__, new_new_n602__, new_new_n603__, new_new_n604__,
    new_new_n605__, new_new_n606__, new_new_n607__, new_new_n608__,
    new_new_n609__, new_new_n610__, new_new_n612__, new_new_n613__,
    new_new_n614__, new_new_n615__, new_new_n616__, new_new_n617__,
    new_new_n618__, new_new_n619__, new_new_n620__, new_new_n621__,
    new_new_n622__, new_new_n623__, new_new_n624__, new_new_n625__,
    new_new_n626__, new_new_n627__, new_new_n628__, new_new_n629__,
    new_new_n630__, new_new_n631__, new_new_n632__, new_new_n633__,
    new_new_n634__, new_new_n635__, new_new_n636__, new_new_n637__,
    new_new_n638__, new_new_n639__, new_new_n640__, new_new_n641__,
    new_new_n642__, new_new_n643__, new_new_n644__, new_new_n645__,
    new_new_n646__, new_new_n647__, new_new_n648__, new_new_n649__,
    new_new_n650__, new_new_n651__, new_new_n652__, new_new_n653__,
    new_new_n654__, new_new_n655__, new_new_n656__, new_new_n657__,
    new_new_n658__, new_new_n659__, new_new_n660__, new_new_n661__,
    new_new_n662__, new_new_n663__, new_new_n664__, new_new_n665__,
    new_new_n666__, new_new_n667__, new_new_n668__, new_new_n669__,
    new_new_n670__, new_new_n671__, new_new_n672__, new_new_n673__,
    new_new_n674__, new_new_n675__, new_new_n676__, new_new_n677__,
    new_new_n678__, new_new_n679__, new_new_n680__, new_new_n681__,
    new_new_n682__, new_new_n683__, new_new_n684__, new_new_n685__,
    new_new_n686__, new_new_n687__, new_new_n688__, new_new_n689__,
    new_new_n691__, new_new_n692__, new_new_n693__, new_new_n694__,
    new_new_n695__, new_new_n696__, new_new_n697__, new_new_n698__,
    new_new_n699__, new_new_n700__, new_new_n701__, new_new_n702__,
    new_new_n703__, new_new_n704__, new_new_n705__, new_new_n706__,
    new_new_n707__, new_new_n708__, new_new_n709__, new_new_n710__,
    new_new_n711__, new_new_n712__, new_new_n713__, new_new_n714__,
    new_new_n715__, new_new_n716__, new_new_n717__, new_new_n718__,
    new_new_n719__, new_new_n720__, new_new_n721__, new_new_n722__,
    new_new_n723__, new_new_n724__, new_new_n725__, new_new_n726__,
    new_new_n727__, new_new_n728__, new_new_n729__, new_new_n730__,
    new_new_n731__, new_new_n732__, new_new_n733__, new_new_n734__,
    new_new_n735__, new_new_n736__, new_new_n737__, new_new_n738__,
    new_new_n739__, new_new_n740__, new_new_n741__, new_new_n742__,
    new_new_n743__, new_new_n744__, new_new_n745__, new_new_n746__,
    new_new_n747__, new_new_n748__, new_new_n749__, new_new_n750__,
    new_new_n751__, new_new_n752__, new_new_n753__, new_new_n754__,
    new_new_n755__, new_new_n756__, new_new_n758__, new_new_n759__,
    new_new_n760__, new_new_n761__, new_new_n762__, new_new_n763__,
    new_new_n764__, new_new_n765__, new_new_n766__, new_new_n767__,
    new_new_n768__, new_new_n769__, new_new_n770__, new_new_n771__,
    new_new_n772__, new_new_n773__, new_new_n774__, new_new_n775__,
    new_new_n776__, new_new_n777__, new_new_n778__, new_new_n779__,
    new_new_n780__, new_new_n781__, new_new_n782__, new_new_n783__,
    new_new_n784__, new_new_n785__, new_new_n786__, new_new_n787__,
    new_new_n788__, new_new_n789__, new_new_n790__, new_new_n791__,
    new_new_n792__, new_new_n793__, new_new_n794__, new_new_n795__,
    new_new_n796__, new_new_n797__, new_new_n798__, new_new_n799__,
    new_new_n800__, new_new_n801__, new_new_n802__, new_new_n803__,
    new_new_n804__, new_new_n805__, new_new_n806__, new_new_n807__,
    new_new_n808__, new_new_n809__, new_new_n810__, new_new_n811__,
    new_new_n812__, new_new_n813__, new_new_n814__, new_new_n815__,
    new_new_n816__, new_new_n817__, new_new_n818__, new_new_n819__,
    new_new_n820__, new_new_n821__, new_new_n822__, new_new_n823__,
    new_new_n824__, new_new_n825__, new_new_n826__, new_new_n827__,
    new_new_n828__, new_new_n829__, new_new_n830__, new_new_n831__,
    new_new_n832__, new_new_n833__, new_new_n834__, new_new_n835__,
    new_new_n836__, new_new_n837__, new_new_n838__, new_new_n839__,
    new_new_n840__, new_new_n841__, new_new_n842__, new_new_n844__,
    new_new_n845__, new_new_n846__, new_new_n847__, new_new_n848__,
    new_new_n849__, new_new_n850__, new_new_n851__, new_new_n852__,
    new_new_n853__, new_new_n854__, new_new_n855__, new_new_n856__,
    new_new_n857__, new_new_n858__, new_new_n859__, new_new_n860__,
    new_new_n861__, new_new_n862__, new_new_n863__, new_new_n864__,
    new_new_n865__, new_new_n866__, new_new_n867__, new_new_n868__,
    new_new_n869__, new_new_n870__, new_new_n871__, new_new_n872__,
    new_new_n873__, new_new_n874__, new_new_n875__, new_new_n876__,
    new_new_n877__, new_new_n878__, new_new_n879__, new_new_n880__,
    new_new_n881__, new_new_n882__, new_new_n883__, new_new_n884__,
    new_new_n885__, new_new_n886__, new_new_n887__, new_new_n888__,
    new_new_n889__, new_new_n890__, new_new_n891__, new_new_n892__,
    new_new_n893__, new_new_n894__, new_new_n895__, new_new_n896__,
    new_new_n897__, new_new_n898__, new_new_n899__, new_new_n900__,
    new_new_n901__, new_new_n902__, new_new_n903__, new_new_n904__,
    new_new_n905__, new_new_n906__, new_new_n907__, new_new_n908__,
    new_new_n909__, new_new_n910__, new_new_n911__, new_new_n912__,
    new_new_n913__, new_new_n914__, new_new_n915__, new_new_n916__,
    new_new_n917__, new_new_n918__, new_new_n919__, new_new_n920__,
    new_new_n921__, new_new_n922__, new_new_n923__, new_new_n924__,
    new_new_n925__, new_new_n926__, new_new_n928__, new_new_n929__,
    new_new_n930__, new_new_n931__, new_new_n932__, new_new_n933__,
    new_new_n934__, new_new_n935__, new_new_n936__, new_new_n937__,
    new_new_n938__, new_new_n939__, new_new_n940__, new_new_n941__,
    new_new_n942__, new_new_n943__, new_new_n944__, new_new_n945__,
    new_new_n946__, new_new_n947__, new_new_n948__, new_new_n949__,
    new_new_n950__, new_new_n951__, new_new_n952__, new_new_n953__,
    new_new_n954__, new_new_n955__, new_new_n956__, new_new_n957__,
    new_new_n958__, new_new_n959__, new_new_n960__, new_new_n961__,
    new_new_n962__, new_new_n963__, new_new_n964__, new_new_n965__,
    new_new_n966__, new_new_n967__, new_new_n968__, new_new_n969__,
    new_new_n970__, new_new_n971__, new_new_n972__, new_new_n973__,
    new_new_n974__, new_new_n975__, new_new_n976__, new_new_n977__,
    new_new_n978__, new_new_n979__, new_new_n980__, new_new_n981__,
    new_new_n982__, new_new_n983__, new_new_n984__, new_new_n985__,
    new_new_n986__, new_new_n987__, new_new_n988__, new_new_n989__,
    new_new_n990__, new_new_n991__, new_new_n992__, new_new_n993__,
    new_new_n994__, new_new_n995__, new_new_n996__, new_new_n997__,
    new_new_n998__, new_new_n999__, new_new_n1000__, new_new_n1001__,
    new_new_n1002__, new_new_n1003__, new_new_n1004__, new_new_n1005__,
    new_new_n1006__, new_new_n1007__, new_new_n1008__, new_new_n1009__,
    new_new_n1010__, new_new_n1011__, new_new_n1012__, new_new_n1013__,
    new_new_n1014__, new_new_n1015__, new_new_n1016__, new_new_n1017__,
    new_new_n1018__, new_new_n1019__, new_new_n1020__, new_new_n1021__,
    new_new_n1022__, new_new_n1023__, new_new_n1024__, new_new_n1025__,
    new_new_n1026__, new_new_n1027__, new_new_n1028__, new_new_n1029__,
    new_new_n1030__, new_new_n1031__, new_new_n1032__, new_new_n1033__,
    new_new_n1034__, new_new_n1036__, new_new_n1037__, new_new_n1038__,
    new_new_n1039__, new_new_n1040__, new_new_n1041__, new_new_n1042__,
    new_new_n1043__, new_new_n1044__, new_new_n1045__, new_new_n1046__,
    new_new_n1047__, new_new_n1048__, new_new_n1049__, new_new_n1050__,
    new_new_n1051__, new_new_n1052__, new_new_n1053__, new_new_n1054__,
    new_new_n1055__, new_new_n1056__, new_new_n1057__, new_new_n1058__,
    new_new_n1059__, new_new_n1060__, new_new_n1061__, new_new_n1062__,
    new_new_n1063__, new_new_n1064__, new_new_n1065__, new_new_n1066__,
    new_new_n1067__, new_new_n1068__, new_new_n1069__, new_new_n1070__,
    new_new_n1071__, new_new_n1072__, new_new_n1073__, new_new_n1074__,
    new_new_n1075__, new_new_n1076__, new_new_n1077__, new_new_n1078__,
    new_new_n1079__, new_new_n1080__, new_new_n1081__, new_new_n1082__,
    new_new_n1083__, new_new_n1084__, new_new_n1085__, new_new_n1086__,
    new_new_n1087__, new_new_n1088__, new_new_n1089__, new_new_n1090__,
    new_new_n1091__, new_new_n1092__, new_new_n1093__, new_new_n1094__,
    new_new_n1095__, new_new_n1096__, new_new_n1097__, new_new_n1098__,
    new_new_n1099__, new_new_n1100__, new_new_n1101__, new_new_n1102__,
    new_new_n1103__, new_new_n1104__, new_new_n1105__, new_new_n1106__,
    new_new_n1107__, new_new_n1108__, new_new_n1109__, new_new_n1110__,
    new_new_n1111__, new_new_n1112__, new_new_n1113__, new_new_n1114__,
    new_new_n1115__, new_new_n1117__, new_new_n1118__, new_new_n1119__,
    new_new_n1120__, new_new_n1121__, new_new_n1122__, new_new_n1123__,
    new_new_n1124__, new_new_n1125__, new_new_n1126__, new_new_n1127__,
    new_new_n1128__, new_new_n1129__, new_new_n1130__, new_new_n1131__,
    new_new_n1132__, new_new_n1133__, new_new_n1134__, new_new_n1135__,
    new_new_n1136__, new_new_n1137__, new_new_n1138__, new_new_n1139__,
    new_new_n1140__, new_new_n1141__, new_new_n1142__, new_new_n1143__,
    new_new_n1144__, new_new_n1145__, new_new_n1146__, new_new_n1147__,
    new_new_n1148__, new_new_n1149__, new_new_n1150__, new_new_n1151__,
    new_new_n1152__, new_new_n1153__, new_new_n1154__, new_new_n1155__,
    new_new_n1156__, new_new_n1157__, new_new_n1158__, new_new_n1159__,
    new_new_n1160__, new_new_n1161__, new_new_n1162__, new_new_n1163__,
    new_new_n1164__, new_new_n1165__, new_new_n1166__, new_new_n1167__,
    new_new_n1168__, new_new_n1169__, new_new_n1170__, new_new_n1171__,
    new_new_n1172__, new_new_n1173__, new_new_n1174__, new_new_n1175__,
    new_new_n1176__, new_new_n1177__, new_new_n1178__, new_new_n1179__,
    new_new_n1180__, new_new_n1181__, new_new_n1182__, new_new_n1183__,
    new_new_n1184__, new_new_n1185__, new_new_n1186__, new_new_n1187__,
    new_new_n1188__, new_new_n1189__, new_new_n1190__, new_new_n1191__,
    new_new_n1192__, new_new_n1193__, new_new_n1194__, new_new_n1195__,
    new_new_n1196__, new_new_n1197__, new_new_n1198__, new_new_n1199__,
    new_new_n1200__, new_new_n1201__, new_new_n1202__, new_new_n1203__,
    new_new_n1204__, new_new_n1205__, new_new_n1206__, new_new_n1207__,
    new_new_n1208__, new_new_n1209__, new_new_n1210__, new_new_n1211__,
    new_new_n1212__, new_new_n1213__, new_new_n1214__, new_new_n1215__,
    new_new_n1216__, new_new_n1217__, new_new_n1218__, new_new_n1219__,
    new_new_n1220__, new_new_n1222__, new_new_n1223__, new_new_n1224__,
    new_new_n1225__, new_new_n1226__, new_new_n1227__, new_new_n1228__,
    new_new_n1229__, new_new_n1230__, new_new_n1231__, new_new_n1232__,
    new_new_n1233__, new_new_n1234__, new_new_n1235__, new_new_n1236__,
    new_new_n1237__, new_new_n1238__, new_new_n1239__, new_new_n1240__,
    new_new_n1241__, new_new_n1242__, new_new_n1243__, new_new_n1244__,
    new_new_n1245__, new_new_n1246__, new_new_n1247__, new_new_n1248__,
    new_new_n1249__, new_new_n1250__, new_new_n1251__, new_new_n1252__,
    new_new_n1253__, new_new_n1254__, new_new_n1255__, new_new_n1256__,
    new_new_n1257__, new_new_n1258__, new_new_n1259__, new_new_n1260__,
    new_new_n1261__, new_new_n1262__, new_new_n1263__, new_new_n1264__,
    new_new_n1265__, new_new_n1266__, new_new_n1267__, new_new_n1268__,
    new_new_n1269__, new_new_n1270__, new_new_n1271__, new_new_n1272__,
    new_new_n1273__, new_new_n1274__, new_new_n1275__, new_new_n1276__,
    new_new_n1277__, new_new_n1278__, new_new_n1279__, new_new_n1280__,
    new_new_n1281__, new_new_n1282__, new_new_n1283__, new_new_n1284__,
    new_new_n1285__, new_new_n1286__, new_new_n1287__, new_new_n1288__,
    new_new_n1289__, new_new_n1290__, new_new_n1291__, new_new_n1292__,
    new_new_n1293__, new_new_n1294__, new_new_n1295__, new_new_n1296__,
    new_new_n1297__, new_new_n1298__, new_new_n1299__, new_new_n1300__,
    new_new_n1301__, new_new_n1302__, new_new_n1303__, new_new_n1304__,
    new_new_n1305__, new_new_n1306__, new_new_n1307__, new_new_n1308__,
    new_new_n1309__, new_new_n1310__, new_new_n1311__, new_new_n1312__,
    new_new_n1313__, new_new_n1314__, new_new_n1315__, new_new_n1316__,
    new_new_n1318__, new_new_n1319__, new_new_n1320__, new_new_n1321__,
    new_new_n1322__, new_new_n1323__, new_new_n1324__, new_new_n1325__,
    new_new_n1326__, new_new_n1327__, new_new_n1328__, new_new_n1329__,
    new_new_n1330__, new_new_n1331__, new_new_n1332__, new_new_n1333__,
    new_new_n1334__, new_new_n1335__, new_new_n1336__, new_new_n1337__,
    new_new_n1338__, new_new_n1339__, new_new_n1340__, new_new_n1341__,
    new_new_n1342__, new_new_n1343__, new_new_n1344__, new_new_n1345__,
    new_new_n1346__, new_new_n1347__, new_new_n1348__, new_new_n1349__,
    new_new_n1350__, new_new_n1351__, new_new_n1352__, new_new_n1353__,
    new_new_n1354__, new_new_n1355__, new_new_n1356__, new_new_n1357__,
    new_new_n1358__, new_new_n1359__, new_new_n1360__, new_new_n1361__,
    new_new_n1362__, new_new_n1363__, new_new_n1364__, new_new_n1365__,
    new_new_n1366__, new_new_n1367__, new_new_n1368__, new_new_n1369__,
    new_new_n1370__, new_new_n1371__, new_new_n1372__, new_new_n1373__,
    new_new_n1374__, new_new_n1375__, new_new_n1376__, new_new_n1377__,
    new_new_n1378__, new_new_n1379__, new_new_n1380__, new_new_n1381__,
    new_new_n1382__, new_new_n1383__, new_new_n1384__, new_new_n1385__,
    new_new_n1386__, new_new_n1387__, new_new_n1388__, new_new_n1389__,
    new_new_n1390__, new_new_n1391__, new_new_n1392__, new_new_n1393__,
    new_new_n1394__, new_new_n1395__, new_new_n1396__, new_new_n1397__,
    new_new_n1398__, new_new_n1399__, new_new_n1400__, new_new_n1401__,
    new_new_n1402__, new_new_n1403__, new_new_n1404__, new_new_n1405__,
    new_new_n1406__, new_new_n1407__, new_new_n1408__, new_new_n1409__,
    new_new_n1410__, new_new_n1411__, new_new_n1412__, new_new_n1413__,
    new_new_n1414__, new_new_n1415__, new_new_n1416__, new_new_n1417__,
    new_new_n1418__, new_new_n1419__, new_new_n1420__, new_new_n1421__,
    new_new_n1422__, new_new_n1423__, new_new_n1424__, new_new_n1425__,
    new_new_n1426__, new_new_n1427__, new_new_n1428__, new_new_n1429__,
    new_new_n1430__, new_new_n1431__, new_new_n1432__, new_new_n1433__,
    new_new_n1435__, new_new_n1436__, new_new_n1437__, new_new_n1438__,
    new_new_n1439__, new_new_n1440__, new_new_n1441__, new_new_n1442__,
    new_new_n1443__, new_new_n1444__, new_new_n1445__, new_new_n1446__,
    new_new_n1447__, new_new_n1448__, new_new_n1449__, new_new_n1450__,
    new_new_n1451__, new_new_n1452__, new_new_n1453__, new_new_n1454__,
    new_new_n1455__, new_new_n1456__, new_new_n1457__, new_new_n1458__,
    new_new_n1459__, new_new_n1460__, new_new_n1461__, new_new_n1462__,
    new_new_n1463__, new_new_n1464__, new_new_n1465__, new_new_n1466__,
    new_new_n1467__, new_new_n1468__, new_new_n1469__, new_new_n1470__,
    new_new_n1471__, new_new_n1472__, new_new_n1473__, new_new_n1474__,
    new_new_n1475__, new_new_n1476__, new_new_n1477__, new_new_n1478__,
    new_new_n1479__, new_new_n1480__, new_new_n1481__, new_new_n1482__,
    new_new_n1483__, new_new_n1484__, new_new_n1485__, new_new_n1486__,
    new_new_n1487__, new_new_n1488__, new_new_n1489__, new_new_n1490__,
    new_new_n1491__, new_new_n1492__, new_new_n1493__, new_new_n1494__,
    new_new_n1495__, new_new_n1496__, new_new_n1497__, new_new_n1498__,
    new_new_n1499__, new_new_n1500__, new_new_n1501__, new_new_n1502__,
    new_new_n1503__, new_new_n1504__, new_new_n1505__, new_new_n1506__,
    new_new_n1507__, new_new_n1508__, new_new_n1509__, new_new_n1510__,
    new_new_n1511__, new_new_n1512__, new_new_n1513__, new_new_n1514__,
    new_new_n1515__, new_new_n1516__, new_new_n1517__, new_new_n1518__,
    new_new_n1519__, new_new_n1520__, new_new_n1521__, new_new_n1522__,
    new_new_n1523__, new_new_n1524__, new_new_n1525__, new_new_n1526__,
    new_new_n1527__, new_new_n1528__, new_new_n1529__, new_new_n1530__,
    new_new_n1531__, new_new_n1532__, new_new_n1533__, new_new_n1535__,
    new_new_n1536__, new_new_n1537__, new_new_n1538__, new_new_n1539__,
    new_new_n1540__, new_new_n1541__, new_new_n1542__, new_new_n1543__,
    new_new_n1544__, new_new_n1545__, new_new_n1546__, new_new_n1547__,
    new_new_n1548__, new_new_n1549__, new_new_n1550__, new_new_n1551__,
    new_new_n1552__, new_new_n1553__, new_new_n1554__, new_new_n1555__,
    new_new_n1556__, new_new_n1557__, new_new_n1558__, new_new_n1559__,
    new_new_n1560__, new_new_n1561__, new_new_n1562__, new_new_n1563__,
    new_new_n1564__, new_new_n1565__, new_new_n1566__, new_new_n1567__,
    new_new_n1568__, new_new_n1569__, new_new_n1570__, new_new_n1571__,
    new_new_n1572__, new_new_n1573__, new_new_n1574__, new_new_n1575__,
    new_new_n1576__, new_new_n1577__, new_new_n1578__, new_new_n1579__,
    new_new_n1580__, new_new_n1581__, new_new_n1582__, new_new_n1583__,
    new_new_n1584__, new_new_n1585__, new_new_n1586__, new_new_n1587__,
    new_new_n1588__, new_new_n1589__, new_new_n1590__, new_new_n1591__,
    new_new_n1592__, new_new_n1593__, new_new_n1594__, new_new_n1595__,
    new_new_n1596__, new_new_n1597__, new_new_n1598__, new_new_n1599__,
    new_new_n1600__, new_new_n1601__, new_new_n1602__, new_new_n1603__,
    new_new_n1604__, new_new_n1605__, new_new_n1606__, new_new_n1607__,
    new_new_n1608__, new_new_n1609__, new_new_n1610__, new_new_n1611__,
    new_new_n1612__, new_new_n1613__, new_new_n1614__, new_new_n1615__,
    new_new_n1616__, new_new_n1617__, new_new_n1618__, new_new_n1619__,
    new_new_n1620__, new_new_n1621__, new_new_n1622__, new_new_n1623__,
    new_new_n1624__, new_new_n1625__, new_new_n1626__, new_new_n1627__,
    new_new_n1628__, new_new_n1629__, new_new_n1630__, new_new_n1631__,
    new_new_n1632__, new_new_n1633__, new_new_n1634__, new_new_n1635__,
    new_new_n1636__, new_new_n1637__, new_new_n1638__, new_new_n1639__,
    new_new_n1640__, new_new_n1641__, new_new_n1642__, new_new_n1643__,
    new_new_n1644__, new_new_n1645__, new_new_n1647__, new_new_n1648__,
    new_new_n1649__, new_new_n1650__, new_new_n1651__, new_new_n1652__,
    new_new_n1653__, new_new_n1654__, new_new_n1655__, new_new_n1656__,
    new_new_n1657__, new_new_n1658__, new_new_n1659__, new_new_n1660__,
    new_new_n1661__, new_new_n1662__, new_new_n1663__, new_new_n1664__,
    new_new_n1665__, new_new_n1666__, new_new_n1667__, new_new_n1668__,
    new_new_n1669__, new_new_n1670__, new_new_n1671__, new_new_n1672__,
    new_new_n1673__, new_new_n1674__, new_new_n1675__, new_new_n1676__,
    new_new_n1677__, new_new_n1678__, new_new_n1679__, new_new_n1680__,
    new_new_n1681__, new_new_n1682__, new_new_n1683__, new_new_n1684__,
    new_new_n1685__, new_new_n1686__, new_new_n1687__, new_new_n1688__,
    new_new_n1689__, new_new_n1690__, new_new_n1691__, new_new_n1692__,
    new_new_n1693__, new_new_n1694__, new_new_n1695__, new_new_n1696__,
    new_new_n1697__, new_new_n1698__, new_new_n1699__, new_new_n1700__,
    new_new_n1701__, new_new_n1702__, new_new_n1703__, new_new_n1704__,
    new_new_n1705__, new_new_n1706__, new_new_n1707__, new_new_n1708__,
    new_new_n1709__, new_new_n1710__, new_new_n1711__, new_new_n1712__,
    new_new_n1713__, new_new_n1714__, new_new_n1715__, new_new_n1716__,
    new_new_n1717__, new_new_n1718__, new_new_n1719__, new_new_n1720__,
    new_new_n1721__, new_new_n1722__, new_new_n1723__, new_new_n1724__,
    new_new_n1725__, new_new_n1726__, new_new_n1727__, new_new_n1728__,
    new_new_n1729__, new_new_n1730__, new_new_n1731__, new_new_n1732__,
    new_new_n1733__, new_new_n1734__, new_new_n1735__, new_new_n1736__,
    new_new_n1737__, new_new_n1738__, new_new_n1739__, new_new_n1740__,
    new_new_n1741__, new_new_n1742__, new_new_n1743__, new_new_n1744__,
    new_new_n1745__, new_new_n1746__, new_new_n1747__, new_new_n1748__,
    new_new_n1749__, new_new_n1750__, new_new_n1751__, new_new_n1752__,
    new_new_n1753__, new_new_n1754__, new_new_n1755__, new_new_n1756__,
    new_new_n1757__, new_new_n1758__, new_new_n1759__, new_new_n1760__,
    new_new_n1761__, new_new_n1762__, new_new_n1763__, new_new_n1764__,
    new_new_n1765__, new_new_n1766__, new_new_n1767__, new_new_n1768__,
    new_new_n1769__, new_new_n1770__, new_new_n1771__, new_new_n1772__,
    new_new_n1773__, new_new_n1774__, new_new_n1776__, new_new_n1777__,
    new_new_n1778__, new_new_n1779__, new_new_n1780__, new_new_n1781__,
    new_new_n1782__, new_new_n1783__, new_new_n1784__, new_new_n1785__,
    new_new_n1786__, new_new_n1787__, new_new_n1788__, new_new_n1789__,
    new_new_n1790__, new_new_n1791__, new_new_n1792__, new_new_n1793__,
    new_new_n1794__, new_new_n1795__, new_new_n1796__, new_new_n1797__,
    new_new_n1798__, new_new_n1799__, new_new_n1800__, new_new_n1801__,
    new_new_n1802__, new_new_n1803__, new_new_n1804__, new_new_n1805__,
    new_new_n1806__, new_new_n1807__, new_new_n1808__, new_new_n1809__,
    new_new_n1810__, new_new_n1811__, new_new_n1812__, new_new_n1813__,
    new_new_n1814__, new_new_n1815__, new_new_n1816__, new_new_n1817__,
    new_new_n1818__, new_new_n1819__, new_new_n1820__, new_new_n1821__,
    new_new_n1822__, new_new_n1823__, new_new_n1824__, new_new_n1825__,
    new_new_n1826__, new_new_n1827__, new_new_n1828__, new_new_n1829__,
    new_new_n1830__, new_new_n1831__, new_new_n1832__, new_new_n1833__,
    new_new_n1834__, new_new_n1835__, new_new_n1836__, new_new_n1837__,
    new_new_n1838__, new_new_n1839__, new_new_n1840__, new_new_n1841__,
    new_new_n1842__, new_new_n1843__, new_new_n1844__, new_new_n1845__,
    new_new_n1846__, new_new_n1847__, new_new_n1848__, new_new_n1849__,
    new_new_n1850__, new_new_n1851__, new_new_n1852__, new_new_n1853__,
    new_new_n1854__, new_new_n1855__, new_new_n1856__, new_new_n1857__,
    new_new_n1858__, new_new_n1859__, new_new_n1860__, new_new_n1861__,
    new_new_n1862__, new_new_n1863__, new_new_n1864__, new_new_n1865__,
    new_new_n1866__, new_new_n1867__, new_new_n1868__, new_new_n1869__,
    new_new_n1870__, new_new_n1871__, new_new_n1872__, new_new_n1873__,
    new_new_n1874__, new_new_n1875__, new_new_n1876__, new_new_n1877__,
    new_new_n1878__, new_new_n1879__, new_new_n1880__, new_new_n1881__,
    new_new_n1882__, new_new_n1883__, new_new_n1884__, new_new_n1885__,
    new_new_n1886__, new_new_n1887__, new_new_n1888__, new_new_n1889__,
    new_new_n1890__, new_new_n1891__, new_new_n1892__, new_new_n1893__,
    new_new_n1894__, new_new_n1895__, new_new_n1897__, new_new_n1898__,
    new_new_n1899__, new_new_n1900__, new_new_n1901__, new_new_n1902__,
    new_new_n1903__, new_new_n1904__, new_new_n1905__, new_new_n1906__,
    new_new_n1907__, new_new_n1908__, new_new_n1909__, new_new_n1910__,
    new_new_n1911__, new_new_n1912__, new_new_n1913__, new_new_n1914__,
    new_new_n1915__, new_new_n1916__, new_new_n1917__, new_new_n1918__,
    new_new_n1919__, new_new_n1920__, new_new_n1921__, new_new_n1922__,
    new_new_n1923__, new_new_n1924__, new_new_n1925__, new_new_n1926__,
    new_new_n1927__, new_new_n1928__, new_new_n1929__, new_new_n1930__,
    new_new_n1931__, new_new_n1932__, new_new_n1933__, new_new_n1934__,
    new_new_n1935__, new_new_n1936__, new_new_n1937__, new_new_n1938__,
    new_new_n1939__, new_new_n1940__, new_new_n1941__, new_new_n1942__,
    new_new_n1943__, new_new_n1944__, new_new_n1945__, new_new_n1946__,
    new_new_n1947__, new_new_n1948__, new_new_n1949__, new_new_n1950__,
    new_new_n1951__, new_new_n1952__, new_new_n1953__, new_new_n1954__,
    new_new_n1955__, new_new_n1956__, new_new_n1957__, new_new_n1958__,
    new_new_n1959__, new_new_n1960__, new_new_n1961__, new_new_n1962__,
    new_new_n1963__, new_new_n1964__, new_new_n1965__, new_new_n1966__,
    new_new_n1967__, new_new_n1968__, new_new_n1969__, new_new_n1970__,
    new_new_n1971__, new_new_n1972__, new_new_n1973__, new_new_n1974__,
    new_new_n1975__, new_new_n1976__, new_new_n1977__, new_new_n1978__,
    new_new_n1979__, new_new_n1980__, new_new_n1981__, new_new_n1982__,
    new_new_n1983__, new_new_n1984__, new_new_n1985__, new_new_n1986__,
    new_new_n1987__, new_new_n1988__, new_new_n1989__, new_new_n1990__,
    new_new_n1991__, new_new_n1992__, new_new_n1993__, new_new_n1994__,
    new_new_n1995__, new_new_n1996__, new_new_n1997__, new_new_n1998__,
    new_new_n1999__, new_new_n2000__, new_new_n2001__, new_new_n2002__,
    new_new_n2003__, new_new_n2004__, new_new_n2005__, new_new_n2006__,
    new_new_n2007__, new_new_n2008__, new_new_n2009__, new_new_n2010__,
    new_new_n2011__, new_new_n2012__, new_new_n2013__, new_new_n2014__,
    new_new_n2015__, new_new_n2016__, new_new_n2017__, new_new_n2018__,
    new_new_n2019__, new_new_n2020__, new_new_n2021__, new_new_n2022__,
    new_new_n2023__, new_new_n2024__, new_new_n2025__, new_new_n2026__,
    new_new_n2027__, new_new_n2028__, new_new_n2029__, new_new_n2030__,
    new_new_n2031__, new_new_n2033__, new_new_n2034__, new_new_n2035__,
    new_new_n2036__, new_new_n2037__, new_new_n2038__, new_new_n2039__,
    new_new_n2040__, new_new_n2041__, new_new_n2042__, new_new_n2043__,
    new_new_n2044__, new_new_n2045__, new_new_n2046__, new_new_n2047__,
    new_new_n2048__, new_new_n2049__, new_new_n2050__, new_new_n2051__,
    new_new_n2052__, new_new_n2053__, new_new_n2054__, new_new_n2055__,
    new_new_n2056__, new_new_n2057__, new_new_n2058__, new_new_n2059__,
    new_new_n2060__, new_new_n2061__, new_new_n2062__, new_new_n2063__,
    new_new_n2064__, new_new_n2065__, new_new_n2066__, new_new_n2067__,
    new_new_n2068__, new_new_n2069__, new_new_n2070__, new_new_n2071__,
    new_new_n2072__, new_new_n2073__, new_new_n2074__, new_new_n2075__,
    new_new_n2076__, new_new_n2077__, new_new_n2078__, new_new_n2079__,
    new_new_n2080__, new_new_n2081__, new_new_n2082__, new_new_n2083__,
    new_new_n2084__, new_new_n2085__, new_new_n2086__, new_new_n2087__,
    new_new_n2088__, new_new_n2089__, new_new_n2090__, new_new_n2091__,
    new_new_n2092__, new_new_n2093__, new_new_n2094__, new_new_n2095__,
    new_new_n2096__, new_new_n2097__, new_new_n2098__, new_new_n2099__,
    new_new_n2100__, new_new_n2101__, new_new_n2102__, new_new_n2103__,
    new_new_n2104__, new_new_n2105__, new_new_n2106__, new_new_n2107__,
    new_new_n2108__, new_new_n2109__, new_new_n2110__, new_new_n2111__,
    new_new_n2112__, new_new_n2113__, new_new_n2114__, new_new_n2115__,
    new_new_n2116__, new_new_n2117__, new_new_n2118__, new_new_n2119__,
    new_new_n2120__, new_new_n2121__, new_new_n2122__, new_new_n2123__,
    new_new_n2124__, new_new_n2125__, new_new_n2126__, new_new_n2127__,
    new_new_n2128__, new_new_n2129__, new_new_n2130__, new_new_n2131__,
    new_new_n2132__, new_new_n2133__, new_new_n2134__, new_new_n2135__,
    new_new_n2136__, new_new_n2137__, new_new_n2138__, new_new_n2139__,
    new_new_n2140__, new_new_n2141__, new_new_n2142__, new_new_n2143__,
    new_new_n2144__, new_new_n2145__, new_new_n2146__, new_new_n2147__,
    new_new_n2148__, new_new_n2149__, new_new_n2150__, new_new_n2151__,
    new_new_n2152__, new_new_n2153__, new_new_n2154__, new_new_n2155__,
    new_new_n2156__, new_new_n2157__, new_new_n2158__, new_new_n2159__,
    new_new_n2160__, new_new_n2161__, new_new_n2162__, new_new_n2163__,
    new_new_n2164__, new_new_n2165__, new_new_n2166__, new_new_n2167__,
    new_new_n2169__, new_new_n2170__, new_new_n2171__, new_new_n2172__,
    new_new_n2173__, new_new_n2174__, new_new_n2175__, new_new_n2176__,
    new_new_n2177__, new_new_n2178__, new_new_n2179__, new_new_n2180__,
    new_new_n2181__, new_new_n2182__, new_new_n2183__, new_new_n2184__,
    new_new_n2185__, new_new_n2186__, new_new_n2187__, new_new_n2188__,
    new_new_n2189__, new_new_n2190__, new_new_n2191__, new_new_n2192__,
    new_new_n2193__, new_new_n2194__, new_new_n2195__, new_new_n2196__,
    new_new_n2197__, new_new_n2198__, new_new_n2199__, new_new_n2200__,
    new_new_n2201__, new_new_n2202__, new_new_n2203__, new_new_n2204__,
    new_new_n2205__, new_new_n2206__, new_new_n2207__, new_new_n2208__,
    new_new_n2209__, new_new_n2210__, new_new_n2211__, new_new_n2212__,
    new_new_n2213__, new_new_n2214__, new_new_n2215__, new_new_n2216__,
    new_new_n2217__, new_new_n2218__, new_new_n2219__, new_new_n2220__,
    new_new_n2221__, new_new_n2222__, new_new_n2223__, new_new_n2224__,
    new_new_n2225__, new_new_n2226__, new_new_n2227__, new_new_n2228__,
    new_new_n2229__, new_new_n2230__, new_new_n2231__, new_new_n2232__,
    new_new_n2233__, new_new_n2234__, new_new_n2235__, new_new_n2236__,
    new_new_n2237__, new_new_n2238__, new_new_n2239__, new_new_n2240__,
    new_new_n2241__, new_new_n2242__, new_new_n2243__, new_new_n2244__,
    new_new_n2245__, new_new_n2246__, new_new_n2247__, new_new_n2248__,
    new_new_n2249__, new_new_n2250__, new_new_n2251__, new_new_n2252__,
    new_new_n2253__, new_new_n2254__, new_new_n2255__, new_new_n2256__,
    new_new_n2257__, new_new_n2258__, new_new_n2259__, new_new_n2260__,
    new_new_n2261__, new_new_n2262__, new_new_n2263__, new_new_n2264__,
    new_new_n2265__, new_new_n2266__, new_new_n2267__, new_new_n2268__,
    new_new_n2269__, new_new_n2270__, new_new_n2271__, new_new_n2272__,
    new_new_n2273__, new_new_n2274__, new_new_n2275__, new_new_n2276__,
    new_new_n2277__, new_new_n2278__, new_new_n2279__, new_new_n2280__,
    new_new_n2281__, new_new_n2282__, new_new_n2283__, new_new_n2284__,
    new_new_n2285__, new_new_n2286__, new_new_n2287__, new_new_n2288__,
    new_new_n2289__, new_new_n2290__, new_new_n2291__, new_new_n2292__,
    new_new_n2293__, new_new_n2294__, new_new_n2295__, new_new_n2296__,
    new_new_n2297__, new_new_n2298__, new_new_n2299__, new_new_n2300__,
    new_new_n2301__, new_new_n2302__, new_new_n2303__, new_new_n2304__,
    new_new_n2305__, new_new_n2306__, new_new_n2307__, new_new_n2308__,
    new_new_n2309__, new_new_n2310__, new_new_n2311__, new_new_n2312__,
    new_new_n2313__, new_new_n2314__, new_new_n2315__, new_new_n2316__,
    new_new_n2317__, new_new_n2319__, new_new_n2320__, new_new_n2321__,
    new_new_n2322__, new_new_n2323__, new_new_n2324__, new_new_n2325__,
    new_new_n2326__, new_new_n2327__, new_new_n2328__, new_new_n2329__,
    new_new_n2330__, new_new_n2331__, new_new_n2332__, new_new_n2333__,
    new_new_n2334__, new_new_n2335__, new_new_n2336__, new_new_n2337__,
    new_new_n2338__, new_new_n2339__, new_new_n2340__, new_new_n2341__,
    new_new_n2342__, new_new_n2343__, new_new_n2344__, new_new_n2345__,
    new_new_n2346__, new_new_n2347__, new_new_n2348__, new_new_n2349__,
    new_new_n2350__, new_new_n2351__, new_new_n2352__, new_new_n2353__,
    new_new_n2354__, new_new_n2355__, new_new_n2356__, new_new_n2357__,
    new_new_n2358__, new_new_n2359__, new_new_n2360__, new_new_n2361__,
    new_new_n2362__, new_new_n2363__, new_new_n2364__, new_new_n2365__,
    new_new_n2366__, new_new_n2367__, new_new_n2368__, new_new_n2369__,
    new_new_n2370__, new_new_n2371__, new_new_n2372__, new_new_n2373__,
    new_new_n2374__, new_new_n2375__, new_new_n2376__, new_new_n2377__,
    new_new_n2378__, new_new_n2379__, new_new_n2380__, new_new_n2381__,
    new_new_n2382__, new_new_n2383__, new_new_n2384__, new_new_n2385__,
    new_new_n2386__, new_new_n2387__, new_new_n2388__, new_new_n2389__,
    new_new_n2390__, new_new_n2391__, new_new_n2392__, new_new_n2393__,
    new_new_n2394__, new_new_n2395__, new_new_n2396__, new_new_n2397__,
    new_new_n2398__, new_new_n2399__, new_new_n2400__, new_new_n2401__,
    new_new_n2402__, new_new_n2403__, new_new_n2404__, new_new_n2405__,
    new_new_n2406__, new_new_n2407__, new_new_n2408__, new_new_n2409__,
    new_new_n2410__, new_new_n2411__, new_new_n2412__, new_new_n2413__,
    new_new_n2414__, new_new_n2415__, new_new_n2416__, new_new_n2417__,
    new_new_n2418__, new_new_n2419__, new_new_n2420__, new_new_n2421__,
    new_new_n2422__, new_new_n2423__, new_new_n2424__, new_new_n2425__,
    new_new_n2426__, new_new_n2427__, new_new_n2428__, new_new_n2429__,
    new_new_n2430__, new_new_n2431__, new_new_n2432__, new_new_n2433__,
    new_new_n2434__, new_new_n2435__, new_new_n2436__, new_new_n2437__,
    new_new_n2438__, new_new_n2439__, new_new_n2440__, new_new_n2441__,
    new_new_n2442__, new_new_n2443__, new_new_n2444__, new_new_n2445__,
    new_new_n2446__, new_new_n2447__, new_new_n2448__, new_new_n2449__,
    new_new_n2450__, new_new_n2451__, new_new_n2452__, new_new_n2453__,
    new_new_n2454__, new_new_n2455__, new_new_n2456__, new_new_n2457__,
    new_new_n2458__, new_new_n2459__, new_new_n2460__, new_new_n2461__,
    new_new_n2463__, new_new_n2464__, new_new_n2465__, new_new_n2466__,
    new_new_n2467__, new_new_n2468__, new_new_n2469__, new_new_n2470__,
    new_new_n2471__, new_new_n2472__, new_new_n2473__, new_new_n2474__,
    new_new_n2475__, new_new_n2476__, new_new_n2477__, new_new_n2478__,
    new_new_n2479__, new_new_n2480__, new_new_n2481__, new_new_n2482__,
    new_new_n2483__, new_new_n2484__, new_new_n2485__, new_new_n2486__,
    new_new_n2487__, new_new_n2488__, new_new_n2489__, new_new_n2490__,
    new_new_n2491__, new_new_n2492__, new_new_n2493__, new_new_n2494__,
    new_new_n2495__, new_new_n2496__, new_new_n2497__, new_new_n2498__,
    new_new_n2499__, new_new_n2500__, new_new_n2501__, new_new_n2502__,
    new_new_n2503__, new_new_n2504__, new_new_n2505__, new_new_n2506__,
    new_new_n2507__, new_new_n2508__, new_new_n2509__, new_new_n2510__,
    new_new_n2511__, new_new_n2512__, new_new_n2513__, new_new_n2514__,
    new_new_n2515__, new_new_n2516__, new_new_n2517__, new_new_n2518__,
    new_new_n2519__, new_new_n2520__, new_new_n2521__, new_new_n2522__,
    new_new_n2523__, new_new_n2524__, new_new_n2525__, new_new_n2526__,
    new_new_n2527__, new_new_n2528__, new_new_n2529__, new_new_n2530__,
    new_new_n2531__, new_new_n2532__, new_new_n2533__, new_new_n2534__,
    new_new_n2535__, new_new_n2536__, new_new_n2537__, new_new_n2538__,
    new_new_n2539__, new_new_n2540__, new_new_n2541__, new_new_n2542__,
    new_new_n2543__, new_new_n2544__, new_new_n2545__, new_new_n2546__,
    new_new_n2547__, new_new_n2548__, new_new_n2549__, new_new_n2550__,
    new_new_n2551__, new_new_n2552__, new_new_n2553__, new_new_n2554__,
    new_new_n2555__, new_new_n2556__, new_new_n2557__, new_new_n2558__,
    new_new_n2559__, new_new_n2560__, new_new_n2561__, new_new_n2562__,
    new_new_n2563__, new_new_n2564__, new_new_n2565__, new_new_n2566__,
    new_new_n2567__, new_new_n2568__, new_new_n2569__, new_new_n2570__,
    new_new_n2571__, new_new_n2572__, new_new_n2573__, new_new_n2574__,
    new_new_n2575__, new_new_n2576__, new_new_n2577__, new_new_n2578__,
    new_new_n2579__, new_new_n2580__, new_new_n2581__, new_new_n2582__,
    new_new_n2583__, new_new_n2584__, new_new_n2585__, new_new_n2586__,
    new_new_n2587__, new_new_n2588__, new_new_n2589__, new_new_n2590__,
    new_new_n2591__, new_new_n2592__, new_new_n2593__, new_new_n2594__,
    new_new_n2595__, new_new_n2596__, new_new_n2597__, new_new_n2598__,
    new_new_n2599__, new_new_n2600__, new_new_n2601__, new_new_n2602__,
    new_new_n2603__, new_new_n2604__, new_new_n2605__, new_new_n2606__,
    new_new_n2607__, new_new_n2608__, new_new_n2609__, new_new_n2610__,
    new_new_n2611__, new_new_n2612__, new_new_n2613__, new_new_n2614__,
    new_new_n2615__, new_new_n2616__, new_new_n2617__, new_new_n2618__,
    new_new_n2619__, new_new_n2621__, new_new_n2622__, new_new_n2623__,
    new_new_n2624__, new_new_n2625__, new_new_n2626__, new_new_n2627__,
    new_new_n2628__, new_new_n2629__, new_new_n2630__, new_new_n2631__,
    new_new_n2632__, new_new_n2633__, new_new_n2634__, new_new_n2635__,
    new_new_n2636__, new_new_n2637__, new_new_n2638__, new_new_n2639__,
    new_new_n2640__, new_new_n2641__, new_new_n2642__, new_new_n2643__,
    new_new_n2644__, new_new_n2645__, new_new_n2646__, new_new_n2647__,
    new_new_n2648__, new_new_n2649__, new_new_n2650__, new_new_n2651__,
    new_new_n2652__, new_new_n2653__, new_new_n2654__, new_new_n2655__,
    new_new_n2656__, new_new_n2657__, new_new_n2658__, new_new_n2659__,
    new_new_n2660__, new_new_n2661__, new_new_n2662__, new_new_n2663__,
    new_new_n2664__, new_new_n2665__, new_new_n2666__, new_new_n2667__,
    new_new_n2668__, new_new_n2669__, new_new_n2670__, new_new_n2671__,
    new_new_n2672__, new_new_n2673__, new_new_n2674__, new_new_n2675__,
    new_new_n2676__, new_new_n2677__, new_new_n2678__, new_new_n2679__,
    new_new_n2680__, new_new_n2681__, new_new_n2682__, new_new_n2683__,
    new_new_n2684__, new_new_n2685__, new_new_n2686__, new_new_n2687__,
    new_new_n2688__, new_new_n2689__, new_new_n2690__, new_new_n2691__,
    new_new_n2692__, new_new_n2693__, new_new_n2694__, new_new_n2695__,
    new_new_n2696__, new_new_n2697__, new_new_n2698__, new_new_n2699__,
    new_new_n2700__, new_new_n2701__, new_new_n2702__, new_new_n2703__,
    new_new_n2704__, new_new_n2705__, new_new_n2706__, new_new_n2707__,
    new_new_n2708__, new_new_n2709__, new_new_n2710__, new_new_n2711__,
    new_new_n2712__, new_new_n2713__, new_new_n2714__, new_new_n2715__,
    new_new_n2716__, new_new_n2717__, new_new_n2718__, new_new_n2719__,
    new_new_n2720__, new_new_n2721__, new_new_n2722__, new_new_n2723__,
    new_new_n2724__, new_new_n2725__, new_new_n2726__, new_new_n2727__,
    new_new_n2728__, new_new_n2729__, new_new_n2730__, new_new_n2731__,
    new_new_n2732__, new_new_n2733__, new_new_n2734__, new_new_n2735__,
    new_new_n2736__, new_new_n2737__, new_new_n2738__, new_new_n2739__,
    new_new_n2740__, new_new_n2741__, new_new_n2742__, new_new_n2743__,
    new_new_n2744__, new_new_n2745__, new_new_n2746__, new_new_n2747__,
    new_new_n2748__, new_new_n2749__, new_new_n2750__, new_new_n2751__,
    new_new_n2752__, new_new_n2753__, new_new_n2754__, new_new_n2755__,
    new_new_n2756__, new_new_n2757__, new_new_n2758__, new_new_n2759__,
    new_new_n2760__, new_new_n2761__, new_new_n2762__, new_new_n2763__,
    new_new_n2764__, new_new_n2765__, new_new_n2766__, new_new_n2767__,
    new_new_n2768__, new_new_n2770__, new_new_n2771__, new_new_n2772__,
    new_new_n2773__, new_new_n2774__, new_new_n2775__, new_new_n2776__,
    new_new_n2777__, new_new_n2778__, new_new_n2779__, new_new_n2780__,
    new_new_n2781__, new_new_n2782__, new_new_n2783__, new_new_n2784__,
    new_new_n2785__, new_new_n2786__, new_new_n2787__, new_new_n2788__,
    new_new_n2789__, new_new_n2790__, new_new_n2791__, new_new_n2792__,
    new_new_n2793__, new_new_n2794__, new_new_n2795__, new_new_n2796__,
    new_new_n2797__, new_new_n2798__, new_new_n2799__, new_new_n2800__,
    new_new_n2801__, new_new_n2802__, new_new_n2803__, new_new_n2804__,
    new_new_n2805__, new_new_n2806__, new_new_n2807__, new_new_n2808__,
    new_new_n2809__, new_new_n2810__, new_new_n2811__, new_new_n2812__,
    new_new_n2813__, new_new_n2814__, new_new_n2815__, new_new_n2816__,
    new_new_n2817__, new_new_n2818__, new_new_n2819__, new_new_n2820__,
    new_new_n2821__, new_new_n2822__, new_new_n2823__, new_new_n2824__,
    new_new_n2825__, new_new_n2826__, new_new_n2827__, new_new_n2828__,
    new_new_n2829__, new_new_n2830__, new_new_n2831__, new_new_n2832__,
    new_new_n2833__, new_new_n2834__, new_new_n2835__, new_new_n2836__,
    new_new_n2837__, new_new_n2838__, new_new_n2839__, new_new_n2840__,
    new_new_n2841__, new_new_n2842__, new_new_n2843__, new_new_n2844__,
    new_new_n2845__, new_new_n2846__, new_new_n2847__, new_new_n2848__,
    new_new_n2849__, new_new_n2850__, new_new_n2851__, new_new_n2852__,
    new_new_n2853__, new_new_n2854__, new_new_n2855__, new_new_n2856__,
    new_new_n2857__, new_new_n2858__, new_new_n2859__, new_new_n2860__,
    new_new_n2861__, new_new_n2862__, new_new_n2863__, new_new_n2864__,
    new_new_n2865__, new_new_n2866__, new_new_n2867__, new_new_n2868__,
    new_new_n2869__, new_new_n2870__, new_new_n2871__, new_new_n2872__,
    new_new_n2873__, new_new_n2874__, new_new_n2875__, new_new_n2876__,
    new_new_n2877__, new_new_n2878__, new_new_n2879__, new_new_n2880__,
    new_new_n2881__, new_new_n2882__, new_new_n2883__, new_new_n2884__,
    new_new_n2885__, new_new_n2886__, new_new_n2887__, new_new_n2888__,
    new_new_n2889__, new_new_n2890__, new_new_n2891__, new_new_n2892__,
    new_new_n2893__, new_new_n2894__, new_new_n2895__, new_new_n2896__,
    new_new_n2897__, new_new_n2898__, new_new_n2899__, new_new_n2900__,
    new_new_n2901__, new_new_n2902__, new_new_n2903__, new_new_n2904__,
    new_new_n2905__, new_new_n2906__, new_new_n2907__, new_new_n2908__,
    new_new_n2909__, new_new_n2910__, new_new_n2911__, new_new_n2912__,
    new_new_n2913__, new_new_n2914__, new_new_n2915__, new_new_n2916__,
    new_new_n2918__, new_new_n2919__, new_new_n2920__, new_new_n2921__,
    new_new_n2922__, new_new_n2923__, new_new_n2924__, new_new_n2925__,
    new_new_n2926__, new_new_n2927__, new_new_n2928__, new_new_n2929__,
    new_new_n2930__, new_new_n2931__, new_new_n2932__, new_new_n2933__,
    new_new_n2934__, new_new_n2935__, new_new_n2936__, new_new_n2937__,
    new_new_n2938__, new_new_n2939__, new_new_n2940__, new_new_n2941__,
    new_new_n2942__, new_new_n2943__, new_new_n2944__, new_new_n2945__,
    new_new_n2946__, new_new_n2947__, new_new_n2948__, new_new_n2949__,
    new_new_n2950__, new_new_n2951__, new_new_n2952__, new_new_n2953__,
    new_new_n2954__, new_new_n2955__, new_new_n2956__, new_new_n2957__,
    new_new_n2958__, new_new_n2959__, new_new_n2960__, new_new_n2961__,
    new_new_n2962__, new_new_n2963__, new_new_n2964__, new_new_n2965__,
    new_new_n2966__, new_new_n2967__, new_new_n2968__, new_new_n2969__,
    new_new_n2970__, new_new_n2971__, new_new_n2972__, new_new_n2973__,
    new_new_n2974__, new_new_n2975__, new_new_n2976__, new_new_n2977__,
    new_new_n2978__, new_new_n2979__, new_new_n2980__, new_new_n2981__,
    new_new_n2982__, new_new_n2983__, new_new_n2984__, new_new_n2985__,
    new_new_n2986__, new_new_n2987__, new_new_n2988__, new_new_n2989__,
    new_new_n2990__, new_new_n2991__, new_new_n2992__, new_new_n2993__,
    new_new_n2994__, new_new_n2995__, new_new_n2996__, new_new_n2997__,
    new_new_n2998__, new_new_n2999__, new_new_n3000__, new_new_n3001__,
    new_new_n3002__, new_new_n3003__, new_new_n3004__, new_new_n3005__,
    new_new_n3006__, new_new_n3007__, new_new_n3008__, new_new_n3009__,
    new_new_n3010__, new_new_n3011__, new_new_n3012__, new_new_n3013__,
    new_new_n3014__, new_new_n3015__, new_new_n3016__, new_new_n3017__,
    new_new_n3018__, new_new_n3019__, new_new_n3020__, new_new_n3021__,
    new_new_n3022__, new_new_n3023__, new_new_n3024__, new_new_n3025__,
    new_new_n3026__, new_new_n3027__, new_new_n3028__, new_new_n3029__,
    new_new_n3030__, new_new_n3031__, new_new_n3032__, new_new_n3033__,
    new_new_n3034__, new_new_n3035__, new_new_n3036__, new_new_n3037__,
    new_new_n3038__, new_new_n3039__, new_new_n3040__, new_new_n3041__,
    new_new_n3042__, new_new_n3043__, new_new_n3044__, new_new_n3045__,
    new_new_n3046__, new_new_n3047__, new_new_n3048__, new_new_n3049__,
    new_new_n3050__, new_new_n3051__, new_new_n3052__, new_new_n3053__,
    new_new_n3054__, new_new_n3055__, new_new_n3056__, new_new_n3057__,
    new_new_n3058__, new_new_n3059__, new_new_n3060__, new_new_n3061__,
    new_new_n3062__, new_new_n3063__, new_new_n3064__, new_new_n3065__,
    new_new_n3066__, new_new_n3067__, new_new_n3068__, new_new_n3069__,
    new_new_n3070__, new_new_n3071__, new_new_n3072__, new_new_n3073__,
    new_new_n3074__, new_new_n3075__, new_new_n3076__, new_new_n3077__,
    new_new_n3078__, new_new_n3079__, new_new_n3080__, new_new_n3081__,
    new_new_n3082__, new_new_n3084__, new_new_n3085__, new_new_n3086__,
    new_new_n3087__, new_new_n3088__, new_new_n3089__, new_new_n3090__,
    new_new_n3091__, new_new_n3092__, new_new_n3093__, new_new_n3094__,
    new_new_n3095__, new_new_n3096__, new_new_n3097__, new_new_n3098__,
    new_new_n3099__, new_new_n3100__, new_new_n3101__, new_new_n3102__,
    new_new_n3103__, new_new_n3104__, new_new_n3105__, new_new_n3106__,
    new_new_n3107__, new_new_n3108__, new_new_n3109__, new_new_n3110__,
    new_new_n3111__, new_new_n3112__, new_new_n3113__, new_new_n3114__,
    new_new_n3115__, new_new_n3116__, new_new_n3117__, new_new_n3118__,
    new_new_n3119__, new_new_n3120__, new_new_n3121__, new_new_n3122__,
    new_new_n3123__, new_new_n3124__, new_new_n3125__, new_new_n3126__,
    new_new_n3127__, new_new_n3128__, new_new_n3129__, new_new_n3130__,
    new_new_n3131__, new_new_n3132__, new_new_n3133__, new_new_n3134__,
    new_new_n3135__, new_new_n3136__, new_new_n3137__, new_new_n3138__,
    new_new_n3139__, new_new_n3140__, new_new_n3141__, new_new_n3142__,
    new_new_n3143__, new_new_n3144__, new_new_n3145__, new_new_n3146__,
    new_new_n3147__, new_new_n3148__, new_new_n3149__, new_new_n3150__,
    new_new_n3151__, new_new_n3152__, new_new_n3153__, new_new_n3154__,
    new_new_n3155__, new_new_n3156__, new_new_n3157__, new_new_n3158__,
    new_new_n3159__, new_new_n3160__, new_new_n3161__, new_new_n3162__,
    new_new_n3163__, new_new_n3164__, new_new_n3165__, new_new_n3166__,
    new_new_n3167__, new_new_n3168__, new_new_n3169__, new_new_n3170__,
    new_new_n3171__, new_new_n3172__, new_new_n3173__, new_new_n3174__,
    new_new_n3175__, new_new_n3176__, new_new_n3177__, new_new_n3178__,
    new_new_n3179__, new_new_n3180__, new_new_n3181__, new_new_n3182__,
    new_new_n3183__, new_new_n3184__, new_new_n3185__, new_new_n3186__,
    new_new_n3187__, new_new_n3188__, new_new_n3189__, new_new_n3190__,
    new_new_n3191__, new_new_n3192__, new_new_n3193__, new_new_n3194__,
    new_new_n3195__, new_new_n3196__, new_new_n3197__, new_new_n3198__,
    new_new_n3199__, new_new_n3200__, new_new_n3201__, new_new_n3202__,
    new_new_n3203__, new_new_n3204__, new_new_n3205__, new_new_n3206__,
    new_new_n3207__, new_new_n3208__, new_new_n3209__, new_new_n3210__,
    new_new_n3211__, new_new_n3212__, new_new_n3213__, new_new_n3214__,
    new_new_n3215__, new_new_n3216__, new_new_n3217__, new_new_n3218__,
    new_new_n3219__, new_new_n3220__, new_new_n3221__, new_new_n3222__,
    new_new_n3223__, new_new_n3224__, new_new_n3225__, new_new_n3226__,
    new_new_n3227__, new_new_n3228__, new_new_n3229__, new_new_n3230__,
    new_new_n3231__, new_new_n3232__, new_new_n3233__, new_new_n3234__,
    new_new_n3235__, new_new_n3236__, new_new_n3237__, new_new_n3238__,
    new_new_n3239__, new_new_n3240__, new_new_n3241__, new_new_n3242__,
    new_new_n3243__, new_new_n3245__, new_new_n3246__, new_new_n3247__,
    new_new_n3248__, new_new_n3249__, new_new_n3250__, new_new_n3251__,
    new_new_n3252__, new_new_n3253__, new_new_n3254__, new_new_n3255__,
    new_new_n3256__, new_new_n3257__, new_new_n3258__, new_new_n3259__,
    new_new_n3260__, new_new_n3261__, new_new_n3262__, new_new_n3263__,
    new_new_n3264__, new_new_n3265__, new_new_n3266__, new_new_n3267__,
    new_new_n3268__, new_new_n3269__, new_new_n3270__, new_new_n3271__,
    new_new_n3272__, new_new_n3273__, new_new_n3274__, new_new_n3275__,
    new_new_n3276__, new_new_n3277__, new_new_n3278__, new_new_n3279__,
    new_new_n3280__, new_new_n3281__, new_new_n3282__, new_new_n3283__,
    new_new_n3284__, new_new_n3285__, new_new_n3286__, new_new_n3287__,
    new_new_n3288__, new_new_n3289__, new_new_n3290__, new_new_n3291__,
    new_new_n3292__, new_new_n3293__, new_new_n3294__, new_new_n3295__,
    new_new_n3296__, new_new_n3297__, new_new_n3298__, new_new_n3299__,
    new_new_n3300__, new_new_n3301__, new_new_n3302__, new_new_n3303__,
    new_new_n3304__, new_new_n3305__, new_new_n3306__, new_new_n3307__,
    new_new_n3308__, new_new_n3309__, new_new_n3310__, new_new_n3311__,
    new_new_n3312__, new_new_n3313__, new_new_n3314__, new_new_n3315__,
    new_new_n3316__, new_new_n3317__, new_new_n3318__, new_new_n3319__,
    new_new_n3320__, new_new_n3321__, new_new_n3322__, new_new_n3323__,
    new_new_n3324__, new_new_n3325__, new_new_n3326__, new_new_n3327__,
    new_new_n3328__, new_new_n3329__, new_new_n3330__, new_new_n3331__,
    new_new_n3332__, new_new_n3333__, new_new_n3334__, new_new_n3335__,
    new_new_n3336__, new_new_n3337__, new_new_n3338__, new_new_n3339__,
    new_new_n3340__, new_new_n3341__, new_new_n3342__, new_new_n3343__,
    new_new_n3344__, new_new_n3345__, new_new_n3346__, new_new_n3347__,
    new_new_n3348__, new_new_n3349__, new_new_n3350__, new_new_n3351__,
    new_new_n3352__, new_new_n3353__, new_new_n3354__, new_new_n3355__,
    new_new_n3356__, new_new_n3357__, new_new_n3358__, new_new_n3359__,
    new_new_n3360__, new_new_n3361__, new_new_n3362__, new_new_n3363__,
    new_new_n3364__, new_new_n3365__, new_new_n3366__, new_new_n3367__,
    new_new_n3368__, new_new_n3369__, new_new_n3370__, new_new_n3371__,
    new_new_n3372__, new_new_n3373__, new_new_n3374__, new_new_n3375__,
    new_new_n3376__, new_new_n3377__, new_new_n3378__, new_new_n3379__,
    new_new_n3380__, new_new_n3381__, new_new_n3382__, new_new_n3383__,
    new_new_n3384__, new_new_n3385__, new_new_n3386__, new_new_n3387__,
    new_new_n3388__, new_new_n3389__, new_new_n3390__, new_new_n3391__,
    new_new_n3392__, new_new_n3393__, new_new_n3394__, new_new_n3395__,
    new_new_n3396__, new_new_n3397__, new_new_n3398__, new_new_n3399__,
    new_new_n3400__, new_new_n3401__, new_new_n3402__, new_new_n3403__,
    new_new_n3404__, new_new_n3405__, new_new_n3406__, new_new_n3407__,
    new_new_n3408__, new_new_n3409__, new_new_n3410__, new_new_n3411__,
    new_new_n3412__, new_new_n3413__, new_new_n3414__, new_new_n3415__,
    new_new_n3416__, new_new_n3417__, new_new_n3418__, new_new_n3419__,
    new_new_n3420__, new_new_n3421__, new_new_n3422__, new_new_n3423__,
    new_new_n3424__, new_new_n3425__, new_new_n3426__, new_new_n3427__,
    new_new_n3428__, new_new_n3429__, new_new_n3430__, new_new_n3431__,
    new_new_n3432__, new_new_n3433__, new_new_n3434__, new_new_n3435__,
    new_new_n3436__, new_new_n3438__, new_new_n3439__, new_new_n3440__,
    new_new_n3441__, new_new_n3442__, new_new_n3443__, new_new_n3444__,
    new_new_n3445__, new_new_n3446__, new_new_n3447__, new_new_n3448__,
    new_new_n3449__, new_new_n3450__, new_new_n3451__, new_new_n3452__,
    new_new_n3453__, new_new_n3454__, new_new_n3455__, new_new_n3456__,
    new_new_n3457__, new_new_n3458__, new_new_n3459__, new_new_n3460__,
    new_new_n3461__, new_new_n3462__, new_new_n3463__, new_new_n3464__,
    new_new_n3465__, new_new_n3466__, new_new_n3467__, new_new_n3468__,
    new_new_n3469__, new_new_n3470__, new_new_n3471__, new_new_n3472__,
    new_new_n3473__, new_new_n3474__, new_new_n3475__, new_new_n3476__,
    new_new_n3477__, new_new_n3478__, new_new_n3479__, new_new_n3480__,
    new_new_n3481__, new_new_n3482__, new_new_n3483__, new_new_n3484__,
    new_new_n3485__, new_new_n3486__, new_new_n3487__, new_new_n3488__,
    new_new_n3489__, new_new_n3490__, new_new_n3491__, new_new_n3492__,
    new_new_n3493__, new_new_n3494__, new_new_n3495__, new_new_n3496__,
    new_new_n3497__, new_new_n3498__, new_new_n3499__, new_new_n3500__,
    new_new_n3501__, new_new_n3502__, new_new_n3503__, new_new_n3504__,
    new_new_n3505__, new_new_n3506__, new_new_n3507__, new_new_n3508__,
    new_new_n3509__, new_new_n3510__, new_new_n3511__, new_new_n3512__,
    new_new_n3513__, new_new_n3514__, new_new_n3515__, new_new_n3516__,
    new_new_n3517__, new_new_n3518__, new_new_n3519__, new_new_n3520__,
    new_new_n3521__, new_new_n3522__, new_new_n3523__, new_new_n3524__,
    new_new_n3525__, new_new_n3526__, new_new_n3527__, new_new_n3528__,
    new_new_n3529__, new_new_n3530__, new_new_n3531__, new_new_n3532__,
    new_new_n3533__, new_new_n3534__, new_new_n3535__, new_new_n3536__,
    new_new_n3537__, new_new_n3538__, new_new_n3539__, new_new_n3540__,
    new_new_n3541__, new_new_n3542__, new_new_n3543__, new_new_n3544__,
    new_new_n3545__, new_new_n3546__, new_new_n3547__, new_new_n3548__,
    new_new_n3549__, new_new_n3550__, new_new_n3551__, new_new_n3552__,
    new_new_n3553__, new_new_n3554__, new_new_n3555__, new_new_n3556__,
    new_new_n3557__, new_new_n3558__, new_new_n3559__, new_new_n3560__,
    new_new_n3561__, new_new_n3562__, new_new_n3563__, new_new_n3564__,
    new_new_n3565__, new_new_n3566__, new_new_n3567__, new_new_n3568__,
    new_new_n3569__, new_new_n3570__, new_new_n3571__, new_new_n3572__,
    new_new_n3573__, new_new_n3574__, new_new_n3575__, new_new_n3576__,
    new_new_n3577__, new_new_n3578__, new_new_n3579__, new_new_n3580__,
    new_new_n3581__, new_new_n3582__, new_new_n3583__, new_new_n3584__,
    new_new_n3585__, new_new_n3586__, new_new_n3587__, new_new_n3588__,
    new_new_n3589__, new_new_n3590__, new_new_n3591__, new_new_n3592__,
    new_new_n3593__, new_new_n3594__, new_new_n3595__, new_new_n3596__,
    new_new_n3597__, new_new_n3598__, new_new_n3599__, new_new_n3600__,
    new_new_n3602__, new_new_n3603__, new_new_n3604__, new_new_n3605__,
    new_new_n3606__, new_new_n3607__, new_new_n3608__, new_new_n3609__,
    new_new_n3610__, new_new_n3611__, new_new_n3612__, new_new_n3613__,
    new_new_n3614__, new_new_n3615__, new_new_n3616__, new_new_n3617__,
    new_new_n3618__, new_new_n3619__, new_new_n3620__, new_new_n3621__,
    new_new_n3622__, new_new_n3623__, new_new_n3624__, new_new_n3625__,
    new_new_n3626__, new_new_n3627__, new_new_n3628__, new_new_n3629__,
    new_new_n3630__, new_new_n3631__, new_new_n3632__, new_new_n3633__,
    new_new_n3634__, new_new_n3635__, new_new_n3636__, new_new_n3637__,
    new_new_n3638__, new_new_n3639__, new_new_n3640__, new_new_n3641__,
    new_new_n3642__, new_new_n3643__, new_new_n3644__, new_new_n3645__,
    new_new_n3646__, new_new_n3647__, new_new_n3648__, new_new_n3649__,
    new_new_n3650__, new_new_n3651__, new_new_n3652__, new_new_n3653__,
    new_new_n3654__, new_new_n3655__, new_new_n3656__, new_new_n3657__,
    new_new_n3658__, new_new_n3659__, new_new_n3660__, new_new_n3661__,
    new_new_n3662__, new_new_n3663__, new_new_n3664__, new_new_n3665__,
    new_new_n3666__, new_new_n3667__, new_new_n3668__, new_new_n3669__,
    new_new_n3670__, new_new_n3671__, new_new_n3672__, new_new_n3673__,
    new_new_n3674__, new_new_n3675__, new_new_n3676__, new_new_n3677__,
    new_new_n3678__, new_new_n3679__, new_new_n3680__, new_new_n3681__,
    new_new_n3682__, new_new_n3683__, new_new_n3684__, new_new_n3685__,
    new_new_n3686__, new_new_n3687__, new_new_n3688__, new_new_n3689__,
    new_new_n3690__, new_new_n3691__, new_new_n3692__, new_new_n3693__,
    new_new_n3694__, new_new_n3695__, new_new_n3696__, new_new_n3697__,
    new_new_n3698__, new_new_n3699__, new_new_n3700__, new_new_n3701__,
    new_new_n3702__, new_new_n3703__, new_new_n3704__, new_new_n3705__,
    new_new_n3706__, new_new_n3707__, new_new_n3708__, new_new_n3709__,
    new_new_n3710__, new_new_n3711__, new_new_n3712__, new_new_n3713__,
    new_new_n3714__, new_new_n3715__, new_new_n3716__, new_new_n3717__,
    new_new_n3718__, new_new_n3719__, new_new_n3720__, new_new_n3721__,
    new_new_n3722__, new_new_n3723__, new_new_n3724__, new_new_n3725__,
    new_new_n3726__, new_new_n3727__, new_new_n3728__, new_new_n3729__,
    new_new_n3730__, new_new_n3731__, new_new_n3732__, new_new_n3733__,
    new_new_n3734__, new_new_n3735__, new_new_n3736__, new_new_n3737__,
    new_new_n3738__, new_new_n3739__, new_new_n3740__, new_new_n3741__,
    new_new_n3742__, new_new_n3743__, new_new_n3744__, new_new_n3745__,
    new_new_n3746__, new_new_n3747__, new_new_n3748__, new_new_n3749__,
    new_new_n3750__, new_new_n3751__, new_new_n3752__, new_new_n3753__,
    new_new_n3754__, new_new_n3755__, new_new_n3756__, new_new_n3757__,
    new_new_n3758__, new_new_n3759__, new_new_n3760__, new_new_n3761__,
    new_new_n3762__, new_new_n3763__, new_new_n3764__, new_new_n3765__,
    new_new_n3766__, new_new_n3767__, new_new_n3768__, new_new_n3769__,
    new_new_n3770__, new_new_n3771__, new_new_n3772__, new_new_n3773__,
    new_new_n3774__, new_new_n3775__, new_new_n3776__, new_new_n3777__,
    new_new_n3778__, new_new_n3779__, new_new_n3780__, new_new_n3781__,
    new_new_n3782__, new_new_n3783__, new_new_n3784__, new_new_n3785__,
    new_new_n3786__, new_new_n3787__, new_new_n3788__, new_new_n3789__,
    new_new_n3790__, new_new_n3791__, new_new_n3792__, new_new_n3793__,
    new_new_n3794__, new_new_n3795__, new_new_n3796__, new_new_n3797__,
    new_new_n3799__, new_new_n3800__, new_new_n3801__, new_new_n3802__,
    new_new_n3803__, new_new_n3804__, new_new_n3805__, new_new_n3806__,
    new_new_n3807__, new_new_n3808__, new_new_n3809__, new_new_n3810__,
    new_new_n3811__, new_new_n3812__, new_new_n3813__, new_new_n3814__,
    new_new_n3815__, new_new_n3816__, new_new_n3817__, new_new_n3818__,
    new_new_n3819__, new_new_n3820__, new_new_n3821__, new_new_n3822__,
    new_new_n3823__, new_new_n3824__, new_new_n3825__, new_new_n3826__,
    new_new_n3827__, new_new_n3828__, new_new_n3829__, new_new_n3830__,
    new_new_n3831__, new_new_n3832__, new_new_n3833__, new_new_n3834__,
    new_new_n3835__, new_new_n3836__, new_new_n3837__, new_new_n3838__,
    new_new_n3839__, new_new_n3840__, new_new_n3841__, new_new_n3842__,
    new_new_n3843__, new_new_n3844__, new_new_n3845__, new_new_n3846__,
    new_new_n3847__, new_new_n3848__, new_new_n3849__, new_new_n3850__,
    new_new_n3851__, new_new_n3852__, new_new_n3853__, new_new_n3854__,
    new_new_n3855__, new_new_n3856__, new_new_n3857__, new_new_n3858__,
    new_new_n3859__, new_new_n3860__, new_new_n3861__, new_new_n3862__,
    new_new_n3863__, new_new_n3864__, new_new_n3865__, new_new_n3866__,
    new_new_n3867__, new_new_n3868__, new_new_n3869__, new_new_n3870__,
    new_new_n3871__, new_new_n3872__, new_new_n3873__, new_new_n3874__,
    new_new_n3875__, new_new_n3876__, new_new_n3877__, new_new_n3878__,
    new_new_n3879__, new_new_n3880__, new_new_n3881__, new_new_n3882__,
    new_new_n3883__, new_new_n3884__, new_new_n3885__, new_new_n3886__,
    new_new_n3887__, new_new_n3888__, new_new_n3889__, new_new_n3890__,
    new_new_n3891__, new_new_n3892__, new_new_n3893__, new_new_n3894__,
    new_new_n3895__, new_new_n3896__, new_new_n3897__, new_new_n3898__,
    new_new_n3899__, new_new_n3900__, new_new_n3901__, new_new_n3902__,
    new_new_n3903__, new_new_n3904__, new_new_n3905__, new_new_n3906__,
    new_new_n3907__, new_new_n3908__, new_new_n3909__, new_new_n3910__,
    new_new_n3911__, new_new_n3912__, new_new_n3913__, new_new_n3914__,
    new_new_n3915__, new_new_n3916__, new_new_n3917__, new_new_n3918__,
    new_new_n3919__, new_new_n3920__, new_new_n3921__, new_new_n3922__,
    new_new_n3923__, new_new_n3924__, new_new_n3925__, new_new_n3926__,
    new_new_n3927__, new_new_n3928__, new_new_n3929__, new_new_n3930__,
    new_new_n3931__, new_new_n3932__, new_new_n3933__, new_new_n3934__,
    new_new_n3935__, new_new_n3936__, new_new_n3937__, new_new_n3938__,
    new_new_n3939__, new_new_n3940__, new_new_n3941__, new_new_n3942__,
    new_new_n3943__, new_new_n3944__, new_new_n3945__, new_new_n3946__,
    new_new_n3947__, new_new_n3948__, new_new_n3949__, new_new_n3950__,
    new_new_n3951__, new_new_n3952__, new_new_n3953__, new_new_n3954__,
    new_new_n3955__, new_new_n3956__, new_new_n3957__, new_new_n3958__,
    new_new_n3959__, new_new_n3960__, new_new_n3961__, new_new_n3962__,
    new_new_n3963__, new_new_n3964__, new_new_n3965__, new_new_n3966__,
    new_new_n3967__, new_new_n3968__, new_new_n3969__, new_new_n3970__,
    new_new_n3971__, new_new_n3972__, new_new_n3973__, new_new_n3974__,
    new_new_n3975__, new_new_n3976__, new_new_n3978__, new_new_n3979__,
    new_new_n3980__, new_new_n3981__, new_new_n3982__, new_new_n3983__,
    new_new_n3984__, new_new_n3985__, new_new_n3986__, new_new_n3987__,
    new_new_n3988__, new_new_n3989__, new_new_n3990__, new_new_n3991__,
    new_new_n3992__, new_new_n3993__, new_new_n3994__, new_new_n3995__,
    new_new_n3996__, new_new_n3997__, new_new_n3998__, new_new_n3999__,
    new_new_n4000__, new_new_n4001__, new_new_n4002__, new_new_n4003__,
    new_new_n4004__, new_new_n4005__, new_new_n4006__, new_new_n4007__,
    new_new_n4008__, new_new_n4009__, new_new_n4010__, new_new_n4011__,
    new_new_n4012__, new_new_n4013__, new_new_n4014__, new_new_n4015__,
    new_new_n4016__, new_new_n4017__, new_new_n4018__, new_new_n4019__,
    new_new_n4020__, new_new_n4021__, new_new_n4022__, new_new_n4023__,
    new_new_n4024__, new_new_n4025__, new_new_n4026__, new_new_n4027__,
    new_new_n4028__, new_new_n4029__, new_new_n4030__, new_new_n4031__,
    new_new_n4032__, new_new_n4033__, new_new_n4034__, new_new_n4035__,
    new_new_n4036__, new_new_n4037__, new_new_n4038__, new_new_n4039__,
    new_new_n4040__, new_new_n4041__, new_new_n4042__, new_new_n4043__,
    new_new_n4044__, new_new_n4045__, new_new_n4046__, new_new_n4047__,
    new_new_n4048__, new_new_n4049__, new_new_n4050__, new_new_n4051__,
    new_new_n4052__, new_new_n4053__, new_new_n4054__, new_new_n4055__,
    new_new_n4056__, new_new_n4057__, new_new_n4058__, new_new_n4059__,
    new_new_n4060__, new_new_n4061__, new_new_n4062__, new_new_n4063__,
    new_new_n4064__, new_new_n4065__, new_new_n4066__, new_new_n4067__,
    new_new_n4068__, new_new_n4069__, new_new_n4070__, new_new_n4071__,
    new_new_n4072__, new_new_n4073__, new_new_n4074__, new_new_n4075__,
    new_new_n4076__, new_new_n4077__, new_new_n4078__, new_new_n4079__,
    new_new_n4080__, new_new_n4081__, new_new_n4082__, new_new_n4083__,
    new_new_n4084__, new_new_n4085__, new_new_n4086__, new_new_n4087__,
    new_new_n4088__, new_new_n4089__, new_new_n4090__, new_new_n4091__,
    new_new_n4092__, new_new_n4093__, new_new_n4094__, new_new_n4095__,
    new_new_n4096__, new_new_n4097__, new_new_n4098__, new_new_n4099__,
    new_new_n4100__, new_new_n4101__, new_new_n4102__, new_new_n4103__,
    new_new_n4104__, new_new_n4105__, new_new_n4106__, new_new_n4107__,
    new_new_n4108__, new_new_n4109__, new_new_n4110__, new_new_n4111__,
    new_new_n4112__, new_new_n4113__, new_new_n4114__, new_new_n4115__,
    new_new_n4116__, new_new_n4117__, new_new_n4118__, new_new_n4119__,
    new_new_n4120__, new_new_n4121__, new_new_n4122__, new_new_n4123__,
    new_new_n4124__, new_new_n4125__, new_new_n4126__, new_new_n4127__,
    new_new_n4128__, new_new_n4129__, new_new_n4130__, new_new_n4131__,
    new_new_n4132__, new_new_n4133__, new_new_n4134__, new_new_n4135__,
    new_new_n4136__, new_new_n4137__, new_new_n4138__, new_new_n4139__,
    new_new_n4140__, new_new_n4141__, new_new_n4142__, new_new_n4143__,
    new_new_n4144__, new_new_n4145__, new_new_n4146__, new_new_n4147__,
    new_new_n4148__, new_new_n4149__, new_new_n4150__, new_new_n4151__,
    new_new_n4152__, new_new_n4153__, new_new_n4154__, new_new_n4155__,
    new_new_n4156__, new_new_n4157__, new_new_n4158__, new_new_n4159__,
    new_new_n4160__, new_new_n4161__, new_new_n4162__, new_new_n4163__,
    new_new_n4164__, new_new_n4165__, new_new_n4166__, new_new_n4167__,
    new_new_n4168__, new_new_n4169__, new_new_n4170__, new_new_n4171__,
    new_new_n4172__, new_new_n4173__, new_new_n4174__, new_new_n4175__,
    new_new_n4176__, new_new_n4177__, new_new_n4178__, new_new_n4180__,
    new_new_n4181__, new_new_n4182__, new_new_n4183__, new_new_n4184__,
    new_new_n4185__, new_new_n4186__, new_new_n4187__, new_new_n4188__,
    new_new_n4189__, new_new_n4190__, new_new_n4191__, new_new_n4192__,
    new_new_n4193__, new_new_n4194__, new_new_n4195__, new_new_n4196__,
    new_new_n4197__, new_new_n4198__, new_new_n4199__, new_new_n4200__,
    new_new_n4201__, new_new_n4202__, new_new_n4203__, new_new_n4204__,
    new_new_n4205__, new_new_n4206__, new_new_n4207__, new_new_n4208__,
    new_new_n4209__, new_new_n4210__, new_new_n4211__, new_new_n4212__,
    new_new_n4213__, new_new_n4214__, new_new_n4215__, new_new_n4216__,
    new_new_n4217__, new_new_n4218__, new_new_n4219__, new_new_n4220__,
    new_new_n4221__, new_new_n4222__, new_new_n4223__, new_new_n4224__,
    new_new_n4225__, new_new_n4226__, new_new_n4227__, new_new_n4228__,
    new_new_n4229__, new_new_n4230__, new_new_n4231__, new_new_n4232__,
    new_new_n4233__, new_new_n4234__, new_new_n4235__, new_new_n4236__,
    new_new_n4237__, new_new_n4238__, new_new_n4239__, new_new_n4240__,
    new_new_n4241__, new_new_n4242__, new_new_n4243__, new_new_n4244__,
    new_new_n4245__, new_new_n4246__, new_new_n4247__, new_new_n4248__,
    new_new_n4249__, new_new_n4250__, new_new_n4251__, new_new_n4252__,
    new_new_n4253__, new_new_n4254__, new_new_n4255__, new_new_n4256__,
    new_new_n4257__, new_new_n4258__, new_new_n4259__, new_new_n4260__,
    new_new_n4261__, new_new_n4262__, new_new_n4263__, new_new_n4264__,
    new_new_n4265__, new_new_n4266__, new_new_n4267__, new_new_n4268__,
    new_new_n4269__, new_new_n4270__, new_new_n4271__, new_new_n4272__,
    new_new_n4273__, new_new_n4274__, new_new_n4275__, new_new_n4276__,
    new_new_n4277__, new_new_n4278__, new_new_n4279__, new_new_n4280__,
    new_new_n4281__, new_new_n4282__, new_new_n4283__, new_new_n4284__,
    new_new_n4285__, new_new_n4286__, new_new_n4287__, new_new_n4288__,
    new_new_n4289__, new_new_n4290__, new_new_n4291__, new_new_n4292__,
    new_new_n4293__, new_new_n4294__, new_new_n4295__, new_new_n4296__,
    new_new_n4297__, new_new_n4298__, new_new_n4299__, new_new_n4300__,
    new_new_n4301__, new_new_n4302__, new_new_n4303__, new_new_n4304__,
    new_new_n4305__, new_new_n4306__, new_new_n4307__, new_new_n4308__,
    new_new_n4309__, new_new_n4310__, new_new_n4311__, new_new_n4312__,
    new_new_n4313__, new_new_n4314__, new_new_n4315__, new_new_n4316__,
    new_new_n4317__, new_new_n4318__, new_new_n4319__, new_new_n4320__,
    new_new_n4321__, new_new_n4322__, new_new_n4323__, new_new_n4324__,
    new_new_n4325__, new_new_n4326__, new_new_n4327__, new_new_n4328__,
    new_new_n4329__, new_new_n4330__, new_new_n4331__, new_new_n4332__,
    new_new_n4333__, new_new_n4334__, new_new_n4335__, new_new_n4336__,
    new_new_n4337__, new_new_n4338__, new_new_n4339__, new_new_n4340__,
    new_new_n4341__, new_new_n4342__, new_new_n4343__, new_new_n4344__,
    new_new_n4345__, new_new_n4346__, new_new_n4347__, new_new_n4348__,
    new_new_n4349__, new_new_n4350__, new_new_n4351__, new_new_n4352__,
    new_new_n4353__, new_new_n4354__, new_new_n4355__, new_new_n4356__,
    new_new_n4357__, new_new_n4358__, new_new_n4359__, new_new_n4360__,
    new_new_n4361__, new_new_n4362__, new_new_n4363__, new_new_n4364__,
    new_new_n4365__, new_new_n4366__, new_new_n4367__, new_new_n4368__,
    new_new_n4369__, new_new_n4370__, new_new_n4372__, new_new_n4373__,
    new_new_n4374__, new_new_n4375__, new_new_n4376__, new_new_n4377__,
    new_new_n4378__, new_new_n4379__, new_new_n4380__, new_new_n4381__,
    new_new_n4382__, new_new_n4383__, new_new_n4384__, new_new_n4385__,
    new_new_n4386__, new_new_n4387__, new_new_n4388__, new_new_n4389__,
    new_new_n4390__, new_new_n4391__, new_new_n4392__, new_new_n4393__,
    new_new_n4394__, new_new_n4395__, new_new_n4396__, new_new_n4397__,
    new_new_n4398__, new_new_n4399__, new_new_n4400__, new_new_n4401__,
    new_new_n4402__, new_new_n4403__, new_new_n4404__, new_new_n4405__,
    new_new_n4406__, new_new_n4407__, new_new_n4408__, new_new_n4409__,
    new_new_n4410__, new_new_n4411__, new_new_n4412__, new_new_n4413__,
    new_new_n4414__, new_new_n4415__, new_new_n4416__, new_new_n4417__,
    new_new_n4418__, new_new_n4419__, new_new_n4420__, new_new_n4421__,
    new_new_n4422__, new_new_n4423__, new_new_n4424__, new_new_n4425__,
    new_new_n4426__, new_new_n4427__, new_new_n4428__, new_new_n4429__,
    new_new_n4430__, new_new_n4431__, new_new_n4432__, new_new_n4433__,
    new_new_n4434__, new_new_n4435__, new_new_n4436__, new_new_n4437__,
    new_new_n4438__, new_new_n4439__, new_new_n4440__, new_new_n4441__,
    new_new_n4442__, new_new_n4443__, new_new_n4444__, new_new_n4445__,
    new_new_n4446__, new_new_n4447__, new_new_n4448__, new_new_n4449__,
    new_new_n4450__, new_new_n4451__, new_new_n4452__, new_new_n4453__,
    new_new_n4454__, new_new_n4455__, new_new_n4456__, new_new_n4457__,
    new_new_n4458__, new_new_n4459__, new_new_n4460__, new_new_n4461__,
    new_new_n4462__, new_new_n4463__, new_new_n4464__, new_new_n4465__,
    new_new_n4466__, new_new_n4467__, new_new_n4468__, new_new_n4469__,
    new_new_n4470__, new_new_n4471__, new_new_n4472__, new_new_n4473__,
    new_new_n4474__, new_new_n4475__, new_new_n4476__, new_new_n4477__,
    new_new_n4478__, new_new_n4479__, new_new_n4480__, new_new_n4481__,
    new_new_n4482__, new_new_n4483__, new_new_n4484__, new_new_n4485__,
    new_new_n4486__, new_new_n4487__, new_new_n4488__, new_new_n4489__,
    new_new_n4490__, new_new_n4491__, new_new_n4492__, new_new_n4493__,
    new_new_n4494__, new_new_n4495__, new_new_n4496__, new_new_n4497__,
    new_new_n4498__, new_new_n4499__, new_new_n4500__, new_new_n4501__,
    new_new_n4502__, new_new_n4503__, new_new_n4504__, new_new_n4505__,
    new_new_n4506__, new_new_n4507__, new_new_n4508__, new_new_n4509__,
    new_new_n4510__, new_new_n4511__, new_new_n4512__, new_new_n4513__,
    new_new_n4514__, new_new_n4515__, new_new_n4516__, new_new_n4517__,
    new_new_n4518__, new_new_n4519__, new_new_n4520__, new_new_n4521__,
    new_new_n4522__, new_new_n4523__, new_new_n4524__, new_new_n4525__,
    new_new_n4526__, new_new_n4527__, new_new_n4528__, new_new_n4529__,
    new_new_n4530__, new_new_n4531__, new_new_n4532__, new_new_n4533__,
    new_new_n4534__, new_new_n4535__, new_new_n4536__, new_new_n4537__,
    new_new_n4538__, new_new_n4539__, new_new_n4540__, new_new_n4541__,
    new_new_n4542__, new_new_n4543__, new_new_n4544__, new_new_n4545__,
    new_new_n4546__, new_new_n4547__, new_new_n4548__, new_new_n4549__,
    new_new_n4550__, new_new_n4551__, new_new_n4552__, new_new_n4553__,
    new_new_n4554__, new_new_n4555__, new_new_n4556__, new_new_n4557__,
    new_new_n4558__, new_new_n4559__, new_new_n4560__, new_new_n4561__,
    new_new_n4562__, new_new_n4563__, new_new_n4564__, new_new_n4565__,
    new_new_n4566__, new_new_n4567__, new_new_n4568__, new_new_n4569__,
    new_new_n4570__, new_new_n4571__, new_new_n4572__, new_new_n4573__,
    new_new_n4574__, new_new_n4575__, new_new_n4576__, new_new_n4577__,
    new_new_n4578__, new_new_n4579__, new_new_n4581__, new_new_n4582__,
    new_new_n4583__, new_new_n4584__, new_new_n4585__, new_new_n4586__,
    new_new_n4587__, new_new_n4588__, new_new_n4589__, new_new_n4590__,
    new_new_n4591__, new_new_n4592__, new_new_n4593__, new_new_n4594__,
    new_new_n4595__, new_new_n4596__, new_new_n4597__, new_new_n4598__,
    new_new_n4599__, new_new_n4600__, new_new_n4601__, new_new_n4602__,
    new_new_n4603__, new_new_n4604__, new_new_n4605__, new_new_n4606__,
    new_new_n4607__, new_new_n4608__, new_new_n4609__, new_new_n4610__,
    new_new_n4611__, new_new_n4612__, new_new_n4613__, new_new_n4614__,
    new_new_n4615__, new_new_n4616__, new_new_n4617__, new_new_n4618__,
    new_new_n4619__, new_new_n4620__, new_new_n4621__, new_new_n4622__,
    new_new_n4623__, new_new_n4624__, new_new_n4625__, new_new_n4626__,
    new_new_n4627__, new_new_n4628__, new_new_n4629__, new_new_n4630__,
    new_new_n4631__, new_new_n4632__, new_new_n4633__, new_new_n4634__,
    new_new_n4635__, new_new_n4636__, new_new_n4637__, new_new_n4638__,
    new_new_n4639__, new_new_n4640__, new_new_n4641__, new_new_n4642__,
    new_new_n4643__, new_new_n4644__, new_new_n4645__, new_new_n4646__,
    new_new_n4647__, new_new_n4648__, new_new_n4649__, new_new_n4650__,
    new_new_n4651__, new_new_n4652__, new_new_n4653__, new_new_n4654__,
    new_new_n4655__, new_new_n4656__, new_new_n4657__, new_new_n4658__,
    new_new_n4659__, new_new_n4660__, new_new_n4661__, new_new_n4662__,
    new_new_n4663__, new_new_n4664__, new_new_n4665__, new_new_n4666__,
    new_new_n4667__, new_new_n4668__, new_new_n4669__, new_new_n4670__,
    new_new_n4671__, new_new_n4672__, new_new_n4673__, new_new_n4674__,
    new_new_n4675__, new_new_n4676__, new_new_n4677__, new_new_n4678__,
    new_new_n4679__, new_new_n4680__, new_new_n4681__, new_new_n4682__,
    new_new_n4683__, new_new_n4684__, new_new_n4685__, new_new_n4686__,
    new_new_n4687__, new_new_n4688__, new_new_n4689__, new_new_n4690__,
    new_new_n4691__, new_new_n4692__, new_new_n4693__, new_new_n4694__,
    new_new_n4695__, new_new_n4696__, new_new_n4697__, new_new_n4698__,
    new_new_n4699__, new_new_n4700__, new_new_n4701__, new_new_n4702__,
    new_new_n4703__, new_new_n4704__, new_new_n4705__, new_new_n4706__,
    new_new_n4707__, new_new_n4708__, new_new_n4709__, new_new_n4710__,
    new_new_n4711__, new_new_n4712__, new_new_n4713__, new_new_n4714__,
    new_new_n4715__, new_new_n4716__, new_new_n4717__, new_new_n4718__,
    new_new_n4719__, new_new_n4720__, new_new_n4721__, new_new_n4722__,
    new_new_n4723__, new_new_n4724__, new_new_n4725__, new_new_n4726__,
    new_new_n4727__, new_new_n4728__, new_new_n4729__, new_new_n4730__,
    new_new_n4731__, new_new_n4732__, new_new_n4733__, new_new_n4734__,
    new_new_n4735__, new_new_n4736__, new_new_n4737__, new_new_n4738__,
    new_new_n4739__, new_new_n4740__, new_new_n4741__, new_new_n4742__,
    new_new_n4743__, new_new_n4744__, new_new_n4745__, new_new_n4746__,
    new_new_n4747__, new_new_n4748__, new_new_n4749__, new_new_n4750__,
    new_new_n4751__, new_new_n4752__, new_new_n4753__, new_new_n4754__,
    new_new_n4755__, new_new_n4756__, new_new_n4757__, new_new_n4758__,
    new_new_n4759__, new_new_n4760__, new_new_n4761__, new_new_n4762__,
    new_new_n4763__, new_new_n4764__, new_new_n4765__, new_new_n4766__,
    new_new_n4767__, new_new_n4768__, new_new_n4769__, new_new_n4770__,
    new_new_n4771__, new_new_n4772__, new_new_n4774__, new_new_n4775__,
    new_new_n4776__, new_new_n4777__, new_new_n4778__, new_new_n4779__,
    new_new_n4780__, new_new_n4781__, new_new_n4782__, new_new_n4783__,
    new_new_n4784__, new_new_n4785__, new_new_n4786__, new_new_n4787__,
    new_new_n4788__, new_new_n4789__, new_new_n4790__, new_new_n4791__,
    new_new_n4792__, new_new_n4793__, new_new_n4794__, new_new_n4795__,
    new_new_n4796__, new_new_n4797__, new_new_n4798__, new_new_n4799__,
    new_new_n4800__, new_new_n4801__, new_new_n4802__, new_new_n4803__,
    new_new_n4804__, new_new_n4805__, new_new_n4806__, new_new_n4807__,
    new_new_n4808__, new_new_n4809__, new_new_n4810__, new_new_n4811__,
    new_new_n4812__, new_new_n4813__, new_new_n4814__, new_new_n4815__,
    new_new_n4816__, new_new_n4817__, new_new_n4818__, new_new_n4819__,
    new_new_n4820__, new_new_n4821__, new_new_n4822__, new_new_n4823__,
    new_new_n4824__, new_new_n4825__, new_new_n4826__, new_new_n4827__,
    new_new_n4828__, new_new_n4829__, new_new_n4830__, new_new_n4831__,
    new_new_n4832__, new_new_n4833__, new_new_n4834__, new_new_n4835__,
    new_new_n4836__, new_new_n4837__, new_new_n4838__, new_new_n4839__,
    new_new_n4840__, new_new_n4841__, new_new_n4842__, new_new_n4843__,
    new_new_n4844__, new_new_n4845__, new_new_n4846__, new_new_n4847__,
    new_new_n4848__, new_new_n4849__, new_new_n4850__, new_new_n4851__,
    new_new_n4852__, new_new_n4853__, new_new_n4854__, new_new_n4855__,
    new_new_n4856__, new_new_n4857__, new_new_n4858__, new_new_n4859__,
    new_new_n4860__, new_new_n4861__, new_new_n4862__, new_new_n4863__,
    new_new_n4864__, new_new_n4865__, new_new_n4866__, new_new_n4867__,
    new_new_n4868__, new_new_n4869__, new_new_n4870__, new_new_n4871__,
    new_new_n4872__, new_new_n4873__, new_new_n4874__, new_new_n4875__,
    new_new_n4876__, new_new_n4877__, new_new_n4878__, new_new_n4879__,
    new_new_n4880__, new_new_n4881__, new_new_n4882__, new_new_n4883__,
    new_new_n4884__, new_new_n4885__, new_new_n4886__, new_new_n4887__,
    new_new_n4888__, new_new_n4889__, new_new_n4890__, new_new_n4891__,
    new_new_n4892__, new_new_n4893__, new_new_n4894__, new_new_n4895__,
    new_new_n4896__, new_new_n4897__, new_new_n4898__, new_new_n4899__,
    new_new_n4900__, new_new_n4901__, new_new_n4902__, new_new_n4903__,
    new_new_n4904__, new_new_n4905__, new_new_n4906__, new_new_n4907__,
    new_new_n4908__, new_new_n4909__, new_new_n4910__, new_new_n4911__,
    new_new_n4912__, new_new_n4913__, new_new_n4914__, new_new_n4915__,
    new_new_n4916__, new_new_n4917__, new_new_n4918__, new_new_n4919__,
    new_new_n4920__, new_new_n4921__, new_new_n4922__, new_new_n4923__,
    new_new_n4924__, new_new_n4925__, new_new_n4926__, new_new_n4927__,
    new_new_n4928__, new_new_n4929__, new_new_n4930__, new_new_n4931__,
    new_new_n4932__, new_new_n4933__, new_new_n4934__, new_new_n4935__,
    new_new_n4936__, new_new_n4937__, new_new_n4938__, new_new_n4939__,
    new_new_n4940__, new_new_n4941__, new_new_n4942__, new_new_n4943__,
    new_new_n4944__, new_new_n4945__, new_new_n4946__, new_new_n4947__,
    new_new_n4948__, new_new_n4949__, new_new_n4950__, new_new_n4951__,
    new_new_n4952__, new_new_n4953__, new_new_n4954__, new_new_n4955__,
    new_new_n4956__, new_new_n4957__, new_new_n4958__, new_new_n4959__,
    new_new_n4960__, new_new_n4961__, new_new_n4962__, new_new_n4963__,
    new_new_n4964__, new_new_n4965__, new_new_n4966__, new_new_n4967__,
    new_new_n4968__, new_new_n4969__, new_new_n4970__, new_new_n4971__,
    new_new_n4972__, new_new_n4973__, new_new_n4974__, new_new_n4975__,
    new_new_n4976__, new_new_n4977__, new_new_n4978__, new_new_n4979__,
    new_new_n4980__, new_new_n4981__, new_new_n4982__, new_new_n4983__,
    new_new_n4984__, new_new_n4985__, new_new_n4986__, new_new_n4987__,
    new_new_n4988__, new_new_n4989__, new_new_n4990__, new_new_n4991__,
    new_new_n4992__, new_new_n4993__, new_new_n4994__, new_new_n4995__,
    new_new_n4996__, new_new_n4997__, new_new_n4998__, new_new_n4999__,
    new_new_n5000__, new_new_n5001__, new_new_n5002__, new_new_n5004__,
    new_new_n5005__, new_new_n5006__, new_new_n5007__, new_new_n5008__,
    new_new_n5009__, new_new_n5010__, new_new_n5011__, new_new_n5012__,
    new_new_n5013__, new_new_n5014__, new_new_n5015__, new_new_n5016__,
    new_new_n5017__, new_new_n5018__, new_new_n5019__, new_new_n5020__,
    new_new_n5021__, new_new_n5022__, new_new_n5023__, new_new_n5024__,
    new_new_n5025__, new_new_n5026__, new_new_n5027__, new_new_n5028__,
    new_new_n5029__, new_new_n5030__, new_new_n5031__, new_new_n5032__,
    new_new_n5033__, new_new_n5034__, new_new_n5035__, new_new_n5036__,
    new_new_n5037__, new_new_n5038__, new_new_n5039__, new_new_n5040__,
    new_new_n5041__, new_new_n5042__, new_new_n5043__, new_new_n5044__,
    new_new_n5045__, new_new_n5046__, new_new_n5047__, new_new_n5048__,
    new_new_n5049__, new_new_n5050__, new_new_n5051__, new_new_n5052__,
    new_new_n5053__, new_new_n5054__, new_new_n5055__, new_new_n5056__,
    new_new_n5057__, new_new_n5058__, new_new_n5059__, new_new_n5060__,
    new_new_n5061__, new_new_n5062__, new_new_n5063__, new_new_n5064__,
    new_new_n5065__, new_new_n5066__, new_new_n5067__, new_new_n5068__,
    new_new_n5069__, new_new_n5070__, new_new_n5071__, new_new_n5072__,
    new_new_n5073__, new_new_n5074__, new_new_n5075__, new_new_n5076__,
    new_new_n5077__, new_new_n5078__, new_new_n5079__, new_new_n5080__,
    new_new_n5081__, new_new_n5082__, new_new_n5083__, new_new_n5084__,
    new_new_n5085__, new_new_n5086__, new_new_n5087__, new_new_n5088__,
    new_new_n5089__, new_new_n5090__, new_new_n5091__, new_new_n5092__,
    new_new_n5093__, new_new_n5094__, new_new_n5095__, new_new_n5096__,
    new_new_n5097__, new_new_n5098__, new_new_n5099__, new_new_n5100__,
    new_new_n5101__, new_new_n5102__, new_new_n5103__, new_new_n5104__,
    new_new_n5105__, new_new_n5106__, new_new_n5107__, new_new_n5108__,
    new_new_n5109__, new_new_n5110__, new_new_n5111__, new_new_n5112__,
    new_new_n5113__, new_new_n5114__, new_new_n5115__, new_new_n5116__,
    new_new_n5117__, new_new_n5118__, new_new_n5119__, new_new_n5120__,
    new_new_n5121__, new_new_n5122__, new_new_n5123__, new_new_n5124__,
    new_new_n5125__, new_new_n5126__, new_new_n5127__, new_new_n5128__,
    new_new_n5129__, new_new_n5130__, new_new_n5131__, new_new_n5132__,
    new_new_n5133__, new_new_n5134__, new_new_n5135__, new_new_n5136__,
    new_new_n5137__, new_new_n5138__, new_new_n5139__, new_new_n5140__,
    new_new_n5141__, new_new_n5142__, new_new_n5143__, new_new_n5144__,
    new_new_n5145__, new_new_n5146__, new_new_n5147__, new_new_n5148__,
    new_new_n5149__, new_new_n5150__, new_new_n5151__, new_new_n5152__,
    new_new_n5153__, new_new_n5154__, new_new_n5155__, new_new_n5156__,
    new_new_n5157__, new_new_n5158__, new_new_n5159__, new_new_n5160__,
    new_new_n5161__, new_new_n5162__, new_new_n5163__, new_new_n5164__,
    new_new_n5165__, new_new_n5166__, new_new_n5167__, new_new_n5168__,
    new_new_n5169__, new_new_n5170__, new_new_n5171__, new_new_n5172__,
    new_new_n5173__, new_new_n5174__, new_new_n5175__, new_new_n5176__,
    new_new_n5177__, new_new_n5178__, new_new_n5179__, new_new_n5180__,
    new_new_n5181__, new_new_n5182__, new_new_n5183__, new_new_n5184__,
    new_new_n5185__, new_new_n5186__, new_new_n5187__, new_new_n5188__,
    new_new_n5189__, new_new_n5190__, new_new_n5191__, new_new_n5192__,
    new_new_n5193__, new_new_n5194__, new_new_n5195__, new_new_n5196__,
    new_new_n5197__, new_new_n5198__, new_new_n5199__, new_new_n5200__,
    new_new_n5201__, new_new_n5202__, new_new_n5203__, new_new_n5204__,
    new_new_n5205__, new_new_n5207__, new_new_n5208__, new_new_n5209__,
    new_new_n5210__, new_new_n5211__, new_new_n5212__, new_new_n5213__,
    new_new_n5214__, new_new_n5215__, new_new_n5216__, new_new_n5217__,
    new_new_n5218__, new_new_n5219__, new_new_n5220__, new_new_n5221__,
    new_new_n5222__, new_new_n5223__, new_new_n5224__, new_new_n5225__,
    new_new_n5226__, new_new_n5227__, new_new_n5228__, new_new_n5229__,
    new_new_n5230__, new_new_n5231__, new_new_n5232__, new_new_n5233__,
    new_new_n5234__, new_new_n5235__, new_new_n5236__, new_new_n5237__,
    new_new_n5238__, new_new_n5239__, new_new_n5240__, new_new_n5241__,
    new_new_n5242__, new_new_n5243__, new_new_n5244__, new_new_n5245__,
    new_new_n5246__, new_new_n5247__, new_new_n5248__, new_new_n5249__,
    new_new_n5250__, new_new_n5251__, new_new_n5252__, new_new_n5253__,
    new_new_n5254__, new_new_n5255__, new_new_n5256__, new_new_n5257__,
    new_new_n5258__, new_new_n5259__, new_new_n5260__, new_new_n5261__,
    new_new_n5262__, new_new_n5263__, new_new_n5264__, new_new_n5265__,
    new_new_n5266__, new_new_n5267__, new_new_n5268__, new_new_n5269__,
    new_new_n5270__, new_new_n5271__, new_new_n5272__, new_new_n5273__,
    new_new_n5274__, new_new_n5275__, new_new_n5276__, new_new_n5277__,
    new_new_n5278__, new_new_n5279__, new_new_n5280__, new_new_n5281__,
    new_new_n5282__, new_new_n5283__, new_new_n5284__, new_new_n5285__,
    new_new_n5286__, new_new_n5287__, new_new_n5288__, new_new_n5289__,
    new_new_n5290__, new_new_n5291__, new_new_n5292__, new_new_n5293__,
    new_new_n5294__, new_new_n5295__, new_new_n5296__, new_new_n5297__,
    new_new_n5298__, new_new_n5299__, new_new_n5300__, new_new_n5301__,
    new_new_n5302__, new_new_n5303__, new_new_n5304__, new_new_n5305__,
    new_new_n5306__, new_new_n5307__, new_new_n5308__, new_new_n5309__,
    new_new_n5310__, new_new_n5311__, new_new_n5312__, new_new_n5313__,
    new_new_n5314__, new_new_n5315__, new_new_n5316__, new_new_n5317__,
    new_new_n5318__, new_new_n5319__, new_new_n5320__, new_new_n5321__,
    new_new_n5322__, new_new_n5323__, new_new_n5324__, new_new_n5325__,
    new_new_n5326__, new_new_n5327__, new_new_n5328__, new_new_n5329__,
    new_new_n5330__, new_new_n5331__, new_new_n5332__, new_new_n5333__,
    new_new_n5334__, new_new_n5335__, new_new_n5336__, new_new_n5337__,
    new_new_n5338__, new_new_n5339__, new_new_n5340__, new_new_n5341__,
    new_new_n5342__, new_new_n5343__, new_new_n5344__, new_new_n5345__,
    new_new_n5346__, new_new_n5347__, new_new_n5348__, new_new_n5349__,
    new_new_n5350__, new_new_n5351__, new_new_n5352__, new_new_n5353__,
    new_new_n5354__, new_new_n5355__, new_new_n5356__, new_new_n5357__,
    new_new_n5358__, new_new_n5359__, new_new_n5360__, new_new_n5361__,
    new_new_n5362__, new_new_n5363__, new_new_n5364__, new_new_n5365__,
    new_new_n5366__, new_new_n5367__, new_new_n5368__, new_new_n5369__,
    new_new_n5370__, new_new_n5371__, new_new_n5372__, new_new_n5373__,
    new_new_n5374__, new_new_n5375__, new_new_n5376__, new_new_n5377__,
    new_new_n5378__, new_new_n5379__, new_new_n5380__, new_new_n5381__,
    new_new_n5382__, new_new_n5383__, new_new_n5384__, new_new_n5385__,
    new_new_n5386__, new_new_n5387__, new_new_n5388__, new_new_n5389__,
    new_new_n5390__, new_new_n5391__, new_new_n5392__, new_new_n5393__,
    new_new_n5394__, new_new_n5395__, new_new_n5396__, new_new_n5397__,
    new_new_n5398__, new_new_n5399__, new_new_n5400__, new_new_n5401__,
    new_new_n5402__, new_new_n5403__, new_new_n5404__, new_new_n5405__,
    new_new_n5406__, new_new_n5407__, new_new_n5408__, new_new_n5409__,
    new_new_n5410__, new_new_n5411__, new_new_n5412__, new_new_n5413__,
    new_new_n5414__, new_new_n5415__, new_new_n5416__, new_new_n5417__,
    new_new_n5418__, new_new_n5419__, new_new_n5420__, new_new_n5421__,
    new_new_n5422__, new_new_n5423__, new_new_n5424__, new_new_n5425__,
    new_new_n5426__, new_new_n5427__, new_new_n5429__, new_new_n5430__,
    new_new_n5431__, new_new_n5432__, new_new_n5433__, new_new_n5434__,
    new_new_n5435__, new_new_n5436__, new_new_n5437__, new_new_n5438__,
    new_new_n5439__, new_new_n5440__, new_new_n5441__, new_new_n5442__,
    new_new_n5443__, new_new_n5444__, new_new_n5445__, new_new_n5446__,
    new_new_n5447__, new_new_n5448__, new_new_n5449__, new_new_n5450__,
    new_new_n5451__, new_new_n5452__, new_new_n5453__, new_new_n5454__,
    new_new_n5455__, new_new_n5456__, new_new_n5457__, new_new_n5458__,
    new_new_n5459__, new_new_n5460__, new_new_n5461__, new_new_n5462__,
    new_new_n5463__, new_new_n5464__, new_new_n5465__, new_new_n5466__,
    new_new_n5467__, new_new_n5468__, new_new_n5469__, new_new_n5470__,
    new_new_n5471__, new_new_n5472__, new_new_n5473__, new_new_n5474__,
    new_new_n5475__, new_new_n5476__, new_new_n5477__, new_new_n5478__,
    new_new_n5479__, new_new_n5480__, new_new_n5481__, new_new_n5482__,
    new_new_n5483__, new_new_n5484__, new_new_n5485__, new_new_n5486__,
    new_new_n5487__, new_new_n5488__, new_new_n5489__, new_new_n5490__,
    new_new_n5491__, new_new_n5492__, new_new_n5493__, new_new_n5494__,
    new_new_n5495__, new_new_n5496__, new_new_n5497__, new_new_n5498__,
    new_new_n5499__, new_new_n5500__, new_new_n5501__, new_new_n5502__,
    new_new_n5503__, new_new_n5504__, new_new_n5505__, new_new_n5506__,
    new_new_n5507__, new_new_n5508__, new_new_n5509__, new_new_n5510__,
    new_new_n5511__, new_new_n5512__, new_new_n5513__, new_new_n5514__,
    new_new_n5515__, new_new_n5516__, new_new_n5517__, new_new_n5518__,
    new_new_n5519__, new_new_n5520__, new_new_n5521__, new_new_n5522__,
    new_new_n5523__, new_new_n5524__, new_new_n5525__, new_new_n5526__,
    new_new_n5527__, new_new_n5528__, new_new_n5529__, new_new_n5530__,
    new_new_n5531__, new_new_n5532__, new_new_n5533__, new_new_n5534__,
    new_new_n5535__, new_new_n5536__, new_new_n5537__, new_new_n5538__,
    new_new_n5539__, new_new_n5540__, new_new_n5541__, new_new_n5542__,
    new_new_n5543__, new_new_n5544__, new_new_n5545__, new_new_n5546__,
    new_new_n5547__, new_new_n5548__, new_new_n5549__, new_new_n5550__,
    new_new_n5551__, new_new_n5552__, new_new_n5553__, new_new_n5554__,
    new_new_n5555__, new_new_n5556__, new_new_n5557__, new_new_n5558__,
    new_new_n5559__, new_new_n5560__, new_new_n5561__, new_new_n5562__,
    new_new_n5563__, new_new_n5564__, new_new_n5565__, new_new_n5566__,
    new_new_n5567__, new_new_n5568__, new_new_n5569__, new_new_n5570__,
    new_new_n5571__, new_new_n5572__, new_new_n5573__, new_new_n5574__,
    new_new_n5575__, new_new_n5576__, new_new_n5577__, new_new_n5578__,
    new_new_n5579__, new_new_n5580__, new_new_n5581__, new_new_n5582__,
    new_new_n5583__, new_new_n5584__, new_new_n5585__, new_new_n5586__,
    new_new_n5587__, new_new_n5588__, new_new_n5589__, new_new_n5590__,
    new_new_n5591__, new_new_n5592__, new_new_n5593__, new_new_n5594__,
    new_new_n5595__, new_new_n5596__, new_new_n5597__, new_new_n5598__,
    new_new_n5599__, new_new_n5600__, new_new_n5601__, new_new_n5602__,
    new_new_n5603__, new_new_n5604__, new_new_n5605__, new_new_n5606__,
    new_new_n5607__, new_new_n5608__, new_new_n5609__, new_new_n5610__,
    new_new_n5611__, new_new_n5612__, new_new_n5613__, new_new_n5614__,
    new_new_n5615__, new_new_n5616__, new_new_n5617__, new_new_n5618__,
    new_new_n5619__, new_new_n5620__, new_new_n5621__, new_new_n5622__,
    new_new_n5623__, new_new_n5624__, new_new_n5625__, new_new_n5626__,
    new_new_n5627__, new_new_n5628__, new_new_n5629__, new_new_n5630__,
    new_new_n5631__, new_new_n5632__, new_new_n5633__, new_new_n5634__,
    new_new_n5635__, new_new_n5636__, new_new_n5637__, new_new_n5638__,
    new_new_n5639__, new_new_n5640__, new_new_n5641__, new_new_n5642__,
    new_new_n5643__, new_new_n5644__, new_new_n5645__, new_new_n5646__,
    new_new_n5648__, new_new_n5649__, new_new_n5650__, new_new_n5651__,
    new_new_n5652__, new_new_n5653__, new_new_n5654__, new_new_n5655__,
    new_new_n5656__, new_new_n5657__, new_new_n5658__, new_new_n5659__,
    new_new_n5660__, new_new_n5661__, new_new_n5662__, new_new_n5663__,
    new_new_n5664__, new_new_n5665__, new_new_n5666__, new_new_n5667__,
    new_new_n5668__, new_new_n5669__, new_new_n5670__, new_new_n5671__,
    new_new_n5672__, new_new_n5673__, new_new_n5674__, new_new_n5675__,
    new_new_n5676__, new_new_n5677__, new_new_n5678__, new_new_n5679__,
    new_new_n5680__, new_new_n5681__, new_new_n5682__, new_new_n5683__,
    new_new_n5684__, new_new_n5685__, new_new_n5686__, new_new_n5687__,
    new_new_n5688__, new_new_n5689__, new_new_n5690__, new_new_n5691__,
    new_new_n5692__, new_new_n5693__, new_new_n5694__, new_new_n5695__,
    new_new_n5696__, new_new_n5697__, new_new_n5698__, new_new_n5699__,
    new_new_n5700__, new_new_n5701__, new_new_n5702__, new_new_n5703__,
    new_new_n5704__, new_new_n5705__, new_new_n5706__, new_new_n5707__,
    new_new_n5708__, new_new_n5709__, new_new_n5710__, new_new_n5711__,
    new_new_n5712__, new_new_n5713__, new_new_n5714__, new_new_n5715__,
    new_new_n5716__, new_new_n5717__, new_new_n5718__, new_new_n5719__,
    new_new_n5720__, new_new_n5721__, new_new_n5722__, new_new_n5723__,
    new_new_n5724__, new_new_n5725__, new_new_n5726__, new_new_n5727__,
    new_new_n5728__, new_new_n5729__, new_new_n5730__, new_new_n5731__,
    new_new_n5732__, new_new_n5733__, new_new_n5734__, new_new_n5735__,
    new_new_n5736__, new_new_n5737__, new_new_n5738__, new_new_n5739__,
    new_new_n5740__, new_new_n5741__, new_new_n5742__, new_new_n5743__,
    new_new_n5744__, new_new_n5745__, new_new_n5746__, new_new_n5747__,
    new_new_n5748__, new_new_n5749__, new_new_n5750__, new_new_n5751__,
    new_new_n5752__, new_new_n5753__, new_new_n5754__, new_new_n5755__,
    new_new_n5756__, new_new_n5757__, new_new_n5758__, new_new_n5759__,
    new_new_n5760__, new_new_n5761__, new_new_n5762__, new_new_n5763__,
    new_new_n5764__, new_new_n5765__, new_new_n5766__, new_new_n5767__,
    new_new_n5768__, new_new_n5769__, new_new_n5770__, new_new_n5771__,
    new_new_n5772__, new_new_n5773__, new_new_n5774__, new_new_n5775__,
    new_new_n5776__, new_new_n5777__, new_new_n5778__, new_new_n5779__,
    new_new_n5780__, new_new_n5781__, new_new_n5782__, new_new_n5783__,
    new_new_n5784__, new_new_n5785__, new_new_n5786__, new_new_n5787__,
    new_new_n5788__, new_new_n5789__, new_new_n5790__, new_new_n5791__,
    new_new_n5792__, new_new_n5793__, new_new_n5794__, new_new_n5795__,
    new_new_n5796__, new_new_n5797__, new_new_n5798__, new_new_n5799__,
    new_new_n5800__, new_new_n5801__, new_new_n5802__, new_new_n5803__,
    new_new_n5804__, new_new_n5805__, new_new_n5806__, new_new_n5807__,
    new_new_n5808__, new_new_n5809__, new_new_n5810__, new_new_n5811__,
    new_new_n5812__, new_new_n5813__, new_new_n5814__, new_new_n5815__,
    new_new_n5816__, new_new_n5817__, new_new_n5818__, new_new_n5819__,
    new_new_n5820__, new_new_n5821__, new_new_n5822__, new_new_n5823__,
    new_new_n5824__, new_new_n5825__, new_new_n5826__, new_new_n5827__,
    new_new_n5828__, new_new_n5829__, new_new_n5830__, new_new_n5831__,
    new_new_n5832__, new_new_n5833__, new_new_n5834__, new_new_n5835__,
    new_new_n5836__, new_new_n5837__, new_new_n5838__, new_new_n5839__,
    new_new_n5840__, new_new_n5841__, new_new_n5842__, new_new_n5843__,
    new_new_n5844__, new_new_n5845__, new_new_n5846__, new_new_n5847__,
    new_new_n5848__, new_new_n5849__, new_new_n5850__, new_new_n5851__,
    new_new_n5852__, new_new_n5853__, new_new_n5854__, new_new_n5855__,
    new_new_n5856__, new_new_n5857__, new_new_n5858__, new_new_n5859__,
    new_new_n5860__, new_new_n5861__, new_new_n5862__, new_new_n5863__,
    new_new_n5864__, new_new_n5865__, new_new_n5866__, new_new_n5867__,
    new_new_n5868__, new_new_n5869__, new_new_n5870__, new_new_n5871__,
    new_new_n5872__, new_new_n5873__, new_new_n5874__, new_new_n5875__,
    new_new_n5876__, new_new_n5877__, new_new_n5878__, new_new_n5879__,
    new_new_n5880__, new_new_n5881__, new_new_n5882__, new_new_n5883__,
    new_new_n5884__, new_new_n5885__, new_new_n5886__, new_new_n5887__,
    new_new_n5888__, new_new_n5890__, new_new_n5891__, new_new_n5892__,
    new_new_n5893__, new_new_n5894__, new_new_n5895__, new_new_n5896__,
    new_new_n5897__, new_new_n5898__, new_new_n5899__, new_new_n5900__,
    new_new_n5901__, new_new_n5902__, new_new_n5903__, new_new_n5904__,
    new_new_n5905__, new_new_n5906__, new_new_n5907__, new_new_n5908__,
    new_new_n5909__, new_new_n5910__, new_new_n5911__, new_new_n5912__,
    new_new_n5913__, new_new_n5914__, new_new_n5915__, new_new_n5916__,
    new_new_n5917__, new_new_n5918__, new_new_n5919__, new_new_n5920__,
    new_new_n5921__, new_new_n5922__, new_new_n5923__, new_new_n5924__,
    new_new_n5925__, new_new_n5926__, new_new_n5927__, new_new_n5928__,
    new_new_n5929__, new_new_n5930__, new_new_n5931__, new_new_n5932__,
    new_new_n5933__, new_new_n5934__, new_new_n5935__, new_new_n5936__,
    new_new_n5937__, new_new_n5938__, new_new_n5939__, new_new_n5940__,
    new_new_n5941__, new_new_n5942__, new_new_n5943__, new_new_n5944__,
    new_new_n5945__, new_new_n5946__, new_new_n5947__, new_new_n5948__,
    new_new_n5949__, new_new_n5950__, new_new_n5951__, new_new_n5952__,
    new_new_n5953__, new_new_n5954__, new_new_n5955__, new_new_n5956__,
    new_new_n5957__, new_new_n5958__, new_new_n5959__, new_new_n5960__,
    new_new_n5961__, new_new_n5962__, new_new_n5963__, new_new_n5964__,
    new_new_n5965__, new_new_n5966__, new_new_n5967__, new_new_n5968__,
    new_new_n5969__, new_new_n5970__, new_new_n5971__, new_new_n5972__,
    new_new_n5973__, new_new_n5974__, new_new_n5975__, new_new_n5976__,
    new_new_n5977__, new_new_n5978__, new_new_n5979__, new_new_n5980__,
    new_new_n5981__, new_new_n5982__, new_new_n5983__, new_new_n5984__,
    new_new_n5985__, new_new_n5986__, new_new_n5987__, new_new_n5988__,
    new_new_n5989__, new_new_n5990__, new_new_n5991__, new_new_n5992__,
    new_new_n5993__, new_new_n5994__, new_new_n5995__, new_new_n5996__,
    new_new_n5997__, new_new_n5998__, new_new_n5999__, new_new_n6000__,
    new_new_n6001__, new_new_n6002__, new_new_n6003__, new_new_n6004__,
    new_new_n6005__, new_new_n6006__, new_new_n6007__, new_new_n6008__,
    new_new_n6009__, new_new_n6010__, new_new_n6011__, new_new_n6012__,
    new_new_n6013__, new_new_n6014__, new_new_n6015__, new_new_n6016__,
    new_new_n6017__, new_new_n6018__, new_new_n6019__, new_new_n6020__,
    new_new_n6021__, new_new_n6022__, new_new_n6023__, new_new_n6024__,
    new_new_n6025__, new_new_n6026__, new_new_n6027__, new_new_n6028__,
    new_new_n6029__, new_new_n6030__, new_new_n6031__, new_new_n6032__,
    new_new_n6033__, new_new_n6034__, new_new_n6035__, new_new_n6036__,
    new_new_n6037__, new_new_n6038__, new_new_n6039__, new_new_n6040__,
    new_new_n6041__, new_new_n6042__, new_new_n6043__, new_new_n6044__,
    new_new_n6045__, new_new_n6046__, new_new_n6047__, new_new_n6048__,
    new_new_n6049__, new_new_n6050__, new_new_n6051__, new_new_n6052__,
    new_new_n6053__, new_new_n6054__, new_new_n6055__, new_new_n6056__,
    new_new_n6057__, new_new_n6058__, new_new_n6059__, new_new_n6060__,
    new_new_n6061__, new_new_n6062__, new_new_n6063__, new_new_n6064__,
    new_new_n6065__, new_new_n6066__, new_new_n6067__, new_new_n6068__,
    new_new_n6069__, new_new_n6070__, new_new_n6071__, new_new_n6072__,
    new_new_n6073__, new_new_n6074__, new_new_n6075__, new_new_n6076__,
    new_new_n6077__, new_new_n6078__, new_new_n6079__, new_new_n6080__,
    new_new_n6081__, new_new_n6082__, new_new_n6083__, new_new_n6084__,
    new_new_n6085__, new_new_n6086__, new_new_n6087__, new_new_n6088__,
    new_new_n6089__, new_new_n6090__, new_new_n6091__, new_new_n6092__,
    new_new_n6093__, new_new_n6094__, new_new_n6095__, new_new_n6096__,
    new_new_n6097__, new_new_n6098__, new_new_n6099__, new_new_n6100__,
    new_new_n6101__, new_new_n6102__, new_new_n6103__, new_new_n6104__,
    new_new_n6105__, new_new_n6106__, new_new_n6107__, new_new_n6108__,
    new_new_n6109__, new_new_n6110__, new_new_n6111__, new_new_n6112__,
    new_new_n6113__, new_new_n6115__, new_new_n6116__, new_new_n6117__,
    new_new_n6118__, new_new_n6119__, new_new_n6120__, new_new_n6121__,
    new_new_n6122__, new_new_n6123__, new_new_n6124__, new_new_n6125__,
    new_new_n6126__, new_new_n6127__, new_new_n6128__, new_new_n6129__,
    new_new_n6130__, new_new_n6131__, new_new_n6132__, new_new_n6133__,
    new_new_n6134__, new_new_n6135__, new_new_n6136__, new_new_n6137__,
    new_new_n6138__, new_new_n6139__, new_new_n6140__, new_new_n6141__,
    new_new_n6142__, new_new_n6143__, new_new_n6144__, new_new_n6145__,
    new_new_n6146__, new_new_n6147__, new_new_n6148__, new_new_n6149__,
    new_new_n6150__, new_new_n6151__, new_new_n6152__, new_new_n6153__,
    new_new_n6154__, new_new_n6155__, new_new_n6156__, new_new_n6157__,
    new_new_n6158__, new_new_n6159__, new_new_n6160__, new_new_n6161__,
    new_new_n6162__, new_new_n6163__, new_new_n6164__, new_new_n6165__,
    new_new_n6166__, new_new_n6167__, new_new_n6168__, new_new_n6169__,
    new_new_n6170__, new_new_n6171__, new_new_n6172__, new_new_n6173__,
    new_new_n6174__, new_new_n6175__, new_new_n6176__, new_new_n6177__,
    new_new_n6178__, new_new_n6179__, new_new_n6180__, new_new_n6181__,
    new_new_n6182__, new_new_n6183__, new_new_n6184__, new_new_n6185__,
    new_new_n6186__, new_new_n6187__, new_new_n6188__, new_new_n6189__,
    new_new_n6190__, new_new_n6191__, new_new_n6192__, new_new_n6193__,
    new_new_n6194__, new_new_n6195__, new_new_n6196__, new_new_n6197__,
    new_new_n6198__, new_new_n6199__, new_new_n6200__, new_new_n6201__,
    new_new_n6202__, new_new_n6203__, new_new_n6204__, new_new_n6205__,
    new_new_n6206__, new_new_n6207__, new_new_n6208__, new_new_n6209__,
    new_new_n6210__, new_new_n6211__, new_new_n6212__, new_new_n6213__,
    new_new_n6214__, new_new_n6215__, new_new_n6216__, new_new_n6217__,
    new_new_n6218__, new_new_n6219__, new_new_n6220__, new_new_n6221__,
    new_new_n6222__, new_new_n6223__, new_new_n6224__, new_new_n6225__,
    new_new_n6226__, new_new_n6227__, new_new_n6228__, new_new_n6229__,
    new_new_n6230__, new_new_n6231__, new_new_n6232__, new_new_n6233__,
    new_new_n6234__, new_new_n6235__, new_new_n6236__, new_new_n6237__,
    new_new_n6238__, new_new_n6239__, new_new_n6240__, new_new_n6241__,
    new_new_n6242__, new_new_n6243__, new_new_n6244__, new_new_n6245__,
    new_new_n6246__, new_new_n6247__, new_new_n6248__, new_new_n6249__,
    new_new_n6250__, new_new_n6251__, new_new_n6252__, new_new_n6253__,
    new_new_n6254__, new_new_n6255__, new_new_n6256__, new_new_n6257__,
    new_new_n6258__, new_new_n6259__, new_new_n6260__, new_new_n6261__,
    new_new_n6262__, new_new_n6263__, new_new_n6264__, new_new_n6265__,
    new_new_n6266__, new_new_n6267__, new_new_n6268__, new_new_n6269__,
    new_new_n6270__, new_new_n6271__, new_new_n6272__, new_new_n6273__,
    new_new_n6274__, new_new_n6275__, new_new_n6276__, new_new_n6277__,
    new_new_n6278__, new_new_n6279__, new_new_n6280__, new_new_n6281__,
    new_new_n6282__, new_new_n6283__, new_new_n6284__, new_new_n6285__,
    new_new_n6286__, new_new_n6287__, new_new_n6288__, new_new_n6289__,
    new_new_n6290__, new_new_n6291__, new_new_n6292__, new_new_n6293__,
    new_new_n6294__, new_new_n6295__, new_new_n6296__, new_new_n6297__,
    new_new_n6298__, new_new_n6299__, new_new_n6300__, new_new_n6301__,
    new_new_n6302__, new_new_n6303__, new_new_n6304__, new_new_n6305__,
    new_new_n6306__, new_new_n6307__, new_new_n6308__, new_new_n6309__,
    new_new_n6310__, new_new_n6311__, new_new_n6312__, new_new_n6313__,
    new_new_n6314__, new_new_n6315__, new_new_n6316__, new_new_n6317__,
    new_new_n6318__, new_new_n6319__, new_new_n6320__, new_new_n6321__,
    new_new_n6322__, new_new_n6323__, new_new_n6324__, new_new_n6325__,
    new_new_n6326__, new_new_n6327__, new_new_n6328__, new_new_n6329__,
    new_new_n6330__, new_new_n6331__, new_new_n6332__, new_new_n6333__,
    new_new_n6334__, new_new_n6335__, new_new_n6336__, new_new_n6337__,
    new_new_n6338__, new_new_n6339__, new_new_n6340__, new_new_n6341__,
    new_new_n6342__, new_new_n6343__, new_new_n6344__, new_new_n6345__,
    new_new_n6346__, new_new_n6347__, new_new_n6348__, new_new_n6349__,
    new_new_n6350__, new_new_n6351__, new_new_n6353__, new_new_n6354__,
    new_new_n6355__, new_new_n6356__, new_new_n6357__, new_new_n6358__,
    new_new_n6359__, new_new_n6360__, new_new_n6361__, new_new_n6362__,
    new_new_n6363__, new_new_n6364__, new_new_n6365__, new_new_n6366__,
    new_new_n6367__, new_new_n6368__, new_new_n6369__, new_new_n6370__,
    new_new_n6371__, new_new_n6372__, new_new_n6373__, new_new_n6374__,
    new_new_n6375__, new_new_n6376__, new_new_n6377__, new_new_n6378__,
    new_new_n6379__, new_new_n6380__, new_new_n6381__, new_new_n6382__,
    new_new_n6383__, new_new_n6384__, new_new_n6385__, new_new_n6386__,
    new_new_n6387__, new_new_n6388__, new_new_n6389__, new_new_n6390__,
    new_new_n6391__, new_new_n6392__, new_new_n6393__, new_new_n6394__,
    new_new_n6395__, new_new_n6396__, new_new_n6397__, new_new_n6398__,
    new_new_n6399__, new_new_n6400__, new_new_n6401__, new_new_n6402__,
    new_new_n6403__, new_new_n6404__, new_new_n6405__, new_new_n6406__,
    new_new_n6407__, new_new_n6408__, new_new_n6409__, new_new_n6410__,
    new_new_n6411__, new_new_n6412__, new_new_n6413__, new_new_n6414__,
    new_new_n6415__, new_new_n6416__, new_new_n6417__, new_new_n6418__,
    new_new_n6419__, new_new_n6420__, new_new_n6421__, new_new_n6422__,
    new_new_n6423__, new_new_n6424__, new_new_n6425__, new_new_n6426__,
    new_new_n6427__, new_new_n6428__, new_new_n6429__, new_new_n6430__,
    new_new_n6431__, new_new_n6432__, new_new_n6433__, new_new_n6434__,
    new_new_n6435__, new_new_n6436__, new_new_n6437__, new_new_n6438__,
    new_new_n6439__, new_new_n6440__, new_new_n6441__, new_new_n6442__,
    new_new_n6443__, new_new_n6444__, new_new_n6445__, new_new_n6446__,
    new_new_n6447__, new_new_n6448__, new_new_n6449__, new_new_n6450__,
    new_new_n6451__, new_new_n6452__, new_new_n6453__, new_new_n6454__,
    new_new_n6455__, new_new_n6456__, new_new_n6457__, new_new_n6458__,
    new_new_n6459__, new_new_n6460__, new_new_n6461__, new_new_n6462__,
    new_new_n6463__, new_new_n6464__, new_new_n6465__, new_new_n6466__,
    new_new_n6467__, new_new_n6468__, new_new_n6469__, new_new_n6470__,
    new_new_n6471__, new_new_n6472__, new_new_n6473__, new_new_n6474__,
    new_new_n6475__, new_new_n6476__, new_new_n6477__, new_new_n6478__,
    new_new_n6479__, new_new_n6480__, new_new_n6481__, new_new_n6482__,
    new_new_n6483__, new_new_n6484__, new_new_n6485__, new_new_n6486__,
    new_new_n6487__, new_new_n6488__, new_new_n6489__, new_new_n6490__,
    new_new_n6491__, new_new_n6492__, new_new_n6493__, new_new_n6494__,
    new_new_n6495__, new_new_n6496__, new_new_n6497__, new_new_n6498__,
    new_new_n6499__, new_new_n6500__, new_new_n6501__, new_new_n6502__,
    new_new_n6503__, new_new_n6504__, new_new_n6505__, new_new_n6506__,
    new_new_n6507__, new_new_n6508__, new_new_n6509__, new_new_n6510__,
    new_new_n6511__, new_new_n6512__, new_new_n6513__, new_new_n6514__,
    new_new_n6515__, new_new_n6516__, new_new_n6517__, new_new_n6518__,
    new_new_n6519__, new_new_n6520__, new_new_n6521__, new_new_n6522__,
    new_new_n6523__, new_new_n6524__, new_new_n6525__, new_new_n6526__,
    new_new_n6527__, new_new_n6528__, new_new_n6529__, new_new_n6530__,
    new_new_n6531__, new_new_n6532__, new_new_n6533__, new_new_n6534__,
    new_new_n6535__, new_new_n6536__, new_new_n6537__, new_new_n6538__,
    new_new_n6539__, new_new_n6540__, new_new_n6541__, new_new_n6542__,
    new_new_n6543__, new_new_n6544__, new_new_n6545__, new_new_n6546__,
    new_new_n6547__, new_new_n6548__, new_new_n6549__, new_new_n6550__,
    new_new_n6551__, new_new_n6552__, new_new_n6553__, new_new_n6554__,
    new_new_n6555__, new_new_n6556__, new_new_n6557__, new_new_n6558__,
    new_new_n6559__, new_new_n6560__, new_new_n6561__, new_new_n6562__,
    new_new_n6563__, new_new_n6564__, new_new_n6565__, new_new_n6566__,
    new_new_n6567__, new_new_n6568__, new_new_n6569__, new_new_n6570__,
    new_new_n6571__, new_new_n6572__, new_new_n6573__, new_new_n6574__,
    new_new_n6575__, new_new_n6576__, new_new_n6577__, new_new_n6578__,
    new_new_n6579__, new_new_n6580__, new_new_n6581__, new_new_n6582__,
    new_new_n6583__, new_new_n6584__, new_new_n6585__, new_new_n6586__,
    new_new_n6587__, new_new_n6588__, new_new_n6589__, new_new_n6590__,
    new_new_n6591__, new_new_n6592__, new_new_n6593__, new_new_n6594__,
    new_new_n6595__, new_new_n6596__, new_new_n6597__, new_new_n6598__,
    new_new_n6599__, new_new_n6600__, new_new_n6601__, new_new_n6602__,
    new_new_n6603__, new_new_n6605__, new_new_n6606__, new_new_n6607__,
    new_new_n6608__, new_new_n6609__, new_new_n6610__, new_new_n6611__,
    new_new_n6612__, new_new_n6613__, new_new_n6614__, new_new_n6615__,
    new_new_n6616__, new_new_n6617__, new_new_n6618__, new_new_n6619__,
    new_new_n6620__, new_new_n6621__, new_new_n6622__, new_new_n6623__,
    new_new_n6624__, new_new_n6625__, new_new_n6626__, new_new_n6627__,
    new_new_n6628__, new_new_n6629__, new_new_n6630__, new_new_n6631__,
    new_new_n6632__, new_new_n6633__, new_new_n6634__, new_new_n6635__,
    new_new_n6636__, new_new_n6637__, new_new_n6638__, new_new_n6639__,
    new_new_n6640__, new_new_n6641__, new_new_n6642__, new_new_n6643__,
    new_new_n6644__, new_new_n6645__, new_new_n6646__, new_new_n6647__,
    new_new_n6648__, new_new_n6649__, new_new_n6650__, new_new_n6651__,
    new_new_n6652__, new_new_n6653__, new_new_n6654__, new_new_n6655__,
    new_new_n6656__, new_new_n6657__, new_new_n6658__, new_new_n6659__,
    new_new_n6660__, new_new_n6661__, new_new_n6662__, new_new_n6663__,
    new_new_n6664__, new_new_n6665__, new_new_n6666__, new_new_n6667__,
    new_new_n6668__, new_new_n6669__, new_new_n6670__, new_new_n6671__,
    new_new_n6672__, new_new_n6673__, new_new_n6674__, new_new_n6675__,
    new_new_n6676__, new_new_n6677__, new_new_n6678__, new_new_n6679__,
    new_new_n6680__, new_new_n6681__, new_new_n6682__, new_new_n6683__,
    new_new_n6684__, new_new_n6685__, new_new_n6686__, new_new_n6687__,
    new_new_n6688__, new_new_n6689__, new_new_n6690__, new_new_n6691__,
    new_new_n6692__, new_new_n6693__, new_new_n6694__, new_new_n6695__,
    new_new_n6696__, new_new_n6697__, new_new_n6698__, new_new_n6699__,
    new_new_n6700__, new_new_n6701__, new_new_n6702__, new_new_n6703__,
    new_new_n6704__, new_new_n6705__, new_new_n6706__, new_new_n6707__,
    new_new_n6708__, new_new_n6709__, new_new_n6710__, new_new_n6711__,
    new_new_n6712__, new_new_n6713__, new_new_n6714__, new_new_n6715__,
    new_new_n6716__, new_new_n6717__, new_new_n6718__, new_new_n6719__,
    new_new_n6720__, new_new_n6721__, new_new_n6722__, new_new_n6723__,
    new_new_n6724__, new_new_n6725__, new_new_n6726__, new_new_n6727__,
    new_new_n6728__, new_new_n6729__, new_new_n6730__, new_new_n6731__,
    new_new_n6732__, new_new_n6733__, new_new_n6734__, new_new_n6735__,
    new_new_n6736__, new_new_n6737__, new_new_n6738__, new_new_n6739__,
    new_new_n6740__, new_new_n6741__, new_new_n6742__, new_new_n6743__,
    new_new_n6744__, new_new_n6745__, new_new_n6746__, new_new_n6747__,
    new_new_n6748__, new_new_n6749__, new_new_n6750__, new_new_n6751__,
    new_new_n6752__, new_new_n6753__, new_new_n6754__, new_new_n6755__,
    new_new_n6756__, new_new_n6757__, new_new_n6758__, new_new_n6759__,
    new_new_n6760__, new_new_n6761__, new_new_n6762__, new_new_n6763__,
    new_new_n6764__, new_new_n6765__, new_new_n6766__, new_new_n6767__,
    new_new_n6768__, new_new_n6769__, new_new_n6770__, new_new_n6771__,
    new_new_n6772__, new_new_n6773__, new_new_n6774__, new_new_n6775__,
    new_new_n6776__, new_new_n6777__, new_new_n6778__, new_new_n6779__,
    new_new_n6780__, new_new_n6781__, new_new_n6782__, new_new_n6783__,
    new_new_n6784__, new_new_n6785__, new_new_n6786__, new_new_n6787__,
    new_new_n6788__, new_new_n6789__, new_new_n6790__, new_new_n6791__,
    new_new_n6792__, new_new_n6793__, new_new_n6794__, new_new_n6795__,
    new_new_n6796__, new_new_n6797__, new_new_n6798__, new_new_n6799__,
    new_new_n6800__, new_new_n6801__, new_new_n6802__, new_new_n6803__,
    new_new_n6804__, new_new_n6805__, new_new_n6806__, new_new_n6807__,
    new_new_n6808__, new_new_n6809__, new_new_n6810__, new_new_n6811__,
    new_new_n6812__, new_new_n6813__, new_new_n6814__, new_new_n6815__,
    new_new_n6816__, new_new_n6817__, new_new_n6818__, new_new_n6819__,
    new_new_n6820__, new_new_n6821__, new_new_n6822__, new_new_n6823__,
    new_new_n6824__, new_new_n6825__, new_new_n6826__, new_new_n6827__,
    new_new_n6828__, new_new_n6829__, new_new_n6830__, new_new_n6831__,
    new_new_n6832__, new_new_n6833__, new_new_n6834__, new_new_n6835__,
    new_new_n6836__, new_new_n6837__, new_new_n6838__, new_new_n6839__,
    new_new_n6840__, new_new_n6841__, new_new_n6842__, new_new_n6843__,
    new_new_n6844__, new_new_n6845__, new_new_n6846__, new_new_n6847__,
    new_new_n6848__, new_new_n6849__, new_new_n6850__, new_new_n6851__,
    new_new_n6853__, new_new_n6854__, new_new_n6855__, new_new_n6856__,
    new_new_n6857__, new_new_n6858__, new_new_n6859__, new_new_n6860__,
    new_new_n6861__, new_new_n6862__, new_new_n6863__, new_new_n6864__,
    new_new_n6865__, new_new_n6866__, new_new_n6867__, new_new_n6868__,
    new_new_n6869__, new_new_n6870__, new_new_n6871__, new_new_n6872__,
    new_new_n6873__, new_new_n6874__, new_new_n6875__, new_new_n6876__,
    new_new_n6877__, new_new_n6878__, new_new_n6879__, new_new_n6880__,
    new_new_n6881__, new_new_n6882__, new_new_n6883__, new_new_n6884__,
    new_new_n6885__, new_new_n6886__, new_new_n6887__, new_new_n6888__,
    new_new_n6889__, new_new_n6890__, new_new_n6891__, new_new_n6892__,
    new_new_n6893__, new_new_n6894__, new_new_n6895__, new_new_n6896__,
    new_new_n6897__, new_new_n6898__, new_new_n6899__, new_new_n6900__,
    new_new_n6901__, new_new_n6902__, new_new_n6903__, new_new_n6904__,
    new_new_n6905__, new_new_n6906__, new_new_n6907__, new_new_n6908__,
    new_new_n6909__, new_new_n6910__, new_new_n6911__, new_new_n6912__,
    new_new_n6913__, new_new_n6914__, new_new_n6915__, new_new_n6916__,
    new_new_n6917__, new_new_n6918__, new_new_n6919__, new_new_n6920__,
    new_new_n6921__, new_new_n6922__, new_new_n6923__, new_new_n6924__,
    new_new_n6925__, new_new_n6926__, new_new_n6927__, new_new_n6928__,
    new_new_n6929__, new_new_n6930__, new_new_n6931__, new_new_n6932__,
    new_new_n6933__, new_new_n6934__, new_new_n6935__, new_new_n6936__,
    new_new_n6937__, new_new_n6938__, new_new_n6939__, new_new_n6940__,
    new_new_n6941__, new_new_n6942__, new_new_n6943__, new_new_n6944__,
    new_new_n6945__, new_new_n6946__, new_new_n6947__, new_new_n6948__,
    new_new_n6949__, new_new_n6950__, new_new_n6951__, new_new_n6952__,
    new_new_n6953__, new_new_n6954__, new_new_n6955__, new_new_n6956__,
    new_new_n6957__, new_new_n6958__, new_new_n6959__, new_new_n6960__,
    new_new_n6961__, new_new_n6962__, new_new_n6963__, new_new_n6964__,
    new_new_n6965__, new_new_n6966__, new_new_n6967__, new_new_n6968__,
    new_new_n6969__, new_new_n6970__, new_new_n6971__, new_new_n6972__,
    new_new_n6973__, new_new_n6974__, new_new_n6975__, new_new_n6976__,
    new_new_n6977__, new_new_n6978__, new_new_n6979__, new_new_n6980__,
    new_new_n6981__, new_new_n6982__, new_new_n6983__, new_new_n6984__,
    new_new_n6985__, new_new_n6986__, new_new_n6987__, new_new_n6988__,
    new_new_n6989__, new_new_n6990__, new_new_n6991__, new_new_n6992__,
    new_new_n6993__, new_new_n6994__, new_new_n6995__, new_new_n6996__,
    new_new_n6997__, new_new_n6998__, new_new_n6999__, new_new_n7000__,
    new_new_n7001__, new_new_n7002__, new_new_n7003__, new_new_n7004__,
    new_new_n7005__, new_new_n7006__, new_new_n7007__, new_new_n7008__,
    new_new_n7009__, new_new_n7010__, new_new_n7011__, new_new_n7012__,
    new_new_n7013__, new_new_n7014__, new_new_n7015__, new_new_n7016__,
    new_new_n7017__, new_new_n7018__, new_new_n7019__, new_new_n7020__,
    new_new_n7021__, new_new_n7022__, new_new_n7023__, new_new_n7024__,
    new_new_n7025__, new_new_n7026__, new_new_n7027__, new_new_n7028__,
    new_new_n7029__, new_new_n7030__, new_new_n7031__, new_new_n7032__,
    new_new_n7033__, new_new_n7034__, new_new_n7035__, new_new_n7036__,
    new_new_n7037__, new_new_n7038__, new_new_n7039__, new_new_n7040__,
    new_new_n7041__, new_new_n7042__, new_new_n7043__, new_new_n7044__,
    new_new_n7045__, new_new_n7046__, new_new_n7047__, new_new_n7048__,
    new_new_n7049__, new_new_n7050__, new_new_n7051__, new_new_n7052__,
    new_new_n7053__, new_new_n7054__, new_new_n7055__, new_new_n7056__,
    new_new_n7057__, new_new_n7058__, new_new_n7059__, new_new_n7060__,
    new_new_n7061__, new_new_n7062__, new_new_n7063__, new_new_n7064__,
    new_new_n7065__, new_new_n7066__, new_new_n7067__, new_new_n7068__,
    new_new_n7069__, new_new_n7070__, new_new_n7071__, new_new_n7072__,
    new_new_n7073__, new_new_n7074__, new_new_n7075__, new_new_n7076__,
    new_new_n7077__, new_new_n7078__, new_new_n7079__, new_new_n7081__,
    new_new_n7082__, new_new_n7083__, new_new_n7084__, new_new_n7085__,
    new_new_n7086__, new_new_n7087__, new_new_n7088__, new_new_n7089__,
    new_new_n7090__, new_new_n7091__, new_new_n7092__, new_new_n7093__,
    new_new_n7094__, new_new_n7095__, new_new_n7096__, new_new_n7097__,
    new_new_n7098__, new_new_n7099__, new_new_n7100__, new_new_n7101__,
    new_new_n7102__, new_new_n7103__, new_new_n7104__, new_new_n7105__,
    new_new_n7106__, new_new_n7107__, new_new_n7108__, new_new_n7109__,
    new_new_n7110__, new_new_n7111__, new_new_n7112__, new_new_n7113__,
    new_new_n7114__, new_new_n7115__, new_new_n7116__, new_new_n7117__,
    new_new_n7118__, new_new_n7119__, new_new_n7120__, new_new_n7121__,
    new_new_n7122__, new_new_n7123__, new_new_n7124__, new_new_n7125__,
    new_new_n7126__, new_new_n7127__, new_new_n7128__, new_new_n7129__,
    new_new_n7130__, new_new_n7131__, new_new_n7132__, new_new_n7133__,
    new_new_n7134__, new_new_n7135__, new_new_n7136__, new_new_n7137__,
    new_new_n7138__, new_new_n7139__, new_new_n7140__, new_new_n7141__,
    new_new_n7142__, new_new_n7143__, new_new_n7144__, new_new_n7145__,
    new_new_n7146__, new_new_n7147__, new_new_n7148__, new_new_n7149__,
    new_new_n7150__, new_new_n7151__, new_new_n7152__, new_new_n7153__,
    new_new_n7154__, new_new_n7155__, new_new_n7156__, new_new_n7157__,
    new_new_n7158__, new_new_n7159__, new_new_n7160__, new_new_n7161__,
    new_new_n7162__, new_new_n7163__, new_new_n7164__, new_new_n7165__,
    new_new_n7166__, new_new_n7167__, new_new_n7168__, new_new_n7169__,
    new_new_n7170__, new_new_n7171__, new_new_n7172__, new_new_n7173__,
    new_new_n7174__, new_new_n7175__, new_new_n7176__, new_new_n7177__,
    new_new_n7178__, new_new_n7179__, new_new_n7180__, new_new_n7181__,
    new_new_n7182__, new_new_n7183__, new_new_n7184__, new_new_n7185__,
    new_new_n7186__, new_new_n7187__, new_new_n7188__, new_new_n7189__,
    new_new_n7190__, new_new_n7191__, new_new_n7192__, new_new_n7193__,
    new_new_n7194__, new_new_n7195__, new_new_n7196__, new_new_n7197__,
    new_new_n7198__, new_new_n7199__, new_new_n7200__, new_new_n7201__,
    new_new_n7202__, new_new_n7203__, new_new_n7204__, new_new_n7205__,
    new_new_n7206__, new_new_n7207__, new_new_n7208__, new_new_n7209__,
    new_new_n7210__, new_new_n7211__, new_new_n7212__, new_new_n7213__,
    new_new_n7214__, new_new_n7215__, new_new_n7216__, new_new_n7217__,
    new_new_n7218__, new_new_n7219__, new_new_n7220__, new_new_n7221__,
    new_new_n7222__, new_new_n7223__, new_new_n7224__, new_new_n7225__,
    new_new_n7226__, new_new_n7227__, new_new_n7228__, new_new_n7229__,
    new_new_n7230__, new_new_n7231__, new_new_n7232__, new_new_n7233__,
    new_new_n7234__, new_new_n7235__, new_new_n7236__, new_new_n7237__,
    new_new_n7238__, new_new_n7239__, new_new_n7240__, new_new_n7241__,
    new_new_n7242__, new_new_n7243__, new_new_n7244__, new_new_n7245__,
    new_new_n7246__, new_new_n7247__, new_new_n7248__, new_new_n7249__,
    new_new_n7250__, new_new_n7251__, new_new_n7252__, new_new_n7253__,
    new_new_n7254__, new_new_n7255__, new_new_n7256__, new_new_n7257__,
    new_new_n7258__, new_new_n7259__, new_new_n7260__, new_new_n7261__,
    new_new_n7262__, new_new_n7263__, new_new_n7264__, new_new_n7265__,
    new_new_n7266__, new_new_n7267__, new_new_n7268__, new_new_n7269__,
    new_new_n7270__, new_new_n7271__, new_new_n7272__, new_new_n7273__,
    new_new_n7274__, new_new_n7275__, new_new_n7276__, new_new_n7277__,
    new_new_n7278__, new_new_n7279__, new_new_n7280__, new_new_n7281__,
    new_new_n7282__, new_new_n7283__, new_new_n7284__, new_new_n7285__,
    new_new_n7286__, new_new_n7287__, new_new_n7288__, new_new_n7289__,
    new_new_n7290__, new_new_n7291__, new_new_n7292__, new_new_n7293__,
    new_new_n7294__, new_new_n7295__, new_new_n7296__, new_new_n7297__,
    new_new_n7298__, new_new_n7299__, new_new_n7300__, new_new_n7301__,
    new_new_n7302__, new_new_n7303__, new_new_n7304__, new_new_n7305__,
    new_new_n7306__, new_new_n7307__, new_new_n7308__, new_new_n7309__,
    new_new_n7310__, new_new_n7311__, new_new_n7312__, new_new_n7313__,
    new_new_n7314__, new_new_n7315__, new_new_n7316__, new_new_n7317__,
    new_new_n7318__, new_new_n7319__, new_new_n7320__, new_new_n7321__,
    new_new_n7322__, new_new_n7323__, new_new_n7324__, new_new_n7325__,
    new_new_n7326__, new_new_n7327__, new_new_n7328__, new_new_n7329__,
    new_new_n7330__, new_new_n7331__, new_new_n7332__, new_new_n7333__,
    new_new_n7334__, new_new_n7335__, new_new_n7336__, new_new_n7337__,
    new_new_n7338__, new_new_n7339__, new_new_n7340__, new_new_n7341__,
    new_new_n7342__, new_new_n7343__, new_new_n7344__, new_new_n7345__,
    new_new_n7346__, new_new_n7347__, new_new_n7348__, new_new_n7349__,
    new_new_n7350__, new_new_n7351__, new_new_n7352__, new_new_n7353__,
    new_new_n7354__, new_new_n7355__, new_new_n7356__, new_new_n7357__,
    new_new_n7358__, new_new_n7359__, new_new_n7360__, new_new_n7361__,
    new_new_n7362__, new_new_n7363__, new_new_n7364__, new_new_n7366__,
    new_new_n7367__, new_new_n7368__, new_new_n7369__, new_new_n7370__,
    new_new_n7371__, new_new_n7372__, new_new_n7373__, new_new_n7374__,
    new_new_n7375__, new_new_n7376__, new_new_n7377__, new_new_n7378__,
    new_new_n7379__, new_new_n7380__, new_new_n7381__, new_new_n7382__,
    new_new_n7383__, new_new_n7384__, new_new_n7385__, new_new_n7386__,
    new_new_n7387__, new_new_n7388__, new_new_n7389__, new_new_n7390__,
    new_new_n7391__, new_new_n7392__, new_new_n7393__, new_new_n7394__,
    new_new_n7395__, new_new_n7396__, new_new_n7397__, new_new_n7398__,
    new_new_n7399__, new_new_n7400__, new_new_n7401__, new_new_n7402__,
    new_new_n7403__, new_new_n7404__, new_new_n7405__, new_new_n7406__,
    new_new_n7407__, new_new_n7408__, new_new_n7409__, new_new_n7410__,
    new_new_n7411__, new_new_n7412__, new_new_n7413__, new_new_n7414__,
    new_new_n7415__, new_new_n7416__, new_new_n7417__, new_new_n7418__,
    new_new_n7419__, new_new_n7420__, new_new_n7421__, new_new_n7422__,
    new_new_n7423__, new_new_n7424__, new_new_n7425__, new_new_n7426__,
    new_new_n7427__, new_new_n7428__, new_new_n7429__, new_new_n7430__,
    new_new_n7431__, new_new_n7432__, new_new_n7433__, new_new_n7434__,
    new_new_n7435__, new_new_n7436__, new_new_n7437__, new_new_n7438__,
    new_new_n7439__, new_new_n7440__, new_new_n7441__, new_new_n7442__,
    new_new_n7443__, new_new_n7444__, new_new_n7445__, new_new_n7446__,
    new_new_n7447__, new_new_n7448__, new_new_n7449__, new_new_n7450__,
    new_new_n7451__, new_new_n7452__, new_new_n7453__, new_new_n7454__,
    new_new_n7455__, new_new_n7456__, new_new_n7457__, new_new_n7458__,
    new_new_n7459__, new_new_n7460__, new_new_n7461__, new_new_n7462__,
    new_new_n7463__, new_new_n7464__, new_new_n7465__, new_new_n7466__,
    new_new_n7467__, new_new_n7468__, new_new_n7469__, new_new_n7470__,
    new_new_n7471__, new_new_n7472__, new_new_n7473__, new_new_n7474__,
    new_new_n7475__, new_new_n7476__, new_new_n7477__, new_new_n7478__,
    new_new_n7479__, new_new_n7480__, new_new_n7481__, new_new_n7482__,
    new_new_n7483__, new_new_n7484__, new_new_n7485__, new_new_n7486__,
    new_new_n7487__, new_new_n7488__, new_new_n7489__, new_new_n7490__,
    new_new_n7491__, new_new_n7492__, new_new_n7493__, new_new_n7494__,
    new_new_n7495__, new_new_n7496__, new_new_n7497__, new_new_n7498__,
    new_new_n7499__, new_new_n7500__, new_new_n7501__, new_new_n7502__,
    new_new_n7503__, new_new_n7504__, new_new_n7505__, new_new_n7506__,
    new_new_n7507__, new_new_n7508__, new_new_n7509__, new_new_n7510__,
    new_new_n7511__, new_new_n7512__, new_new_n7513__, new_new_n7514__,
    new_new_n7515__, new_new_n7516__, new_new_n7517__, new_new_n7518__,
    new_new_n7519__, new_new_n7520__, new_new_n7521__, new_new_n7522__,
    new_new_n7523__, new_new_n7524__, new_new_n7525__, new_new_n7526__,
    new_new_n7527__, new_new_n7528__, new_new_n7529__, new_new_n7530__,
    new_new_n7531__, new_new_n7532__, new_new_n7533__, new_new_n7534__,
    new_new_n7535__, new_new_n7536__, new_new_n7537__, new_new_n7538__,
    new_new_n7539__, new_new_n7540__, new_new_n7541__, new_new_n7542__,
    new_new_n7543__, new_new_n7544__, new_new_n7545__, new_new_n7546__,
    new_new_n7547__, new_new_n7548__, new_new_n7549__, new_new_n7550__,
    new_new_n7551__, new_new_n7552__, new_new_n7553__, new_new_n7554__,
    new_new_n7555__, new_new_n7556__, new_new_n7557__, new_new_n7558__,
    new_new_n7559__, new_new_n7560__, new_new_n7561__, new_new_n7562__,
    new_new_n7563__, new_new_n7564__, new_new_n7565__, new_new_n7566__,
    new_new_n7567__, new_new_n7568__, new_new_n7569__, new_new_n7570__,
    new_new_n7571__, new_new_n7572__, new_new_n7573__, new_new_n7574__,
    new_new_n7575__, new_new_n7576__, new_new_n7577__, new_new_n7578__,
    new_new_n7579__, new_new_n7580__, new_new_n7581__, new_new_n7582__,
    new_new_n7583__, new_new_n7584__, new_new_n7585__, new_new_n7586__,
    new_new_n7587__, new_new_n7588__, new_new_n7589__, new_new_n7590__,
    new_new_n7591__, new_new_n7592__, new_new_n7593__, new_new_n7594__,
    new_new_n7595__, new_new_n7596__, new_new_n7597__, new_new_n7598__,
    new_new_n7599__, new_new_n7600__, new_new_n7601__, new_new_n7602__,
    new_new_n7603__, new_new_n7604__, new_new_n7605__, new_new_n7606__,
    new_new_n7607__, new_new_n7608__, new_new_n7609__, new_new_n7610__,
    new_new_n7611__, new_new_n7612__, new_new_n7613__, new_new_n7614__,
    new_new_n7615__, new_new_n7616__, new_new_n7617__, new_new_n7618__,
    new_new_n7619__, new_new_n7620__, new_new_n7621__, new_new_n7622__,
    new_new_n7623__, new_new_n7624__, new_new_n7626__, new_new_n7627__,
    new_new_n7628__, new_new_n7629__, new_new_n7630__, new_new_n7631__,
    new_new_n7632__, new_new_n7633__, new_new_n7634__, new_new_n7635__,
    new_new_n7636__, new_new_n7637__, new_new_n7638__, new_new_n7639__,
    new_new_n7640__, new_new_n7641__, new_new_n7642__, new_new_n7643__,
    new_new_n7644__, new_new_n7645__, new_new_n7646__, new_new_n7647__,
    new_new_n7648__, new_new_n7649__, new_new_n7650__, new_new_n7651__,
    new_new_n7652__, new_new_n7653__, new_new_n7654__, new_new_n7655__,
    new_new_n7656__, new_new_n7657__, new_new_n7658__, new_new_n7659__,
    new_new_n7660__, new_new_n7661__, new_new_n7662__, new_new_n7663__,
    new_new_n7664__, new_new_n7665__, new_new_n7666__, new_new_n7667__,
    new_new_n7668__, new_new_n7669__, new_new_n7670__, new_new_n7671__,
    new_new_n7672__, new_new_n7673__, new_new_n7674__, new_new_n7675__,
    new_new_n7676__, new_new_n7677__, new_new_n7678__, new_new_n7679__,
    new_new_n7680__, new_new_n7681__, new_new_n7682__, new_new_n7683__,
    new_new_n7684__, new_new_n7685__, new_new_n7686__, new_new_n7687__,
    new_new_n7688__, new_new_n7689__, new_new_n7690__, new_new_n7691__,
    new_new_n7692__, new_new_n7693__, new_new_n7694__, new_new_n7695__,
    new_new_n7696__, new_new_n7697__, new_new_n7698__, new_new_n7699__,
    new_new_n7700__, new_new_n7701__, new_new_n7702__, new_new_n7703__,
    new_new_n7704__, new_new_n7705__, new_new_n7706__, new_new_n7707__,
    new_new_n7708__, new_new_n7709__, new_new_n7710__, new_new_n7711__,
    new_new_n7712__, new_new_n7713__, new_new_n7714__, new_new_n7715__,
    new_new_n7716__, new_new_n7717__, new_new_n7718__, new_new_n7719__,
    new_new_n7720__, new_new_n7721__, new_new_n7722__, new_new_n7723__,
    new_new_n7724__, new_new_n7725__, new_new_n7726__, new_new_n7727__,
    new_new_n7728__, new_new_n7729__, new_new_n7730__, new_new_n7731__,
    new_new_n7732__, new_new_n7733__, new_new_n7734__, new_new_n7735__,
    new_new_n7736__, new_new_n7737__, new_new_n7738__, new_new_n7739__,
    new_new_n7740__, new_new_n7741__, new_new_n7742__, new_new_n7743__,
    new_new_n7744__, new_new_n7745__, new_new_n7746__, new_new_n7747__,
    new_new_n7748__, new_new_n7749__, new_new_n7750__, new_new_n7751__,
    new_new_n7752__, new_new_n7753__, new_new_n7754__, new_new_n7755__,
    new_new_n7756__, new_new_n7757__, new_new_n7758__, new_new_n7759__,
    new_new_n7760__, new_new_n7761__, new_new_n7762__, new_new_n7763__,
    new_new_n7764__, new_new_n7765__, new_new_n7766__, new_new_n7767__,
    new_new_n7768__, new_new_n7769__, new_new_n7770__, new_new_n7771__,
    new_new_n7772__, new_new_n7773__, new_new_n7774__, new_new_n7775__,
    new_new_n7776__, new_new_n7777__, new_new_n7778__, new_new_n7779__,
    new_new_n7780__, new_new_n7781__, new_new_n7782__, new_new_n7783__,
    new_new_n7784__, new_new_n7785__, new_new_n7786__, new_new_n7787__,
    new_new_n7788__, new_new_n7789__, new_new_n7790__, new_new_n7791__,
    new_new_n7792__, new_new_n7793__, new_new_n7794__, new_new_n7795__,
    new_new_n7796__, new_new_n7797__, new_new_n7798__, new_new_n7799__,
    new_new_n7800__, new_new_n7801__, new_new_n7802__, new_new_n7803__,
    new_new_n7804__, new_new_n7805__, new_new_n7806__, new_new_n7807__,
    new_new_n7808__, new_new_n7809__, new_new_n7810__, new_new_n7811__,
    new_new_n7812__, new_new_n7813__, new_new_n7814__, new_new_n7815__,
    new_new_n7816__, new_new_n7817__, new_new_n7818__, new_new_n7819__,
    new_new_n7820__, new_new_n7821__, new_new_n7822__, new_new_n7823__,
    new_new_n7824__, new_new_n7825__, new_new_n7826__, new_new_n7827__,
    new_new_n7828__, new_new_n7829__, new_new_n7830__, new_new_n7831__,
    new_new_n7832__, new_new_n7833__, new_new_n7834__, new_new_n7835__,
    new_new_n7836__, new_new_n7837__, new_new_n7838__, new_new_n7839__,
    new_new_n7840__, new_new_n7841__, new_new_n7842__, new_new_n7843__,
    new_new_n7844__, new_new_n7845__, new_new_n7846__, new_new_n7847__,
    new_new_n7848__, new_new_n7849__, new_new_n7850__, new_new_n7851__,
    new_new_n7852__, new_new_n7853__, new_new_n7854__, new_new_n7855__,
    new_new_n7856__, new_new_n7857__, new_new_n7858__, new_new_n7859__,
    new_new_n7860__, new_new_n7861__, new_new_n7862__, new_new_n7863__,
    new_new_n7864__, new_new_n7865__, new_new_n7866__, new_new_n7867__,
    new_new_n7868__, new_new_n7869__, new_new_n7870__, new_new_n7871__,
    new_new_n7872__, new_new_n7873__, new_new_n7874__, new_new_n7875__,
    new_new_n7876__, new_new_n7877__, new_new_n7878__, new_new_n7879__,
    new_new_n7880__, new_new_n7881__, new_new_n7882__, new_new_n7884__,
    new_new_n7885__, new_new_n7886__, new_new_n7887__, new_new_n7888__,
    new_new_n7889__, new_new_n7890__, new_new_n7891__, new_new_n7892__,
    new_new_n7893__, new_new_n7894__, new_new_n7895__, new_new_n7896__,
    new_new_n7897__, new_new_n7898__, new_new_n7899__, new_new_n7900__,
    new_new_n7901__, new_new_n7902__, new_new_n7903__, new_new_n7904__,
    new_new_n7905__, new_new_n7906__, new_new_n7907__, new_new_n7908__,
    new_new_n7909__, new_new_n7910__, new_new_n7911__, new_new_n7912__,
    new_new_n7913__, new_new_n7914__, new_new_n7915__, new_new_n7916__,
    new_new_n7917__, new_new_n7918__, new_new_n7919__, new_new_n7920__,
    new_new_n7921__, new_new_n7922__, new_new_n7923__, new_new_n7924__,
    new_new_n7925__, new_new_n7926__, new_new_n7927__, new_new_n7928__,
    new_new_n7929__, new_new_n7930__, new_new_n7931__, new_new_n7932__,
    new_new_n7933__, new_new_n7934__, new_new_n7935__, new_new_n7936__,
    new_new_n7937__, new_new_n7938__, new_new_n7939__, new_new_n7940__,
    new_new_n7941__, new_new_n7942__, new_new_n7943__, new_new_n7944__,
    new_new_n7945__, new_new_n7946__, new_new_n7947__, new_new_n7948__,
    new_new_n7949__, new_new_n7950__, new_new_n7951__, new_new_n7952__,
    new_new_n7953__, new_new_n7954__, new_new_n7955__, new_new_n7956__,
    new_new_n7957__, new_new_n7958__, new_new_n7959__, new_new_n7960__,
    new_new_n7961__, new_new_n7962__, new_new_n7963__, new_new_n7964__,
    new_new_n7965__, new_new_n7966__, new_new_n7967__, new_new_n7968__,
    new_new_n7969__, new_new_n7970__, new_new_n7971__, new_new_n7972__,
    new_new_n7973__, new_new_n7974__, new_new_n7975__, new_new_n7976__,
    new_new_n7977__, new_new_n7978__, new_new_n7979__, new_new_n7980__,
    new_new_n7981__, new_new_n7982__, new_new_n7983__, new_new_n7984__,
    new_new_n7985__, new_new_n7986__, new_new_n7987__, new_new_n7988__,
    new_new_n7989__, new_new_n7990__, new_new_n7991__, new_new_n7992__,
    new_new_n7993__, new_new_n7994__, new_new_n7995__, new_new_n7996__,
    new_new_n7997__, new_new_n7998__, new_new_n7999__, new_new_n8000__,
    new_new_n8001__, new_new_n8002__, new_new_n8003__, new_new_n8004__,
    new_new_n8005__, new_new_n8006__, new_new_n8007__, new_new_n8008__,
    new_new_n8009__, new_new_n8010__, new_new_n8011__, new_new_n8012__,
    new_new_n8013__, new_new_n8014__, new_new_n8015__, new_new_n8016__,
    new_new_n8017__, new_new_n8018__, new_new_n8019__, new_new_n8020__,
    new_new_n8021__, new_new_n8022__, new_new_n8023__, new_new_n8024__,
    new_new_n8025__, new_new_n8026__, new_new_n8027__, new_new_n8028__,
    new_new_n8029__, new_new_n8030__, new_new_n8031__, new_new_n8032__,
    new_new_n8033__, new_new_n8034__, new_new_n8035__, new_new_n8036__,
    new_new_n8037__, new_new_n8038__, new_new_n8039__, new_new_n8040__,
    new_new_n8041__, new_new_n8042__, new_new_n8043__, new_new_n8044__,
    new_new_n8045__, new_new_n8046__, new_new_n8047__, new_new_n8048__,
    new_new_n8049__, new_new_n8050__, new_new_n8051__, new_new_n8052__,
    new_new_n8053__, new_new_n8054__, new_new_n8055__, new_new_n8056__,
    new_new_n8057__, new_new_n8058__, new_new_n8059__, new_new_n8060__,
    new_new_n8061__, new_new_n8062__, new_new_n8063__, new_new_n8064__,
    new_new_n8065__, new_new_n8066__, new_new_n8067__, new_new_n8068__,
    new_new_n8069__, new_new_n8070__, new_new_n8071__, new_new_n8072__,
    new_new_n8073__, new_new_n8074__, new_new_n8075__, new_new_n8076__,
    new_new_n8077__, new_new_n8078__, new_new_n8079__, new_new_n8080__,
    new_new_n8081__, new_new_n8082__, new_new_n8083__, new_new_n8084__,
    new_new_n8085__, new_new_n8086__, new_new_n8087__, new_new_n8088__,
    new_new_n8089__, new_new_n8090__, new_new_n8091__, new_new_n8092__,
    new_new_n8093__, new_new_n8094__, new_new_n8095__, new_new_n8096__,
    new_new_n8097__, new_new_n8098__, new_new_n8099__, new_new_n8100__,
    new_new_n8101__, new_new_n8102__, new_new_n8103__, new_new_n8104__,
    new_new_n8105__, new_new_n8106__, new_new_n8107__, new_new_n8108__,
    new_new_n8109__, new_new_n8110__, new_new_n8111__, new_new_n8112__,
    new_new_n8113__, new_new_n8114__, new_new_n8115__, new_new_n8116__,
    new_new_n8117__, new_new_n8118__, new_new_n8119__, new_new_n8120__,
    new_new_n8121__, new_new_n8122__, new_new_n8123__, new_new_n8124__,
    new_new_n8125__, new_new_n8126__, new_new_n8127__, new_new_n8128__,
    new_new_n8129__, new_new_n8130__, new_new_n8131__, new_new_n8132__,
    new_new_n8133__, new_new_n8134__, new_new_n8136__, new_new_n8137__,
    new_new_n8138__, new_new_n8139__, new_new_n8140__, new_new_n8141__,
    new_new_n8142__, new_new_n8143__, new_new_n8144__, new_new_n8145__,
    new_new_n8146__, new_new_n8147__, new_new_n8148__, new_new_n8149__,
    new_new_n8150__, new_new_n8151__, new_new_n8152__, new_new_n8153__,
    new_new_n8154__, new_new_n8155__, new_new_n8156__, new_new_n8157__,
    new_new_n8158__, new_new_n8159__, new_new_n8160__, new_new_n8161__,
    new_new_n8162__, new_new_n8163__, new_new_n8164__, new_new_n8165__,
    new_new_n8166__, new_new_n8167__, new_new_n8168__, new_new_n8169__,
    new_new_n8170__, new_new_n8171__, new_new_n8172__, new_new_n8173__,
    new_new_n8174__, new_new_n8175__, new_new_n8176__, new_new_n8177__,
    new_new_n8178__, new_new_n8179__, new_new_n8180__, new_new_n8181__,
    new_new_n8182__, new_new_n8183__, new_new_n8184__, new_new_n8185__,
    new_new_n8186__, new_new_n8187__, new_new_n8188__, new_new_n8189__,
    new_new_n8190__, new_new_n8191__, new_new_n8192__, new_new_n8193__,
    new_new_n8194__, new_new_n8195__, new_new_n8196__, new_new_n8197__,
    new_new_n8198__, new_new_n8199__, new_new_n8200__, new_new_n8201__,
    new_new_n8202__, new_new_n8203__, new_new_n8204__, new_new_n8205__,
    new_new_n8206__, new_new_n8207__, new_new_n8208__, new_new_n8209__,
    new_new_n8210__, new_new_n8211__, new_new_n8212__, new_new_n8213__,
    new_new_n8214__, new_new_n8215__, new_new_n8216__, new_new_n8217__,
    new_new_n8218__, new_new_n8219__, new_new_n8220__, new_new_n8221__,
    new_new_n8222__, new_new_n8223__, new_new_n8224__, new_new_n8225__,
    new_new_n8226__, new_new_n8227__, new_new_n8228__, new_new_n8229__,
    new_new_n8230__, new_new_n8231__, new_new_n8232__, new_new_n8233__,
    new_new_n8234__, new_new_n8235__, new_new_n8236__, new_new_n8237__,
    new_new_n8238__, new_new_n8239__, new_new_n8240__, new_new_n8241__,
    new_new_n8242__, new_new_n8243__, new_new_n8244__, new_new_n8245__,
    new_new_n8246__, new_new_n8247__, new_new_n8248__, new_new_n8249__,
    new_new_n8250__, new_new_n8251__, new_new_n8252__, new_new_n8253__,
    new_new_n8254__, new_new_n8255__, new_new_n8256__, new_new_n8257__,
    new_new_n8258__, new_new_n8259__, new_new_n8260__, new_new_n8261__,
    new_new_n8262__, new_new_n8263__, new_new_n8264__, new_new_n8265__,
    new_new_n8266__, new_new_n8267__, new_new_n8268__, new_new_n8269__,
    new_new_n8270__, new_new_n8271__, new_new_n8272__, new_new_n8273__,
    new_new_n8274__, new_new_n8275__, new_new_n8276__, new_new_n8277__,
    new_new_n8278__, new_new_n8279__, new_new_n8280__, new_new_n8281__,
    new_new_n8282__, new_new_n8283__, new_new_n8284__, new_new_n8285__,
    new_new_n8286__, new_new_n8287__, new_new_n8288__, new_new_n8289__,
    new_new_n8290__, new_new_n8291__, new_new_n8292__, new_new_n8293__,
    new_new_n8294__, new_new_n8295__, new_new_n8296__, new_new_n8297__,
    new_new_n8298__, new_new_n8299__, new_new_n8300__, new_new_n8301__,
    new_new_n8302__, new_new_n8303__, new_new_n8304__, new_new_n8305__,
    new_new_n8306__, new_new_n8307__, new_new_n8308__, new_new_n8309__,
    new_new_n8310__, new_new_n8311__, new_new_n8312__, new_new_n8313__,
    new_new_n8314__, new_new_n8315__, new_new_n8316__, new_new_n8317__,
    new_new_n8318__, new_new_n8319__, new_new_n8320__, new_new_n8321__,
    new_new_n8322__, new_new_n8323__, new_new_n8324__, new_new_n8325__,
    new_new_n8326__, new_new_n8327__, new_new_n8328__, new_new_n8329__,
    new_new_n8330__, new_new_n8331__, new_new_n8332__, new_new_n8333__,
    new_new_n8334__, new_new_n8335__, new_new_n8336__, new_new_n8337__,
    new_new_n8338__, new_new_n8339__, new_new_n8340__, new_new_n8341__,
    new_new_n8342__, new_new_n8343__, new_new_n8344__, new_new_n8345__,
    new_new_n8346__, new_new_n8347__, new_new_n8348__, new_new_n8349__,
    new_new_n8350__, new_new_n8351__, new_new_n8352__, new_new_n8353__,
    new_new_n8354__, new_new_n8355__, new_new_n8356__, new_new_n8357__,
    new_new_n8358__, new_new_n8359__, new_new_n8360__, new_new_n8361__,
    new_new_n8362__, new_new_n8363__, new_new_n8364__, new_new_n8365__,
    new_new_n8366__, new_new_n8367__, new_new_n8368__, new_new_n8369__,
    new_new_n8370__, new_new_n8371__, new_new_n8372__, new_new_n8373__,
    new_new_n8374__, new_new_n8375__, new_new_n8376__, new_new_n8377__,
    new_new_n8378__, new_new_n8379__, new_new_n8380__, new_new_n8381__,
    new_new_n8382__, new_new_n8383__, new_new_n8384__, new_new_n8385__,
    new_new_n8386__, new_new_n8387__, new_new_n8388__, new_new_n8389__,
    new_new_n8390__, new_new_n8391__, new_new_n8392__, new_new_n8393__,
    new_new_n8394__, new_new_n8395__, new_new_n8397__, new_new_n8398__,
    new_new_n8399__, new_new_n8400__, new_new_n8401__, new_new_n8402__,
    new_new_n8403__, new_new_n8404__, new_new_n8405__, new_new_n8406__,
    new_new_n8407__, new_new_n8408__, new_new_n8409__, new_new_n8410__,
    new_new_n8411__, new_new_n8412__, new_new_n8413__, new_new_n8414__,
    new_new_n8415__, new_new_n8416__, new_new_n8417__, new_new_n8418__,
    new_new_n8419__, new_new_n8420__, new_new_n8421__, new_new_n8422__,
    new_new_n8423__, new_new_n8424__, new_new_n8425__, new_new_n8426__,
    new_new_n8427__, new_new_n8428__, new_new_n8429__, new_new_n8430__,
    new_new_n8431__, new_new_n8432__, new_new_n8433__, new_new_n8434__,
    new_new_n8435__, new_new_n8436__, new_new_n8437__, new_new_n8438__,
    new_new_n8439__, new_new_n8440__, new_new_n8441__, new_new_n8442__,
    new_new_n8443__, new_new_n8444__, new_new_n8445__, new_new_n8446__,
    new_new_n8447__, new_new_n8448__, new_new_n8449__, new_new_n8450__,
    new_new_n8451__, new_new_n8452__, new_new_n8453__, new_new_n8454__,
    new_new_n8455__, new_new_n8456__, new_new_n8457__, new_new_n8458__,
    new_new_n8459__, new_new_n8460__, new_new_n8461__, new_new_n8462__,
    new_new_n8463__, new_new_n8464__, new_new_n8465__, new_new_n8466__,
    new_new_n8467__, new_new_n8468__, new_new_n8469__, new_new_n8470__,
    new_new_n8471__, new_new_n8472__, new_new_n8473__, new_new_n8474__,
    new_new_n8475__, new_new_n8476__, new_new_n8477__, new_new_n8478__,
    new_new_n8479__, new_new_n8480__, new_new_n8481__, new_new_n8482__,
    new_new_n8483__, new_new_n8484__, new_new_n8485__, new_new_n8486__,
    new_new_n8487__, new_new_n8488__, new_new_n8489__, new_new_n8490__,
    new_new_n8491__, new_new_n8492__, new_new_n8493__, new_new_n8494__,
    new_new_n8495__, new_new_n8496__, new_new_n8497__, new_new_n8498__,
    new_new_n8499__, new_new_n8500__, new_new_n8501__, new_new_n8502__,
    new_new_n8503__, new_new_n8504__, new_new_n8505__, new_new_n8506__,
    new_new_n8507__, new_new_n8508__, new_new_n8509__, new_new_n8510__,
    new_new_n8511__, new_new_n8512__, new_new_n8513__, new_new_n8514__,
    new_new_n8515__, new_new_n8516__, new_new_n8517__, new_new_n8518__,
    new_new_n8519__, new_new_n8520__, new_new_n8521__, new_new_n8522__,
    new_new_n8523__, new_new_n8524__, new_new_n8525__, new_new_n8526__,
    new_new_n8527__, new_new_n8528__, new_new_n8529__, new_new_n8530__,
    new_new_n8531__, new_new_n8532__, new_new_n8533__, new_new_n8534__,
    new_new_n8535__, new_new_n8536__, new_new_n8537__, new_new_n8538__,
    new_new_n8539__, new_new_n8540__, new_new_n8541__, new_new_n8542__,
    new_new_n8543__, new_new_n8544__, new_new_n8545__, new_new_n8546__,
    new_new_n8547__, new_new_n8548__, new_new_n8549__, new_new_n8550__,
    new_new_n8551__, new_new_n8552__, new_new_n8553__, new_new_n8554__,
    new_new_n8555__, new_new_n8556__, new_new_n8557__, new_new_n8558__,
    new_new_n8559__, new_new_n8560__, new_new_n8561__, new_new_n8562__,
    new_new_n8563__, new_new_n8564__, new_new_n8565__, new_new_n8566__,
    new_new_n8567__, new_new_n8568__, new_new_n8569__, new_new_n8570__,
    new_new_n8571__, new_new_n8572__, new_new_n8573__, new_new_n8574__,
    new_new_n8575__, new_new_n8576__, new_new_n8577__, new_new_n8578__,
    new_new_n8579__, new_new_n8580__, new_new_n8581__, new_new_n8582__,
    new_new_n8583__, new_new_n8584__, new_new_n8585__, new_new_n8586__,
    new_new_n8587__, new_new_n8588__, new_new_n8589__, new_new_n8590__,
    new_new_n8591__, new_new_n8592__, new_new_n8593__, new_new_n8594__,
    new_new_n8595__, new_new_n8596__, new_new_n8597__, new_new_n8598__,
    new_new_n8599__, new_new_n8600__, new_new_n8601__, new_new_n8602__,
    new_new_n8603__, new_new_n8604__, new_new_n8605__, new_new_n8606__,
    new_new_n8607__, new_new_n8608__, new_new_n8609__, new_new_n8610__,
    new_new_n8611__, new_new_n8612__, new_new_n8613__, new_new_n8614__,
    new_new_n8615__, new_new_n8616__, new_new_n8617__, new_new_n8618__,
    new_new_n8619__, new_new_n8620__, new_new_n8621__, new_new_n8622__,
    new_new_n8623__, new_new_n8624__, new_new_n8625__, new_new_n8626__,
    new_new_n8627__, new_new_n8628__, new_new_n8629__, new_new_n8630__,
    new_new_n8631__, new_new_n8632__, new_new_n8633__, new_new_n8634__,
    new_new_n8635__, new_new_n8636__, new_new_n8637__, new_new_n8638__,
    new_new_n8639__, new_new_n8640__, new_new_n8641__, new_new_n8642__,
    new_new_n8643__, new_new_n8644__, new_new_n8645__, new_new_n8646__,
    new_new_n8647__, new_new_n8648__, new_new_n8649__, new_new_n8650__,
    new_new_n8651__, new_new_n8652__, new_new_n8653__, new_new_n8654__,
    new_new_n8655__, new_new_n8656__, new_new_n8657__, new_new_n8658__,
    new_new_n8659__, new_new_n8660__, new_new_n8661__, new_new_n8662__,
    new_new_n8663__, new_new_n8664__, new_new_n8665__, new_new_n8666__,
    new_new_n8667__, new_new_n8668__, new_new_n8669__, new_new_n8670__,
    new_new_n8671__, new_new_n8672__, new_new_n8673__, new_new_n8674__,
    new_new_n8675__, new_new_n8676__, new_new_n8677__, new_new_n8678__,
    new_new_n8680__, new_new_n8681__, new_new_n8682__, new_new_n8683__,
    new_new_n8684__, new_new_n8685__, new_new_n8686__, new_new_n8687__,
    new_new_n8688__, new_new_n8689__, new_new_n8690__, new_new_n8691__,
    new_new_n8692__, new_new_n8693__, new_new_n8694__, new_new_n8695__,
    new_new_n8696__, new_new_n8697__, new_new_n8698__, new_new_n8699__,
    new_new_n8700__, new_new_n8701__, new_new_n8702__, new_new_n8703__,
    new_new_n8704__, new_new_n8705__, new_new_n8706__, new_new_n8707__,
    new_new_n8708__, new_new_n8709__, new_new_n8710__, new_new_n8711__,
    new_new_n8712__, new_new_n8713__, new_new_n8714__, new_new_n8715__,
    new_new_n8716__, new_new_n8717__, new_new_n8718__, new_new_n8719__,
    new_new_n8720__, new_new_n8721__, new_new_n8722__, new_new_n8723__,
    new_new_n8724__, new_new_n8725__, new_new_n8726__, new_new_n8727__,
    new_new_n8728__, new_new_n8729__, new_new_n8730__, new_new_n8731__,
    new_new_n8732__, new_new_n8733__, new_new_n8734__, new_new_n8735__,
    new_new_n8736__, new_new_n8737__, new_new_n8738__, new_new_n8739__,
    new_new_n8740__, new_new_n8741__, new_new_n8742__, new_new_n8743__,
    new_new_n8744__, new_new_n8745__, new_new_n8746__, new_new_n8747__,
    new_new_n8748__, new_new_n8749__, new_new_n8750__, new_new_n8751__,
    new_new_n8752__, new_new_n8753__, new_new_n8754__, new_new_n8755__,
    new_new_n8756__, new_new_n8757__, new_new_n8758__, new_new_n8759__,
    new_new_n8760__, new_new_n8761__, new_new_n8762__, new_new_n8763__,
    new_new_n8764__, new_new_n8765__, new_new_n8766__, new_new_n8767__,
    new_new_n8768__, new_new_n8769__, new_new_n8770__, new_new_n8771__,
    new_new_n8772__, new_new_n8773__, new_new_n8774__, new_new_n8775__,
    new_new_n8776__, new_new_n8777__, new_new_n8778__, new_new_n8779__,
    new_new_n8780__, new_new_n8781__, new_new_n8782__, new_new_n8783__,
    new_new_n8784__, new_new_n8785__, new_new_n8786__, new_new_n8787__,
    new_new_n8788__, new_new_n8789__, new_new_n8790__, new_new_n8791__,
    new_new_n8792__, new_new_n8793__, new_new_n8794__, new_new_n8795__,
    new_new_n8796__, new_new_n8797__, new_new_n8798__, new_new_n8799__,
    new_new_n8800__, new_new_n8801__, new_new_n8802__, new_new_n8803__,
    new_new_n8804__, new_new_n8805__, new_new_n8806__, new_new_n8807__,
    new_new_n8808__, new_new_n8809__, new_new_n8810__, new_new_n8811__,
    new_new_n8812__, new_new_n8813__, new_new_n8814__, new_new_n8815__,
    new_new_n8816__, new_new_n8817__, new_new_n8818__, new_new_n8819__,
    new_new_n8820__, new_new_n8821__, new_new_n8822__, new_new_n8823__,
    new_new_n8824__, new_new_n8825__, new_new_n8826__, new_new_n8827__,
    new_new_n8828__, new_new_n8829__, new_new_n8830__, new_new_n8831__,
    new_new_n8832__, new_new_n8833__, new_new_n8834__, new_new_n8835__,
    new_new_n8836__, new_new_n8837__, new_new_n8838__, new_new_n8839__,
    new_new_n8840__, new_new_n8841__, new_new_n8842__, new_new_n8843__,
    new_new_n8844__, new_new_n8845__, new_new_n8846__, new_new_n8847__,
    new_new_n8848__, new_new_n8849__, new_new_n8850__, new_new_n8851__,
    new_new_n8852__, new_new_n8853__, new_new_n8854__, new_new_n8855__,
    new_new_n8856__, new_new_n8857__, new_new_n8858__, new_new_n8859__,
    new_new_n8860__, new_new_n8861__, new_new_n8862__, new_new_n8863__,
    new_new_n8864__, new_new_n8865__, new_new_n8866__, new_new_n8867__,
    new_new_n8868__, new_new_n8869__, new_new_n8870__, new_new_n8871__,
    new_new_n8872__, new_new_n8873__, new_new_n8874__, new_new_n8875__,
    new_new_n8876__, new_new_n8877__, new_new_n8878__, new_new_n8879__,
    new_new_n8880__, new_new_n8881__, new_new_n8882__, new_new_n8883__,
    new_new_n8884__, new_new_n8885__, new_new_n8886__, new_new_n8887__,
    new_new_n8888__, new_new_n8889__, new_new_n8890__, new_new_n8891__,
    new_new_n8892__, new_new_n8893__, new_new_n8894__, new_new_n8895__,
    new_new_n8896__, new_new_n8897__, new_new_n8898__, new_new_n8899__,
    new_new_n8900__, new_new_n8901__, new_new_n8902__, new_new_n8903__,
    new_new_n8904__, new_new_n8905__, new_new_n8906__, new_new_n8907__,
    new_new_n8908__, new_new_n8909__, new_new_n8910__, new_new_n8911__,
    new_new_n8912__, new_new_n8913__, new_new_n8914__, new_new_n8915__,
    new_new_n8916__, new_new_n8917__, new_new_n8918__, new_new_n8919__,
    new_new_n8920__, new_new_n8921__, new_new_n8922__, new_new_n8923__,
    new_new_n8924__, new_new_n8925__, new_new_n8926__, new_new_n8927__,
    new_new_n8928__, new_new_n8929__, new_new_n8930__, new_new_n8931__,
    new_new_n8932__, new_new_n8933__, new_new_n8934__, new_new_n8935__,
    new_new_n8936__, new_new_n8937__, new_new_n8938__, new_new_n8939__,
    new_new_n8940__, new_new_n8941__, new_new_n8942__, new_new_n8943__,
    new_new_n8944__, new_new_n8945__, new_new_n8946__, new_new_n8947__,
    new_new_n8948__, new_new_n8949__, new_new_n8950__, new_new_n8951__,
    new_new_n8952__, new_new_n8953__, new_new_n8954__, new_new_n8955__,
    new_new_n8956__, new_new_n8957__, new_new_n8958__, new_new_n8959__,
    new_new_n8960__, new_new_n8961__, new_new_n8962__, new_new_n8963__,
    new_new_n8964__, new_new_n8965__, new_new_n8966__, new_new_n8967__,
    new_new_n8968__, new_new_n8969__, new_new_n8970__, new_new_n8971__,
    new_new_n8972__, new_new_n8973__, new_new_n8974__, new_new_n8975__,
    new_new_n8977__, new_new_n8978__, new_new_n8979__, new_new_n8980__,
    new_new_n8981__, new_new_n8982__, new_new_n8983__, new_new_n8984__,
    new_new_n8985__, new_new_n8986__, new_new_n8987__, new_new_n8988__,
    new_new_n8989__, new_new_n8990__, new_new_n8991__, new_new_n8992__,
    new_new_n8993__, new_new_n8994__, new_new_n8995__, new_new_n8996__,
    new_new_n8997__, new_new_n8998__, new_new_n8999__, new_new_n9000__,
    new_new_n9001__, new_new_n9002__, new_new_n9003__, new_new_n9004__,
    new_new_n9005__, new_new_n9006__, new_new_n9007__, new_new_n9008__,
    new_new_n9009__, new_new_n9010__, new_new_n9011__, new_new_n9012__,
    new_new_n9013__, new_new_n9014__, new_new_n9015__, new_new_n9016__,
    new_new_n9017__, new_new_n9018__, new_new_n9019__, new_new_n9020__,
    new_new_n9021__, new_new_n9022__, new_new_n9023__, new_new_n9024__,
    new_new_n9025__, new_new_n9026__, new_new_n9027__, new_new_n9028__,
    new_new_n9029__, new_new_n9030__, new_new_n9031__, new_new_n9032__,
    new_new_n9033__, new_new_n9034__, new_new_n9035__, new_new_n9036__,
    new_new_n9037__, new_new_n9038__, new_new_n9039__, new_new_n9040__,
    new_new_n9041__, new_new_n9042__, new_new_n9043__, new_new_n9044__,
    new_new_n9045__, new_new_n9046__, new_new_n9047__, new_new_n9048__,
    new_new_n9049__, new_new_n9050__, new_new_n9051__, new_new_n9052__,
    new_new_n9053__, new_new_n9054__, new_new_n9055__, new_new_n9056__,
    new_new_n9057__, new_new_n9058__, new_new_n9059__, new_new_n9060__,
    new_new_n9061__, new_new_n9062__, new_new_n9063__, new_new_n9064__,
    new_new_n9065__, new_new_n9066__, new_new_n9067__, new_new_n9068__,
    new_new_n9069__, new_new_n9070__, new_new_n9071__, new_new_n9072__,
    new_new_n9073__, new_new_n9074__, new_new_n9075__, new_new_n9076__,
    new_new_n9077__, new_new_n9078__, new_new_n9079__, new_new_n9080__,
    new_new_n9081__, new_new_n9082__, new_new_n9083__, new_new_n9084__,
    new_new_n9085__, new_new_n9086__, new_new_n9087__, new_new_n9088__,
    new_new_n9089__, new_new_n9090__, new_new_n9091__, new_new_n9092__,
    new_new_n9093__, new_new_n9094__, new_new_n9095__, new_new_n9096__,
    new_new_n9097__, new_new_n9098__, new_new_n9099__, new_new_n9100__,
    new_new_n9101__, new_new_n9102__, new_new_n9103__, new_new_n9104__,
    new_new_n9105__, new_new_n9106__, new_new_n9107__, new_new_n9108__,
    new_new_n9109__, new_new_n9110__, new_new_n9111__, new_new_n9112__,
    new_new_n9113__, new_new_n9114__, new_new_n9115__, new_new_n9116__,
    new_new_n9117__, new_new_n9118__, new_new_n9119__, new_new_n9120__,
    new_new_n9121__, new_new_n9122__, new_new_n9123__, new_new_n9124__,
    new_new_n9125__, new_new_n9126__, new_new_n9127__, new_new_n9128__,
    new_new_n9129__, new_new_n9130__, new_new_n9131__, new_new_n9132__,
    new_new_n9133__, new_new_n9134__, new_new_n9135__, new_new_n9136__,
    new_new_n9137__, new_new_n9138__, new_new_n9139__, new_new_n9140__,
    new_new_n9141__, new_new_n9142__, new_new_n9143__, new_new_n9144__,
    new_new_n9145__, new_new_n9146__, new_new_n9147__, new_new_n9148__,
    new_new_n9149__, new_new_n9150__, new_new_n9151__, new_new_n9152__,
    new_new_n9153__, new_new_n9154__, new_new_n9155__, new_new_n9156__,
    new_new_n9157__, new_new_n9158__, new_new_n9159__, new_new_n9160__,
    new_new_n9161__, new_new_n9162__, new_new_n9163__, new_new_n9164__,
    new_new_n9165__, new_new_n9166__, new_new_n9167__, new_new_n9168__,
    new_new_n9169__, new_new_n9170__, new_new_n9171__, new_new_n9172__,
    new_new_n9173__, new_new_n9174__, new_new_n9175__, new_new_n9176__,
    new_new_n9177__, new_new_n9178__, new_new_n9179__, new_new_n9180__,
    new_new_n9181__, new_new_n9182__, new_new_n9183__, new_new_n9184__,
    new_new_n9185__, new_new_n9186__, new_new_n9187__, new_new_n9188__,
    new_new_n9189__, new_new_n9190__, new_new_n9191__, new_new_n9192__,
    new_new_n9193__, new_new_n9194__, new_new_n9195__, new_new_n9196__,
    new_new_n9197__, new_new_n9198__, new_new_n9199__, new_new_n9200__,
    new_new_n9201__, new_new_n9202__, new_new_n9203__, new_new_n9204__,
    new_new_n9205__, new_new_n9206__, new_new_n9207__, new_new_n9208__,
    new_new_n9209__, new_new_n9210__, new_new_n9211__, new_new_n9212__,
    new_new_n9213__, new_new_n9214__, new_new_n9215__, new_new_n9216__,
    new_new_n9217__, new_new_n9218__, new_new_n9219__, new_new_n9220__,
    new_new_n9221__, new_new_n9222__, new_new_n9223__, new_new_n9224__,
    new_new_n9225__, new_new_n9226__, new_new_n9227__, new_new_n9228__,
    new_new_n9229__, new_new_n9230__, new_new_n9231__, new_new_n9232__,
    new_new_n9233__, new_new_n9234__, new_new_n9235__, new_new_n9236__,
    new_new_n9237__, new_new_n9238__, new_new_n9239__, new_new_n9240__,
    new_new_n9241__, new_new_n9242__, new_new_n9243__, new_new_n9244__,
    new_new_n9245__, new_new_n9246__, new_new_n9247__, new_new_n9248__,
    new_new_n9249__, new_new_n9250__, new_new_n9251__, new_new_n9252__,
    new_new_n9253__, new_new_n9254__, new_new_n9255__, new_new_n9256__,
    new_new_n9258__, new_new_n9259__, new_new_n9260__, new_new_n9261__,
    new_new_n9262__, new_new_n9263__, new_new_n9264__, new_new_n9265__,
    new_new_n9266__, new_new_n9267__, new_new_n9268__, new_new_n9269__,
    new_new_n9270__, new_new_n9271__, new_new_n9272__, new_new_n9273__,
    new_new_n9274__, new_new_n9275__, new_new_n9276__, new_new_n9277__,
    new_new_n9278__, new_new_n9279__, new_new_n9280__, new_new_n9281__,
    new_new_n9282__, new_new_n9283__, new_new_n9284__, new_new_n9285__,
    new_new_n9286__, new_new_n9287__, new_new_n9288__, new_new_n9289__,
    new_new_n9290__, new_new_n9291__, new_new_n9292__, new_new_n9293__,
    new_new_n9294__, new_new_n9295__, new_new_n9296__, new_new_n9297__,
    new_new_n9298__, new_new_n9299__, new_new_n9300__, new_new_n9301__,
    new_new_n9302__, new_new_n9303__, new_new_n9304__, new_new_n9305__,
    new_new_n9306__, new_new_n9307__, new_new_n9308__, new_new_n9309__,
    new_new_n9310__, new_new_n9311__, new_new_n9312__, new_new_n9313__,
    new_new_n9314__, new_new_n9315__, new_new_n9316__, new_new_n9317__,
    new_new_n9318__, new_new_n9319__, new_new_n9320__, new_new_n9321__,
    new_new_n9322__, new_new_n9323__, new_new_n9324__, new_new_n9325__,
    new_new_n9326__, new_new_n9327__, new_new_n9328__, new_new_n9329__,
    new_new_n9330__, new_new_n9331__, new_new_n9332__, new_new_n9333__,
    new_new_n9334__, new_new_n9335__, new_new_n9336__, new_new_n9337__,
    new_new_n9338__, new_new_n9339__, new_new_n9340__, new_new_n9341__,
    new_new_n9342__, new_new_n9343__, new_new_n9344__, new_new_n9345__,
    new_new_n9346__, new_new_n9347__, new_new_n9348__, new_new_n9349__,
    new_new_n9350__, new_new_n9351__, new_new_n9352__, new_new_n9353__,
    new_new_n9354__, new_new_n9355__, new_new_n9356__, new_new_n9357__,
    new_new_n9358__, new_new_n9359__, new_new_n9360__, new_new_n9361__,
    new_new_n9362__, new_new_n9363__, new_new_n9364__, new_new_n9365__,
    new_new_n9366__, new_new_n9367__, new_new_n9368__, new_new_n9369__,
    new_new_n9370__, new_new_n9371__, new_new_n9372__, new_new_n9373__,
    new_new_n9374__, new_new_n9375__, new_new_n9376__, new_new_n9377__,
    new_new_n9378__, new_new_n9379__, new_new_n9380__, new_new_n9381__,
    new_new_n9382__, new_new_n9383__, new_new_n9384__, new_new_n9385__,
    new_new_n9386__, new_new_n9387__, new_new_n9388__, new_new_n9389__,
    new_new_n9390__, new_new_n9391__, new_new_n9392__, new_new_n9393__,
    new_new_n9394__, new_new_n9395__, new_new_n9396__, new_new_n9397__,
    new_new_n9398__, new_new_n9399__, new_new_n9400__, new_new_n9401__,
    new_new_n9402__, new_new_n9403__, new_new_n9404__, new_new_n9405__,
    new_new_n9406__, new_new_n9407__, new_new_n9408__, new_new_n9409__,
    new_new_n9410__, new_new_n9411__, new_new_n9412__, new_new_n9413__,
    new_new_n9414__, new_new_n9415__, new_new_n9416__, new_new_n9417__,
    new_new_n9418__, new_new_n9419__, new_new_n9420__, new_new_n9421__,
    new_new_n9422__, new_new_n9423__, new_new_n9424__, new_new_n9425__,
    new_new_n9426__, new_new_n9427__, new_new_n9428__, new_new_n9429__,
    new_new_n9430__, new_new_n9431__, new_new_n9432__, new_new_n9433__,
    new_new_n9434__, new_new_n9435__, new_new_n9436__, new_new_n9437__,
    new_new_n9438__, new_new_n9439__, new_new_n9440__, new_new_n9441__,
    new_new_n9442__, new_new_n9443__, new_new_n9444__, new_new_n9445__,
    new_new_n9446__, new_new_n9447__, new_new_n9448__, new_new_n9449__,
    new_new_n9450__, new_new_n9451__, new_new_n9452__, new_new_n9453__,
    new_new_n9454__, new_new_n9455__, new_new_n9456__, new_new_n9457__,
    new_new_n9458__, new_new_n9459__, new_new_n9460__, new_new_n9461__,
    new_new_n9462__, new_new_n9463__, new_new_n9464__, new_new_n9465__,
    new_new_n9466__, new_new_n9467__, new_new_n9468__, new_new_n9469__,
    new_new_n9470__, new_new_n9471__, new_new_n9472__, new_new_n9473__,
    new_new_n9474__, new_new_n9475__, new_new_n9476__, new_new_n9477__,
    new_new_n9478__, new_new_n9479__, new_new_n9480__, new_new_n9481__,
    new_new_n9482__, new_new_n9483__, new_new_n9484__, new_new_n9485__,
    new_new_n9486__, new_new_n9487__, new_new_n9488__, new_new_n9489__,
    new_new_n9490__, new_new_n9491__, new_new_n9492__, new_new_n9493__,
    new_new_n9494__, new_new_n9495__, new_new_n9496__, new_new_n9497__,
    new_new_n9498__, new_new_n9499__, new_new_n9500__, new_new_n9501__,
    new_new_n9502__, new_new_n9503__, new_new_n9504__, new_new_n9505__,
    new_new_n9506__, new_new_n9507__, new_new_n9508__, new_new_n9509__,
    new_new_n9510__, new_new_n9511__, new_new_n9512__, new_new_n9513__,
    new_new_n9514__, new_new_n9515__, new_new_n9516__, new_new_n9517__,
    new_new_n9518__, new_new_n9519__, new_new_n9520__, new_new_n9521__,
    new_new_n9522__, new_new_n9523__, new_new_n9524__, new_new_n9525__,
    new_new_n9526__, new_new_n9527__, new_new_n9528__, new_new_n9529__,
    new_new_n9530__, new_new_n9531__, new_new_n9532__, new_new_n9533__,
    new_new_n9534__, new_new_n9535__, new_new_n9536__, new_new_n9537__,
    new_new_n9538__, new_new_n9539__, new_new_n9540__, new_new_n9541__,
    new_new_n9542__, new_new_n9543__, new_new_n9544__, new_new_n9545__,
    new_new_n9546__, new_new_n9547__, new_new_n9548__, new_new_n9549__,
    new_new_n9550__, new_new_n9551__, new_new_n9552__, new_new_n9553__,
    new_new_n9554__, new_new_n9555__, new_new_n9556__, new_new_n9557__,
    new_new_n9558__, new_new_n9559__, new_new_n9560__, new_new_n9562__,
    new_new_n9563__, new_new_n9564__, new_new_n9565__, new_new_n9566__,
    new_new_n9567__, new_new_n9568__, new_new_n9569__, new_new_n9570__,
    new_new_n9571__, new_new_n9572__, new_new_n9573__, new_new_n9574__,
    new_new_n9575__, new_new_n9576__, new_new_n9577__, new_new_n9578__,
    new_new_n9579__, new_new_n9580__, new_new_n9581__, new_new_n9582__,
    new_new_n9583__, new_new_n9584__, new_new_n9585__, new_new_n9586__,
    new_new_n9587__, new_new_n9588__, new_new_n9589__, new_new_n9590__,
    new_new_n9591__, new_new_n9592__, new_new_n9593__, new_new_n9594__,
    new_new_n9595__, new_new_n9596__, new_new_n9597__, new_new_n9598__,
    new_new_n9599__, new_new_n9600__, new_new_n9601__, new_new_n9602__,
    new_new_n9603__, new_new_n9604__, new_new_n9605__, new_new_n9606__,
    new_new_n9607__, new_new_n9608__, new_new_n9609__, new_new_n9610__,
    new_new_n9611__, new_new_n9612__, new_new_n9613__, new_new_n9614__,
    new_new_n9615__, new_new_n9616__, new_new_n9617__, new_new_n9618__,
    new_new_n9619__, new_new_n9620__, new_new_n9621__, new_new_n9622__,
    new_new_n9623__, new_new_n9624__, new_new_n9625__, new_new_n9626__,
    new_new_n9627__, new_new_n9628__, new_new_n9629__, new_new_n9630__,
    new_new_n9631__, new_new_n9632__, new_new_n9633__, new_new_n9634__,
    new_new_n9635__, new_new_n9636__, new_new_n9637__, new_new_n9638__,
    new_new_n9639__, new_new_n9640__, new_new_n9641__, new_new_n9642__,
    new_new_n9643__, new_new_n9644__, new_new_n9645__, new_new_n9646__,
    new_new_n9647__, new_new_n9648__, new_new_n9649__, new_new_n9650__,
    new_new_n9651__, new_new_n9652__, new_new_n9653__, new_new_n9654__,
    new_new_n9655__, new_new_n9656__, new_new_n9657__, new_new_n9658__,
    new_new_n9659__, new_new_n9660__, new_new_n9661__, new_new_n9662__,
    new_new_n9663__, new_new_n9664__, new_new_n9665__, new_new_n9666__,
    new_new_n9667__, new_new_n9668__, new_new_n9669__, new_new_n9670__,
    new_new_n9671__, new_new_n9672__, new_new_n9673__, new_new_n9674__,
    new_new_n9675__, new_new_n9676__, new_new_n9677__, new_new_n9678__,
    new_new_n9679__, new_new_n9680__, new_new_n9681__, new_new_n9682__,
    new_new_n9683__, new_new_n9684__, new_new_n9685__, new_new_n9686__,
    new_new_n9687__, new_new_n9688__, new_new_n9689__, new_new_n9690__,
    new_new_n9691__, new_new_n9692__, new_new_n9693__, new_new_n9694__,
    new_new_n9695__, new_new_n9696__, new_new_n9697__, new_new_n9698__,
    new_new_n9699__, new_new_n9700__, new_new_n9701__, new_new_n9702__,
    new_new_n9703__, new_new_n9704__, new_new_n9705__, new_new_n9706__,
    new_new_n9707__, new_new_n9708__, new_new_n9709__, new_new_n9710__,
    new_new_n9711__, new_new_n9712__, new_new_n9713__, new_new_n9714__,
    new_new_n9715__, new_new_n9716__, new_new_n9717__, new_new_n9718__,
    new_new_n9719__, new_new_n9720__, new_new_n9721__, new_new_n9722__,
    new_new_n9723__, new_new_n9724__, new_new_n9725__, new_new_n9726__,
    new_new_n9727__, new_new_n9728__, new_new_n9729__, new_new_n9730__,
    new_new_n9731__, new_new_n9732__, new_new_n9733__, new_new_n9734__,
    new_new_n9735__, new_new_n9736__, new_new_n9737__, new_new_n9738__,
    new_new_n9739__, new_new_n9740__, new_new_n9741__, new_new_n9742__,
    new_new_n9743__, new_new_n9744__, new_new_n9745__, new_new_n9746__,
    new_new_n9747__, new_new_n9748__, new_new_n9749__, new_new_n9750__,
    new_new_n9751__, new_new_n9752__, new_new_n9753__, new_new_n9754__,
    new_new_n9755__, new_new_n9756__, new_new_n9757__, new_new_n9758__,
    new_new_n9759__, new_new_n9760__, new_new_n9761__, new_new_n9762__,
    new_new_n9763__, new_new_n9764__, new_new_n9765__, new_new_n9766__,
    new_new_n9767__, new_new_n9768__, new_new_n9769__, new_new_n9770__,
    new_new_n9771__, new_new_n9772__, new_new_n9773__, new_new_n9774__,
    new_new_n9775__, new_new_n9776__, new_new_n9777__, new_new_n9778__,
    new_new_n9779__, new_new_n9780__, new_new_n9781__, new_new_n9782__,
    new_new_n9783__, new_new_n9784__, new_new_n9785__, new_new_n9786__,
    new_new_n9787__, new_new_n9788__, new_new_n9789__, new_new_n9790__,
    new_new_n9791__, new_new_n9792__, new_new_n9793__, new_new_n9794__,
    new_new_n9795__, new_new_n9796__, new_new_n9797__, new_new_n9798__,
    new_new_n9799__, new_new_n9800__, new_new_n9801__, new_new_n9802__,
    new_new_n9803__, new_new_n9804__, new_new_n9805__, new_new_n9806__,
    new_new_n9807__, new_new_n9808__, new_new_n9809__, new_new_n9810__,
    new_new_n9811__, new_new_n9812__, new_new_n9813__, new_new_n9814__,
    new_new_n9815__, new_new_n9816__, new_new_n9817__, new_new_n9818__,
    new_new_n9819__, new_new_n9820__, new_new_n9821__, new_new_n9822__,
    new_new_n9823__, new_new_n9824__, new_new_n9825__, new_new_n9826__,
    new_new_n9827__, new_new_n9828__, new_new_n9829__, new_new_n9830__,
    new_new_n9831__, new_new_n9832__, new_new_n9833__, new_new_n9834__,
    new_new_n9835__, new_new_n9836__, new_new_n9837__, new_new_n9838__,
    new_new_n9839__, new_new_n9840__, new_new_n9841__, new_new_n9842__,
    new_new_n9843__, new_new_n9845__, new_new_n9846__, new_new_n9847__,
    new_new_n9848__, new_new_n9849__, new_new_n9850__, new_new_n9851__,
    new_new_n9852__, new_new_n9853__, new_new_n9854__, new_new_n9855__,
    new_new_n9856__, new_new_n9857__, new_new_n9858__, new_new_n9859__,
    new_new_n9860__, new_new_n9861__, new_new_n9862__, new_new_n9863__,
    new_new_n9864__, new_new_n9865__, new_new_n9866__, new_new_n9867__,
    new_new_n9868__, new_new_n9869__, new_new_n9870__, new_new_n9871__,
    new_new_n9872__, new_new_n9873__, new_new_n9874__, new_new_n9875__,
    new_new_n9876__, new_new_n9877__, new_new_n9878__, new_new_n9879__,
    new_new_n9880__, new_new_n9881__, new_new_n9882__, new_new_n9883__,
    new_new_n9884__, new_new_n9885__, new_new_n9886__, new_new_n9887__,
    new_new_n9888__, new_new_n9889__, new_new_n9890__, new_new_n9891__,
    new_new_n9892__, new_new_n9893__, new_new_n9894__, new_new_n9895__,
    new_new_n9896__, new_new_n9897__, new_new_n9898__, new_new_n9899__,
    new_new_n9900__, new_new_n9901__, new_new_n9902__, new_new_n9903__,
    new_new_n9904__, new_new_n9905__, new_new_n9906__, new_new_n9907__,
    new_new_n9908__, new_new_n9909__, new_new_n9910__, new_new_n9911__,
    new_new_n9912__, new_new_n9913__, new_new_n9914__, new_new_n9915__,
    new_new_n9916__, new_new_n9917__, new_new_n9918__, new_new_n9919__,
    new_new_n9920__, new_new_n9921__, new_new_n9922__, new_new_n9923__,
    new_new_n9924__, new_new_n9925__, new_new_n9926__, new_new_n9927__,
    new_new_n9928__, new_new_n9929__, new_new_n9930__, new_new_n9931__,
    new_new_n9932__, new_new_n9933__, new_new_n9934__, new_new_n9935__,
    new_new_n9936__, new_new_n9937__, new_new_n9938__, new_new_n9939__,
    new_new_n9940__, new_new_n9941__, new_new_n9942__, new_new_n9943__,
    new_new_n9944__, new_new_n9945__, new_new_n9946__, new_new_n9947__,
    new_new_n9948__, new_new_n9949__, new_new_n9950__, new_new_n9951__,
    new_new_n9952__, new_new_n9953__, new_new_n9954__, new_new_n9955__,
    new_new_n9956__, new_new_n9957__, new_new_n9958__, new_new_n9959__,
    new_new_n9960__, new_new_n9961__, new_new_n9962__, new_new_n9963__,
    new_new_n9964__, new_new_n9965__, new_new_n9966__, new_new_n9967__,
    new_new_n9968__, new_new_n9969__, new_new_n9970__, new_new_n9971__,
    new_new_n9972__, new_new_n9973__, new_new_n9974__, new_new_n9975__,
    new_new_n9976__, new_new_n9977__, new_new_n9978__, new_new_n9979__,
    new_new_n9980__, new_new_n9981__, new_new_n9982__, new_new_n9983__,
    new_new_n9984__, new_new_n9985__, new_new_n9986__, new_new_n9987__,
    new_new_n9988__, new_new_n9989__, new_new_n9990__, new_new_n9991__,
    new_new_n9992__, new_new_n9993__, new_new_n9994__, new_new_n9995__,
    new_new_n9996__, new_new_n9997__, new_new_n9998__, new_new_n9999__,
    new_new_n10000__, new_new_n10001__, new_new_n10002__, new_new_n10003__,
    new_new_n10004__, new_new_n10005__, new_new_n10006__, new_new_n10007__,
    new_new_n10008__, new_new_n10009__, new_new_n10010__, new_new_n10011__,
    new_new_n10012__, new_new_n10013__, new_new_n10014__, new_new_n10015__,
    new_new_n10016__, new_new_n10017__, new_new_n10018__, new_new_n10019__,
    new_new_n10020__, new_new_n10021__, new_new_n10022__, new_new_n10023__,
    new_new_n10024__, new_new_n10025__, new_new_n10026__, new_new_n10027__,
    new_new_n10028__, new_new_n10029__, new_new_n10030__, new_new_n10031__,
    new_new_n10032__, new_new_n10033__, new_new_n10034__, new_new_n10035__,
    new_new_n10036__, new_new_n10037__, new_new_n10038__, new_new_n10039__,
    new_new_n10040__, new_new_n10041__, new_new_n10042__, new_new_n10043__,
    new_new_n10044__, new_new_n10045__, new_new_n10046__, new_new_n10047__,
    new_new_n10048__, new_new_n10049__, new_new_n10050__, new_new_n10051__,
    new_new_n10052__, new_new_n10053__, new_new_n10054__, new_new_n10055__,
    new_new_n10056__, new_new_n10057__, new_new_n10058__, new_new_n10059__,
    new_new_n10060__, new_new_n10061__, new_new_n10062__, new_new_n10063__,
    new_new_n10064__, new_new_n10065__, new_new_n10066__, new_new_n10067__,
    new_new_n10068__, new_new_n10069__, new_new_n10070__, new_new_n10071__,
    new_new_n10072__, new_new_n10073__, new_new_n10074__, new_new_n10075__,
    new_new_n10076__, new_new_n10077__, new_new_n10078__, new_new_n10079__,
    new_new_n10080__, new_new_n10081__, new_new_n10082__, new_new_n10083__,
    new_new_n10084__, new_new_n10085__, new_new_n10086__, new_new_n10087__,
    new_new_n10088__, new_new_n10089__, new_new_n10090__, new_new_n10091__,
    new_new_n10092__, new_new_n10093__, new_new_n10094__, new_new_n10095__,
    new_new_n10096__, new_new_n10097__, new_new_n10098__, new_new_n10099__,
    new_new_n10100__, new_new_n10101__, new_new_n10102__, new_new_n10103__,
    new_new_n10104__, new_new_n10105__, new_new_n10106__, new_new_n10107__,
    new_new_n10108__, new_new_n10109__, new_new_n10110__, new_new_n10111__,
    new_new_n10112__, new_new_n10113__, new_new_n10114__, new_new_n10115__,
    new_new_n10116__, new_new_n10117__, new_new_n10118__, new_new_n10119__,
    new_new_n10120__, new_new_n10121__, new_new_n10122__, new_new_n10123__,
    new_new_n10124__, new_new_n10125__, new_new_n10126__, new_new_n10127__,
    new_new_n10128__, new_new_n10129__, new_new_n10130__, new_new_n10132__,
    new_new_n10133__, new_new_n10134__, new_new_n10135__, new_new_n10136__,
    new_new_n10137__, new_new_n10138__, new_new_n10139__, new_new_n10140__,
    new_new_n10141__, new_new_n10142__, new_new_n10143__, new_new_n10144__,
    new_new_n10145__, new_new_n10146__, new_new_n10147__, new_new_n10148__,
    new_new_n10149__, new_new_n10150__, new_new_n10151__, new_new_n10152__,
    new_new_n10153__, new_new_n10154__, new_new_n10155__, new_new_n10156__,
    new_new_n10157__, new_new_n10158__, new_new_n10159__, new_new_n10160__,
    new_new_n10161__, new_new_n10162__, new_new_n10163__, new_new_n10164__,
    new_new_n10165__, new_new_n10166__, new_new_n10167__, new_new_n10168__,
    new_new_n10169__, new_new_n10170__, new_new_n10171__, new_new_n10172__,
    new_new_n10173__, new_new_n10174__, new_new_n10175__, new_new_n10176__,
    new_new_n10177__, new_new_n10178__, new_new_n10179__, new_new_n10180__,
    new_new_n10181__, new_new_n10182__, new_new_n10183__, new_new_n10184__,
    new_new_n10185__, new_new_n10186__, new_new_n10187__, new_new_n10188__,
    new_new_n10189__, new_new_n10190__, new_new_n10191__, new_new_n10192__,
    new_new_n10193__, new_new_n10194__, new_new_n10195__, new_new_n10196__,
    new_new_n10197__, new_new_n10198__, new_new_n10199__, new_new_n10200__,
    new_new_n10201__, new_new_n10202__, new_new_n10203__, new_new_n10204__,
    new_new_n10205__, new_new_n10206__, new_new_n10207__, new_new_n10208__,
    new_new_n10209__, new_new_n10210__, new_new_n10211__, new_new_n10212__,
    new_new_n10213__, new_new_n10214__, new_new_n10215__, new_new_n10216__,
    new_new_n10217__, new_new_n10218__, new_new_n10219__, new_new_n10220__,
    new_new_n10221__, new_new_n10222__, new_new_n10223__, new_new_n10224__,
    new_new_n10225__, new_new_n10226__, new_new_n10227__, new_new_n10228__,
    new_new_n10229__, new_new_n10230__, new_new_n10231__, new_new_n10232__,
    new_new_n10233__, new_new_n10234__, new_new_n10235__, new_new_n10236__,
    new_new_n10237__, new_new_n10238__, new_new_n10239__, new_new_n10240__,
    new_new_n10241__, new_new_n10242__, new_new_n10243__, new_new_n10244__,
    new_new_n10245__, new_new_n10246__, new_new_n10247__, new_new_n10248__,
    new_new_n10249__, new_new_n10250__, new_new_n10251__, new_new_n10252__,
    new_new_n10253__, new_new_n10254__, new_new_n10255__, new_new_n10256__,
    new_new_n10257__, new_new_n10258__, new_new_n10259__, new_new_n10260__,
    new_new_n10261__, new_new_n10262__, new_new_n10263__, new_new_n10264__,
    new_new_n10265__, new_new_n10266__, new_new_n10267__, new_new_n10268__,
    new_new_n10269__, new_new_n10270__, new_new_n10271__, new_new_n10272__,
    new_new_n10273__, new_new_n10274__, new_new_n10275__, new_new_n10276__,
    new_new_n10277__, new_new_n10278__, new_new_n10279__, new_new_n10280__,
    new_new_n10281__, new_new_n10282__, new_new_n10283__, new_new_n10284__,
    new_new_n10285__, new_new_n10286__, new_new_n10287__, new_new_n10288__,
    new_new_n10289__, new_new_n10290__, new_new_n10291__, new_new_n10292__,
    new_new_n10293__, new_new_n10294__, new_new_n10295__, new_new_n10296__,
    new_new_n10297__, new_new_n10298__, new_new_n10299__, new_new_n10300__,
    new_new_n10301__, new_new_n10302__, new_new_n10303__, new_new_n10304__,
    new_new_n10305__, new_new_n10306__, new_new_n10307__, new_new_n10308__,
    new_new_n10309__, new_new_n10310__, new_new_n10311__, new_new_n10312__,
    new_new_n10313__, new_new_n10314__, new_new_n10315__, new_new_n10316__,
    new_new_n10317__, new_new_n10318__, new_new_n10319__, new_new_n10320__,
    new_new_n10321__, new_new_n10322__, new_new_n10323__, new_new_n10324__,
    new_new_n10325__, new_new_n10326__, new_new_n10327__, new_new_n10328__,
    new_new_n10329__, new_new_n10330__, new_new_n10331__, new_new_n10332__,
    new_new_n10333__, new_new_n10334__, new_new_n10335__, new_new_n10336__,
    new_new_n10337__, new_new_n10338__, new_new_n10339__, new_new_n10340__,
    new_new_n10341__, new_new_n10342__, new_new_n10343__, new_new_n10344__,
    new_new_n10345__, new_new_n10346__, new_new_n10347__, new_new_n10348__,
    new_new_n10349__, new_new_n10350__, new_new_n10351__, new_new_n10352__,
    new_new_n10353__, new_new_n10354__, new_new_n10355__, new_new_n10356__,
    new_new_n10357__, new_new_n10358__, new_new_n10359__, new_new_n10360__,
    new_new_n10361__, new_new_n10362__, new_new_n10363__, new_new_n10364__,
    new_new_n10365__, new_new_n10366__, new_new_n10367__, new_new_n10368__,
    new_new_n10369__, new_new_n10370__, new_new_n10371__, new_new_n10372__,
    new_new_n10373__, new_new_n10374__, new_new_n10375__, new_new_n10376__,
    new_new_n10377__, new_new_n10378__, new_new_n10379__, new_new_n10380__,
    new_new_n10381__, new_new_n10382__, new_new_n10383__, new_new_n10384__,
    new_new_n10385__, new_new_n10386__, new_new_n10387__, new_new_n10388__,
    new_new_n10389__, new_new_n10390__, new_new_n10391__, new_new_n10392__,
    new_new_n10393__, new_new_n10394__, new_new_n10395__, new_new_n10396__,
    new_new_n10397__, new_new_n10398__, new_new_n10399__, new_new_n10400__,
    new_new_n10401__, new_new_n10402__, new_new_n10403__, new_new_n10404__,
    new_new_n10405__, new_new_n10406__, new_new_n10407__, new_new_n10408__,
    new_new_n10409__, new_new_n10410__, new_new_n10411__, new_new_n10412__,
    new_new_n10413__, new_new_n10414__, new_new_n10415__, new_new_n10416__,
    new_new_n10417__, new_new_n10418__, new_new_n10419__, new_new_n10420__,
    new_new_n10421__, new_new_n10422__, new_new_n10423__, new_new_n10424__,
    new_new_n10425__, new_new_n10426__, new_new_n10427__, new_new_n10428__,
    new_new_n10429__, new_new_n10430__, new_new_n10431__, new_new_n10432__,
    new_new_n10433__, new_new_n10434__, new_new_n10435__, new_new_n10436__,
    new_new_n10437__, new_new_n10438__, new_new_n10439__, new_new_n10440__,
    new_new_n10441__, new_new_n10442__, new_new_n10443__, new_new_n10444__,
    new_new_n10445__, new_new_n10446__, new_new_n10447__, new_new_n10449__,
    new_new_n10450__, new_new_n10451__, new_new_n10452__, new_new_n10453__,
    new_new_n10454__, new_new_n10455__, new_new_n10456__, new_new_n10457__,
    new_new_n10458__, new_new_n10459__, new_new_n10460__, new_new_n10461__,
    new_new_n10462__, new_new_n10463__, new_new_n10464__, new_new_n10465__,
    new_new_n10466__, new_new_n10467__, new_new_n10468__, new_new_n10469__,
    new_new_n10470__, new_new_n10471__, new_new_n10472__, new_new_n10473__,
    new_new_n10474__, new_new_n10475__, new_new_n10476__, new_new_n10477__,
    new_new_n10478__, new_new_n10479__, new_new_n10480__, new_new_n10481__,
    new_new_n10482__, new_new_n10483__, new_new_n10484__, new_new_n10485__,
    new_new_n10486__, new_new_n10487__, new_new_n10488__, new_new_n10489__,
    new_new_n10490__, new_new_n10491__, new_new_n10492__, new_new_n10493__,
    new_new_n10494__, new_new_n10495__, new_new_n10496__, new_new_n10497__,
    new_new_n10498__, new_new_n10499__, new_new_n10500__, new_new_n10501__,
    new_new_n10502__, new_new_n10503__, new_new_n10504__, new_new_n10505__,
    new_new_n10506__, new_new_n10507__, new_new_n10508__, new_new_n10509__,
    new_new_n10510__, new_new_n10511__, new_new_n10512__, new_new_n10513__,
    new_new_n10514__, new_new_n10515__, new_new_n10516__, new_new_n10517__,
    new_new_n10518__, new_new_n10519__, new_new_n10520__, new_new_n10521__,
    new_new_n10522__, new_new_n10523__, new_new_n10524__, new_new_n10525__,
    new_new_n10526__, new_new_n10527__, new_new_n10528__, new_new_n10529__,
    new_new_n10530__, new_new_n10531__, new_new_n10532__, new_new_n10533__,
    new_new_n10534__, new_new_n10535__, new_new_n10536__, new_new_n10537__,
    new_new_n10538__, new_new_n10539__, new_new_n10540__, new_new_n10541__,
    new_new_n10542__, new_new_n10543__, new_new_n10544__, new_new_n10545__,
    new_new_n10546__, new_new_n10547__, new_new_n10548__, new_new_n10549__,
    new_new_n10550__, new_new_n10551__, new_new_n10552__, new_new_n10553__,
    new_new_n10554__, new_new_n10555__, new_new_n10556__, new_new_n10557__,
    new_new_n10558__, new_new_n10559__, new_new_n10560__, new_new_n10561__,
    new_new_n10562__, new_new_n10563__, new_new_n10564__, new_new_n10565__,
    new_new_n10566__, new_new_n10567__, new_new_n10568__, new_new_n10569__,
    new_new_n10570__, new_new_n10571__, new_new_n10572__, new_new_n10573__,
    new_new_n10574__, new_new_n10575__, new_new_n10576__, new_new_n10577__,
    new_new_n10578__, new_new_n10579__, new_new_n10580__, new_new_n10581__,
    new_new_n10582__, new_new_n10583__, new_new_n10584__, new_new_n10585__,
    new_new_n10586__, new_new_n10587__, new_new_n10588__, new_new_n10589__,
    new_new_n10590__, new_new_n10591__, new_new_n10592__, new_new_n10593__,
    new_new_n10594__, new_new_n10595__, new_new_n10596__, new_new_n10597__,
    new_new_n10598__, new_new_n10599__, new_new_n10600__, new_new_n10601__,
    new_new_n10602__, new_new_n10603__, new_new_n10604__, new_new_n10605__,
    new_new_n10606__, new_new_n10607__, new_new_n10608__, new_new_n10609__,
    new_new_n10610__, new_new_n10611__, new_new_n10612__, new_new_n10613__,
    new_new_n10614__, new_new_n10615__, new_new_n10616__, new_new_n10617__,
    new_new_n10618__, new_new_n10619__, new_new_n10620__, new_new_n10621__,
    new_new_n10622__, new_new_n10623__, new_new_n10624__, new_new_n10625__,
    new_new_n10626__, new_new_n10627__, new_new_n10628__, new_new_n10629__,
    new_new_n10630__, new_new_n10631__, new_new_n10632__, new_new_n10633__,
    new_new_n10634__, new_new_n10635__, new_new_n10636__, new_new_n10637__,
    new_new_n10638__, new_new_n10639__, new_new_n10640__, new_new_n10641__,
    new_new_n10642__, new_new_n10643__, new_new_n10644__, new_new_n10645__,
    new_new_n10646__, new_new_n10647__, new_new_n10648__, new_new_n10649__,
    new_new_n10650__, new_new_n10651__, new_new_n10652__, new_new_n10653__,
    new_new_n10654__, new_new_n10655__, new_new_n10656__, new_new_n10657__,
    new_new_n10658__, new_new_n10659__, new_new_n10660__, new_new_n10661__,
    new_new_n10662__, new_new_n10663__, new_new_n10664__, new_new_n10665__,
    new_new_n10666__, new_new_n10667__, new_new_n10668__, new_new_n10669__,
    new_new_n10670__, new_new_n10671__, new_new_n10672__, new_new_n10673__,
    new_new_n10674__, new_new_n10675__, new_new_n10676__, new_new_n10677__,
    new_new_n10678__, new_new_n10679__, new_new_n10680__, new_new_n10681__,
    new_new_n10682__, new_new_n10683__, new_new_n10684__, new_new_n10685__,
    new_new_n10686__, new_new_n10687__, new_new_n10688__, new_new_n10689__,
    new_new_n10690__, new_new_n10691__, new_new_n10692__, new_new_n10693__,
    new_new_n10694__, new_new_n10695__, new_new_n10696__, new_new_n10697__,
    new_new_n10698__, new_new_n10699__, new_new_n10700__, new_new_n10701__,
    new_new_n10702__, new_new_n10703__, new_new_n10704__, new_new_n10705__,
    new_new_n10706__, new_new_n10707__, new_new_n10708__, new_new_n10709__,
    new_new_n10710__, new_new_n10711__, new_new_n10712__, new_new_n10713__,
    new_new_n10714__, new_new_n10715__, new_new_n10716__, new_new_n10717__,
    new_new_n10718__, new_new_n10719__, new_new_n10720__, new_new_n10721__,
    new_new_n10722__, new_new_n10723__, new_new_n10724__, new_new_n10725__,
    new_new_n10726__, new_new_n10727__, new_new_n10728__, new_new_n10729__,
    new_new_n10730__, new_new_n10731__, new_new_n10732__, new_new_n10733__,
    new_new_n10734__, new_new_n10735__, new_new_n10736__, new_new_n10737__,
    new_new_n10738__, new_new_n10739__, new_new_n10740__, new_new_n10741__,
    new_new_n10742__, new_new_n10743__, new_new_n10744__, new_new_n10745__,
    new_new_n10746__, new_new_n10747__, new_new_n10748__, new_new_n10750__,
    new_new_n10751__, new_new_n10752__, new_new_n10753__, new_new_n10754__,
    new_new_n10755__, new_new_n10756__, new_new_n10757__, new_new_n10758__,
    new_new_n10759__, new_new_n10760__, new_new_n10761__, new_new_n10762__,
    new_new_n10763__, new_new_n10764__, new_new_n10765__, new_new_n10766__,
    new_new_n10767__, new_new_n10768__, new_new_n10769__, new_new_n10770__,
    new_new_n10771__, new_new_n10772__, new_new_n10773__, new_new_n10774__,
    new_new_n10775__, new_new_n10776__, new_new_n10777__, new_new_n10778__,
    new_new_n10779__, new_new_n10780__, new_new_n10781__, new_new_n10782__,
    new_new_n10783__, new_new_n10784__, new_new_n10785__, new_new_n10786__,
    new_new_n10787__, new_new_n10788__, new_new_n10789__, new_new_n10790__,
    new_new_n10791__, new_new_n10792__, new_new_n10793__, new_new_n10794__,
    new_new_n10795__, new_new_n10796__, new_new_n10797__, new_new_n10798__,
    new_new_n10799__, new_new_n10800__, new_new_n10801__, new_new_n10802__,
    new_new_n10803__, new_new_n10804__, new_new_n10805__, new_new_n10806__,
    new_new_n10807__, new_new_n10808__, new_new_n10809__, new_new_n10810__,
    new_new_n10811__, new_new_n10812__, new_new_n10813__, new_new_n10814__,
    new_new_n10815__, new_new_n10816__, new_new_n10817__, new_new_n10818__,
    new_new_n10819__, new_new_n10820__, new_new_n10821__, new_new_n10822__,
    new_new_n10823__, new_new_n10824__, new_new_n10825__, new_new_n10826__,
    new_new_n10827__, new_new_n10828__, new_new_n10829__, new_new_n10830__,
    new_new_n10831__, new_new_n10832__, new_new_n10833__, new_new_n10834__,
    new_new_n10835__, new_new_n10836__, new_new_n10837__, new_new_n10838__,
    new_new_n10839__, new_new_n10840__, new_new_n10841__, new_new_n10842__,
    new_new_n10843__, new_new_n10844__, new_new_n10845__, new_new_n10846__,
    new_new_n10847__, new_new_n10848__, new_new_n10849__, new_new_n10850__,
    new_new_n10851__, new_new_n10852__, new_new_n10853__, new_new_n10854__,
    new_new_n10855__, new_new_n10856__, new_new_n10857__, new_new_n10858__,
    new_new_n10859__, new_new_n10860__, new_new_n10861__, new_new_n10862__,
    new_new_n10863__, new_new_n10864__, new_new_n10865__, new_new_n10866__,
    new_new_n10867__, new_new_n10868__, new_new_n10869__, new_new_n10870__,
    new_new_n10871__, new_new_n10872__, new_new_n10873__, new_new_n10874__,
    new_new_n10875__, new_new_n10876__, new_new_n10877__, new_new_n10878__,
    new_new_n10879__, new_new_n10880__, new_new_n10881__, new_new_n10882__,
    new_new_n10883__, new_new_n10884__, new_new_n10885__, new_new_n10886__,
    new_new_n10887__, new_new_n10888__, new_new_n10889__, new_new_n10890__,
    new_new_n10891__, new_new_n10892__, new_new_n10893__, new_new_n10894__,
    new_new_n10895__, new_new_n10896__, new_new_n10897__, new_new_n10898__,
    new_new_n10899__, new_new_n10900__, new_new_n10901__, new_new_n10902__,
    new_new_n10903__, new_new_n10904__, new_new_n10905__, new_new_n10906__,
    new_new_n10907__, new_new_n10908__, new_new_n10909__, new_new_n10910__,
    new_new_n10911__, new_new_n10912__, new_new_n10913__, new_new_n10914__,
    new_new_n10915__, new_new_n10916__, new_new_n10917__, new_new_n10918__,
    new_new_n10919__, new_new_n10920__, new_new_n10921__, new_new_n10922__,
    new_new_n10923__, new_new_n10924__, new_new_n10925__, new_new_n10926__,
    new_new_n10927__, new_new_n10928__, new_new_n10929__, new_new_n10930__,
    new_new_n10931__, new_new_n10932__, new_new_n10933__, new_new_n10934__,
    new_new_n10935__, new_new_n10936__, new_new_n10937__, new_new_n10938__,
    new_new_n10939__, new_new_n10940__, new_new_n10941__, new_new_n10942__,
    new_new_n10943__, new_new_n10944__, new_new_n10945__, new_new_n10946__,
    new_new_n10947__, new_new_n10948__, new_new_n10949__, new_new_n10950__,
    new_new_n10951__, new_new_n10952__, new_new_n10953__, new_new_n10954__,
    new_new_n10955__, new_new_n10956__, new_new_n10957__, new_new_n10958__,
    new_new_n10959__, new_new_n10960__, new_new_n10961__, new_new_n10962__,
    new_new_n10963__, new_new_n10964__, new_new_n10965__, new_new_n10966__,
    new_new_n10967__, new_new_n10968__, new_new_n10969__, new_new_n10970__,
    new_new_n10971__, new_new_n10972__, new_new_n10973__, new_new_n10974__,
    new_new_n10975__, new_new_n10976__, new_new_n10977__, new_new_n10978__,
    new_new_n10979__, new_new_n10980__, new_new_n10981__, new_new_n10982__,
    new_new_n10983__, new_new_n10984__, new_new_n10985__, new_new_n10986__,
    new_new_n10987__, new_new_n10988__, new_new_n10989__, new_new_n10990__,
    new_new_n10991__, new_new_n10992__, new_new_n10993__, new_new_n10994__,
    new_new_n10995__, new_new_n10996__, new_new_n10997__, new_new_n10998__,
    new_new_n10999__, new_new_n11000__, new_new_n11001__, new_new_n11002__,
    new_new_n11003__, new_new_n11004__, new_new_n11005__, new_new_n11006__,
    new_new_n11007__, new_new_n11008__, new_new_n11009__, new_new_n11010__,
    new_new_n11011__, new_new_n11012__, new_new_n11013__, new_new_n11014__,
    new_new_n11015__, new_new_n11016__, new_new_n11017__, new_new_n11018__,
    new_new_n11019__, new_new_n11020__, new_new_n11021__, new_new_n11022__,
    new_new_n11023__, new_new_n11024__, new_new_n11025__, new_new_n11026__,
    new_new_n11027__, new_new_n11028__, new_new_n11029__, new_new_n11030__,
    new_new_n11031__, new_new_n11032__, new_new_n11033__, new_new_n11034__,
    new_new_n11035__, new_new_n11036__, new_new_n11037__, new_new_n11038__,
    new_new_n11039__, new_new_n11040__, new_new_n11041__, new_new_n11042__,
    new_new_n11043__, new_new_n11044__, new_new_n11045__, new_new_n11046__,
    new_new_n11047__, new_new_n11048__, new_new_n11049__, new_new_n11050__,
    new_new_n11052__, new_new_n11053__, new_new_n11054__, new_new_n11055__,
    new_new_n11056__, new_new_n11057__, new_new_n11058__, new_new_n11059__,
    new_new_n11060__, new_new_n11061__, new_new_n11062__, new_new_n11063__,
    new_new_n11064__, new_new_n11065__, new_new_n11066__, new_new_n11067__,
    new_new_n11068__, new_new_n11069__, new_new_n11070__, new_new_n11071__,
    new_new_n11072__, new_new_n11073__, new_new_n11074__, new_new_n11075__,
    new_new_n11076__, new_new_n11077__, new_new_n11078__, new_new_n11079__,
    new_new_n11080__, new_new_n11081__, new_new_n11082__, new_new_n11083__,
    new_new_n11084__, new_new_n11085__, new_new_n11086__, new_new_n11087__,
    new_new_n11088__, new_new_n11089__, new_new_n11090__, new_new_n11091__,
    new_new_n11092__, new_new_n11093__, new_new_n11094__, new_new_n11095__,
    new_new_n11096__, new_new_n11097__, new_new_n11098__, new_new_n11099__,
    new_new_n11100__, new_new_n11101__, new_new_n11102__, new_new_n11103__,
    new_new_n11104__, new_new_n11105__, new_new_n11106__, new_new_n11107__,
    new_new_n11108__, new_new_n11109__, new_new_n11110__, new_new_n11111__,
    new_new_n11112__, new_new_n11113__, new_new_n11114__, new_new_n11115__,
    new_new_n11116__, new_new_n11117__, new_new_n11118__, new_new_n11119__,
    new_new_n11120__, new_new_n11121__, new_new_n11122__, new_new_n11123__,
    new_new_n11124__, new_new_n11125__, new_new_n11126__, new_new_n11127__,
    new_new_n11128__, new_new_n11129__, new_new_n11130__, new_new_n11131__,
    new_new_n11132__, new_new_n11133__, new_new_n11134__, new_new_n11135__,
    new_new_n11136__, new_new_n11137__, new_new_n11138__, new_new_n11139__,
    new_new_n11140__, new_new_n11141__, new_new_n11142__, new_new_n11143__,
    new_new_n11144__, new_new_n11145__, new_new_n11146__, new_new_n11147__,
    new_new_n11148__, new_new_n11149__, new_new_n11150__, new_new_n11151__,
    new_new_n11152__, new_new_n11153__, new_new_n11154__, new_new_n11155__,
    new_new_n11156__, new_new_n11157__, new_new_n11158__, new_new_n11159__,
    new_new_n11160__, new_new_n11161__, new_new_n11162__, new_new_n11163__,
    new_new_n11164__, new_new_n11165__, new_new_n11166__, new_new_n11167__,
    new_new_n11168__, new_new_n11169__, new_new_n11170__, new_new_n11171__,
    new_new_n11172__, new_new_n11173__, new_new_n11174__, new_new_n11175__,
    new_new_n11176__, new_new_n11177__, new_new_n11178__, new_new_n11179__,
    new_new_n11180__, new_new_n11181__, new_new_n11182__, new_new_n11183__,
    new_new_n11184__, new_new_n11185__, new_new_n11186__, new_new_n11187__,
    new_new_n11188__, new_new_n11189__, new_new_n11190__, new_new_n11191__,
    new_new_n11192__, new_new_n11193__, new_new_n11194__, new_new_n11195__,
    new_new_n11196__, new_new_n11197__, new_new_n11198__, new_new_n11199__,
    new_new_n11200__, new_new_n11201__, new_new_n11202__, new_new_n11203__,
    new_new_n11204__, new_new_n11205__, new_new_n11206__, new_new_n11207__,
    new_new_n11208__, new_new_n11209__, new_new_n11210__, new_new_n11211__,
    new_new_n11212__, new_new_n11213__, new_new_n11214__, new_new_n11215__,
    new_new_n11216__, new_new_n11217__, new_new_n11218__, new_new_n11219__,
    new_new_n11220__, new_new_n11221__, new_new_n11222__, new_new_n11223__,
    new_new_n11224__, new_new_n11225__, new_new_n11226__, new_new_n11227__,
    new_new_n11228__, new_new_n11229__, new_new_n11230__, new_new_n11231__,
    new_new_n11232__, new_new_n11233__, new_new_n11234__, new_new_n11235__,
    new_new_n11236__, new_new_n11237__, new_new_n11238__, new_new_n11239__,
    new_new_n11240__, new_new_n11241__, new_new_n11242__, new_new_n11243__,
    new_new_n11244__, new_new_n11245__, new_new_n11246__, new_new_n11247__,
    new_new_n11248__, new_new_n11249__, new_new_n11250__, new_new_n11251__,
    new_new_n11252__, new_new_n11253__, new_new_n11254__, new_new_n11255__,
    new_new_n11256__, new_new_n11257__, new_new_n11258__, new_new_n11259__,
    new_new_n11260__, new_new_n11261__, new_new_n11262__, new_new_n11263__,
    new_new_n11264__, new_new_n11265__, new_new_n11266__, new_new_n11267__,
    new_new_n11268__, new_new_n11269__, new_new_n11270__, new_new_n11271__,
    new_new_n11272__, new_new_n11273__, new_new_n11274__, new_new_n11275__,
    new_new_n11276__, new_new_n11277__, new_new_n11278__, new_new_n11279__,
    new_new_n11280__, new_new_n11281__, new_new_n11282__, new_new_n11283__,
    new_new_n11284__, new_new_n11285__, new_new_n11286__, new_new_n11287__,
    new_new_n11288__, new_new_n11289__, new_new_n11290__, new_new_n11291__,
    new_new_n11292__, new_new_n11293__, new_new_n11294__, new_new_n11295__,
    new_new_n11296__, new_new_n11297__, new_new_n11298__, new_new_n11299__,
    new_new_n11300__, new_new_n11301__, new_new_n11302__, new_new_n11303__,
    new_new_n11304__, new_new_n11305__, new_new_n11306__, new_new_n11307__,
    new_new_n11308__, new_new_n11309__, new_new_n11310__, new_new_n11311__,
    new_new_n11312__, new_new_n11313__, new_new_n11314__, new_new_n11315__,
    new_new_n11316__, new_new_n11317__, new_new_n11318__, new_new_n11319__,
    new_new_n11320__, new_new_n11321__, new_new_n11322__, new_new_n11324__,
    new_new_n11325__, new_new_n11326__, new_new_n11327__, new_new_n11328__,
    new_new_n11329__, new_new_n11330__, new_new_n11331__, new_new_n11332__,
    new_new_n11333__, new_new_n11334__, new_new_n11335__, new_new_n11336__,
    new_new_n11337__, new_new_n11338__, new_new_n11339__, new_new_n11340__,
    new_new_n11341__, new_new_n11342__, new_new_n11343__, new_new_n11344__,
    new_new_n11345__, new_new_n11346__, new_new_n11347__, new_new_n11348__,
    new_new_n11349__, new_new_n11350__, new_new_n11351__, new_new_n11352__,
    new_new_n11353__, new_new_n11354__, new_new_n11355__, new_new_n11356__,
    new_new_n11357__, new_new_n11358__, new_new_n11359__, new_new_n11360__,
    new_new_n11361__, new_new_n11362__, new_new_n11363__, new_new_n11364__,
    new_new_n11365__, new_new_n11366__, new_new_n11367__, new_new_n11368__,
    new_new_n11369__, new_new_n11370__, new_new_n11371__, new_new_n11372__,
    new_new_n11373__, new_new_n11374__, new_new_n11375__, new_new_n11376__,
    new_new_n11377__, new_new_n11378__, new_new_n11379__, new_new_n11380__,
    new_new_n11381__, new_new_n11382__, new_new_n11383__, new_new_n11384__,
    new_new_n11385__, new_new_n11386__, new_new_n11387__, new_new_n11388__,
    new_new_n11389__, new_new_n11390__, new_new_n11391__, new_new_n11392__,
    new_new_n11393__, new_new_n11394__, new_new_n11395__, new_new_n11396__,
    new_new_n11397__, new_new_n11398__, new_new_n11399__, new_new_n11400__,
    new_new_n11401__, new_new_n11402__, new_new_n11403__, new_new_n11404__,
    new_new_n11405__, new_new_n11406__, new_new_n11407__, new_new_n11408__,
    new_new_n11409__, new_new_n11410__, new_new_n11411__, new_new_n11412__,
    new_new_n11413__, new_new_n11414__, new_new_n11415__, new_new_n11416__,
    new_new_n11417__, new_new_n11418__, new_new_n11419__, new_new_n11420__,
    new_new_n11421__, new_new_n11422__, new_new_n11423__, new_new_n11424__,
    new_new_n11425__, new_new_n11426__, new_new_n11427__, new_new_n11428__,
    new_new_n11429__, new_new_n11430__, new_new_n11431__, new_new_n11432__,
    new_new_n11433__, new_new_n11434__, new_new_n11435__, new_new_n11436__,
    new_new_n11437__, new_new_n11438__, new_new_n11439__, new_new_n11440__,
    new_new_n11441__, new_new_n11442__, new_new_n11443__, new_new_n11444__,
    new_new_n11445__, new_new_n11446__, new_new_n11447__, new_new_n11448__,
    new_new_n11449__, new_new_n11450__, new_new_n11451__, new_new_n11452__,
    new_new_n11453__, new_new_n11454__, new_new_n11455__, new_new_n11456__,
    new_new_n11457__, new_new_n11458__, new_new_n11459__, new_new_n11460__,
    new_new_n11461__, new_new_n11462__, new_new_n11463__, new_new_n11464__,
    new_new_n11465__, new_new_n11466__, new_new_n11467__, new_new_n11468__,
    new_new_n11469__, new_new_n11470__, new_new_n11471__, new_new_n11472__,
    new_new_n11473__, new_new_n11474__, new_new_n11475__, new_new_n11476__,
    new_new_n11477__, new_new_n11478__, new_new_n11479__, new_new_n11480__,
    new_new_n11481__, new_new_n11482__, new_new_n11483__, new_new_n11484__,
    new_new_n11485__, new_new_n11486__, new_new_n11487__, new_new_n11488__,
    new_new_n11489__, new_new_n11490__, new_new_n11491__, new_new_n11492__,
    new_new_n11493__, new_new_n11494__, new_new_n11495__, new_new_n11496__,
    new_new_n11497__, new_new_n11498__, new_new_n11499__, new_new_n11500__,
    new_new_n11501__, new_new_n11502__, new_new_n11503__, new_new_n11504__,
    new_new_n11505__, new_new_n11506__, new_new_n11507__, new_new_n11508__,
    new_new_n11509__, new_new_n11510__, new_new_n11511__, new_new_n11512__,
    new_new_n11513__, new_new_n11514__, new_new_n11515__, new_new_n11516__,
    new_new_n11517__, new_new_n11518__, new_new_n11519__, new_new_n11520__,
    new_new_n11521__, new_new_n11522__, new_new_n11523__, new_new_n11524__,
    new_new_n11525__, new_new_n11526__, new_new_n11527__, new_new_n11528__,
    new_new_n11529__, new_new_n11530__, new_new_n11531__, new_new_n11532__,
    new_new_n11533__, new_new_n11534__, new_new_n11535__, new_new_n11536__,
    new_new_n11537__, new_new_n11538__, new_new_n11539__, new_new_n11540__,
    new_new_n11541__, new_new_n11542__, new_new_n11543__, new_new_n11544__,
    new_new_n11545__, new_new_n11546__, new_new_n11547__, new_new_n11548__,
    new_new_n11549__, new_new_n11550__, new_new_n11551__, new_new_n11552__,
    new_new_n11553__, new_new_n11554__, new_new_n11555__, new_new_n11556__,
    new_new_n11557__, new_new_n11558__, new_new_n11559__, new_new_n11560__,
    new_new_n11561__, new_new_n11562__, new_new_n11563__, new_new_n11564__,
    new_new_n11565__, new_new_n11566__, new_new_n11567__, new_new_n11568__,
    new_new_n11569__, new_new_n11570__, new_new_n11571__, new_new_n11572__,
    new_new_n11573__, new_new_n11574__, new_new_n11575__, new_new_n11576__,
    new_new_n11577__, new_new_n11578__, new_new_n11579__, new_new_n11580__,
    new_new_n11581__, new_new_n11582__, new_new_n11583__, new_new_n11584__,
    new_new_n11585__, new_new_n11586__, new_new_n11587__, new_new_n11588__,
    new_new_n11589__, new_new_n11590__, new_new_n11591__, new_new_n11592__,
    new_new_n11593__, new_new_n11595__, new_new_n11596__, new_new_n11597__,
    new_new_n11598__, new_new_n11599__, new_new_n11600__, new_new_n11601__,
    new_new_n11602__, new_new_n11603__, new_new_n11604__, new_new_n11605__,
    new_new_n11606__, new_new_n11607__, new_new_n11608__, new_new_n11609__,
    new_new_n11610__, new_new_n11611__, new_new_n11612__, new_new_n11613__,
    new_new_n11614__, new_new_n11615__, new_new_n11616__, new_new_n11617__,
    new_new_n11618__, new_new_n11619__, new_new_n11620__, new_new_n11621__,
    new_new_n11622__, new_new_n11623__, new_new_n11624__, new_new_n11625__,
    new_new_n11626__, new_new_n11627__, new_new_n11628__, new_new_n11629__,
    new_new_n11630__, new_new_n11631__, new_new_n11632__, new_new_n11633__,
    new_new_n11634__, new_new_n11635__, new_new_n11636__, new_new_n11637__,
    new_new_n11638__, new_new_n11639__, new_new_n11640__, new_new_n11641__,
    new_new_n11642__, new_new_n11643__, new_new_n11644__, new_new_n11645__,
    new_new_n11646__, new_new_n11647__, new_new_n11648__, new_new_n11649__,
    new_new_n11650__, new_new_n11651__, new_new_n11652__, new_new_n11653__,
    new_new_n11654__, new_new_n11655__, new_new_n11656__, new_new_n11657__,
    new_new_n11658__, new_new_n11659__, new_new_n11660__, new_new_n11661__,
    new_new_n11662__, new_new_n11663__, new_new_n11664__, new_new_n11665__,
    new_new_n11666__, new_new_n11667__, new_new_n11668__, new_new_n11669__,
    new_new_n11670__, new_new_n11671__, new_new_n11672__, new_new_n11673__,
    new_new_n11674__, new_new_n11675__, new_new_n11676__, new_new_n11677__,
    new_new_n11678__, new_new_n11679__, new_new_n11680__, new_new_n11681__,
    new_new_n11682__, new_new_n11683__, new_new_n11684__, new_new_n11685__,
    new_new_n11686__, new_new_n11687__, new_new_n11688__, new_new_n11689__,
    new_new_n11690__, new_new_n11691__, new_new_n11692__, new_new_n11693__,
    new_new_n11694__, new_new_n11695__, new_new_n11696__, new_new_n11697__,
    new_new_n11698__, new_new_n11699__, new_new_n11700__, new_new_n11701__,
    new_new_n11702__, new_new_n11703__, new_new_n11704__, new_new_n11705__,
    new_new_n11706__, new_new_n11707__, new_new_n11708__, new_new_n11709__,
    new_new_n11710__, new_new_n11711__, new_new_n11712__, new_new_n11713__,
    new_new_n11714__, new_new_n11715__, new_new_n11716__, new_new_n11717__,
    new_new_n11718__, new_new_n11719__, new_new_n11720__, new_new_n11721__,
    new_new_n11722__, new_new_n11723__, new_new_n11724__, new_new_n11725__,
    new_new_n11726__, new_new_n11727__, new_new_n11728__, new_new_n11729__,
    new_new_n11730__, new_new_n11731__, new_new_n11732__, new_new_n11733__,
    new_new_n11734__, new_new_n11735__, new_new_n11736__, new_new_n11737__,
    new_new_n11738__, new_new_n11739__, new_new_n11740__, new_new_n11741__,
    new_new_n11742__, new_new_n11743__, new_new_n11744__, new_new_n11745__,
    new_new_n11746__, new_new_n11747__, new_new_n11748__, new_new_n11749__,
    new_new_n11750__, new_new_n11751__, new_new_n11752__, new_new_n11753__,
    new_new_n11754__, new_new_n11755__, new_new_n11756__, new_new_n11757__,
    new_new_n11758__, new_new_n11759__, new_new_n11760__, new_new_n11761__,
    new_new_n11762__, new_new_n11763__, new_new_n11764__, new_new_n11765__,
    new_new_n11766__, new_new_n11767__, new_new_n11768__, new_new_n11769__,
    new_new_n11770__, new_new_n11771__, new_new_n11772__, new_new_n11773__,
    new_new_n11774__, new_new_n11775__, new_new_n11776__, new_new_n11777__,
    new_new_n11778__, new_new_n11779__, new_new_n11780__, new_new_n11781__,
    new_new_n11782__, new_new_n11783__, new_new_n11784__, new_new_n11785__,
    new_new_n11786__, new_new_n11787__, new_new_n11788__, new_new_n11789__,
    new_new_n11790__, new_new_n11791__, new_new_n11792__, new_new_n11793__,
    new_new_n11794__, new_new_n11795__, new_new_n11796__, new_new_n11797__,
    new_new_n11798__, new_new_n11799__, new_new_n11800__, new_new_n11801__,
    new_new_n11802__, new_new_n11803__, new_new_n11804__, new_new_n11805__,
    new_new_n11806__, new_new_n11807__, new_new_n11808__, new_new_n11809__,
    new_new_n11810__, new_new_n11811__, new_new_n11812__, new_new_n11813__,
    new_new_n11814__, new_new_n11815__, new_new_n11816__, new_new_n11817__,
    new_new_n11818__, new_new_n11819__, new_new_n11820__, new_new_n11821__,
    new_new_n11822__, new_new_n11823__, new_new_n11824__, new_new_n11825__,
    new_new_n11826__, new_new_n11827__, new_new_n11828__, new_new_n11829__,
    new_new_n11830__, new_new_n11831__, new_new_n11832__, new_new_n11833__,
    new_new_n11834__, new_new_n11835__, new_new_n11836__, new_new_n11837__,
    new_new_n11838__, new_new_n11839__, new_new_n11840__, new_new_n11841__,
    new_new_n11842__, new_new_n11843__, new_new_n11844__, new_new_n11845__,
    new_new_n11846__, new_new_n11847__, new_new_n11848__, new_new_n11849__,
    new_new_n11850__, new_new_n11851__, new_new_n11852__, new_new_n11853__,
    new_new_n11854__, new_new_n11855__, new_new_n11856__, new_new_n11857__,
    new_new_n11858__, new_new_n11859__, new_new_n11860__, new_new_n11861__,
    new_new_n11862__, new_new_n11863__, new_new_n11864__, new_new_n11865__,
    new_new_n11866__, new_new_n11867__, new_new_n11868__, new_new_n11869__,
    new_new_n11870__, new_new_n11871__, new_new_n11872__, new_new_n11873__,
    new_new_n11874__, new_new_n11875__, new_new_n11876__, new_new_n11878__,
    new_new_n11879__, new_new_n11880__, new_new_n11881__, new_new_n11882__,
    new_new_n11883__, new_new_n11884__, new_new_n11885__, new_new_n11886__,
    new_new_n11887__, new_new_n11888__, new_new_n11889__, new_new_n11890__,
    new_new_n11891__, new_new_n11892__, new_new_n11893__, new_new_n11894__,
    new_new_n11895__, new_new_n11896__, new_new_n11897__, new_new_n11898__,
    new_new_n11899__, new_new_n11900__, new_new_n11901__, new_new_n11902__,
    new_new_n11903__, new_new_n11904__, new_new_n11905__, new_new_n11906__,
    new_new_n11907__, new_new_n11908__, new_new_n11909__, new_new_n11910__,
    new_new_n11911__, new_new_n11912__, new_new_n11913__, new_new_n11914__,
    new_new_n11915__, new_new_n11916__, new_new_n11917__, new_new_n11918__,
    new_new_n11919__, new_new_n11920__, new_new_n11921__, new_new_n11922__,
    new_new_n11923__, new_new_n11924__, new_new_n11925__, new_new_n11926__,
    new_new_n11927__, new_new_n11928__, new_new_n11929__, new_new_n11930__,
    new_new_n11931__, new_new_n11932__, new_new_n11933__, new_new_n11934__,
    new_new_n11935__, new_new_n11936__, new_new_n11937__, new_new_n11938__,
    new_new_n11939__, new_new_n11940__, new_new_n11941__, new_new_n11942__,
    new_new_n11943__, new_new_n11944__, new_new_n11945__, new_new_n11946__,
    new_new_n11947__, new_new_n11948__, new_new_n11949__, new_new_n11950__,
    new_new_n11951__, new_new_n11952__, new_new_n11953__, new_new_n11954__,
    new_new_n11955__, new_new_n11956__, new_new_n11957__, new_new_n11958__,
    new_new_n11959__, new_new_n11960__, new_new_n11961__, new_new_n11962__,
    new_new_n11963__, new_new_n11964__, new_new_n11965__, new_new_n11966__,
    new_new_n11967__, new_new_n11968__, new_new_n11969__, new_new_n11970__,
    new_new_n11971__, new_new_n11972__, new_new_n11973__, new_new_n11974__,
    new_new_n11975__, new_new_n11976__, new_new_n11977__, new_new_n11978__,
    new_new_n11979__, new_new_n11980__, new_new_n11981__, new_new_n11982__,
    new_new_n11983__, new_new_n11984__, new_new_n11985__, new_new_n11986__,
    new_new_n11987__, new_new_n11988__, new_new_n11989__, new_new_n11990__,
    new_new_n11991__, new_new_n11992__, new_new_n11993__, new_new_n11994__,
    new_new_n11995__, new_new_n11996__, new_new_n11997__, new_new_n11998__,
    new_new_n11999__, new_new_n12000__, new_new_n12001__, new_new_n12002__,
    new_new_n12003__, new_new_n12004__, new_new_n12005__, new_new_n12006__,
    new_new_n12007__, new_new_n12008__, new_new_n12009__, new_new_n12010__,
    new_new_n12011__, new_new_n12012__, new_new_n12013__, new_new_n12014__,
    new_new_n12015__, new_new_n12016__, new_new_n12017__, new_new_n12018__,
    new_new_n12019__, new_new_n12020__, new_new_n12021__, new_new_n12022__,
    new_new_n12023__, new_new_n12024__, new_new_n12025__, new_new_n12026__,
    new_new_n12027__, new_new_n12028__, new_new_n12029__, new_new_n12030__,
    new_new_n12031__, new_new_n12032__, new_new_n12033__, new_new_n12034__,
    new_new_n12035__, new_new_n12036__, new_new_n12037__, new_new_n12038__,
    new_new_n12039__, new_new_n12040__, new_new_n12041__, new_new_n12042__,
    new_new_n12043__, new_new_n12044__, new_new_n12045__, new_new_n12046__,
    new_new_n12047__, new_new_n12048__, new_new_n12049__, new_new_n12050__,
    new_new_n12051__, new_new_n12052__, new_new_n12053__, new_new_n12054__,
    new_new_n12055__, new_new_n12056__, new_new_n12057__, new_new_n12058__,
    new_new_n12059__, new_new_n12060__, new_new_n12061__, new_new_n12062__,
    new_new_n12063__, new_new_n12064__, new_new_n12065__, new_new_n12066__,
    new_new_n12067__, new_new_n12068__, new_new_n12069__, new_new_n12070__,
    new_new_n12071__, new_new_n12072__, new_new_n12073__, new_new_n12074__,
    new_new_n12075__, new_new_n12076__, new_new_n12077__, new_new_n12078__,
    new_new_n12079__, new_new_n12080__, new_new_n12081__, new_new_n12082__,
    new_new_n12083__, new_new_n12084__, new_new_n12085__, new_new_n12086__,
    new_new_n12087__, new_new_n12088__, new_new_n12089__, new_new_n12090__,
    new_new_n12091__, new_new_n12092__, new_new_n12093__, new_new_n12094__,
    new_new_n12095__, new_new_n12096__, new_new_n12097__, new_new_n12098__,
    new_new_n12099__, new_new_n12100__, new_new_n12101__, new_new_n12102__,
    new_new_n12103__, new_new_n12104__, new_new_n12105__, new_new_n12106__,
    new_new_n12107__, new_new_n12108__, new_new_n12109__, new_new_n12110__,
    new_new_n12111__, new_new_n12112__, new_new_n12113__, new_new_n12114__,
    new_new_n12115__, new_new_n12116__, new_new_n12117__, new_new_n12118__,
    new_new_n12119__, new_new_n12120__, new_new_n12121__, new_new_n12122__,
    new_new_n12123__, new_new_n12124__, new_new_n12125__, new_new_n12126__,
    new_new_n12127__, new_new_n12128__, new_new_n12129__, new_new_n12130__,
    new_new_n12131__, new_new_n12132__, new_new_n12133__, new_new_n12134__,
    new_new_n12135__, new_new_n12136__, new_new_n12137__, new_new_n12138__,
    new_new_n12139__, new_new_n12140__, new_new_n12141__, new_new_n12142__,
    new_new_n12143__, new_new_n12144__, new_new_n12145__, new_new_n12146__,
    new_new_n12147__, new_new_n12148__, new_new_n12149__, new_new_n12150__,
    new_new_n12152__, new_new_n12153__, new_new_n12154__, new_new_n12155__,
    new_new_n12156__, new_new_n12157__, new_new_n12158__, new_new_n12159__,
    new_new_n12160__, new_new_n12161__, new_new_n12162__, new_new_n12163__,
    new_new_n12164__, new_new_n12165__, new_new_n12166__, new_new_n12167__,
    new_new_n12168__, new_new_n12169__, new_new_n12170__, new_new_n12171__,
    new_new_n12172__, new_new_n12173__, new_new_n12174__, new_new_n12175__,
    new_new_n12176__, new_new_n12177__, new_new_n12178__, new_new_n12179__,
    new_new_n12180__, new_new_n12181__, new_new_n12182__, new_new_n12183__,
    new_new_n12184__, new_new_n12185__, new_new_n12186__, new_new_n12187__,
    new_new_n12188__, new_new_n12189__, new_new_n12190__, new_new_n12191__,
    new_new_n12192__, new_new_n12193__, new_new_n12194__, new_new_n12195__,
    new_new_n12196__, new_new_n12197__, new_new_n12198__, new_new_n12199__,
    new_new_n12200__, new_new_n12201__, new_new_n12202__, new_new_n12203__,
    new_new_n12204__, new_new_n12205__, new_new_n12206__, new_new_n12207__,
    new_new_n12208__, new_new_n12209__, new_new_n12210__, new_new_n12211__,
    new_new_n12212__, new_new_n12213__, new_new_n12214__, new_new_n12215__,
    new_new_n12216__, new_new_n12217__, new_new_n12218__, new_new_n12219__,
    new_new_n12220__, new_new_n12221__, new_new_n12222__, new_new_n12223__,
    new_new_n12224__, new_new_n12225__, new_new_n12226__, new_new_n12227__,
    new_new_n12228__, new_new_n12229__, new_new_n12230__, new_new_n12231__,
    new_new_n12232__, new_new_n12233__, new_new_n12234__, new_new_n12235__,
    new_new_n12236__, new_new_n12237__, new_new_n12238__, new_new_n12239__,
    new_new_n12240__, new_new_n12241__, new_new_n12242__, new_new_n12243__,
    new_new_n12244__, new_new_n12245__, new_new_n12246__, new_new_n12247__,
    new_new_n12248__, new_new_n12249__, new_new_n12250__, new_new_n12251__,
    new_new_n12252__, new_new_n12253__, new_new_n12254__, new_new_n12255__,
    new_new_n12256__, new_new_n12257__, new_new_n12258__, new_new_n12259__,
    new_new_n12260__, new_new_n12261__, new_new_n12262__, new_new_n12263__,
    new_new_n12264__, new_new_n12265__, new_new_n12266__, new_new_n12267__,
    new_new_n12268__, new_new_n12269__, new_new_n12270__, new_new_n12271__,
    new_new_n12272__, new_new_n12273__, new_new_n12274__, new_new_n12275__,
    new_new_n12276__, new_new_n12277__, new_new_n12278__, new_new_n12279__,
    new_new_n12280__, new_new_n12281__, new_new_n12282__, new_new_n12283__,
    new_new_n12284__, new_new_n12285__, new_new_n12286__, new_new_n12287__,
    new_new_n12288__, new_new_n12289__, new_new_n12290__, new_new_n12291__,
    new_new_n12292__, new_new_n12293__, new_new_n12294__, new_new_n12295__,
    new_new_n12296__, new_new_n12297__, new_new_n12298__, new_new_n12299__,
    new_new_n12300__, new_new_n12301__, new_new_n12302__, new_new_n12303__,
    new_new_n12304__, new_new_n12305__, new_new_n12306__, new_new_n12307__,
    new_new_n12308__, new_new_n12309__, new_new_n12310__, new_new_n12311__,
    new_new_n12312__, new_new_n12313__, new_new_n12314__, new_new_n12315__,
    new_new_n12316__, new_new_n12317__, new_new_n12318__, new_new_n12319__,
    new_new_n12320__, new_new_n12321__, new_new_n12322__, new_new_n12323__,
    new_new_n12324__, new_new_n12325__, new_new_n12326__, new_new_n12327__,
    new_new_n12328__, new_new_n12329__, new_new_n12330__, new_new_n12331__,
    new_new_n12332__, new_new_n12333__, new_new_n12334__, new_new_n12335__,
    new_new_n12336__, new_new_n12337__, new_new_n12338__, new_new_n12339__,
    new_new_n12340__, new_new_n12341__, new_new_n12342__, new_new_n12343__,
    new_new_n12344__, new_new_n12345__, new_new_n12346__, new_new_n12347__,
    new_new_n12348__, new_new_n12349__, new_new_n12350__, new_new_n12351__,
    new_new_n12352__, new_new_n12353__, new_new_n12354__, new_new_n12355__,
    new_new_n12356__, new_new_n12357__, new_new_n12358__, new_new_n12359__,
    new_new_n12360__, new_new_n12361__, new_new_n12362__, new_new_n12363__,
    new_new_n12364__, new_new_n12365__, new_new_n12366__, new_new_n12367__,
    new_new_n12368__, new_new_n12369__, new_new_n12370__, new_new_n12371__,
    new_new_n12372__, new_new_n12373__, new_new_n12374__, new_new_n12375__,
    new_new_n12376__, new_new_n12377__, new_new_n12378__, new_new_n12379__,
    new_new_n12380__, new_new_n12381__, new_new_n12382__, new_new_n12383__,
    new_new_n12384__, new_new_n12385__, new_new_n12386__, new_new_n12387__,
    new_new_n12388__, new_new_n12389__, new_new_n12390__, new_new_n12391__,
    new_new_n12392__, new_new_n12393__, new_new_n12394__, new_new_n12395__,
    new_new_n12396__, new_new_n12397__, new_new_n12398__, new_new_n12399__,
    new_new_n12400__, new_new_n12401__, new_new_n12402__, new_new_n12403__,
    new_new_n12404__, new_new_n12405__, new_new_n12406__, new_new_n12407__,
    new_new_n12409__, new_new_n12410__, new_new_n12411__, new_new_n12412__,
    new_new_n12413__, new_new_n12414__, new_new_n12415__, new_new_n12416__,
    new_new_n12417__, new_new_n12418__, new_new_n12419__, new_new_n12420__,
    new_new_n12421__, new_new_n12422__, new_new_n12423__, new_new_n12424__,
    new_new_n12425__, new_new_n12426__, new_new_n12427__, new_new_n12428__,
    new_new_n12429__, new_new_n12430__, new_new_n12431__, new_new_n12432__,
    new_new_n12433__, new_new_n12434__, new_new_n12435__, new_new_n12436__,
    new_new_n12437__, new_new_n12438__, new_new_n12439__, new_new_n12440__,
    new_new_n12441__, new_new_n12442__, new_new_n12443__, new_new_n12444__,
    new_new_n12445__, new_new_n12446__, new_new_n12447__, new_new_n12448__,
    new_new_n12449__, new_new_n12450__, new_new_n12451__, new_new_n12452__,
    new_new_n12453__, new_new_n12454__, new_new_n12455__, new_new_n12456__,
    new_new_n12457__, new_new_n12458__, new_new_n12459__, new_new_n12460__,
    new_new_n12461__, new_new_n12462__, new_new_n12463__, new_new_n12464__,
    new_new_n12465__, new_new_n12466__, new_new_n12467__, new_new_n12468__,
    new_new_n12469__, new_new_n12470__, new_new_n12471__, new_new_n12472__,
    new_new_n12473__, new_new_n12474__, new_new_n12475__, new_new_n12476__,
    new_new_n12477__, new_new_n12478__, new_new_n12479__, new_new_n12480__,
    new_new_n12481__, new_new_n12482__, new_new_n12483__, new_new_n12484__,
    new_new_n12485__, new_new_n12486__, new_new_n12487__, new_new_n12488__,
    new_new_n12489__, new_new_n12490__, new_new_n12491__, new_new_n12492__,
    new_new_n12493__, new_new_n12494__, new_new_n12495__, new_new_n12496__,
    new_new_n12497__, new_new_n12498__, new_new_n12499__, new_new_n12500__,
    new_new_n12501__, new_new_n12502__, new_new_n12503__, new_new_n12504__,
    new_new_n12505__, new_new_n12506__, new_new_n12507__, new_new_n12508__,
    new_new_n12509__, new_new_n12510__, new_new_n12511__, new_new_n12512__,
    new_new_n12513__, new_new_n12514__, new_new_n12515__, new_new_n12516__,
    new_new_n12517__, new_new_n12518__, new_new_n12519__, new_new_n12520__,
    new_new_n12521__, new_new_n12522__, new_new_n12523__, new_new_n12524__,
    new_new_n12525__, new_new_n12526__, new_new_n12527__, new_new_n12528__,
    new_new_n12529__, new_new_n12530__, new_new_n12531__, new_new_n12532__,
    new_new_n12533__, new_new_n12534__, new_new_n12535__, new_new_n12536__,
    new_new_n12537__, new_new_n12538__, new_new_n12539__, new_new_n12540__,
    new_new_n12541__, new_new_n12542__, new_new_n12543__, new_new_n12544__,
    new_new_n12545__, new_new_n12546__, new_new_n12547__, new_new_n12548__,
    new_new_n12549__, new_new_n12550__, new_new_n12551__, new_new_n12552__,
    new_new_n12553__, new_new_n12554__, new_new_n12555__, new_new_n12556__,
    new_new_n12557__, new_new_n12558__, new_new_n12559__, new_new_n12560__,
    new_new_n12561__, new_new_n12562__, new_new_n12563__, new_new_n12564__,
    new_new_n12565__, new_new_n12566__, new_new_n12567__, new_new_n12568__,
    new_new_n12569__, new_new_n12570__, new_new_n12571__, new_new_n12572__,
    new_new_n12573__, new_new_n12574__, new_new_n12575__, new_new_n12576__,
    new_new_n12577__, new_new_n12578__, new_new_n12579__, new_new_n12580__,
    new_new_n12581__, new_new_n12582__, new_new_n12583__, new_new_n12584__,
    new_new_n12585__, new_new_n12586__, new_new_n12587__, new_new_n12588__,
    new_new_n12589__, new_new_n12590__, new_new_n12591__, new_new_n12592__,
    new_new_n12593__, new_new_n12594__, new_new_n12595__, new_new_n12596__,
    new_new_n12597__, new_new_n12598__, new_new_n12599__, new_new_n12600__,
    new_new_n12601__, new_new_n12602__, new_new_n12603__, new_new_n12604__,
    new_new_n12605__, new_new_n12606__, new_new_n12607__, new_new_n12608__,
    new_new_n12609__, new_new_n12610__, new_new_n12611__, new_new_n12612__,
    new_new_n12613__, new_new_n12614__, new_new_n12615__, new_new_n12616__,
    new_new_n12617__, new_new_n12618__, new_new_n12619__, new_new_n12620__,
    new_new_n12621__, new_new_n12622__, new_new_n12623__, new_new_n12624__,
    new_new_n12625__, new_new_n12626__, new_new_n12627__, new_new_n12628__,
    new_new_n12629__, new_new_n12630__, new_new_n12631__, new_new_n12632__,
    new_new_n12633__, new_new_n12634__, new_new_n12635__, new_new_n12636__,
    new_new_n12637__, new_new_n12638__, new_new_n12639__, new_new_n12640__,
    new_new_n12641__, new_new_n12642__, new_new_n12643__, new_new_n12644__,
    new_new_n12645__, new_new_n12646__, new_new_n12647__, new_new_n12648__,
    new_new_n12649__, new_new_n12650__, new_new_n12651__, new_new_n12652__,
    new_new_n12653__, new_new_n12654__, new_new_n12655__, new_new_n12656__,
    new_new_n12657__, new_new_n12658__, new_new_n12659__, new_new_n12660__,
    new_new_n12661__, new_new_n12662__, new_new_n12663__, new_new_n12664__,
    new_new_n12665__, new_new_n12666__, new_new_n12667__, new_new_n12668__,
    new_new_n12669__, new_new_n12670__, new_new_n12671__, new_new_n12672__,
    new_new_n12673__, new_new_n12674__, new_new_n12675__, new_new_n12676__,
    new_new_n12677__, new_new_n12678__, new_new_n12679__, new_new_n12680__,
    new_new_n12682__, new_new_n12683__, new_new_n12684__, new_new_n12685__,
    new_new_n12686__, new_new_n12687__, new_new_n12688__, new_new_n12689__,
    new_new_n12690__, new_new_n12691__, new_new_n12692__, new_new_n12693__,
    new_new_n12694__, new_new_n12695__, new_new_n12696__, new_new_n12697__,
    new_new_n12698__, new_new_n12699__, new_new_n12700__, new_new_n12701__,
    new_new_n12702__, new_new_n12703__, new_new_n12704__, new_new_n12705__,
    new_new_n12706__, new_new_n12707__, new_new_n12708__, new_new_n12709__,
    new_new_n12710__, new_new_n12711__, new_new_n12712__, new_new_n12713__,
    new_new_n12714__, new_new_n12715__, new_new_n12716__, new_new_n12717__,
    new_new_n12718__, new_new_n12719__, new_new_n12720__, new_new_n12721__,
    new_new_n12722__, new_new_n12723__, new_new_n12724__, new_new_n12725__,
    new_new_n12726__, new_new_n12727__, new_new_n12728__, new_new_n12729__,
    new_new_n12730__, new_new_n12731__, new_new_n12732__, new_new_n12733__,
    new_new_n12734__, new_new_n12735__, new_new_n12736__, new_new_n12737__,
    new_new_n12738__, new_new_n12739__, new_new_n12740__, new_new_n12741__,
    new_new_n12742__, new_new_n12743__, new_new_n12744__, new_new_n12745__,
    new_new_n12746__, new_new_n12747__, new_new_n12748__, new_new_n12749__,
    new_new_n12750__, new_new_n12751__, new_new_n12752__, new_new_n12753__,
    new_new_n12754__, new_new_n12755__, new_new_n12756__, new_new_n12757__,
    new_new_n12758__, new_new_n12759__, new_new_n12760__, new_new_n12761__,
    new_new_n12762__, new_new_n12763__, new_new_n12764__, new_new_n12765__,
    new_new_n12766__, new_new_n12767__, new_new_n12768__, new_new_n12769__,
    new_new_n12770__, new_new_n12771__, new_new_n12772__, new_new_n12773__,
    new_new_n12774__, new_new_n12775__, new_new_n12776__, new_new_n12777__,
    new_new_n12778__, new_new_n12779__, new_new_n12780__, new_new_n12781__,
    new_new_n12782__, new_new_n12783__, new_new_n12784__, new_new_n12785__,
    new_new_n12786__, new_new_n12787__, new_new_n12788__, new_new_n12789__,
    new_new_n12790__, new_new_n12791__, new_new_n12792__, new_new_n12793__,
    new_new_n12794__, new_new_n12795__, new_new_n12796__, new_new_n12797__,
    new_new_n12798__, new_new_n12799__, new_new_n12800__, new_new_n12801__,
    new_new_n12802__, new_new_n12803__, new_new_n12804__, new_new_n12805__,
    new_new_n12806__, new_new_n12807__, new_new_n12808__, new_new_n12809__,
    new_new_n12810__, new_new_n12811__, new_new_n12812__, new_new_n12813__,
    new_new_n12814__, new_new_n12815__, new_new_n12816__, new_new_n12817__,
    new_new_n12818__, new_new_n12819__, new_new_n12820__, new_new_n12821__,
    new_new_n12822__, new_new_n12823__, new_new_n12824__, new_new_n12825__,
    new_new_n12826__, new_new_n12827__, new_new_n12828__, new_new_n12829__,
    new_new_n12830__, new_new_n12831__, new_new_n12832__, new_new_n12833__,
    new_new_n12834__, new_new_n12835__, new_new_n12836__, new_new_n12837__,
    new_new_n12838__, new_new_n12839__, new_new_n12840__, new_new_n12841__,
    new_new_n12842__, new_new_n12843__, new_new_n12844__, new_new_n12845__,
    new_new_n12846__, new_new_n12847__, new_new_n12848__, new_new_n12849__,
    new_new_n12850__, new_new_n12851__, new_new_n12852__, new_new_n12853__,
    new_new_n12854__, new_new_n12855__, new_new_n12856__, new_new_n12857__,
    new_new_n12858__, new_new_n12859__, new_new_n12860__, new_new_n12861__,
    new_new_n12862__, new_new_n12863__, new_new_n12864__, new_new_n12865__,
    new_new_n12866__, new_new_n12867__, new_new_n12868__, new_new_n12869__,
    new_new_n12870__, new_new_n12871__, new_new_n12872__, new_new_n12873__,
    new_new_n12874__, new_new_n12875__, new_new_n12876__, new_new_n12877__,
    new_new_n12878__, new_new_n12879__, new_new_n12880__, new_new_n12881__,
    new_new_n12882__, new_new_n12883__, new_new_n12884__, new_new_n12885__,
    new_new_n12886__, new_new_n12887__, new_new_n12888__, new_new_n12889__,
    new_new_n12890__, new_new_n12891__, new_new_n12892__, new_new_n12893__,
    new_new_n12894__, new_new_n12895__, new_new_n12896__, new_new_n12897__,
    new_new_n12898__, new_new_n12899__, new_new_n12900__, new_new_n12901__,
    new_new_n12902__, new_new_n12903__, new_new_n12904__, new_new_n12905__,
    new_new_n12906__, new_new_n12907__, new_new_n12908__, new_new_n12909__,
    new_new_n12910__, new_new_n12911__, new_new_n12912__, new_new_n12913__,
    new_new_n12914__, new_new_n12915__, new_new_n12916__, new_new_n12917__,
    new_new_n12918__, new_new_n12919__, new_new_n12920__, new_new_n12921__,
    new_new_n12922__, new_new_n12923__, new_new_n12924__, new_new_n12925__,
    new_new_n12926__, new_new_n12927__, new_new_n12928__, new_new_n12929__,
    new_new_n12930__, new_new_n12931__, new_new_n12932__, new_new_n12933__,
    new_new_n12934__, new_new_n12935__, new_new_n12936__, new_new_n12937__,
    new_new_n12939__, new_new_n12940__, new_new_n12941__, new_new_n12942__,
    new_new_n12943__, new_new_n12944__, new_new_n12945__, new_new_n12946__,
    new_new_n12947__, new_new_n12948__, new_new_n12949__, new_new_n12950__,
    new_new_n12951__, new_new_n12952__, new_new_n12953__, new_new_n12954__,
    new_new_n12955__, new_new_n12956__, new_new_n12957__, new_new_n12958__,
    new_new_n12959__, new_new_n12960__, new_new_n12961__, new_new_n12962__,
    new_new_n12963__, new_new_n12964__, new_new_n12965__, new_new_n12966__,
    new_new_n12967__, new_new_n12968__, new_new_n12969__, new_new_n12970__,
    new_new_n12971__, new_new_n12972__, new_new_n12973__, new_new_n12974__,
    new_new_n12975__, new_new_n12976__, new_new_n12977__, new_new_n12978__,
    new_new_n12979__, new_new_n12980__, new_new_n12981__, new_new_n12982__,
    new_new_n12983__, new_new_n12984__, new_new_n12985__, new_new_n12986__,
    new_new_n12987__, new_new_n12988__, new_new_n12989__, new_new_n12990__,
    new_new_n12991__, new_new_n12992__, new_new_n12993__, new_new_n12994__,
    new_new_n12995__, new_new_n12996__, new_new_n12997__, new_new_n12998__,
    new_new_n12999__, new_new_n13000__, new_new_n13001__, new_new_n13002__,
    new_new_n13003__, new_new_n13004__, new_new_n13005__, new_new_n13006__,
    new_new_n13007__, new_new_n13008__, new_new_n13009__, new_new_n13010__,
    new_new_n13011__, new_new_n13012__, new_new_n13013__, new_new_n13014__,
    new_new_n13015__, new_new_n13016__, new_new_n13017__, new_new_n13018__,
    new_new_n13019__, new_new_n13020__, new_new_n13021__, new_new_n13022__,
    new_new_n13023__, new_new_n13024__, new_new_n13025__, new_new_n13026__,
    new_new_n13027__, new_new_n13028__, new_new_n13029__, new_new_n13030__,
    new_new_n13031__, new_new_n13032__, new_new_n13033__, new_new_n13034__,
    new_new_n13035__, new_new_n13036__, new_new_n13037__, new_new_n13038__,
    new_new_n13039__, new_new_n13040__, new_new_n13041__, new_new_n13042__,
    new_new_n13043__, new_new_n13044__, new_new_n13045__, new_new_n13046__,
    new_new_n13047__, new_new_n13048__, new_new_n13049__, new_new_n13050__,
    new_new_n13051__, new_new_n13052__, new_new_n13053__, new_new_n13054__,
    new_new_n13055__, new_new_n13056__, new_new_n13057__, new_new_n13058__,
    new_new_n13059__, new_new_n13060__, new_new_n13061__, new_new_n13062__,
    new_new_n13063__, new_new_n13064__, new_new_n13065__, new_new_n13066__,
    new_new_n13067__, new_new_n13068__, new_new_n13069__, new_new_n13070__,
    new_new_n13071__, new_new_n13072__, new_new_n13073__, new_new_n13074__,
    new_new_n13075__, new_new_n13076__, new_new_n13077__, new_new_n13078__,
    new_new_n13079__, new_new_n13080__, new_new_n13081__, new_new_n13082__,
    new_new_n13083__, new_new_n13084__, new_new_n13085__, new_new_n13086__,
    new_new_n13087__, new_new_n13088__, new_new_n13089__, new_new_n13090__,
    new_new_n13091__, new_new_n13092__, new_new_n13093__, new_new_n13094__,
    new_new_n13095__, new_new_n13096__, new_new_n13097__, new_new_n13098__,
    new_new_n13099__, new_new_n13100__, new_new_n13101__, new_new_n13102__,
    new_new_n13103__, new_new_n13104__, new_new_n13105__, new_new_n13106__,
    new_new_n13107__, new_new_n13108__, new_new_n13109__, new_new_n13110__,
    new_new_n13111__, new_new_n13112__, new_new_n13113__, new_new_n13114__,
    new_new_n13115__, new_new_n13116__, new_new_n13117__, new_new_n13118__,
    new_new_n13119__, new_new_n13120__, new_new_n13121__, new_new_n13122__,
    new_new_n13123__, new_new_n13124__, new_new_n13125__, new_new_n13126__,
    new_new_n13127__, new_new_n13128__, new_new_n13129__, new_new_n13130__,
    new_new_n13131__, new_new_n13132__, new_new_n13133__, new_new_n13134__,
    new_new_n13135__, new_new_n13136__, new_new_n13137__, new_new_n13138__,
    new_new_n13139__, new_new_n13140__, new_new_n13141__, new_new_n13142__,
    new_new_n13143__, new_new_n13144__, new_new_n13145__, new_new_n13146__,
    new_new_n13147__, new_new_n13148__, new_new_n13149__, new_new_n13150__,
    new_new_n13151__, new_new_n13152__, new_new_n13153__, new_new_n13154__,
    new_new_n13155__, new_new_n13156__, new_new_n13157__, new_new_n13158__,
    new_new_n13159__, new_new_n13160__, new_new_n13161__, new_new_n13162__,
    new_new_n13163__, new_new_n13164__, new_new_n13165__, new_new_n13166__,
    new_new_n13167__, new_new_n13168__, new_new_n13169__, new_new_n13170__,
    new_new_n13171__, new_new_n13172__, new_new_n13173__, new_new_n13174__,
    new_new_n13175__, new_new_n13176__, new_new_n13177__, new_new_n13178__,
    new_new_n13179__, new_new_n13180__, new_new_n13181__, new_new_n13182__,
    new_new_n13183__, new_new_n13184__, new_new_n13185__, new_new_n13186__,
    new_new_n13187__, new_new_n13188__, new_new_n13189__, new_new_n13190__,
    new_new_n13191__, new_new_n13192__, new_new_n13193__, new_new_n13194__,
    new_new_n13195__, new_new_n13196__, new_new_n13197__, new_new_n13198__,
    new_new_n13199__, new_new_n13200__, new_new_n13201__, new_new_n13202__,
    new_new_n13203__, new_new_n13204__, new_new_n13205__, new_new_n13206__,
    new_new_n13207__, new_new_n13208__, new_new_n13209__, new_new_n13211__,
    new_new_n13212__, new_new_n13213__, new_new_n13214__, new_new_n13215__,
    new_new_n13216__, new_new_n13217__, new_new_n13218__, new_new_n13219__,
    new_new_n13220__, new_new_n13221__, new_new_n13222__, new_new_n13223__,
    new_new_n13224__, new_new_n13225__, new_new_n13226__, new_new_n13227__,
    new_new_n13228__, new_new_n13229__, new_new_n13230__, new_new_n13231__,
    new_new_n13232__, new_new_n13233__, new_new_n13234__, new_new_n13235__,
    new_new_n13236__, new_new_n13237__, new_new_n13238__, new_new_n13239__,
    new_new_n13240__, new_new_n13241__, new_new_n13242__, new_new_n13243__,
    new_new_n13244__, new_new_n13245__, new_new_n13246__, new_new_n13247__,
    new_new_n13248__, new_new_n13249__, new_new_n13250__, new_new_n13251__,
    new_new_n13252__, new_new_n13253__, new_new_n13254__, new_new_n13255__,
    new_new_n13256__, new_new_n13257__, new_new_n13258__, new_new_n13259__,
    new_new_n13260__, new_new_n13261__, new_new_n13262__, new_new_n13263__,
    new_new_n13264__, new_new_n13265__, new_new_n13266__, new_new_n13267__,
    new_new_n13268__, new_new_n13269__, new_new_n13270__, new_new_n13271__,
    new_new_n13272__, new_new_n13273__, new_new_n13274__, new_new_n13275__,
    new_new_n13276__, new_new_n13277__, new_new_n13278__, new_new_n13279__,
    new_new_n13280__, new_new_n13281__, new_new_n13282__, new_new_n13283__,
    new_new_n13284__, new_new_n13285__, new_new_n13286__, new_new_n13287__,
    new_new_n13288__, new_new_n13289__, new_new_n13290__, new_new_n13291__,
    new_new_n13292__, new_new_n13293__, new_new_n13294__, new_new_n13295__,
    new_new_n13296__, new_new_n13297__, new_new_n13298__, new_new_n13299__,
    new_new_n13300__, new_new_n13301__, new_new_n13302__, new_new_n13303__,
    new_new_n13304__, new_new_n13305__, new_new_n13306__, new_new_n13307__,
    new_new_n13308__, new_new_n13309__, new_new_n13310__, new_new_n13311__,
    new_new_n13312__, new_new_n13313__, new_new_n13314__, new_new_n13315__,
    new_new_n13316__, new_new_n13317__, new_new_n13318__, new_new_n13319__,
    new_new_n13320__, new_new_n13321__, new_new_n13322__, new_new_n13323__,
    new_new_n13324__, new_new_n13325__, new_new_n13326__, new_new_n13327__,
    new_new_n13328__, new_new_n13329__, new_new_n13330__, new_new_n13331__,
    new_new_n13332__, new_new_n13333__, new_new_n13334__, new_new_n13335__,
    new_new_n13336__, new_new_n13337__, new_new_n13338__, new_new_n13339__,
    new_new_n13340__, new_new_n13341__, new_new_n13342__, new_new_n13343__,
    new_new_n13344__, new_new_n13345__, new_new_n13346__, new_new_n13347__,
    new_new_n13348__, new_new_n13349__, new_new_n13350__, new_new_n13351__,
    new_new_n13352__, new_new_n13353__, new_new_n13354__, new_new_n13355__,
    new_new_n13356__, new_new_n13357__, new_new_n13358__, new_new_n13359__,
    new_new_n13360__, new_new_n13361__, new_new_n13362__, new_new_n13363__,
    new_new_n13364__, new_new_n13365__, new_new_n13366__, new_new_n13367__,
    new_new_n13368__, new_new_n13369__, new_new_n13370__, new_new_n13371__,
    new_new_n13372__, new_new_n13373__, new_new_n13374__, new_new_n13375__,
    new_new_n13376__, new_new_n13377__, new_new_n13378__, new_new_n13379__,
    new_new_n13380__, new_new_n13381__, new_new_n13382__, new_new_n13383__,
    new_new_n13384__, new_new_n13385__, new_new_n13386__, new_new_n13387__,
    new_new_n13388__, new_new_n13389__, new_new_n13390__, new_new_n13391__,
    new_new_n13392__, new_new_n13393__, new_new_n13394__, new_new_n13395__,
    new_new_n13396__, new_new_n13397__, new_new_n13398__, new_new_n13399__,
    new_new_n13400__, new_new_n13401__, new_new_n13402__, new_new_n13403__,
    new_new_n13404__, new_new_n13405__, new_new_n13406__, new_new_n13407__,
    new_new_n13408__, new_new_n13409__, new_new_n13410__, new_new_n13411__,
    new_new_n13412__, new_new_n13413__, new_new_n13414__, new_new_n13415__,
    new_new_n13416__, new_new_n13417__, new_new_n13418__, new_new_n13419__,
    new_new_n13420__, new_new_n13421__, new_new_n13422__, new_new_n13423__,
    new_new_n13424__, new_new_n13425__, new_new_n13426__, new_new_n13427__,
    new_new_n13428__, new_new_n13429__, new_new_n13430__, new_new_n13431__,
    new_new_n13432__, new_new_n13433__, new_new_n13434__, new_new_n13435__,
    new_new_n13436__, new_new_n13437__, new_new_n13438__, new_new_n13439__,
    new_new_n13440__, new_new_n13441__, new_new_n13443__, new_new_n13444__,
    new_new_n13445__, new_new_n13446__, new_new_n13447__, new_new_n13448__,
    new_new_n13449__, new_new_n13450__, new_new_n13451__, new_new_n13452__,
    new_new_n13453__, new_new_n13454__, new_new_n13455__, new_new_n13456__,
    new_new_n13457__, new_new_n13458__, new_new_n13459__, new_new_n13460__,
    new_new_n13461__, new_new_n13462__, new_new_n13463__, new_new_n13464__,
    new_new_n13465__, new_new_n13466__, new_new_n13467__, new_new_n13468__,
    new_new_n13469__, new_new_n13470__, new_new_n13471__, new_new_n13472__,
    new_new_n13473__, new_new_n13474__, new_new_n13475__, new_new_n13476__,
    new_new_n13477__, new_new_n13478__, new_new_n13479__, new_new_n13480__,
    new_new_n13481__, new_new_n13482__, new_new_n13483__, new_new_n13484__,
    new_new_n13485__, new_new_n13486__, new_new_n13487__, new_new_n13488__,
    new_new_n13489__, new_new_n13490__, new_new_n13491__, new_new_n13492__,
    new_new_n13493__, new_new_n13494__, new_new_n13495__, new_new_n13496__,
    new_new_n13497__, new_new_n13498__, new_new_n13499__, new_new_n13500__,
    new_new_n13501__, new_new_n13502__, new_new_n13503__, new_new_n13504__,
    new_new_n13505__, new_new_n13506__, new_new_n13507__, new_new_n13508__,
    new_new_n13509__, new_new_n13510__, new_new_n13511__, new_new_n13512__,
    new_new_n13513__, new_new_n13514__, new_new_n13515__, new_new_n13516__,
    new_new_n13517__, new_new_n13518__, new_new_n13519__, new_new_n13520__,
    new_new_n13521__, new_new_n13522__, new_new_n13523__, new_new_n13524__,
    new_new_n13525__, new_new_n13526__, new_new_n13527__, new_new_n13528__,
    new_new_n13529__, new_new_n13530__, new_new_n13531__, new_new_n13532__,
    new_new_n13533__, new_new_n13534__, new_new_n13535__, new_new_n13536__,
    new_new_n13537__, new_new_n13538__, new_new_n13539__, new_new_n13540__,
    new_new_n13541__, new_new_n13542__, new_new_n13543__, new_new_n13544__,
    new_new_n13545__, new_new_n13546__, new_new_n13547__, new_new_n13548__,
    new_new_n13549__, new_new_n13550__, new_new_n13551__, new_new_n13552__,
    new_new_n13553__, new_new_n13554__, new_new_n13555__, new_new_n13556__,
    new_new_n13557__, new_new_n13558__, new_new_n13559__, new_new_n13560__,
    new_new_n13561__, new_new_n13562__, new_new_n13563__, new_new_n13564__,
    new_new_n13565__, new_new_n13566__, new_new_n13567__, new_new_n13568__,
    new_new_n13569__, new_new_n13570__, new_new_n13571__, new_new_n13572__,
    new_new_n13573__, new_new_n13574__, new_new_n13575__, new_new_n13576__,
    new_new_n13577__, new_new_n13578__, new_new_n13579__, new_new_n13580__,
    new_new_n13581__, new_new_n13582__, new_new_n13583__, new_new_n13584__,
    new_new_n13585__, new_new_n13586__, new_new_n13587__, new_new_n13588__,
    new_new_n13589__, new_new_n13590__, new_new_n13591__, new_new_n13592__,
    new_new_n13593__, new_new_n13594__, new_new_n13595__, new_new_n13596__,
    new_new_n13597__, new_new_n13598__, new_new_n13599__, new_new_n13600__,
    new_new_n13601__, new_new_n13602__, new_new_n13603__, new_new_n13604__,
    new_new_n13605__, new_new_n13606__, new_new_n13607__, new_new_n13608__,
    new_new_n13609__, new_new_n13610__, new_new_n13611__, new_new_n13612__,
    new_new_n13613__, new_new_n13614__, new_new_n13615__, new_new_n13616__,
    new_new_n13617__, new_new_n13618__, new_new_n13619__, new_new_n13620__,
    new_new_n13621__, new_new_n13622__, new_new_n13623__, new_new_n13624__,
    new_new_n13625__, new_new_n13626__, new_new_n13627__, new_new_n13628__,
    new_new_n13629__, new_new_n13630__, new_new_n13631__, new_new_n13632__,
    new_new_n13633__, new_new_n13634__, new_new_n13635__, new_new_n13636__,
    new_new_n13637__, new_new_n13638__, new_new_n13639__, new_new_n13640__,
    new_new_n13641__, new_new_n13642__, new_new_n13643__, new_new_n13644__,
    new_new_n13645__, new_new_n13646__, new_new_n13647__, new_new_n13648__,
    new_new_n13649__, new_new_n13650__, new_new_n13651__, new_new_n13652__,
    new_new_n13653__, new_new_n13654__, new_new_n13655__, new_new_n13656__,
    new_new_n13657__, new_new_n13658__, new_new_n13659__, new_new_n13660__,
    new_new_n13661__, new_new_n13662__, new_new_n13663__, new_new_n13664__,
    new_new_n13665__, new_new_n13666__, new_new_n13667__, new_new_n13668__,
    new_new_n13669__, new_new_n13670__, new_new_n13671__, new_new_n13672__,
    new_new_n13673__, new_new_n13674__, new_new_n13675__, new_new_n13676__,
    new_new_n13677__, new_new_n13678__, new_new_n13679__, new_new_n13680__,
    new_new_n13681__, new_new_n13682__, new_new_n13683__, new_new_n13684__,
    new_new_n13685__, new_new_n13686__, new_new_n13687__, new_new_n13688__,
    new_new_n13689__, new_new_n13690__, new_new_n13691__, new_new_n13692__,
    new_new_n13693__, new_new_n13694__, new_new_n13695__, new_new_n13696__,
    new_new_n13697__, new_new_n13698__, new_new_n13699__, new_new_n13700__,
    new_new_n13701__, new_new_n13702__, new_new_n13703__, new_new_n13704__,
    new_new_n13705__, new_new_n13706__, new_new_n13707__, new_new_n13708__,
    new_new_n13710__, new_new_n13711__, new_new_n13712__, new_new_n13713__,
    new_new_n13714__, new_new_n13715__, new_new_n13716__, new_new_n13717__,
    new_new_n13718__, new_new_n13719__, new_new_n13720__, new_new_n13721__,
    new_new_n13722__, new_new_n13723__, new_new_n13724__, new_new_n13725__,
    new_new_n13726__, new_new_n13727__, new_new_n13728__, new_new_n13729__,
    new_new_n13730__, new_new_n13731__, new_new_n13732__, new_new_n13733__,
    new_new_n13734__, new_new_n13735__, new_new_n13736__, new_new_n13737__,
    new_new_n13738__, new_new_n13739__, new_new_n13740__, new_new_n13741__,
    new_new_n13742__, new_new_n13743__, new_new_n13744__, new_new_n13745__,
    new_new_n13746__, new_new_n13747__, new_new_n13748__, new_new_n13749__,
    new_new_n13750__, new_new_n13751__, new_new_n13752__, new_new_n13753__,
    new_new_n13754__, new_new_n13755__, new_new_n13756__, new_new_n13757__,
    new_new_n13758__, new_new_n13759__, new_new_n13760__, new_new_n13761__,
    new_new_n13762__, new_new_n13763__, new_new_n13764__, new_new_n13765__,
    new_new_n13766__, new_new_n13767__, new_new_n13768__, new_new_n13769__,
    new_new_n13770__, new_new_n13771__, new_new_n13772__, new_new_n13773__,
    new_new_n13774__, new_new_n13775__, new_new_n13776__, new_new_n13777__,
    new_new_n13778__, new_new_n13779__, new_new_n13780__, new_new_n13781__,
    new_new_n13782__, new_new_n13783__, new_new_n13784__, new_new_n13785__,
    new_new_n13786__, new_new_n13787__, new_new_n13788__, new_new_n13789__,
    new_new_n13790__, new_new_n13791__, new_new_n13792__, new_new_n13793__,
    new_new_n13794__, new_new_n13795__, new_new_n13796__, new_new_n13797__,
    new_new_n13798__, new_new_n13799__, new_new_n13800__, new_new_n13801__,
    new_new_n13802__, new_new_n13803__, new_new_n13804__, new_new_n13805__,
    new_new_n13806__, new_new_n13807__, new_new_n13808__, new_new_n13809__,
    new_new_n13810__, new_new_n13811__, new_new_n13812__, new_new_n13813__,
    new_new_n13814__, new_new_n13815__, new_new_n13816__, new_new_n13817__,
    new_new_n13818__, new_new_n13819__, new_new_n13820__, new_new_n13821__,
    new_new_n13822__, new_new_n13823__, new_new_n13824__, new_new_n13825__,
    new_new_n13826__, new_new_n13827__, new_new_n13828__, new_new_n13829__,
    new_new_n13830__, new_new_n13831__, new_new_n13832__, new_new_n13833__,
    new_new_n13834__, new_new_n13835__, new_new_n13836__, new_new_n13837__,
    new_new_n13838__, new_new_n13839__, new_new_n13840__, new_new_n13841__,
    new_new_n13842__, new_new_n13843__, new_new_n13844__, new_new_n13845__,
    new_new_n13846__, new_new_n13847__, new_new_n13848__, new_new_n13849__,
    new_new_n13850__, new_new_n13851__, new_new_n13852__, new_new_n13853__,
    new_new_n13854__, new_new_n13855__, new_new_n13856__, new_new_n13857__,
    new_new_n13858__, new_new_n13859__, new_new_n13860__, new_new_n13861__,
    new_new_n13862__, new_new_n13863__, new_new_n13864__, new_new_n13865__,
    new_new_n13866__, new_new_n13867__, new_new_n13868__, new_new_n13869__,
    new_new_n13870__, new_new_n13871__, new_new_n13872__, new_new_n13873__,
    new_new_n13874__, new_new_n13875__, new_new_n13876__, new_new_n13877__,
    new_new_n13878__, new_new_n13879__, new_new_n13880__, new_new_n13881__,
    new_new_n13882__, new_new_n13883__, new_new_n13884__, new_new_n13885__,
    new_new_n13886__, new_new_n13887__, new_new_n13888__, new_new_n13889__,
    new_new_n13890__, new_new_n13891__, new_new_n13892__, new_new_n13893__,
    new_new_n13894__, new_new_n13895__, new_new_n13896__, new_new_n13897__,
    new_new_n13898__, new_new_n13899__, new_new_n13900__, new_new_n13901__,
    new_new_n13902__, new_new_n13903__, new_new_n13904__, new_new_n13905__,
    new_new_n13906__, new_new_n13907__, new_new_n13908__, new_new_n13909__,
    new_new_n13910__, new_new_n13911__, new_new_n13912__, new_new_n13913__,
    new_new_n13914__, new_new_n13915__, new_new_n13916__, new_new_n13917__,
    new_new_n13918__, new_new_n13919__, new_new_n13920__, new_new_n13921__,
    new_new_n13922__, new_new_n13923__, new_new_n13924__, new_new_n13925__,
    new_new_n13926__, new_new_n13927__, new_new_n13928__, new_new_n13929__,
    new_new_n13930__, new_new_n13931__, new_new_n13932__, new_new_n13933__,
    new_new_n13934__, new_new_n13935__, new_new_n13936__, new_new_n13937__,
    new_new_n13938__, new_new_n13939__, new_new_n13940__, new_new_n13941__,
    new_new_n13942__, new_new_n13943__, new_new_n13944__, new_new_n13945__,
    new_new_n13946__, new_new_n13947__, new_new_n13948__, new_new_n13949__,
    new_new_n13951__, new_new_n13952__, new_new_n13953__, new_new_n13954__,
    new_new_n13955__, new_new_n13956__, new_new_n13957__, new_new_n13958__,
    new_new_n13959__, new_new_n13960__, new_new_n13961__, new_new_n13962__,
    new_new_n13963__, new_new_n13964__, new_new_n13965__, new_new_n13966__,
    new_new_n13967__, new_new_n13968__, new_new_n13969__, new_new_n13970__,
    new_new_n13971__, new_new_n13972__, new_new_n13973__, new_new_n13974__,
    new_new_n13975__, new_new_n13976__, new_new_n13977__, new_new_n13978__,
    new_new_n13979__, new_new_n13980__, new_new_n13981__, new_new_n13982__,
    new_new_n13983__, new_new_n13984__, new_new_n13985__, new_new_n13986__,
    new_new_n13987__, new_new_n13988__, new_new_n13989__, new_new_n13990__,
    new_new_n13991__, new_new_n13992__, new_new_n13993__, new_new_n13994__,
    new_new_n13995__, new_new_n13996__, new_new_n13997__, new_new_n13998__,
    new_new_n13999__, new_new_n14000__, new_new_n14001__, new_new_n14002__,
    new_new_n14003__, new_new_n14004__, new_new_n14005__, new_new_n14006__,
    new_new_n14007__, new_new_n14008__, new_new_n14009__, new_new_n14010__,
    new_new_n14011__, new_new_n14012__, new_new_n14013__, new_new_n14014__,
    new_new_n14015__, new_new_n14016__, new_new_n14017__, new_new_n14018__,
    new_new_n14019__, new_new_n14020__, new_new_n14021__, new_new_n14022__,
    new_new_n14023__, new_new_n14024__, new_new_n14025__, new_new_n14026__,
    new_new_n14027__, new_new_n14028__, new_new_n14029__, new_new_n14030__,
    new_new_n14031__, new_new_n14032__, new_new_n14033__, new_new_n14034__,
    new_new_n14035__, new_new_n14036__, new_new_n14037__, new_new_n14038__,
    new_new_n14039__, new_new_n14040__, new_new_n14041__, new_new_n14042__,
    new_new_n14043__, new_new_n14044__, new_new_n14045__, new_new_n14046__,
    new_new_n14047__, new_new_n14048__, new_new_n14049__, new_new_n14050__,
    new_new_n14051__, new_new_n14052__, new_new_n14053__, new_new_n14054__,
    new_new_n14055__, new_new_n14056__, new_new_n14057__, new_new_n14058__,
    new_new_n14059__, new_new_n14060__, new_new_n14061__, new_new_n14062__,
    new_new_n14063__, new_new_n14064__, new_new_n14065__, new_new_n14066__,
    new_new_n14067__, new_new_n14068__, new_new_n14069__, new_new_n14070__,
    new_new_n14071__, new_new_n14072__, new_new_n14073__, new_new_n14074__,
    new_new_n14075__, new_new_n14076__, new_new_n14077__, new_new_n14078__,
    new_new_n14079__, new_new_n14080__, new_new_n14081__, new_new_n14082__,
    new_new_n14083__, new_new_n14084__, new_new_n14085__, new_new_n14086__,
    new_new_n14087__, new_new_n14088__, new_new_n14089__, new_new_n14090__,
    new_new_n14091__, new_new_n14092__, new_new_n14093__, new_new_n14094__,
    new_new_n14095__, new_new_n14096__, new_new_n14097__, new_new_n14098__,
    new_new_n14099__, new_new_n14100__, new_new_n14101__, new_new_n14102__,
    new_new_n14103__, new_new_n14104__, new_new_n14105__, new_new_n14106__,
    new_new_n14107__, new_new_n14108__, new_new_n14109__, new_new_n14110__,
    new_new_n14111__, new_new_n14112__, new_new_n14113__, new_new_n14114__,
    new_new_n14115__, new_new_n14116__, new_new_n14117__, new_new_n14118__,
    new_new_n14119__, new_new_n14120__, new_new_n14121__, new_new_n14122__,
    new_new_n14123__, new_new_n14124__, new_new_n14125__, new_new_n14126__,
    new_new_n14127__, new_new_n14128__, new_new_n14129__, new_new_n14130__,
    new_new_n14131__, new_new_n14132__, new_new_n14133__, new_new_n14134__,
    new_new_n14135__, new_new_n14136__, new_new_n14137__, new_new_n14138__,
    new_new_n14139__, new_new_n14140__, new_new_n14141__, new_new_n14142__,
    new_new_n14143__, new_new_n14144__, new_new_n14145__, new_new_n14146__,
    new_new_n14147__, new_new_n14148__, new_new_n14149__, new_new_n14150__,
    new_new_n14151__, new_new_n14152__, new_new_n14153__, new_new_n14154__,
    new_new_n14155__, new_new_n14156__, new_new_n14157__, new_new_n14158__,
    new_new_n14159__, new_new_n14160__, new_new_n14161__, new_new_n14162__,
    new_new_n14163__, new_new_n14164__, new_new_n14165__, new_new_n14166__,
    new_new_n14167__, new_new_n14168__, new_new_n14169__, new_new_n14170__,
    new_new_n14171__, new_new_n14172__, new_new_n14173__, new_new_n14174__,
    new_new_n14175__, new_new_n14176__, new_new_n14177__, new_new_n14178__,
    new_new_n14179__, new_new_n14180__, new_new_n14181__, new_new_n14182__,
    new_new_n14183__, new_new_n14184__, new_new_n14185__, new_new_n14186__,
    new_new_n14187__, new_new_n14188__, new_new_n14189__, new_new_n14190__,
    new_new_n14191__, new_new_n14192__, new_new_n14193__, new_new_n14194__,
    new_new_n14195__, new_new_n14196__, new_new_n14198__, new_new_n14199__,
    new_new_n14200__, new_new_n14201__, new_new_n14202__, new_new_n14203__,
    new_new_n14204__, new_new_n14205__, new_new_n14206__, new_new_n14207__,
    new_new_n14208__, new_new_n14209__, new_new_n14210__, new_new_n14211__,
    new_new_n14212__, new_new_n14213__, new_new_n14214__, new_new_n14215__,
    new_new_n14216__, new_new_n14217__, new_new_n14218__, new_new_n14219__,
    new_new_n14220__, new_new_n14221__, new_new_n14222__, new_new_n14223__,
    new_new_n14224__, new_new_n14225__, new_new_n14226__, new_new_n14227__,
    new_new_n14228__, new_new_n14229__, new_new_n14230__, new_new_n14231__,
    new_new_n14232__, new_new_n14233__, new_new_n14234__, new_new_n14235__,
    new_new_n14236__, new_new_n14237__, new_new_n14238__, new_new_n14239__,
    new_new_n14240__, new_new_n14241__, new_new_n14242__, new_new_n14243__,
    new_new_n14244__, new_new_n14245__, new_new_n14246__, new_new_n14247__,
    new_new_n14248__, new_new_n14249__, new_new_n14250__, new_new_n14251__,
    new_new_n14252__, new_new_n14253__, new_new_n14254__, new_new_n14255__,
    new_new_n14256__, new_new_n14257__, new_new_n14258__, new_new_n14259__,
    new_new_n14260__, new_new_n14261__, new_new_n14262__, new_new_n14263__,
    new_new_n14264__, new_new_n14265__, new_new_n14266__, new_new_n14267__,
    new_new_n14268__, new_new_n14269__, new_new_n14270__, new_new_n14271__,
    new_new_n14272__, new_new_n14273__, new_new_n14274__, new_new_n14275__,
    new_new_n14276__, new_new_n14277__, new_new_n14278__, new_new_n14279__,
    new_new_n14280__, new_new_n14281__, new_new_n14282__, new_new_n14283__,
    new_new_n14284__, new_new_n14285__, new_new_n14286__, new_new_n14287__,
    new_new_n14288__, new_new_n14289__, new_new_n14290__, new_new_n14291__,
    new_new_n14292__, new_new_n14293__, new_new_n14294__, new_new_n14295__,
    new_new_n14296__, new_new_n14297__, new_new_n14298__, new_new_n14299__,
    new_new_n14300__, new_new_n14301__, new_new_n14302__, new_new_n14303__,
    new_new_n14304__, new_new_n14305__, new_new_n14306__, new_new_n14307__,
    new_new_n14308__, new_new_n14309__, new_new_n14310__, new_new_n14311__,
    new_new_n14312__, new_new_n14313__, new_new_n14314__, new_new_n14315__,
    new_new_n14316__, new_new_n14317__, new_new_n14318__, new_new_n14319__,
    new_new_n14320__, new_new_n14321__, new_new_n14322__, new_new_n14323__,
    new_new_n14324__, new_new_n14325__, new_new_n14326__, new_new_n14327__,
    new_new_n14328__, new_new_n14329__, new_new_n14330__, new_new_n14331__,
    new_new_n14332__, new_new_n14333__, new_new_n14334__, new_new_n14335__,
    new_new_n14336__, new_new_n14337__, new_new_n14338__, new_new_n14339__,
    new_new_n14340__, new_new_n14341__, new_new_n14342__, new_new_n14343__,
    new_new_n14344__, new_new_n14345__, new_new_n14346__, new_new_n14347__,
    new_new_n14348__, new_new_n14349__, new_new_n14350__, new_new_n14351__,
    new_new_n14352__, new_new_n14353__, new_new_n14354__, new_new_n14355__,
    new_new_n14356__, new_new_n14357__, new_new_n14358__, new_new_n14359__,
    new_new_n14360__, new_new_n14361__, new_new_n14362__, new_new_n14363__,
    new_new_n14364__, new_new_n14365__, new_new_n14366__, new_new_n14367__,
    new_new_n14368__, new_new_n14369__, new_new_n14370__, new_new_n14371__,
    new_new_n14372__, new_new_n14373__, new_new_n14374__, new_new_n14375__,
    new_new_n14376__, new_new_n14377__, new_new_n14378__, new_new_n14379__,
    new_new_n14380__, new_new_n14381__, new_new_n14382__, new_new_n14383__,
    new_new_n14384__, new_new_n14385__, new_new_n14386__, new_new_n14387__,
    new_new_n14388__, new_new_n14389__, new_new_n14390__, new_new_n14391__,
    new_new_n14392__, new_new_n14393__, new_new_n14394__, new_new_n14395__,
    new_new_n14396__, new_new_n14397__, new_new_n14398__, new_new_n14399__,
    new_new_n14400__, new_new_n14401__, new_new_n14402__, new_new_n14403__,
    new_new_n14404__, new_new_n14405__, new_new_n14406__, new_new_n14407__,
    new_new_n14408__, new_new_n14409__, new_new_n14410__, new_new_n14411__,
    new_new_n14412__, new_new_n14413__, new_new_n14414__, new_new_n14415__,
    new_new_n14416__, new_new_n14417__, new_new_n14418__, new_new_n14419__,
    new_new_n14420__, new_new_n14422__, new_new_n14423__, new_new_n14424__,
    new_new_n14425__, new_new_n14426__, new_new_n14427__, new_new_n14428__,
    new_new_n14429__, new_new_n14430__, new_new_n14431__, new_new_n14432__,
    new_new_n14433__, new_new_n14434__, new_new_n14435__, new_new_n14436__,
    new_new_n14437__, new_new_n14438__, new_new_n14439__, new_new_n14440__,
    new_new_n14441__, new_new_n14442__, new_new_n14443__, new_new_n14444__,
    new_new_n14445__, new_new_n14446__, new_new_n14447__, new_new_n14448__,
    new_new_n14449__, new_new_n14450__, new_new_n14451__, new_new_n14452__,
    new_new_n14453__, new_new_n14454__, new_new_n14455__, new_new_n14456__,
    new_new_n14457__, new_new_n14458__, new_new_n14459__, new_new_n14460__,
    new_new_n14461__, new_new_n14462__, new_new_n14463__, new_new_n14464__,
    new_new_n14465__, new_new_n14466__, new_new_n14467__, new_new_n14468__,
    new_new_n14469__, new_new_n14470__, new_new_n14471__, new_new_n14472__,
    new_new_n14473__, new_new_n14474__, new_new_n14475__, new_new_n14476__,
    new_new_n14477__, new_new_n14478__, new_new_n14479__, new_new_n14480__,
    new_new_n14481__, new_new_n14482__, new_new_n14483__, new_new_n14484__,
    new_new_n14485__, new_new_n14486__, new_new_n14487__, new_new_n14488__,
    new_new_n14489__, new_new_n14490__, new_new_n14491__, new_new_n14492__,
    new_new_n14493__, new_new_n14494__, new_new_n14495__, new_new_n14496__,
    new_new_n14497__, new_new_n14498__, new_new_n14499__, new_new_n14500__,
    new_new_n14501__, new_new_n14502__, new_new_n14503__, new_new_n14504__,
    new_new_n14505__, new_new_n14506__, new_new_n14507__, new_new_n14508__,
    new_new_n14509__, new_new_n14510__, new_new_n14511__, new_new_n14512__,
    new_new_n14513__, new_new_n14514__, new_new_n14515__, new_new_n14516__,
    new_new_n14517__, new_new_n14518__, new_new_n14519__, new_new_n14520__,
    new_new_n14521__, new_new_n14522__, new_new_n14523__, new_new_n14524__,
    new_new_n14525__, new_new_n14526__, new_new_n14527__, new_new_n14528__,
    new_new_n14529__, new_new_n14530__, new_new_n14531__, new_new_n14532__,
    new_new_n14533__, new_new_n14534__, new_new_n14535__, new_new_n14536__,
    new_new_n14537__, new_new_n14538__, new_new_n14539__, new_new_n14540__,
    new_new_n14541__, new_new_n14542__, new_new_n14543__, new_new_n14544__,
    new_new_n14545__, new_new_n14546__, new_new_n14547__, new_new_n14548__,
    new_new_n14549__, new_new_n14550__, new_new_n14551__, new_new_n14552__,
    new_new_n14553__, new_new_n14554__, new_new_n14555__, new_new_n14556__,
    new_new_n14557__, new_new_n14558__, new_new_n14559__, new_new_n14560__,
    new_new_n14561__, new_new_n14562__, new_new_n14563__, new_new_n14564__,
    new_new_n14565__, new_new_n14566__, new_new_n14567__, new_new_n14568__,
    new_new_n14569__, new_new_n14570__, new_new_n14571__, new_new_n14572__,
    new_new_n14573__, new_new_n14574__, new_new_n14575__, new_new_n14576__,
    new_new_n14577__, new_new_n14578__, new_new_n14579__, new_new_n14580__,
    new_new_n14581__, new_new_n14582__, new_new_n14583__, new_new_n14584__,
    new_new_n14585__, new_new_n14586__, new_new_n14587__, new_new_n14588__,
    new_new_n14589__, new_new_n14590__, new_new_n14591__, new_new_n14592__,
    new_new_n14593__, new_new_n14594__, new_new_n14595__, new_new_n14596__,
    new_new_n14597__, new_new_n14598__, new_new_n14599__, new_new_n14600__,
    new_new_n14601__, new_new_n14602__, new_new_n14603__, new_new_n14604__,
    new_new_n14605__, new_new_n14606__, new_new_n14607__, new_new_n14608__,
    new_new_n14609__, new_new_n14610__, new_new_n14611__, new_new_n14612__,
    new_new_n14613__, new_new_n14614__, new_new_n14615__, new_new_n14616__,
    new_new_n14617__, new_new_n14618__, new_new_n14619__, new_new_n14620__,
    new_new_n14621__, new_new_n14622__, new_new_n14623__, new_new_n14624__,
    new_new_n14625__, new_new_n14626__, new_new_n14627__, new_new_n14628__,
    new_new_n14630__, new_new_n14631__, new_new_n14632__, new_new_n14633__,
    new_new_n14634__, new_new_n14635__, new_new_n14636__, new_new_n14637__,
    new_new_n14638__, new_new_n14639__, new_new_n14640__, new_new_n14641__,
    new_new_n14642__, new_new_n14643__, new_new_n14644__, new_new_n14645__,
    new_new_n14646__, new_new_n14647__, new_new_n14648__, new_new_n14649__,
    new_new_n14650__, new_new_n14651__, new_new_n14652__, new_new_n14653__,
    new_new_n14654__, new_new_n14655__, new_new_n14656__, new_new_n14657__,
    new_new_n14658__, new_new_n14659__, new_new_n14660__, new_new_n14661__,
    new_new_n14662__, new_new_n14663__, new_new_n14664__, new_new_n14665__,
    new_new_n14666__, new_new_n14667__, new_new_n14668__, new_new_n14669__,
    new_new_n14670__, new_new_n14671__, new_new_n14672__, new_new_n14673__,
    new_new_n14674__, new_new_n14675__, new_new_n14676__, new_new_n14677__,
    new_new_n14678__, new_new_n14679__, new_new_n14680__, new_new_n14681__,
    new_new_n14682__, new_new_n14683__, new_new_n14684__, new_new_n14685__,
    new_new_n14686__, new_new_n14687__, new_new_n14688__, new_new_n14689__,
    new_new_n14690__, new_new_n14691__, new_new_n14692__, new_new_n14693__,
    new_new_n14694__, new_new_n14695__, new_new_n14696__, new_new_n14697__,
    new_new_n14698__, new_new_n14699__, new_new_n14700__, new_new_n14701__,
    new_new_n14702__, new_new_n14703__, new_new_n14704__, new_new_n14705__,
    new_new_n14706__, new_new_n14707__, new_new_n14708__, new_new_n14709__,
    new_new_n14710__, new_new_n14711__, new_new_n14712__, new_new_n14713__,
    new_new_n14714__, new_new_n14715__, new_new_n14716__, new_new_n14717__,
    new_new_n14718__, new_new_n14719__, new_new_n14720__, new_new_n14721__,
    new_new_n14722__, new_new_n14723__, new_new_n14724__, new_new_n14725__,
    new_new_n14726__, new_new_n14727__, new_new_n14728__, new_new_n14729__,
    new_new_n14730__, new_new_n14731__, new_new_n14732__, new_new_n14733__,
    new_new_n14734__, new_new_n14735__, new_new_n14736__, new_new_n14737__,
    new_new_n14738__, new_new_n14739__, new_new_n14740__, new_new_n14741__,
    new_new_n14742__, new_new_n14743__, new_new_n14744__, new_new_n14745__,
    new_new_n14746__, new_new_n14747__, new_new_n14748__, new_new_n14749__,
    new_new_n14750__, new_new_n14751__, new_new_n14752__, new_new_n14753__,
    new_new_n14754__, new_new_n14755__, new_new_n14756__, new_new_n14757__,
    new_new_n14758__, new_new_n14759__, new_new_n14760__, new_new_n14761__,
    new_new_n14762__, new_new_n14763__, new_new_n14764__, new_new_n14765__,
    new_new_n14766__, new_new_n14767__, new_new_n14768__, new_new_n14769__,
    new_new_n14770__, new_new_n14771__, new_new_n14772__, new_new_n14773__,
    new_new_n14774__, new_new_n14775__, new_new_n14776__, new_new_n14777__,
    new_new_n14778__, new_new_n14779__, new_new_n14780__, new_new_n14781__,
    new_new_n14782__, new_new_n14783__, new_new_n14784__, new_new_n14785__,
    new_new_n14786__, new_new_n14787__, new_new_n14788__, new_new_n14789__,
    new_new_n14790__, new_new_n14791__, new_new_n14792__, new_new_n14793__,
    new_new_n14794__, new_new_n14795__, new_new_n14796__, new_new_n14797__,
    new_new_n14798__, new_new_n14799__, new_new_n14800__, new_new_n14801__,
    new_new_n14802__, new_new_n14803__, new_new_n14804__, new_new_n14805__,
    new_new_n14806__, new_new_n14807__, new_new_n14808__, new_new_n14809__,
    new_new_n14810__, new_new_n14811__, new_new_n14812__, new_new_n14813__,
    new_new_n14814__, new_new_n14815__, new_new_n14816__, new_new_n14817__,
    new_new_n14818__, new_new_n14819__, new_new_n14820__, new_new_n14821__,
    new_new_n14822__, new_new_n14823__, new_new_n14824__, new_new_n14825__,
    new_new_n14826__, new_new_n14827__, new_new_n14828__, new_new_n14829__,
    new_new_n14830__, new_new_n14831__, new_new_n14832__, new_new_n14833__,
    new_new_n14834__, new_new_n14835__, new_new_n14836__, new_new_n14837__,
    new_new_n14838__, new_new_n14839__, new_new_n14840__, new_new_n14841__,
    new_new_n14842__, new_new_n14843__, new_new_n14844__, new_new_n14845__,
    new_new_n14846__, new_new_n14847__, new_new_n14848__, new_new_n14849__,
    new_new_n14850__, new_new_n14851__, new_new_n14852__, new_new_n14853__,
    new_new_n14854__, new_new_n14855__, new_new_n14857__, new_new_n14858__,
    new_new_n14859__, new_new_n14860__, new_new_n14861__, new_new_n14862__,
    new_new_n14863__, new_new_n14864__, new_new_n14865__, new_new_n14866__,
    new_new_n14867__, new_new_n14868__, new_new_n14869__, new_new_n14870__,
    new_new_n14871__, new_new_n14872__, new_new_n14873__, new_new_n14874__,
    new_new_n14875__, new_new_n14876__, new_new_n14877__, new_new_n14878__,
    new_new_n14879__, new_new_n14880__, new_new_n14881__, new_new_n14882__,
    new_new_n14883__, new_new_n14884__, new_new_n14885__, new_new_n14886__,
    new_new_n14887__, new_new_n14888__, new_new_n14889__, new_new_n14890__,
    new_new_n14891__, new_new_n14892__, new_new_n14893__, new_new_n14894__,
    new_new_n14895__, new_new_n14896__, new_new_n14897__, new_new_n14898__,
    new_new_n14899__, new_new_n14900__, new_new_n14901__, new_new_n14902__,
    new_new_n14903__, new_new_n14904__, new_new_n14905__, new_new_n14906__,
    new_new_n14907__, new_new_n14908__, new_new_n14909__, new_new_n14910__,
    new_new_n14911__, new_new_n14912__, new_new_n14913__, new_new_n14914__,
    new_new_n14915__, new_new_n14916__, new_new_n14917__, new_new_n14918__,
    new_new_n14919__, new_new_n14920__, new_new_n14921__, new_new_n14922__,
    new_new_n14923__, new_new_n14924__, new_new_n14925__, new_new_n14926__,
    new_new_n14927__, new_new_n14928__, new_new_n14929__, new_new_n14930__,
    new_new_n14931__, new_new_n14932__, new_new_n14933__, new_new_n14934__,
    new_new_n14935__, new_new_n14936__, new_new_n14937__, new_new_n14938__,
    new_new_n14939__, new_new_n14940__, new_new_n14941__, new_new_n14942__,
    new_new_n14943__, new_new_n14944__, new_new_n14945__, new_new_n14946__,
    new_new_n14947__, new_new_n14948__, new_new_n14949__, new_new_n14950__,
    new_new_n14951__, new_new_n14952__, new_new_n14953__, new_new_n14954__,
    new_new_n14955__, new_new_n14956__, new_new_n14957__, new_new_n14958__,
    new_new_n14959__, new_new_n14960__, new_new_n14961__, new_new_n14962__,
    new_new_n14963__, new_new_n14964__, new_new_n14965__, new_new_n14966__,
    new_new_n14967__, new_new_n14968__, new_new_n14969__, new_new_n14970__,
    new_new_n14971__, new_new_n14972__, new_new_n14973__, new_new_n14974__,
    new_new_n14975__, new_new_n14976__, new_new_n14977__, new_new_n14978__,
    new_new_n14979__, new_new_n14980__, new_new_n14981__, new_new_n14982__,
    new_new_n14983__, new_new_n14984__, new_new_n14985__, new_new_n14986__,
    new_new_n14987__, new_new_n14988__, new_new_n14989__, new_new_n14990__,
    new_new_n14991__, new_new_n14992__, new_new_n14993__, new_new_n14994__,
    new_new_n14995__, new_new_n14996__, new_new_n14997__, new_new_n14998__,
    new_new_n14999__, new_new_n15000__, new_new_n15001__, new_new_n15002__,
    new_new_n15003__, new_new_n15004__, new_new_n15005__, new_new_n15006__,
    new_new_n15007__, new_new_n15008__, new_new_n15009__, new_new_n15010__,
    new_new_n15011__, new_new_n15012__, new_new_n15013__, new_new_n15014__,
    new_new_n15015__, new_new_n15016__, new_new_n15017__, new_new_n15018__,
    new_new_n15019__, new_new_n15020__, new_new_n15021__, new_new_n15022__,
    new_new_n15023__, new_new_n15024__, new_new_n15025__, new_new_n15026__,
    new_new_n15027__, new_new_n15028__, new_new_n15029__, new_new_n15030__,
    new_new_n15031__, new_new_n15032__, new_new_n15033__, new_new_n15034__,
    new_new_n15035__, new_new_n15036__, new_new_n15037__, new_new_n15038__,
    new_new_n15039__, new_new_n15040__, new_new_n15041__, new_new_n15042__,
    new_new_n15043__, new_new_n15044__, new_new_n15045__, new_new_n15046__,
    new_new_n15047__, new_new_n15048__, new_new_n15049__, new_new_n15050__,
    new_new_n15051__, new_new_n15052__, new_new_n15053__, new_new_n15054__,
    new_new_n15055__, new_new_n15056__, new_new_n15057__, new_new_n15058__,
    new_new_n15059__, new_new_n15060__, new_new_n15061__, new_new_n15062__,
    new_new_n15063__, new_new_n15064__, new_new_n15065__, new_new_n15066__,
    new_new_n15067__, new_new_n15068__, new_new_n15069__, new_new_n15070__,
    new_new_n15071__, new_new_n15072__, new_new_n15073__, new_new_n15074__,
    new_new_n15075__, new_new_n15076__, new_new_n15077__, new_new_n15078__,
    new_new_n15079__, new_new_n15080__, new_new_n15081__, new_new_n15082__,
    new_new_n15083__, new_new_n15084__, new_new_n15085__, new_new_n15086__,
    new_new_n15087__, new_new_n15088__, new_new_n15089__, new_new_n15090__,
    new_new_n15091__, new_new_n15092__, new_new_n15093__, new_new_n15095__,
    new_new_n15096__, new_new_n15097__, new_new_n15098__, new_new_n15099__,
    new_new_n15100__, new_new_n15101__, new_new_n15102__, new_new_n15103__,
    new_new_n15104__, new_new_n15105__, new_new_n15106__, new_new_n15107__,
    new_new_n15108__, new_new_n15109__, new_new_n15110__, new_new_n15111__,
    new_new_n15112__, new_new_n15113__, new_new_n15114__, new_new_n15115__,
    new_new_n15116__, new_new_n15117__, new_new_n15118__, new_new_n15119__,
    new_new_n15120__, new_new_n15121__, new_new_n15122__, new_new_n15123__,
    new_new_n15124__, new_new_n15125__, new_new_n15126__, new_new_n15127__,
    new_new_n15128__, new_new_n15129__, new_new_n15130__, new_new_n15131__,
    new_new_n15132__, new_new_n15133__, new_new_n15134__, new_new_n15135__,
    new_new_n15136__, new_new_n15137__, new_new_n15138__, new_new_n15139__,
    new_new_n15140__, new_new_n15141__, new_new_n15142__, new_new_n15143__,
    new_new_n15144__, new_new_n15145__, new_new_n15146__, new_new_n15147__,
    new_new_n15148__, new_new_n15149__, new_new_n15150__, new_new_n15151__,
    new_new_n15152__, new_new_n15153__, new_new_n15154__, new_new_n15155__,
    new_new_n15156__, new_new_n15157__, new_new_n15158__, new_new_n15159__,
    new_new_n15160__, new_new_n15161__, new_new_n15162__, new_new_n15163__,
    new_new_n15164__, new_new_n15165__, new_new_n15166__, new_new_n15167__,
    new_new_n15168__, new_new_n15169__, new_new_n15170__, new_new_n15171__,
    new_new_n15172__, new_new_n15173__, new_new_n15174__, new_new_n15175__,
    new_new_n15176__, new_new_n15177__, new_new_n15178__, new_new_n15179__,
    new_new_n15180__, new_new_n15181__, new_new_n15182__, new_new_n15183__,
    new_new_n15184__, new_new_n15185__, new_new_n15186__, new_new_n15187__,
    new_new_n15188__, new_new_n15189__, new_new_n15190__, new_new_n15191__,
    new_new_n15192__, new_new_n15193__, new_new_n15194__, new_new_n15195__,
    new_new_n15196__, new_new_n15197__, new_new_n15198__, new_new_n15199__,
    new_new_n15200__, new_new_n15201__, new_new_n15202__, new_new_n15203__,
    new_new_n15204__, new_new_n15205__, new_new_n15206__, new_new_n15207__,
    new_new_n15208__, new_new_n15209__, new_new_n15210__, new_new_n15211__,
    new_new_n15212__, new_new_n15213__, new_new_n15214__, new_new_n15215__,
    new_new_n15216__, new_new_n15217__, new_new_n15218__, new_new_n15219__,
    new_new_n15220__, new_new_n15221__, new_new_n15222__, new_new_n15223__,
    new_new_n15224__, new_new_n15225__, new_new_n15226__, new_new_n15227__,
    new_new_n15228__, new_new_n15229__, new_new_n15230__, new_new_n15231__,
    new_new_n15232__, new_new_n15233__, new_new_n15234__, new_new_n15235__,
    new_new_n15236__, new_new_n15237__, new_new_n15238__, new_new_n15239__,
    new_new_n15240__, new_new_n15241__, new_new_n15242__, new_new_n15243__,
    new_new_n15244__, new_new_n15245__, new_new_n15246__, new_new_n15247__,
    new_new_n15248__, new_new_n15249__, new_new_n15250__, new_new_n15251__,
    new_new_n15252__, new_new_n15253__, new_new_n15254__, new_new_n15255__,
    new_new_n15256__, new_new_n15257__, new_new_n15258__, new_new_n15259__,
    new_new_n15260__, new_new_n15261__, new_new_n15262__, new_new_n15263__,
    new_new_n15264__, new_new_n15265__, new_new_n15266__, new_new_n15267__,
    new_new_n15268__, new_new_n15269__, new_new_n15270__, new_new_n15271__,
    new_new_n15272__, new_new_n15273__, new_new_n15274__, new_new_n15275__,
    new_new_n15276__, new_new_n15277__, new_new_n15278__, new_new_n15279__,
    new_new_n15280__, new_new_n15281__, new_new_n15282__, new_new_n15283__,
    new_new_n15284__, new_new_n15285__, new_new_n15286__, new_new_n15287__,
    new_new_n15288__, new_new_n15289__, new_new_n15290__, new_new_n15291__,
    new_new_n15292__, new_new_n15293__, new_new_n15294__, new_new_n15295__,
    new_new_n15296__, new_new_n15297__, new_new_n15298__, new_new_n15299__,
    new_new_n15300__, new_new_n15301__, new_new_n15302__, new_new_n15303__,
    new_new_n15304__, new_new_n15305__, new_new_n15306__, new_new_n15307__,
    new_new_n15308__, new_new_n15309__, new_new_n15310__, new_new_n15311__,
    new_new_n15312__, new_new_n15313__, new_new_n15314__, new_new_n15316__,
    new_new_n15317__, new_new_n15318__, new_new_n15319__, new_new_n15320__,
    new_new_n15321__, new_new_n15322__, new_new_n15323__, new_new_n15324__,
    new_new_n15325__, new_new_n15326__, new_new_n15327__, new_new_n15328__,
    new_new_n15329__, new_new_n15330__, new_new_n15331__, new_new_n15332__,
    new_new_n15333__, new_new_n15334__, new_new_n15335__, new_new_n15336__,
    new_new_n15337__, new_new_n15338__, new_new_n15339__, new_new_n15340__,
    new_new_n15341__, new_new_n15342__, new_new_n15343__, new_new_n15344__,
    new_new_n15345__, new_new_n15346__, new_new_n15347__, new_new_n15348__,
    new_new_n15349__, new_new_n15350__, new_new_n15351__, new_new_n15352__,
    new_new_n15353__, new_new_n15354__, new_new_n15355__, new_new_n15356__,
    new_new_n15357__, new_new_n15358__, new_new_n15359__, new_new_n15360__,
    new_new_n15361__, new_new_n15362__, new_new_n15363__, new_new_n15364__,
    new_new_n15365__, new_new_n15366__, new_new_n15367__, new_new_n15368__,
    new_new_n15369__, new_new_n15370__, new_new_n15371__, new_new_n15372__,
    new_new_n15373__, new_new_n15374__, new_new_n15375__, new_new_n15376__,
    new_new_n15377__, new_new_n15378__, new_new_n15379__, new_new_n15380__,
    new_new_n15381__, new_new_n15382__, new_new_n15383__, new_new_n15384__,
    new_new_n15385__, new_new_n15386__, new_new_n15387__, new_new_n15388__,
    new_new_n15389__, new_new_n15390__, new_new_n15391__, new_new_n15392__,
    new_new_n15393__, new_new_n15394__, new_new_n15395__, new_new_n15396__,
    new_new_n15397__, new_new_n15398__, new_new_n15399__, new_new_n15400__,
    new_new_n15401__, new_new_n15402__, new_new_n15403__, new_new_n15404__,
    new_new_n15405__, new_new_n15406__, new_new_n15407__, new_new_n15408__,
    new_new_n15409__, new_new_n15410__, new_new_n15411__, new_new_n15412__,
    new_new_n15413__, new_new_n15414__, new_new_n15415__, new_new_n15416__,
    new_new_n15417__, new_new_n15418__, new_new_n15419__, new_new_n15420__,
    new_new_n15421__, new_new_n15422__, new_new_n15423__, new_new_n15424__,
    new_new_n15425__, new_new_n15426__, new_new_n15427__, new_new_n15428__,
    new_new_n15429__, new_new_n15430__, new_new_n15431__, new_new_n15432__,
    new_new_n15433__, new_new_n15434__, new_new_n15435__, new_new_n15436__,
    new_new_n15437__, new_new_n15438__, new_new_n15439__, new_new_n15440__,
    new_new_n15441__, new_new_n15442__, new_new_n15443__, new_new_n15444__,
    new_new_n15445__, new_new_n15446__, new_new_n15447__, new_new_n15448__,
    new_new_n15449__, new_new_n15450__, new_new_n15451__, new_new_n15452__,
    new_new_n15453__, new_new_n15454__, new_new_n15455__, new_new_n15456__,
    new_new_n15457__, new_new_n15458__, new_new_n15459__, new_new_n15460__,
    new_new_n15461__, new_new_n15462__, new_new_n15463__, new_new_n15464__,
    new_new_n15465__, new_new_n15466__, new_new_n15467__, new_new_n15468__,
    new_new_n15469__, new_new_n15470__, new_new_n15471__, new_new_n15472__,
    new_new_n15473__, new_new_n15474__, new_new_n15475__, new_new_n15476__,
    new_new_n15477__, new_new_n15478__, new_new_n15479__, new_new_n15480__,
    new_new_n15481__, new_new_n15482__, new_new_n15483__, new_new_n15484__,
    new_new_n15485__, new_new_n15486__, new_new_n15487__, new_new_n15488__,
    new_new_n15489__, new_new_n15490__, new_new_n15491__, new_new_n15492__,
    new_new_n15493__, new_new_n15494__, new_new_n15495__, new_new_n15496__,
    new_new_n15497__, new_new_n15498__, new_new_n15499__, new_new_n15500__,
    new_new_n15501__, new_new_n15502__, new_new_n15503__, new_new_n15504__,
    new_new_n15505__, new_new_n15506__, new_new_n15507__, new_new_n15508__,
    new_new_n15509__, new_new_n15510__, new_new_n15511__, new_new_n15512__,
    new_new_n15514__, new_new_n15515__, new_new_n15516__, new_new_n15517__,
    new_new_n15518__, new_new_n15519__, new_new_n15520__, new_new_n15521__,
    new_new_n15522__, new_new_n15523__, new_new_n15524__, new_new_n15525__,
    new_new_n15526__, new_new_n15527__, new_new_n15528__, new_new_n15529__,
    new_new_n15530__, new_new_n15531__, new_new_n15532__, new_new_n15533__,
    new_new_n15534__, new_new_n15535__, new_new_n15536__, new_new_n15537__,
    new_new_n15538__, new_new_n15539__, new_new_n15540__, new_new_n15541__,
    new_new_n15542__, new_new_n15543__, new_new_n15544__, new_new_n15545__,
    new_new_n15546__, new_new_n15547__, new_new_n15548__, new_new_n15549__,
    new_new_n15550__, new_new_n15551__, new_new_n15552__, new_new_n15553__,
    new_new_n15554__, new_new_n15555__, new_new_n15556__, new_new_n15557__,
    new_new_n15558__, new_new_n15559__, new_new_n15560__, new_new_n15561__,
    new_new_n15562__, new_new_n15563__, new_new_n15564__, new_new_n15565__,
    new_new_n15566__, new_new_n15567__, new_new_n15568__, new_new_n15569__,
    new_new_n15570__, new_new_n15571__, new_new_n15572__, new_new_n15573__,
    new_new_n15574__, new_new_n15575__, new_new_n15576__, new_new_n15577__,
    new_new_n15578__, new_new_n15579__, new_new_n15580__, new_new_n15581__,
    new_new_n15582__, new_new_n15583__, new_new_n15584__, new_new_n15585__,
    new_new_n15586__, new_new_n15587__, new_new_n15588__, new_new_n15589__,
    new_new_n15590__, new_new_n15591__, new_new_n15592__, new_new_n15593__,
    new_new_n15594__, new_new_n15595__, new_new_n15596__, new_new_n15597__,
    new_new_n15598__, new_new_n15599__, new_new_n15600__, new_new_n15601__,
    new_new_n15602__, new_new_n15603__, new_new_n15604__, new_new_n15605__,
    new_new_n15606__, new_new_n15607__, new_new_n15608__, new_new_n15609__,
    new_new_n15610__, new_new_n15611__, new_new_n15612__, new_new_n15613__,
    new_new_n15614__, new_new_n15615__, new_new_n15616__, new_new_n15617__,
    new_new_n15618__, new_new_n15619__, new_new_n15620__, new_new_n15621__,
    new_new_n15622__, new_new_n15623__, new_new_n15624__, new_new_n15625__,
    new_new_n15626__, new_new_n15627__, new_new_n15628__, new_new_n15629__,
    new_new_n15630__, new_new_n15631__, new_new_n15632__, new_new_n15633__,
    new_new_n15634__, new_new_n15635__, new_new_n15636__, new_new_n15637__,
    new_new_n15638__, new_new_n15639__, new_new_n15640__, new_new_n15641__,
    new_new_n15642__, new_new_n15643__, new_new_n15644__, new_new_n15645__,
    new_new_n15646__, new_new_n15647__, new_new_n15648__, new_new_n15649__,
    new_new_n15650__, new_new_n15651__, new_new_n15652__, new_new_n15653__,
    new_new_n15654__, new_new_n15655__, new_new_n15656__, new_new_n15657__,
    new_new_n15658__, new_new_n15659__, new_new_n15660__, new_new_n15661__,
    new_new_n15662__, new_new_n15663__, new_new_n15664__, new_new_n15665__,
    new_new_n15666__, new_new_n15667__, new_new_n15668__, new_new_n15669__,
    new_new_n15670__, new_new_n15671__, new_new_n15672__, new_new_n15673__,
    new_new_n15674__, new_new_n15675__, new_new_n15676__, new_new_n15677__,
    new_new_n15678__, new_new_n15679__, new_new_n15680__, new_new_n15681__,
    new_new_n15682__, new_new_n15683__, new_new_n15684__, new_new_n15685__,
    new_new_n15686__, new_new_n15687__, new_new_n15688__, new_new_n15689__,
    new_new_n15690__, new_new_n15691__, new_new_n15692__, new_new_n15693__,
    new_new_n15694__, new_new_n15695__, new_new_n15696__, new_new_n15697__,
    new_new_n15698__, new_new_n15699__, new_new_n15700__, new_new_n15701__,
    new_new_n15703__, new_new_n15704__, new_new_n15705__, new_new_n15706__,
    new_new_n15707__, new_new_n15708__, new_new_n15709__, new_new_n15710__,
    new_new_n15711__, new_new_n15712__, new_new_n15713__, new_new_n15714__,
    new_new_n15715__, new_new_n15716__, new_new_n15717__, new_new_n15718__,
    new_new_n15719__, new_new_n15720__, new_new_n15721__, new_new_n15722__,
    new_new_n15723__, new_new_n15724__, new_new_n15725__, new_new_n15726__,
    new_new_n15727__, new_new_n15728__, new_new_n15729__, new_new_n15730__,
    new_new_n15731__, new_new_n15732__, new_new_n15733__, new_new_n15734__,
    new_new_n15735__, new_new_n15736__, new_new_n15737__, new_new_n15738__,
    new_new_n15739__, new_new_n15740__, new_new_n15741__, new_new_n15742__,
    new_new_n15743__, new_new_n15744__, new_new_n15745__, new_new_n15746__,
    new_new_n15747__, new_new_n15748__, new_new_n15749__, new_new_n15750__,
    new_new_n15751__, new_new_n15752__, new_new_n15753__, new_new_n15754__,
    new_new_n15755__, new_new_n15756__, new_new_n15757__, new_new_n15758__,
    new_new_n15759__, new_new_n15760__, new_new_n15761__, new_new_n15762__,
    new_new_n15763__, new_new_n15764__, new_new_n15765__, new_new_n15766__,
    new_new_n15767__, new_new_n15768__, new_new_n15769__, new_new_n15770__,
    new_new_n15771__, new_new_n15772__, new_new_n15773__, new_new_n15774__,
    new_new_n15775__, new_new_n15776__, new_new_n15777__, new_new_n15778__,
    new_new_n15779__, new_new_n15780__, new_new_n15781__, new_new_n15782__,
    new_new_n15783__, new_new_n15784__, new_new_n15785__, new_new_n15786__,
    new_new_n15787__, new_new_n15788__, new_new_n15789__, new_new_n15790__,
    new_new_n15791__, new_new_n15792__, new_new_n15793__, new_new_n15794__,
    new_new_n15795__, new_new_n15796__, new_new_n15797__, new_new_n15798__,
    new_new_n15799__, new_new_n15800__, new_new_n15801__, new_new_n15802__,
    new_new_n15803__, new_new_n15804__, new_new_n15805__, new_new_n15806__,
    new_new_n15807__, new_new_n15808__, new_new_n15809__, new_new_n15810__,
    new_new_n15811__, new_new_n15812__, new_new_n15813__, new_new_n15814__,
    new_new_n15815__, new_new_n15816__, new_new_n15817__, new_new_n15818__,
    new_new_n15819__, new_new_n15820__, new_new_n15821__, new_new_n15822__,
    new_new_n15823__, new_new_n15824__, new_new_n15825__, new_new_n15826__,
    new_new_n15827__, new_new_n15828__, new_new_n15829__, new_new_n15830__,
    new_new_n15831__, new_new_n15832__, new_new_n15833__, new_new_n15834__,
    new_new_n15835__, new_new_n15836__, new_new_n15837__, new_new_n15838__,
    new_new_n15839__, new_new_n15840__, new_new_n15841__, new_new_n15842__,
    new_new_n15843__, new_new_n15844__, new_new_n15845__, new_new_n15846__,
    new_new_n15847__, new_new_n15848__, new_new_n15849__, new_new_n15850__,
    new_new_n15851__, new_new_n15852__, new_new_n15853__, new_new_n15854__,
    new_new_n15855__, new_new_n15856__, new_new_n15857__, new_new_n15858__,
    new_new_n15859__, new_new_n15860__, new_new_n15861__, new_new_n15862__,
    new_new_n15863__, new_new_n15864__, new_new_n15865__, new_new_n15866__,
    new_new_n15867__, new_new_n15868__, new_new_n15869__, new_new_n15870__,
    new_new_n15871__, new_new_n15872__, new_new_n15873__, new_new_n15874__,
    new_new_n15875__, new_new_n15876__, new_new_n15877__, new_new_n15878__,
    new_new_n15879__, new_new_n15880__, new_new_n15881__, new_new_n15882__,
    new_new_n15883__, new_new_n15884__, new_new_n15885__, new_new_n15886__,
    new_new_n15887__, new_new_n15888__, new_new_n15889__, new_new_n15890__,
    new_new_n15891__, new_new_n15892__, new_new_n15893__, new_new_n15894__,
    new_new_n15895__, new_new_n15896__, new_new_n15897__, new_new_n15898__,
    new_new_n15899__, new_new_n15900__, new_new_n15901__, new_new_n15902__,
    new_new_n15903__, new_new_n15904__, new_new_n15905__, new_new_n15906__,
    new_new_n15907__, new_new_n15908__, new_new_n15909__, new_new_n15910__,
    new_new_n15911__, new_new_n15912__, new_new_n15913__, new_new_n15914__,
    new_new_n15916__, new_new_n15917__, new_new_n15918__, new_new_n15919__,
    new_new_n15920__, new_new_n15921__, new_new_n15922__, new_new_n15923__,
    new_new_n15924__, new_new_n15925__, new_new_n15926__, new_new_n15927__,
    new_new_n15928__, new_new_n15929__, new_new_n15930__, new_new_n15931__,
    new_new_n15932__, new_new_n15933__, new_new_n15934__, new_new_n15935__,
    new_new_n15936__, new_new_n15937__, new_new_n15938__, new_new_n15939__,
    new_new_n15940__, new_new_n15941__, new_new_n15942__, new_new_n15943__,
    new_new_n15944__, new_new_n15945__, new_new_n15946__, new_new_n15947__,
    new_new_n15948__, new_new_n15949__, new_new_n15950__, new_new_n15951__,
    new_new_n15952__, new_new_n15953__, new_new_n15954__, new_new_n15955__,
    new_new_n15956__, new_new_n15957__, new_new_n15958__, new_new_n15959__,
    new_new_n15960__, new_new_n15961__, new_new_n15962__, new_new_n15963__,
    new_new_n15964__, new_new_n15965__, new_new_n15966__, new_new_n15967__,
    new_new_n15968__, new_new_n15969__, new_new_n15970__, new_new_n15971__,
    new_new_n15972__, new_new_n15973__, new_new_n15974__, new_new_n15975__,
    new_new_n15976__, new_new_n15977__, new_new_n15978__, new_new_n15979__,
    new_new_n15980__, new_new_n15981__, new_new_n15982__, new_new_n15983__,
    new_new_n15984__, new_new_n15985__, new_new_n15986__, new_new_n15987__,
    new_new_n15988__, new_new_n15989__, new_new_n15990__, new_new_n15991__,
    new_new_n15992__, new_new_n15993__, new_new_n15994__, new_new_n15995__,
    new_new_n15996__, new_new_n15997__, new_new_n15998__, new_new_n15999__,
    new_new_n16000__, new_new_n16001__, new_new_n16002__, new_new_n16003__,
    new_new_n16004__, new_new_n16005__, new_new_n16006__, new_new_n16007__,
    new_new_n16008__, new_new_n16009__, new_new_n16010__, new_new_n16011__,
    new_new_n16012__, new_new_n16013__, new_new_n16014__, new_new_n16015__,
    new_new_n16016__, new_new_n16017__, new_new_n16018__, new_new_n16019__,
    new_new_n16020__, new_new_n16021__, new_new_n16022__, new_new_n16023__,
    new_new_n16024__, new_new_n16025__, new_new_n16026__, new_new_n16027__,
    new_new_n16028__, new_new_n16029__, new_new_n16030__, new_new_n16031__,
    new_new_n16032__, new_new_n16033__, new_new_n16034__, new_new_n16035__,
    new_new_n16036__, new_new_n16037__, new_new_n16038__, new_new_n16039__,
    new_new_n16040__, new_new_n16041__, new_new_n16042__, new_new_n16043__,
    new_new_n16044__, new_new_n16045__, new_new_n16046__, new_new_n16047__,
    new_new_n16048__, new_new_n16049__, new_new_n16050__, new_new_n16051__,
    new_new_n16052__, new_new_n16053__, new_new_n16054__, new_new_n16055__,
    new_new_n16056__, new_new_n16057__, new_new_n16058__, new_new_n16059__,
    new_new_n16060__, new_new_n16061__, new_new_n16062__, new_new_n16063__,
    new_new_n16064__, new_new_n16065__, new_new_n16066__, new_new_n16067__,
    new_new_n16068__, new_new_n16069__, new_new_n16070__, new_new_n16071__,
    new_new_n16072__, new_new_n16073__, new_new_n16074__, new_new_n16075__,
    new_new_n16076__, new_new_n16077__, new_new_n16078__, new_new_n16079__,
    new_new_n16080__, new_new_n16081__, new_new_n16082__, new_new_n16083__,
    new_new_n16084__, new_new_n16085__, new_new_n16086__, new_new_n16087__,
    new_new_n16088__, new_new_n16089__, new_new_n16090__, new_new_n16091__,
    new_new_n16092__, new_new_n16093__, new_new_n16094__, new_new_n16095__,
    new_new_n16096__, new_new_n16097__, new_new_n16098__, new_new_n16099__,
    new_new_n16100__, new_new_n16101__, new_new_n16102__, new_new_n16103__,
    new_new_n16104__, new_new_n16105__, new_new_n16106__, new_new_n16107__,
    new_new_n16108__, new_new_n16109__, new_new_n16110__, new_new_n16111__,
    new_new_n16112__, new_new_n16113__, new_new_n16114__, new_new_n16115__,
    new_new_n16116__, new_new_n16117__, new_new_n16118__, new_new_n16119__,
    new_new_n16120__, new_new_n16121__, new_new_n16122__, new_new_n16123__,
    new_new_n16124__, new_new_n16125__, new_new_n16126__, new_new_n16127__,
    new_new_n16128__, new_new_n16129__, new_new_n16130__, new_new_n16131__,
    new_new_n16132__, new_new_n16133__, new_new_n16134__, new_new_n16136__,
    new_new_n16137__, new_new_n16138__, new_new_n16139__, new_new_n16140__,
    new_new_n16141__, new_new_n16142__, new_new_n16143__, new_new_n16144__,
    new_new_n16145__, new_new_n16146__, new_new_n16147__, new_new_n16148__,
    new_new_n16149__, new_new_n16150__, new_new_n16151__, new_new_n16152__,
    new_new_n16153__, new_new_n16154__, new_new_n16155__, new_new_n16156__,
    new_new_n16157__, new_new_n16158__, new_new_n16159__, new_new_n16160__,
    new_new_n16161__, new_new_n16162__, new_new_n16163__, new_new_n16164__,
    new_new_n16165__, new_new_n16166__, new_new_n16167__, new_new_n16168__,
    new_new_n16169__, new_new_n16170__, new_new_n16171__, new_new_n16172__,
    new_new_n16173__, new_new_n16174__, new_new_n16175__, new_new_n16176__,
    new_new_n16177__, new_new_n16178__, new_new_n16179__, new_new_n16180__,
    new_new_n16181__, new_new_n16182__, new_new_n16183__, new_new_n16184__,
    new_new_n16185__, new_new_n16186__, new_new_n16187__, new_new_n16188__,
    new_new_n16189__, new_new_n16190__, new_new_n16191__, new_new_n16192__,
    new_new_n16193__, new_new_n16194__, new_new_n16195__, new_new_n16196__,
    new_new_n16197__, new_new_n16198__, new_new_n16199__, new_new_n16200__,
    new_new_n16201__, new_new_n16202__, new_new_n16203__, new_new_n16204__,
    new_new_n16205__, new_new_n16206__, new_new_n16207__, new_new_n16208__,
    new_new_n16209__, new_new_n16210__, new_new_n16211__, new_new_n16212__,
    new_new_n16213__, new_new_n16214__, new_new_n16215__, new_new_n16216__,
    new_new_n16217__, new_new_n16218__, new_new_n16219__, new_new_n16220__,
    new_new_n16221__, new_new_n16222__, new_new_n16223__, new_new_n16224__,
    new_new_n16225__, new_new_n16226__, new_new_n16227__, new_new_n16228__,
    new_new_n16229__, new_new_n16230__, new_new_n16231__, new_new_n16232__,
    new_new_n16233__, new_new_n16234__, new_new_n16235__, new_new_n16236__,
    new_new_n16237__, new_new_n16238__, new_new_n16239__, new_new_n16240__,
    new_new_n16241__, new_new_n16242__, new_new_n16243__, new_new_n16244__,
    new_new_n16245__, new_new_n16246__, new_new_n16247__, new_new_n16248__,
    new_new_n16249__, new_new_n16250__, new_new_n16251__, new_new_n16252__,
    new_new_n16253__, new_new_n16254__, new_new_n16255__, new_new_n16256__,
    new_new_n16257__, new_new_n16258__, new_new_n16259__, new_new_n16260__,
    new_new_n16261__, new_new_n16262__, new_new_n16263__, new_new_n16264__,
    new_new_n16265__, new_new_n16266__, new_new_n16267__, new_new_n16268__,
    new_new_n16269__, new_new_n16270__, new_new_n16271__, new_new_n16272__,
    new_new_n16273__, new_new_n16274__, new_new_n16275__, new_new_n16276__,
    new_new_n16277__, new_new_n16278__, new_new_n16279__, new_new_n16280__,
    new_new_n16281__, new_new_n16282__, new_new_n16283__, new_new_n16284__,
    new_new_n16285__, new_new_n16286__, new_new_n16287__, new_new_n16288__,
    new_new_n16289__, new_new_n16290__, new_new_n16291__, new_new_n16292__,
    new_new_n16293__, new_new_n16294__, new_new_n16295__, new_new_n16296__,
    new_new_n16297__, new_new_n16298__, new_new_n16299__, new_new_n16300__,
    new_new_n16301__, new_new_n16302__, new_new_n16303__, new_new_n16304__,
    new_new_n16305__, new_new_n16306__, new_new_n16307__, new_new_n16308__,
    new_new_n16309__, new_new_n16310__, new_new_n16311__, new_new_n16312__,
    new_new_n16313__, new_new_n16314__, new_new_n16315__, new_new_n16316__,
    new_new_n16317__, new_new_n16318__, new_new_n16319__, new_new_n16320__,
    new_new_n16321__, new_new_n16322__, new_new_n16323__, new_new_n16324__,
    new_new_n16325__, new_new_n16326__, new_new_n16327__, new_new_n16328__,
    new_new_n16329__, new_new_n16330__, new_new_n16331__, new_new_n16332__,
    new_new_n16333__, new_new_n16334__, new_new_n16336__, new_new_n16337__,
    new_new_n16338__, new_new_n16339__, new_new_n16340__, new_new_n16341__,
    new_new_n16342__, new_new_n16343__, new_new_n16344__, new_new_n16345__,
    new_new_n16346__, new_new_n16347__, new_new_n16348__, new_new_n16349__,
    new_new_n16350__, new_new_n16351__, new_new_n16352__, new_new_n16353__,
    new_new_n16354__, new_new_n16355__, new_new_n16356__, new_new_n16357__,
    new_new_n16358__, new_new_n16359__, new_new_n16360__, new_new_n16361__,
    new_new_n16362__, new_new_n16363__, new_new_n16364__, new_new_n16365__,
    new_new_n16366__, new_new_n16367__, new_new_n16368__, new_new_n16369__,
    new_new_n16370__, new_new_n16371__, new_new_n16372__, new_new_n16373__,
    new_new_n16374__, new_new_n16375__, new_new_n16376__, new_new_n16377__,
    new_new_n16378__, new_new_n16379__, new_new_n16380__, new_new_n16381__,
    new_new_n16382__, new_new_n16383__, new_new_n16384__, new_new_n16385__,
    new_new_n16386__, new_new_n16387__, new_new_n16388__, new_new_n16389__,
    new_new_n16390__, new_new_n16391__, new_new_n16392__, new_new_n16393__,
    new_new_n16394__, new_new_n16395__, new_new_n16396__, new_new_n16397__,
    new_new_n16398__, new_new_n16399__, new_new_n16400__, new_new_n16401__,
    new_new_n16402__, new_new_n16403__, new_new_n16404__, new_new_n16405__,
    new_new_n16406__, new_new_n16407__, new_new_n16408__, new_new_n16409__,
    new_new_n16410__, new_new_n16411__, new_new_n16412__, new_new_n16413__,
    new_new_n16414__, new_new_n16415__, new_new_n16416__, new_new_n16417__,
    new_new_n16418__, new_new_n16419__, new_new_n16420__, new_new_n16421__,
    new_new_n16422__, new_new_n16423__, new_new_n16424__, new_new_n16425__,
    new_new_n16426__, new_new_n16427__, new_new_n16428__, new_new_n16429__,
    new_new_n16430__, new_new_n16431__, new_new_n16432__, new_new_n16433__,
    new_new_n16434__, new_new_n16435__, new_new_n16436__, new_new_n16437__,
    new_new_n16438__, new_new_n16439__, new_new_n16440__, new_new_n16441__,
    new_new_n16442__, new_new_n16443__, new_new_n16444__, new_new_n16445__,
    new_new_n16446__, new_new_n16447__, new_new_n16448__, new_new_n16449__,
    new_new_n16450__, new_new_n16451__, new_new_n16452__, new_new_n16453__,
    new_new_n16454__, new_new_n16455__, new_new_n16456__, new_new_n16457__,
    new_new_n16458__, new_new_n16459__, new_new_n16460__, new_new_n16461__,
    new_new_n16462__, new_new_n16463__, new_new_n16464__, new_new_n16465__,
    new_new_n16466__, new_new_n16467__, new_new_n16468__, new_new_n16469__,
    new_new_n16470__, new_new_n16471__, new_new_n16472__, new_new_n16473__,
    new_new_n16474__, new_new_n16475__, new_new_n16476__, new_new_n16477__,
    new_new_n16478__, new_new_n16479__, new_new_n16480__, new_new_n16481__,
    new_new_n16482__, new_new_n16483__, new_new_n16484__, new_new_n16485__,
    new_new_n16486__, new_new_n16487__, new_new_n16488__, new_new_n16489__,
    new_new_n16490__, new_new_n16491__, new_new_n16492__, new_new_n16493__,
    new_new_n16494__, new_new_n16495__, new_new_n16496__, new_new_n16497__,
    new_new_n16498__, new_new_n16499__, new_new_n16500__, new_new_n16501__,
    new_new_n16502__, new_new_n16503__, new_new_n16504__, new_new_n16505__,
    new_new_n16506__, new_new_n16507__, new_new_n16508__, new_new_n16509__,
    new_new_n16510__, new_new_n16511__, new_new_n16513__, new_new_n16514__,
    new_new_n16515__, new_new_n16516__, new_new_n16517__, new_new_n16518__,
    new_new_n16519__, new_new_n16520__, new_new_n16521__, new_new_n16522__,
    new_new_n16523__, new_new_n16524__, new_new_n16525__, new_new_n16526__,
    new_new_n16527__, new_new_n16528__, new_new_n16529__, new_new_n16530__,
    new_new_n16531__, new_new_n16532__, new_new_n16533__, new_new_n16534__,
    new_new_n16535__, new_new_n16536__, new_new_n16537__, new_new_n16538__,
    new_new_n16539__, new_new_n16540__, new_new_n16541__, new_new_n16542__,
    new_new_n16543__, new_new_n16544__, new_new_n16545__, new_new_n16546__,
    new_new_n16547__, new_new_n16548__, new_new_n16549__, new_new_n16550__,
    new_new_n16551__, new_new_n16552__, new_new_n16553__, new_new_n16554__,
    new_new_n16555__, new_new_n16556__, new_new_n16557__, new_new_n16558__,
    new_new_n16559__, new_new_n16560__, new_new_n16561__, new_new_n16562__,
    new_new_n16563__, new_new_n16564__, new_new_n16565__, new_new_n16566__,
    new_new_n16567__, new_new_n16568__, new_new_n16569__, new_new_n16570__,
    new_new_n16571__, new_new_n16572__, new_new_n16573__, new_new_n16574__,
    new_new_n16575__, new_new_n16576__, new_new_n16577__, new_new_n16578__,
    new_new_n16579__, new_new_n16580__, new_new_n16581__, new_new_n16582__,
    new_new_n16583__, new_new_n16584__, new_new_n16585__, new_new_n16586__,
    new_new_n16587__, new_new_n16588__, new_new_n16589__, new_new_n16590__,
    new_new_n16591__, new_new_n16592__, new_new_n16593__, new_new_n16594__,
    new_new_n16595__, new_new_n16596__, new_new_n16597__, new_new_n16598__,
    new_new_n16599__, new_new_n16600__, new_new_n16601__, new_new_n16602__,
    new_new_n16603__, new_new_n16604__, new_new_n16605__, new_new_n16606__,
    new_new_n16607__, new_new_n16608__, new_new_n16609__, new_new_n16610__,
    new_new_n16611__, new_new_n16612__, new_new_n16613__, new_new_n16614__,
    new_new_n16615__, new_new_n16616__, new_new_n16617__, new_new_n16618__,
    new_new_n16619__, new_new_n16620__, new_new_n16621__, new_new_n16622__,
    new_new_n16623__, new_new_n16624__, new_new_n16625__, new_new_n16626__,
    new_new_n16627__, new_new_n16628__, new_new_n16629__, new_new_n16630__,
    new_new_n16631__, new_new_n16632__, new_new_n16633__, new_new_n16634__,
    new_new_n16635__, new_new_n16636__, new_new_n16637__, new_new_n16638__,
    new_new_n16639__, new_new_n16640__, new_new_n16641__, new_new_n16642__,
    new_new_n16643__, new_new_n16644__, new_new_n16645__, new_new_n16646__,
    new_new_n16647__, new_new_n16648__, new_new_n16649__, new_new_n16650__,
    new_new_n16651__, new_new_n16652__, new_new_n16653__, new_new_n16654__,
    new_new_n16655__, new_new_n16656__, new_new_n16657__, new_new_n16658__,
    new_new_n16659__, new_new_n16660__, new_new_n16661__, new_new_n16662__,
    new_new_n16663__, new_new_n16664__, new_new_n16665__, new_new_n16666__,
    new_new_n16667__, new_new_n16668__, new_new_n16669__, new_new_n16670__,
    new_new_n16671__, new_new_n16672__, new_new_n16673__, new_new_n16674__,
    new_new_n16675__, new_new_n16676__, new_new_n16677__, new_new_n16678__,
    new_new_n16679__, new_new_n16680__, new_new_n16681__, new_new_n16682__,
    new_new_n16683__, new_new_n16684__, new_new_n16685__, new_new_n16686__,
    new_new_n16687__, new_new_n16689__, new_new_n16690__, new_new_n16691__,
    new_new_n16692__, new_new_n16693__, new_new_n16694__, new_new_n16695__,
    new_new_n16696__, new_new_n16697__, new_new_n16698__, new_new_n16699__,
    new_new_n16700__, new_new_n16701__, new_new_n16702__, new_new_n16703__,
    new_new_n16704__, new_new_n16705__, new_new_n16706__, new_new_n16707__,
    new_new_n16708__, new_new_n16709__, new_new_n16710__, new_new_n16711__,
    new_new_n16712__, new_new_n16713__, new_new_n16714__, new_new_n16715__,
    new_new_n16716__, new_new_n16717__, new_new_n16718__, new_new_n16719__,
    new_new_n16720__, new_new_n16721__, new_new_n16722__, new_new_n16723__,
    new_new_n16724__, new_new_n16725__, new_new_n16726__, new_new_n16727__,
    new_new_n16728__, new_new_n16729__, new_new_n16730__, new_new_n16731__,
    new_new_n16732__, new_new_n16733__, new_new_n16734__, new_new_n16735__,
    new_new_n16736__, new_new_n16737__, new_new_n16738__, new_new_n16739__,
    new_new_n16740__, new_new_n16741__, new_new_n16742__, new_new_n16743__,
    new_new_n16744__, new_new_n16745__, new_new_n16746__, new_new_n16747__,
    new_new_n16748__, new_new_n16749__, new_new_n16750__, new_new_n16751__,
    new_new_n16752__, new_new_n16753__, new_new_n16754__, new_new_n16755__,
    new_new_n16756__, new_new_n16757__, new_new_n16758__, new_new_n16759__,
    new_new_n16760__, new_new_n16761__, new_new_n16762__, new_new_n16763__,
    new_new_n16764__, new_new_n16765__, new_new_n16766__, new_new_n16767__,
    new_new_n16768__, new_new_n16769__, new_new_n16770__, new_new_n16771__,
    new_new_n16772__, new_new_n16773__, new_new_n16774__, new_new_n16775__,
    new_new_n16776__, new_new_n16777__, new_new_n16778__, new_new_n16779__,
    new_new_n16780__, new_new_n16781__, new_new_n16782__, new_new_n16783__,
    new_new_n16784__, new_new_n16785__, new_new_n16786__, new_new_n16787__,
    new_new_n16788__, new_new_n16789__, new_new_n16790__, new_new_n16791__,
    new_new_n16792__, new_new_n16793__, new_new_n16794__, new_new_n16795__,
    new_new_n16796__, new_new_n16797__, new_new_n16798__, new_new_n16799__,
    new_new_n16800__, new_new_n16801__, new_new_n16802__, new_new_n16803__,
    new_new_n16804__, new_new_n16805__, new_new_n16806__, new_new_n16807__,
    new_new_n16808__, new_new_n16809__, new_new_n16810__, new_new_n16811__,
    new_new_n16812__, new_new_n16813__, new_new_n16814__, new_new_n16815__,
    new_new_n16816__, new_new_n16817__, new_new_n16818__, new_new_n16819__,
    new_new_n16820__, new_new_n16821__, new_new_n16822__, new_new_n16823__,
    new_new_n16824__, new_new_n16825__, new_new_n16826__, new_new_n16827__,
    new_new_n16828__, new_new_n16829__, new_new_n16830__, new_new_n16831__,
    new_new_n16832__, new_new_n16833__, new_new_n16834__, new_new_n16835__,
    new_new_n16836__, new_new_n16837__, new_new_n16838__, new_new_n16839__,
    new_new_n16840__, new_new_n16841__, new_new_n16842__, new_new_n16843__,
    new_new_n16844__, new_new_n16845__, new_new_n16846__, new_new_n16847__,
    new_new_n16848__, new_new_n16849__, new_new_n16850__, new_new_n16851__,
    new_new_n16852__, new_new_n16853__, new_new_n16854__, new_new_n16855__,
    new_new_n16857__, new_new_n16858__, new_new_n16859__, new_new_n16860__,
    new_new_n16861__, new_new_n16862__, new_new_n16863__, new_new_n16864__,
    new_new_n16865__, new_new_n16866__, new_new_n16867__, new_new_n16868__,
    new_new_n16869__, new_new_n16870__, new_new_n16871__, new_new_n16872__,
    new_new_n16873__, new_new_n16874__, new_new_n16875__, new_new_n16876__,
    new_new_n16877__, new_new_n16878__, new_new_n16879__, new_new_n16880__,
    new_new_n16881__, new_new_n16882__, new_new_n16883__, new_new_n16884__,
    new_new_n16885__, new_new_n16886__, new_new_n16887__, new_new_n16888__,
    new_new_n16889__, new_new_n16890__, new_new_n16891__, new_new_n16892__,
    new_new_n16893__, new_new_n16894__, new_new_n16895__, new_new_n16896__,
    new_new_n16897__, new_new_n16898__, new_new_n16899__, new_new_n16900__,
    new_new_n16901__, new_new_n16902__, new_new_n16903__, new_new_n16904__,
    new_new_n16905__, new_new_n16906__, new_new_n16907__, new_new_n16908__,
    new_new_n16909__, new_new_n16910__, new_new_n16911__, new_new_n16912__,
    new_new_n16913__, new_new_n16914__, new_new_n16915__, new_new_n16916__,
    new_new_n16917__, new_new_n16918__, new_new_n16919__, new_new_n16920__,
    new_new_n16921__, new_new_n16922__, new_new_n16923__, new_new_n16924__,
    new_new_n16925__, new_new_n16926__, new_new_n16927__, new_new_n16928__,
    new_new_n16929__, new_new_n16930__, new_new_n16931__, new_new_n16932__,
    new_new_n16933__, new_new_n16934__, new_new_n16935__, new_new_n16936__,
    new_new_n16937__, new_new_n16938__, new_new_n16939__, new_new_n16940__,
    new_new_n16941__, new_new_n16942__, new_new_n16943__, new_new_n16944__,
    new_new_n16945__, new_new_n16946__, new_new_n16947__, new_new_n16948__,
    new_new_n16949__, new_new_n16950__, new_new_n16951__, new_new_n16952__,
    new_new_n16953__, new_new_n16954__, new_new_n16955__, new_new_n16956__,
    new_new_n16957__, new_new_n16958__, new_new_n16959__, new_new_n16960__,
    new_new_n16961__, new_new_n16962__, new_new_n16963__, new_new_n16964__,
    new_new_n16965__, new_new_n16966__, new_new_n16967__, new_new_n16968__,
    new_new_n16969__, new_new_n16970__, new_new_n16971__, new_new_n16972__,
    new_new_n16973__, new_new_n16974__, new_new_n16975__, new_new_n16976__,
    new_new_n16977__, new_new_n16978__, new_new_n16979__, new_new_n16980__,
    new_new_n16981__, new_new_n16982__, new_new_n16983__, new_new_n16984__,
    new_new_n16985__, new_new_n16986__, new_new_n16987__, new_new_n16988__,
    new_new_n16989__, new_new_n16990__, new_new_n16991__, new_new_n16992__,
    new_new_n16993__, new_new_n16994__, new_new_n16995__, new_new_n16996__,
    new_new_n16997__, new_new_n16998__, new_new_n16999__, new_new_n17000__,
    new_new_n17001__, new_new_n17002__, new_new_n17003__, new_new_n17004__,
    new_new_n17005__, new_new_n17006__, new_new_n17007__, new_new_n17008__,
    new_new_n17009__, new_new_n17010__, new_new_n17011__, new_new_n17012__,
    new_new_n17013__, new_new_n17014__, new_new_n17015__, new_new_n17016__,
    new_new_n17017__, new_new_n17018__, new_new_n17019__, new_new_n17020__,
    new_new_n17021__, new_new_n17022__, new_new_n17023__, new_new_n17024__,
    new_new_n17025__, new_new_n17026__, new_new_n17027__, new_new_n17028__,
    new_new_n17029__, new_new_n17030__, new_new_n17031__, new_new_n17032__,
    new_new_n17033__, new_new_n17034__, new_new_n17035__, new_new_n17036__,
    new_new_n17037__, new_new_n17038__, new_new_n17040__, new_new_n17041__,
    new_new_n17042__, new_new_n17043__, new_new_n17044__, new_new_n17045__,
    new_new_n17046__, new_new_n17047__, new_new_n17048__, new_new_n17049__,
    new_new_n17050__, new_new_n17051__, new_new_n17052__, new_new_n17053__,
    new_new_n17054__, new_new_n17055__, new_new_n17056__, new_new_n17057__,
    new_new_n17058__, new_new_n17059__, new_new_n17060__, new_new_n17061__,
    new_new_n17062__, new_new_n17063__, new_new_n17064__, new_new_n17065__,
    new_new_n17066__, new_new_n17067__, new_new_n17068__, new_new_n17069__,
    new_new_n17070__, new_new_n17071__, new_new_n17072__, new_new_n17073__,
    new_new_n17074__, new_new_n17075__, new_new_n17076__, new_new_n17077__,
    new_new_n17078__, new_new_n17079__, new_new_n17080__, new_new_n17081__,
    new_new_n17082__, new_new_n17083__, new_new_n17084__, new_new_n17085__,
    new_new_n17086__, new_new_n17087__, new_new_n17088__, new_new_n17089__,
    new_new_n17090__, new_new_n17091__, new_new_n17092__, new_new_n17093__,
    new_new_n17094__, new_new_n17095__, new_new_n17096__, new_new_n17097__,
    new_new_n17098__, new_new_n17099__, new_new_n17100__, new_new_n17101__,
    new_new_n17102__, new_new_n17103__, new_new_n17104__, new_new_n17105__,
    new_new_n17106__, new_new_n17107__, new_new_n17108__, new_new_n17109__,
    new_new_n17110__, new_new_n17111__, new_new_n17112__, new_new_n17113__,
    new_new_n17114__, new_new_n17115__, new_new_n17116__, new_new_n17117__,
    new_new_n17118__, new_new_n17119__, new_new_n17120__, new_new_n17121__,
    new_new_n17122__, new_new_n17123__, new_new_n17124__, new_new_n17125__,
    new_new_n17126__, new_new_n17127__, new_new_n17128__, new_new_n17129__,
    new_new_n17130__, new_new_n17131__, new_new_n17132__, new_new_n17133__,
    new_new_n17134__, new_new_n17135__, new_new_n17136__, new_new_n17137__,
    new_new_n17138__, new_new_n17139__, new_new_n17140__, new_new_n17141__,
    new_new_n17142__, new_new_n17143__, new_new_n17144__, new_new_n17145__,
    new_new_n17146__, new_new_n17147__, new_new_n17148__, new_new_n17149__,
    new_new_n17150__, new_new_n17151__, new_new_n17152__, new_new_n17153__,
    new_new_n17154__, new_new_n17155__, new_new_n17156__, new_new_n17157__,
    new_new_n17158__, new_new_n17159__, new_new_n17160__, new_new_n17161__,
    new_new_n17162__, new_new_n17163__, new_new_n17164__, new_new_n17165__,
    new_new_n17166__, new_new_n17167__, new_new_n17168__, new_new_n17169__,
    new_new_n17170__, new_new_n17171__, new_new_n17172__, new_new_n17173__,
    new_new_n17174__, new_new_n17175__, new_new_n17176__, new_new_n17177__,
    new_new_n17178__, new_new_n17179__, new_new_n17180__, new_new_n17181__,
    new_new_n17182__, new_new_n17183__, new_new_n17184__, new_new_n17185__,
    new_new_n17186__, new_new_n17187__, new_new_n17188__, new_new_n17189__,
    new_new_n17190__, new_new_n17191__, new_new_n17192__, new_new_n17193__,
    new_new_n17194__, new_new_n17195__, new_new_n17197__, new_new_n17198__,
    new_new_n17199__, new_new_n17200__, new_new_n17201__, new_new_n17202__,
    new_new_n17203__, new_new_n17204__, new_new_n17205__, new_new_n17206__,
    new_new_n17207__, new_new_n17208__, new_new_n17209__, new_new_n17210__,
    new_new_n17211__, new_new_n17212__, new_new_n17213__, new_new_n17214__,
    new_new_n17215__, new_new_n17216__, new_new_n17217__, new_new_n17218__,
    new_new_n17219__, new_new_n17220__, new_new_n17221__, new_new_n17222__,
    new_new_n17223__, new_new_n17224__, new_new_n17225__, new_new_n17226__,
    new_new_n17227__, new_new_n17228__, new_new_n17229__, new_new_n17230__,
    new_new_n17231__, new_new_n17232__, new_new_n17233__, new_new_n17234__,
    new_new_n17235__, new_new_n17236__, new_new_n17237__, new_new_n17238__,
    new_new_n17239__, new_new_n17240__, new_new_n17241__, new_new_n17242__,
    new_new_n17243__, new_new_n17244__, new_new_n17245__, new_new_n17246__,
    new_new_n17247__, new_new_n17248__, new_new_n17249__, new_new_n17250__,
    new_new_n17251__, new_new_n17252__, new_new_n17253__, new_new_n17254__,
    new_new_n17255__, new_new_n17256__, new_new_n17257__, new_new_n17258__,
    new_new_n17259__, new_new_n17260__, new_new_n17261__, new_new_n17262__,
    new_new_n17263__, new_new_n17264__, new_new_n17265__, new_new_n17266__,
    new_new_n17267__, new_new_n17268__, new_new_n17269__, new_new_n17270__,
    new_new_n17271__, new_new_n17272__, new_new_n17273__, new_new_n17274__,
    new_new_n17275__, new_new_n17276__, new_new_n17277__, new_new_n17278__,
    new_new_n17279__, new_new_n17280__, new_new_n17281__, new_new_n17282__,
    new_new_n17283__, new_new_n17284__, new_new_n17285__, new_new_n17286__,
    new_new_n17287__, new_new_n17288__, new_new_n17289__, new_new_n17290__,
    new_new_n17291__, new_new_n17292__, new_new_n17293__, new_new_n17294__,
    new_new_n17295__, new_new_n17296__, new_new_n17297__, new_new_n17298__,
    new_new_n17299__, new_new_n17300__, new_new_n17301__, new_new_n17302__,
    new_new_n17303__, new_new_n17304__, new_new_n17305__, new_new_n17306__,
    new_new_n17307__, new_new_n17308__, new_new_n17309__, new_new_n17310__,
    new_new_n17311__, new_new_n17312__, new_new_n17313__, new_new_n17314__,
    new_new_n17315__, new_new_n17316__, new_new_n17317__, new_new_n17318__,
    new_new_n17319__, new_new_n17320__, new_new_n17321__, new_new_n17322__,
    new_new_n17323__, new_new_n17324__, new_new_n17325__, new_new_n17326__,
    new_new_n17327__, new_new_n17328__, new_new_n17329__, new_new_n17330__,
    new_new_n17331__, new_new_n17332__, new_new_n17333__, new_new_n17334__,
    new_new_n17335__, new_new_n17336__, new_new_n17337__, new_new_n17338__,
    new_new_n17339__, new_new_n17340__, new_new_n17341__, new_new_n17342__,
    new_new_n17343__, new_new_n17344__, new_new_n17345__, new_new_n17346__,
    new_new_n17347__, new_new_n17348__, new_new_n17349__, new_new_n17350__,
    new_new_n17351__, new_new_n17352__, new_new_n17353__, new_new_n17354__,
    new_new_n17355__, new_new_n17356__, new_new_n17357__, new_new_n17358__,
    new_new_n17359__, new_new_n17360__, new_new_n17361__, new_new_n17362__,
    new_new_n17363__, new_new_n17364__, new_new_n17365__, new_new_n17367__,
    new_new_n17368__, new_new_n17369__, new_new_n17370__, new_new_n17371__,
    new_new_n17372__, new_new_n17373__, new_new_n17374__, new_new_n17375__,
    new_new_n17376__, new_new_n17377__, new_new_n17378__, new_new_n17379__,
    new_new_n17380__, new_new_n17381__, new_new_n17382__, new_new_n17383__,
    new_new_n17384__, new_new_n17385__, new_new_n17386__, new_new_n17387__,
    new_new_n17388__, new_new_n17389__, new_new_n17390__, new_new_n17391__,
    new_new_n17392__, new_new_n17393__, new_new_n17394__, new_new_n17395__,
    new_new_n17396__, new_new_n17397__, new_new_n17398__, new_new_n17399__,
    new_new_n17400__, new_new_n17401__, new_new_n17402__, new_new_n17403__,
    new_new_n17404__, new_new_n17405__, new_new_n17406__, new_new_n17407__,
    new_new_n17408__, new_new_n17409__, new_new_n17410__, new_new_n17411__,
    new_new_n17412__, new_new_n17413__, new_new_n17414__, new_new_n17415__,
    new_new_n17416__, new_new_n17417__, new_new_n17418__, new_new_n17419__,
    new_new_n17420__, new_new_n17421__, new_new_n17422__, new_new_n17423__,
    new_new_n17424__, new_new_n17425__, new_new_n17426__, new_new_n17427__,
    new_new_n17428__, new_new_n17429__, new_new_n17430__, new_new_n17431__,
    new_new_n17432__, new_new_n17433__, new_new_n17434__, new_new_n17435__,
    new_new_n17436__, new_new_n17437__, new_new_n17438__, new_new_n17439__,
    new_new_n17440__, new_new_n17441__, new_new_n17442__, new_new_n17443__,
    new_new_n17444__, new_new_n17445__, new_new_n17446__, new_new_n17447__,
    new_new_n17448__, new_new_n17449__, new_new_n17450__, new_new_n17451__,
    new_new_n17452__, new_new_n17453__, new_new_n17454__, new_new_n17455__,
    new_new_n17456__, new_new_n17457__, new_new_n17458__, new_new_n17459__,
    new_new_n17460__, new_new_n17461__, new_new_n17462__, new_new_n17463__,
    new_new_n17464__, new_new_n17465__, new_new_n17466__, new_new_n17467__,
    new_new_n17468__, new_new_n17469__, new_new_n17470__, new_new_n17471__,
    new_new_n17472__, new_new_n17473__, new_new_n17474__, new_new_n17475__,
    new_new_n17476__, new_new_n17477__, new_new_n17478__, new_new_n17479__,
    new_new_n17480__, new_new_n17481__, new_new_n17482__, new_new_n17483__,
    new_new_n17484__, new_new_n17485__, new_new_n17486__, new_new_n17487__,
    new_new_n17488__, new_new_n17489__, new_new_n17490__, new_new_n17491__,
    new_new_n17492__, new_new_n17493__, new_new_n17494__, new_new_n17495__,
    new_new_n17496__, new_new_n17497__, new_new_n17498__, new_new_n17499__,
    new_new_n17500__, new_new_n17501__, new_new_n17502__, new_new_n17503__,
    new_new_n17504__, new_new_n17505__, new_new_n17506__, new_new_n17507__,
    new_new_n17508__, new_new_n17509__, new_new_n17510__, new_new_n17511__,
    new_new_n17512__, new_new_n17513__, new_new_n17514__, new_new_n17515__,
    new_new_n17516__, new_new_n17517__, new_new_n17518__, new_new_n17519__,
    new_new_n17520__, new_new_n17522__, new_new_n17523__, new_new_n17524__,
    new_new_n17525__, new_new_n17526__, new_new_n17527__, new_new_n17528__,
    new_new_n17529__, new_new_n17530__, new_new_n17531__, new_new_n17532__,
    new_new_n17533__, new_new_n17534__, new_new_n17535__, new_new_n17536__,
    new_new_n17537__, new_new_n17538__, new_new_n17539__, new_new_n17540__,
    new_new_n17541__, new_new_n17542__, new_new_n17543__, new_new_n17544__,
    new_new_n17545__, new_new_n17546__, new_new_n17547__, new_new_n17548__,
    new_new_n17549__, new_new_n17550__, new_new_n17551__, new_new_n17552__,
    new_new_n17553__, new_new_n17554__, new_new_n17555__, new_new_n17556__,
    new_new_n17557__, new_new_n17558__, new_new_n17559__, new_new_n17560__,
    new_new_n17561__, new_new_n17562__, new_new_n17563__, new_new_n17564__,
    new_new_n17565__, new_new_n17566__, new_new_n17567__, new_new_n17568__,
    new_new_n17569__, new_new_n17570__, new_new_n17571__, new_new_n17572__,
    new_new_n17573__, new_new_n17574__, new_new_n17575__, new_new_n17576__,
    new_new_n17577__, new_new_n17578__, new_new_n17579__, new_new_n17580__,
    new_new_n17581__, new_new_n17582__, new_new_n17583__, new_new_n17584__,
    new_new_n17585__, new_new_n17586__, new_new_n17587__, new_new_n17588__,
    new_new_n17589__, new_new_n17590__, new_new_n17591__, new_new_n17592__,
    new_new_n17593__, new_new_n17594__, new_new_n17595__, new_new_n17596__,
    new_new_n17597__, new_new_n17598__, new_new_n17599__, new_new_n17600__,
    new_new_n17601__, new_new_n17602__, new_new_n17603__, new_new_n17604__,
    new_new_n17605__, new_new_n17606__, new_new_n17607__, new_new_n17608__,
    new_new_n17609__, new_new_n17610__, new_new_n17611__, new_new_n17612__,
    new_new_n17613__, new_new_n17614__, new_new_n17615__, new_new_n17616__,
    new_new_n17617__, new_new_n17618__, new_new_n17619__, new_new_n17620__,
    new_new_n17621__, new_new_n17622__, new_new_n17623__, new_new_n17624__,
    new_new_n17625__, new_new_n17626__, new_new_n17627__, new_new_n17628__,
    new_new_n17629__, new_new_n17630__, new_new_n17631__, new_new_n17632__,
    new_new_n17633__, new_new_n17634__, new_new_n17635__, new_new_n17636__,
    new_new_n17637__, new_new_n17638__, new_new_n17639__, new_new_n17640__,
    new_new_n17641__, new_new_n17642__, new_new_n17643__, new_new_n17644__,
    new_new_n17645__, new_new_n17646__, new_new_n17647__, new_new_n17648__,
    new_new_n17649__, new_new_n17650__, new_new_n17651__, new_new_n17652__,
    new_new_n17653__, new_new_n17654__, new_new_n17655__, new_new_n17656__,
    new_new_n17657__, new_new_n17658__, new_new_n17659__, new_new_n17660__,
    new_new_n17661__, new_new_n17662__, new_new_n17663__, new_new_n17664__,
    new_new_n17665__, new_new_n17667__, new_new_n17668__, new_new_n17669__,
    new_new_n17670__, new_new_n17671__, new_new_n17672__, new_new_n17673__,
    new_new_n17674__, new_new_n17675__, new_new_n17676__, new_new_n17677__,
    new_new_n17678__, new_new_n17679__, new_new_n17680__, new_new_n17681__,
    new_new_n17682__, new_new_n17683__, new_new_n17684__, new_new_n17685__,
    new_new_n17686__, new_new_n17687__, new_new_n17688__, new_new_n17689__,
    new_new_n17690__, new_new_n17691__, new_new_n17692__, new_new_n17693__,
    new_new_n17694__, new_new_n17695__, new_new_n17696__, new_new_n17697__,
    new_new_n17698__, new_new_n17699__, new_new_n17700__, new_new_n17701__,
    new_new_n17702__, new_new_n17703__, new_new_n17704__, new_new_n17705__,
    new_new_n17706__, new_new_n17707__, new_new_n17708__, new_new_n17709__,
    new_new_n17710__, new_new_n17711__, new_new_n17712__, new_new_n17713__,
    new_new_n17714__, new_new_n17715__, new_new_n17716__, new_new_n17717__,
    new_new_n17718__, new_new_n17719__, new_new_n17720__, new_new_n17721__,
    new_new_n17722__, new_new_n17723__, new_new_n17724__, new_new_n17725__,
    new_new_n17726__, new_new_n17727__, new_new_n17728__, new_new_n17729__,
    new_new_n17730__, new_new_n17731__, new_new_n17732__, new_new_n17733__,
    new_new_n17734__, new_new_n17735__, new_new_n17736__, new_new_n17737__,
    new_new_n17738__, new_new_n17739__, new_new_n17740__, new_new_n17741__,
    new_new_n17742__, new_new_n17743__, new_new_n17744__, new_new_n17745__,
    new_new_n17746__, new_new_n17747__, new_new_n17748__, new_new_n17749__,
    new_new_n17750__, new_new_n17751__, new_new_n17752__, new_new_n17753__,
    new_new_n17754__, new_new_n17755__, new_new_n17756__, new_new_n17757__,
    new_new_n17758__, new_new_n17759__, new_new_n17760__, new_new_n17761__,
    new_new_n17762__, new_new_n17763__, new_new_n17764__, new_new_n17765__,
    new_new_n17766__, new_new_n17767__, new_new_n17768__, new_new_n17769__,
    new_new_n17770__, new_new_n17771__, new_new_n17772__, new_new_n17773__,
    new_new_n17774__, new_new_n17775__, new_new_n17776__, new_new_n17777__,
    new_new_n17778__, new_new_n17779__, new_new_n17780__, new_new_n17781__,
    new_new_n17782__, new_new_n17783__, new_new_n17784__, new_new_n17785__,
    new_new_n17786__, new_new_n17787__, new_new_n17788__, new_new_n17789__,
    new_new_n17790__, new_new_n17791__, new_new_n17792__, new_new_n17793__,
    new_new_n17794__, new_new_n17795__, new_new_n17796__, new_new_n17797__,
    new_new_n17798__, new_new_n17799__, new_new_n17800__, new_new_n17801__,
    new_new_n17802__, new_new_n17803__, new_new_n17804__, new_new_n17805__,
    new_new_n17806__, new_new_n17807__, new_new_n17808__, new_new_n17809__,
    new_new_n17810__, new_new_n17811__, new_new_n17812__, new_new_n17813__,
    new_new_n17814__, new_new_n17815__, new_new_n17817__, new_new_n17818__,
    new_new_n17819__, new_new_n17820__, new_new_n17821__, new_new_n17822__,
    new_new_n17823__, new_new_n17824__, new_new_n17825__, new_new_n17826__,
    new_new_n17827__, new_new_n17828__, new_new_n17829__, new_new_n17830__,
    new_new_n17831__, new_new_n17832__, new_new_n17833__, new_new_n17834__,
    new_new_n17835__, new_new_n17836__, new_new_n17837__, new_new_n17838__,
    new_new_n17839__, new_new_n17840__, new_new_n17841__, new_new_n17842__,
    new_new_n17843__, new_new_n17844__, new_new_n17845__, new_new_n17846__,
    new_new_n17847__, new_new_n17848__, new_new_n17849__, new_new_n17850__,
    new_new_n17851__, new_new_n17852__, new_new_n17853__, new_new_n17854__,
    new_new_n17855__, new_new_n17856__, new_new_n17857__, new_new_n17858__,
    new_new_n17859__, new_new_n17860__, new_new_n17861__, new_new_n17862__,
    new_new_n17863__, new_new_n17864__, new_new_n17865__, new_new_n17866__,
    new_new_n17867__, new_new_n17868__, new_new_n17869__, new_new_n17870__,
    new_new_n17871__, new_new_n17872__, new_new_n17873__, new_new_n17874__,
    new_new_n17875__, new_new_n17876__, new_new_n17877__, new_new_n17878__,
    new_new_n17879__, new_new_n17880__, new_new_n17881__, new_new_n17882__,
    new_new_n17883__, new_new_n17884__, new_new_n17885__, new_new_n17886__,
    new_new_n17887__, new_new_n17888__, new_new_n17889__, new_new_n17890__,
    new_new_n17891__, new_new_n17892__, new_new_n17893__, new_new_n17894__,
    new_new_n17895__, new_new_n17896__, new_new_n17897__, new_new_n17898__,
    new_new_n17899__, new_new_n17900__, new_new_n17901__, new_new_n17902__,
    new_new_n17903__, new_new_n17904__, new_new_n17905__, new_new_n17906__,
    new_new_n17907__, new_new_n17908__, new_new_n17909__, new_new_n17910__,
    new_new_n17911__, new_new_n17912__, new_new_n17913__, new_new_n17914__,
    new_new_n17915__, new_new_n17916__, new_new_n17917__, new_new_n17918__,
    new_new_n17919__, new_new_n17920__, new_new_n17921__, new_new_n17922__,
    new_new_n17923__, new_new_n17924__, new_new_n17925__, new_new_n17926__,
    new_new_n17927__, new_new_n17928__, new_new_n17929__, new_new_n17930__,
    new_new_n17931__, new_new_n17932__, new_new_n17933__, new_new_n17934__,
    new_new_n17935__, new_new_n17936__, new_new_n17937__, new_new_n17938__,
    new_new_n17939__, new_new_n17940__, new_new_n17941__, new_new_n17942__,
    new_new_n17943__, new_new_n17944__, new_new_n17945__, new_new_n17946__,
    new_new_n17947__, new_new_n17948__, new_new_n17949__, new_new_n17950__,
    new_new_n17951__, new_new_n17952__, new_new_n17953__, new_new_n17954__,
    new_new_n17955__, new_new_n17956__, new_new_n17957__, new_new_n17958__,
    new_new_n17959__, new_new_n17960__, new_new_n17961__, new_new_n17962__,
    new_new_n17963__, new_new_n17965__, new_new_n17966__, new_new_n17967__,
    new_new_n17968__, new_new_n17969__, new_new_n17970__, new_new_n17971__,
    new_new_n17972__, new_new_n17973__, new_new_n17974__, new_new_n17975__,
    new_new_n17976__, new_new_n17977__, new_new_n17978__, new_new_n17979__,
    new_new_n17980__, new_new_n17981__, new_new_n17982__, new_new_n17983__,
    new_new_n17984__, new_new_n17985__, new_new_n17986__, new_new_n17987__,
    new_new_n17988__, new_new_n17989__, new_new_n17990__, new_new_n17991__,
    new_new_n17992__, new_new_n17993__, new_new_n17994__, new_new_n17995__,
    new_new_n17996__, new_new_n17997__, new_new_n17998__, new_new_n17999__,
    new_new_n18000__, new_new_n18001__, new_new_n18002__, new_new_n18003__,
    new_new_n18004__, new_new_n18005__, new_new_n18006__, new_new_n18007__,
    new_new_n18008__, new_new_n18009__, new_new_n18010__, new_new_n18011__,
    new_new_n18012__, new_new_n18013__, new_new_n18014__, new_new_n18015__,
    new_new_n18016__, new_new_n18017__, new_new_n18018__, new_new_n18019__,
    new_new_n18020__, new_new_n18021__, new_new_n18022__, new_new_n18023__,
    new_new_n18024__, new_new_n18025__, new_new_n18026__, new_new_n18027__,
    new_new_n18028__, new_new_n18029__, new_new_n18030__, new_new_n18031__,
    new_new_n18032__, new_new_n18033__, new_new_n18034__, new_new_n18035__,
    new_new_n18036__, new_new_n18037__, new_new_n18038__, new_new_n18039__,
    new_new_n18040__, new_new_n18041__, new_new_n18042__, new_new_n18043__,
    new_new_n18044__, new_new_n18045__, new_new_n18046__, new_new_n18047__,
    new_new_n18048__, new_new_n18049__, new_new_n18050__, new_new_n18051__,
    new_new_n18052__, new_new_n18053__, new_new_n18054__, new_new_n18055__,
    new_new_n18056__, new_new_n18057__, new_new_n18058__, new_new_n18059__,
    new_new_n18060__, new_new_n18061__, new_new_n18062__, new_new_n18063__,
    new_new_n18064__, new_new_n18065__, new_new_n18066__, new_new_n18067__,
    new_new_n18068__, new_new_n18069__, new_new_n18070__, new_new_n18071__,
    new_new_n18072__, new_new_n18073__, new_new_n18074__, new_new_n18075__,
    new_new_n18076__, new_new_n18077__, new_new_n18078__, new_new_n18079__,
    new_new_n18080__, new_new_n18081__, new_new_n18082__, new_new_n18083__,
    new_new_n18084__, new_new_n18085__, new_new_n18086__, new_new_n18087__,
    new_new_n18088__, new_new_n18089__, new_new_n18090__, new_new_n18091__,
    new_new_n18093__, new_new_n18094__, new_new_n18095__, new_new_n18096__,
    new_new_n18097__, new_new_n18098__, new_new_n18099__, new_new_n18100__,
    new_new_n18101__, new_new_n18102__, new_new_n18103__, new_new_n18104__,
    new_new_n18105__, new_new_n18106__, new_new_n18107__, new_new_n18108__,
    new_new_n18109__, new_new_n18110__, new_new_n18111__, new_new_n18112__,
    new_new_n18113__, new_new_n18114__, new_new_n18115__, new_new_n18116__,
    new_new_n18117__, new_new_n18118__, new_new_n18119__, new_new_n18120__,
    new_new_n18121__, new_new_n18122__, new_new_n18123__, new_new_n18124__,
    new_new_n18125__, new_new_n18126__, new_new_n18127__, new_new_n18128__,
    new_new_n18129__, new_new_n18130__, new_new_n18131__, new_new_n18132__,
    new_new_n18133__, new_new_n18134__, new_new_n18135__, new_new_n18136__,
    new_new_n18137__, new_new_n18138__, new_new_n18139__, new_new_n18140__,
    new_new_n18141__, new_new_n18142__, new_new_n18143__, new_new_n18144__,
    new_new_n18145__, new_new_n18146__, new_new_n18147__, new_new_n18148__,
    new_new_n18149__, new_new_n18150__, new_new_n18151__, new_new_n18152__,
    new_new_n18153__, new_new_n18154__, new_new_n18155__, new_new_n18156__,
    new_new_n18157__, new_new_n18158__, new_new_n18159__, new_new_n18160__,
    new_new_n18161__, new_new_n18162__, new_new_n18163__, new_new_n18164__,
    new_new_n18165__, new_new_n18166__, new_new_n18167__, new_new_n18168__,
    new_new_n18169__, new_new_n18170__, new_new_n18171__, new_new_n18172__,
    new_new_n18173__, new_new_n18174__, new_new_n18175__, new_new_n18176__,
    new_new_n18177__, new_new_n18178__, new_new_n18179__, new_new_n18180__,
    new_new_n18181__, new_new_n18182__, new_new_n18183__, new_new_n18184__,
    new_new_n18185__, new_new_n18186__, new_new_n18187__, new_new_n18188__,
    new_new_n18189__, new_new_n18190__, new_new_n18191__, new_new_n18192__,
    new_new_n18193__, new_new_n18194__, new_new_n18195__, new_new_n18196__,
    new_new_n18197__, new_new_n18198__, new_new_n18199__, new_new_n18200__,
    new_new_n18201__, new_new_n18202__, new_new_n18203__, new_new_n18204__,
    new_new_n18205__, new_new_n18206__, new_new_n18207__, new_new_n18208__,
    new_new_n18209__, new_new_n18210__, new_new_n18211__, new_new_n18212__,
    new_new_n18213__, new_new_n18214__, new_new_n18215__, new_new_n18216__,
    new_new_n18217__, new_new_n18218__, new_new_n18219__, new_new_n18220__,
    new_new_n18221__, new_new_n18222__, new_new_n18223__, new_new_n18224__,
    new_new_n18225__, new_new_n18226__, new_new_n18227__, new_new_n18228__,
    new_new_n18229__, new_new_n18230__, new_new_n18231__, new_new_n18232__,
    new_new_n18233__, new_new_n18234__, new_new_n18235__, new_new_n18236__,
    new_new_n18237__, new_new_n18239__, new_new_n18240__, new_new_n18241__,
    new_new_n18242__, new_new_n18243__, new_new_n18244__, new_new_n18245__,
    new_new_n18246__, new_new_n18247__, new_new_n18248__, new_new_n18249__,
    new_new_n18250__, new_new_n18251__, new_new_n18252__, new_new_n18253__,
    new_new_n18254__, new_new_n18255__, new_new_n18256__, new_new_n18257__,
    new_new_n18258__, new_new_n18259__, new_new_n18260__, new_new_n18261__,
    new_new_n18262__, new_new_n18263__, new_new_n18264__, new_new_n18265__,
    new_new_n18266__, new_new_n18267__, new_new_n18268__, new_new_n18269__,
    new_new_n18270__, new_new_n18271__, new_new_n18272__, new_new_n18273__,
    new_new_n18274__, new_new_n18275__, new_new_n18276__, new_new_n18277__,
    new_new_n18278__, new_new_n18279__, new_new_n18280__, new_new_n18281__,
    new_new_n18282__, new_new_n18283__, new_new_n18284__, new_new_n18285__,
    new_new_n18286__, new_new_n18287__, new_new_n18288__, new_new_n18289__,
    new_new_n18290__, new_new_n18291__, new_new_n18292__, new_new_n18293__,
    new_new_n18294__, new_new_n18295__, new_new_n18296__, new_new_n18297__,
    new_new_n18298__, new_new_n18299__, new_new_n18300__, new_new_n18301__,
    new_new_n18302__, new_new_n18303__, new_new_n18304__, new_new_n18305__,
    new_new_n18306__, new_new_n18307__, new_new_n18308__, new_new_n18309__,
    new_new_n18310__, new_new_n18311__, new_new_n18312__, new_new_n18313__,
    new_new_n18314__, new_new_n18315__, new_new_n18316__, new_new_n18317__,
    new_new_n18318__, new_new_n18319__, new_new_n18320__, new_new_n18321__,
    new_new_n18322__, new_new_n18323__, new_new_n18324__, new_new_n18325__,
    new_new_n18326__, new_new_n18327__, new_new_n18328__, new_new_n18329__,
    new_new_n18330__, new_new_n18331__, new_new_n18332__, new_new_n18333__,
    new_new_n18334__, new_new_n18335__, new_new_n18336__, new_new_n18337__,
    new_new_n18338__, new_new_n18339__, new_new_n18340__, new_new_n18341__,
    new_new_n18342__, new_new_n18343__, new_new_n18344__, new_new_n18345__,
    new_new_n18346__, new_new_n18347__, new_new_n18348__, new_new_n18349__,
    new_new_n18350__, new_new_n18351__, new_new_n18352__, new_new_n18353__,
    new_new_n18354__, new_new_n18355__, new_new_n18356__, new_new_n18357__,
    new_new_n18358__, new_new_n18359__, new_new_n18360__, new_new_n18362__,
    new_new_n18363__, new_new_n18364__, new_new_n18365__, new_new_n18366__,
    new_new_n18367__, new_new_n18368__, new_new_n18369__, new_new_n18370__,
    new_new_n18371__, new_new_n18372__, new_new_n18373__, new_new_n18374__,
    new_new_n18375__, new_new_n18376__, new_new_n18377__, new_new_n18378__,
    new_new_n18379__, new_new_n18380__, new_new_n18381__, new_new_n18382__,
    new_new_n18383__, new_new_n18384__, new_new_n18385__, new_new_n18386__,
    new_new_n18387__, new_new_n18388__, new_new_n18389__, new_new_n18390__,
    new_new_n18391__, new_new_n18392__, new_new_n18393__, new_new_n18394__,
    new_new_n18395__, new_new_n18396__, new_new_n18397__, new_new_n18398__,
    new_new_n18399__, new_new_n18400__, new_new_n18401__, new_new_n18402__,
    new_new_n18403__, new_new_n18404__, new_new_n18405__, new_new_n18406__,
    new_new_n18407__, new_new_n18408__, new_new_n18409__, new_new_n18410__,
    new_new_n18411__, new_new_n18412__, new_new_n18413__, new_new_n18414__,
    new_new_n18415__, new_new_n18416__, new_new_n18417__, new_new_n18418__,
    new_new_n18419__, new_new_n18420__, new_new_n18421__, new_new_n18422__,
    new_new_n18423__, new_new_n18424__, new_new_n18425__, new_new_n18426__,
    new_new_n18427__, new_new_n18428__, new_new_n18429__, new_new_n18430__,
    new_new_n18431__, new_new_n18432__, new_new_n18433__, new_new_n18434__,
    new_new_n18435__, new_new_n18436__, new_new_n18437__, new_new_n18438__,
    new_new_n18439__, new_new_n18440__, new_new_n18441__, new_new_n18442__,
    new_new_n18443__, new_new_n18444__, new_new_n18445__, new_new_n18446__,
    new_new_n18447__, new_new_n18448__, new_new_n18449__, new_new_n18450__,
    new_new_n18451__, new_new_n18452__, new_new_n18453__, new_new_n18454__,
    new_new_n18455__, new_new_n18456__, new_new_n18457__, new_new_n18458__,
    new_new_n18459__, new_new_n18460__, new_new_n18461__, new_new_n18462__,
    new_new_n18463__, new_new_n18464__, new_new_n18465__, new_new_n18466__,
    new_new_n18467__, new_new_n18468__, new_new_n18469__, new_new_n18470__,
    new_new_n18471__, new_new_n18472__, new_new_n18473__, new_new_n18474__,
    new_new_n18475__, new_new_n18476__, new_new_n18477__, new_new_n18478__,
    new_new_n18479__, new_new_n18480__, new_new_n18481__, new_new_n18482__,
    new_new_n18483__, new_new_n18484__, new_new_n18485__, new_new_n18486__,
    new_new_n18487__, new_new_n18488__, new_new_n18489__, new_new_n18490__,
    new_new_n18491__, new_new_n18492__, new_new_n18494__, new_new_n18495__,
    new_new_n18496__, new_new_n18497__, new_new_n18498__, new_new_n18499__,
    new_new_n18500__, new_new_n18501__, new_new_n18502__, new_new_n18503__,
    new_new_n18504__, new_new_n18505__, new_new_n18506__, new_new_n18507__,
    new_new_n18508__, new_new_n18509__, new_new_n18510__, new_new_n18511__,
    new_new_n18512__, new_new_n18513__, new_new_n18514__, new_new_n18515__,
    new_new_n18516__, new_new_n18517__, new_new_n18518__, new_new_n18519__,
    new_new_n18520__, new_new_n18521__, new_new_n18522__, new_new_n18523__,
    new_new_n18524__, new_new_n18525__, new_new_n18526__, new_new_n18527__,
    new_new_n18528__, new_new_n18529__, new_new_n18530__, new_new_n18531__,
    new_new_n18532__, new_new_n18533__, new_new_n18534__, new_new_n18535__,
    new_new_n18536__, new_new_n18537__, new_new_n18538__, new_new_n18539__,
    new_new_n18540__, new_new_n18541__, new_new_n18542__, new_new_n18543__,
    new_new_n18544__, new_new_n18545__, new_new_n18546__, new_new_n18547__,
    new_new_n18548__, new_new_n18549__, new_new_n18550__, new_new_n18551__,
    new_new_n18552__, new_new_n18553__, new_new_n18554__, new_new_n18555__,
    new_new_n18556__, new_new_n18557__, new_new_n18558__, new_new_n18559__,
    new_new_n18560__, new_new_n18561__, new_new_n18562__, new_new_n18563__,
    new_new_n18564__, new_new_n18565__, new_new_n18566__, new_new_n18567__,
    new_new_n18568__, new_new_n18569__, new_new_n18570__, new_new_n18571__,
    new_new_n18572__, new_new_n18573__, new_new_n18574__, new_new_n18575__,
    new_new_n18576__, new_new_n18577__, new_new_n18578__, new_new_n18579__,
    new_new_n18580__, new_new_n18581__, new_new_n18582__, new_new_n18583__,
    new_new_n18584__, new_new_n18585__, new_new_n18586__, new_new_n18587__,
    new_new_n18588__, new_new_n18589__, new_new_n18590__, new_new_n18591__,
    new_new_n18592__, new_new_n18593__, new_new_n18594__, new_new_n18595__,
    new_new_n18596__, new_new_n18597__, new_new_n18598__, new_new_n18599__,
    new_new_n18600__, new_new_n18601__, new_new_n18602__, new_new_n18603__,
    new_new_n18604__, new_new_n18605__, new_new_n18606__, new_new_n18607__,
    new_new_n18608__, new_new_n18609__, new_new_n18610__, new_new_n18611__,
    new_new_n18613__, new_new_n18614__, new_new_n18615__, new_new_n18616__,
    new_new_n18617__, new_new_n18618__, new_new_n18619__, new_new_n18620__,
    new_new_n18621__, new_new_n18622__, new_new_n18623__, new_new_n18624__,
    new_new_n18625__, new_new_n18626__, new_new_n18627__, new_new_n18628__,
    new_new_n18629__, new_new_n18630__, new_new_n18631__, new_new_n18632__,
    new_new_n18633__, new_new_n18634__, new_new_n18635__, new_new_n18636__,
    new_new_n18637__, new_new_n18638__, new_new_n18639__, new_new_n18640__,
    new_new_n18641__, new_new_n18642__, new_new_n18643__, new_new_n18644__,
    new_new_n18645__, new_new_n18646__, new_new_n18647__, new_new_n18648__,
    new_new_n18649__, new_new_n18650__, new_new_n18651__, new_new_n18652__,
    new_new_n18653__, new_new_n18654__, new_new_n18655__, new_new_n18656__,
    new_new_n18657__, new_new_n18658__, new_new_n18659__, new_new_n18660__,
    new_new_n18661__, new_new_n18662__, new_new_n18663__, new_new_n18664__,
    new_new_n18665__, new_new_n18666__, new_new_n18667__, new_new_n18668__,
    new_new_n18669__, new_new_n18670__, new_new_n18671__, new_new_n18672__,
    new_new_n18673__, new_new_n18674__, new_new_n18675__, new_new_n18676__,
    new_new_n18677__, new_new_n18678__, new_new_n18679__, new_new_n18680__,
    new_new_n18681__, new_new_n18682__, new_new_n18683__, new_new_n18684__,
    new_new_n18685__, new_new_n18686__, new_new_n18687__, new_new_n18688__,
    new_new_n18689__, new_new_n18690__, new_new_n18691__, new_new_n18692__,
    new_new_n18693__, new_new_n18694__, new_new_n18695__, new_new_n18696__,
    new_new_n18697__, new_new_n18698__, new_new_n18699__, new_new_n18700__,
    new_new_n18701__, new_new_n18702__, new_new_n18703__, new_new_n18704__,
    new_new_n18705__, new_new_n18706__, new_new_n18707__, new_new_n18708__,
    new_new_n18709__, new_new_n18710__, new_new_n18711__, new_new_n18712__,
    new_new_n18713__, new_new_n18714__, new_new_n18715__, new_new_n18716__,
    new_new_n18717__, new_new_n18718__, new_new_n18719__, new_new_n18720__,
    new_new_n18721__, new_new_n18722__, new_new_n18723__, new_new_n18725__,
    new_new_n18726__, new_new_n18727__, new_new_n18728__, new_new_n18729__,
    new_new_n18730__, new_new_n18731__, new_new_n18732__, new_new_n18733__,
    new_new_n18734__, new_new_n18735__, new_new_n18736__, new_new_n18737__,
    new_new_n18738__, new_new_n18739__, new_new_n18740__, new_new_n18741__,
    new_new_n18742__, new_new_n18743__, new_new_n18744__, new_new_n18745__,
    new_new_n18746__, new_new_n18747__, new_new_n18748__, new_new_n18749__,
    new_new_n18750__, new_new_n18751__, new_new_n18752__, new_new_n18753__,
    new_new_n18754__, new_new_n18755__, new_new_n18756__, new_new_n18757__,
    new_new_n18758__, new_new_n18759__, new_new_n18760__, new_new_n18761__,
    new_new_n18762__, new_new_n18763__, new_new_n18764__, new_new_n18765__,
    new_new_n18766__, new_new_n18767__, new_new_n18768__, new_new_n18769__,
    new_new_n18770__, new_new_n18771__, new_new_n18772__, new_new_n18773__,
    new_new_n18774__, new_new_n18775__, new_new_n18776__, new_new_n18777__,
    new_new_n18778__, new_new_n18779__, new_new_n18780__, new_new_n18781__,
    new_new_n18782__, new_new_n18783__, new_new_n18784__, new_new_n18785__,
    new_new_n18786__, new_new_n18787__, new_new_n18788__, new_new_n18789__,
    new_new_n18790__, new_new_n18791__, new_new_n18792__, new_new_n18793__,
    new_new_n18794__, new_new_n18795__, new_new_n18796__, new_new_n18797__,
    new_new_n18798__, new_new_n18799__, new_new_n18800__, new_new_n18801__,
    new_new_n18802__, new_new_n18803__, new_new_n18804__, new_new_n18805__,
    new_new_n18806__, new_new_n18807__, new_new_n18808__, new_new_n18809__,
    new_new_n18810__, new_new_n18811__, new_new_n18812__, new_new_n18813__,
    new_new_n18814__, new_new_n18815__, new_new_n18816__, new_new_n18817__,
    new_new_n18818__, new_new_n18819__, new_new_n18820__, new_new_n18821__,
    new_new_n18822__, new_new_n18823__, new_new_n18824__, new_new_n18825__,
    new_new_n18826__, new_new_n18827__, new_new_n18828__, new_new_n18829__,
    new_new_n18830__, new_new_n18831__, new_new_n18832__, new_new_n18833__,
    new_new_n18834__, new_new_n18835__, new_new_n18836__, new_new_n18837__,
    new_new_n18838__, new_new_n18839__, new_new_n18840__, new_new_n18841__,
    new_new_n18842__, new_new_n18843__, new_new_n18844__, new_new_n18845__,
    new_new_n18846__, new_new_n18847__, new_new_n18848__, new_new_n18849__,
    new_new_n18850__, new_new_n18852__, new_new_n18853__, new_new_n18854__,
    new_new_n18855__, new_new_n18856__, new_new_n18857__, new_new_n18858__,
    new_new_n18859__, new_new_n18860__, new_new_n18861__, new_new_n18862__,
    new_new_n18863__, new_new_n18864__, new_new_n18865__, new_new_n18866__,
    new_new_n18867__, new_new_n18868__, new_new_n18869__, new_new_n18870__,
    new_new_n18871__, new_new_n18872__, new_new_n18873__, new_new_n18874__,
    new_new_n18875__, new_new_n18876__, new_new_n18877__, new_new_n18878__,
    new_new_n18879__, new_new_n18880__, new_new_n18881__, new_new_n18882__,
    new_new_n18883__, new_new_n18884__, new_new_n18885__, new_new_n18886__,
    new_new_n18887__, new_new_n18888__, new_new_n18889__, new_new_n18890__,
    new_new_n18891__, new_new_n18892__, new_new_n18893__, new_new_n18894__,
    new_new_n18895__, new_new_n18896__, new_new_n18897__, new_new_n18898__,
    new_new_n18899__, new_new_n18900__, new_new_n18901__, new_new_n18902__,
    new_new_n18903__, new_new_n18904__, new_new_n18905__, new_new_n18906__,
    new_new_n18907__, new_new_n18908__, new_new_n18909__, new_new_n18910__,
    new_new_n18911__, new_new_n18912__, new_new_n18913__, new_new_n18914__,
    new_new_n18915__, new_new_n18916__, new_new_n18917__, new_new_n18918__,
    new_new_n18919__, new_new_n18920__, new_new_n18921__, new_new_n18922__,
    new_new_n18923__, new_new_n18924__, new_new_n18925__, new_new_n18926__,
    new_new_n18927__, new_new_n18928__, new_new_n18929__, new_new_n18930__,
    new_new_n18931__, new_new_n18932__, new_new_n18933__, new_new_n18934__,
    new_new_n18935__, new_new_n18936__, new_new_n18937__, new_new_n18938__,
    new_new_n18939__, new_new_n18940__, new_new_n18941__, new_new_n18942__,
    new_new_n18943__, new_new_n18944__, new_new_n18945__, new_new_n18946__,
    new_new_n18947__, new_new_n18948__, new_new_n18949__, new_new_n18950__,
    new_new_n18951__, new_new_n18952__, new_new_n18953__, new_new_n18954__,
    new_new_n18955__, new_new_n18956__, new_new_n18957__, new_new_n18958__,
    new_new_n18959__, new_new_n18960__, new_new_n18961__, new_new_n18962__,
    new_new_n18963__, new_new_n18965__, new_new_n18966__, new_new_n18967__,
    new_new_n18968__, new_new_n18969__, new_new_n18970__, new_new_n18971__,
    new_new_n18972__, new_new_n18973__, new_new_n18974__, new_new_n18975__,
    new_new_n18976__, new_new_n18977__, new_new_n18978__, new_new_n18979__,
    new_new_n18980__, new_new_n18981__, new_new_n18982__, new_new_n18983__,
    new_new_n18984__, new_new_n18985__, new_new_n18986__, new_new_n18987__,
    new_new_n18988__, new_new_n18989__, new_new_n18990__, new_new_n18991__,
    new_new_n18992__, new_new_n18993__, new_new_n18994__, new_new_n18995__,
    new_new_n18996__, new_new_n18997__, new_new_n18998__, new_new_n18999__,
    new_new_n19000__, new_new_n19001__, new_new_n19002__, new_new_n19003__,
    new_new_n19004__, new_new_n19005__, new_new_n19006__, new_new_n19007__,
    new_new_n19008__, new_new_n19009__, new_new_n19010__, new_new_n19011__,
    new_new_n19012__, new_new_n19013__, new_new_n19014__, new_new_n19015__,
    new_new_n19016__, new_new_n19017__, new_new_n19018__, new_new_n19019__,
    new_new_n19020__, new_new_n19021__, new_new_n19022__, new_new_n19023__,
    new_new_n19024__, new_new_n19025__, new_new_n19026__, new_new_n19027__,
    new_new_n19028__, new_new_n19029__, new_new_n19030__, new_new_n19031__,
    new_new_n19032__, new_new_n19033__, new_new_n19034__, new_new_n19035__,
    new_new_n19036__, new_new_n19037__, new_new_n19038__, new_new_n19039__,
    new_new_n19040__, new_new_n19041__, new_new_n19042__, new_new_n19043__,
    new_new_n19044__, new_new_n19045__, new_new_n19046__, new_new_n19047__,
    new_new_n19048__, new_new_n19049__, new_new_n19050__, new_new_n19051__,
    new_new_n19052__, new_new_n19054__, new_new_n19055__, new_new_n19056__,
    new_new_n19057__, new_new_n19058__, new_new_n19059__, new_new_n19060__,
    new_new_n19061__, new_new_n19062__, new_new_n19063__, new_new_n19064__,
    new_new_n19065__, new_new_n19066__, new_new_n19067__, new_new_n19068__,
    new_new_n19069__, new_new_n19070__, new_new_n19071__, new_new_n19072__,
    new_new_n19073__, new_new_n19074__, new_new_n19075__, new_new_n19076__,
    new_new_n19077__, new_new_n19078__, new_new_n19079__, new_new_n19080__,
    new_new_n19081__, new_new_n19082__, new_new_n19083__, new_new_n19084__,
    new_new_n19085__, new_new_n19086__, new_new_n19087__, new_new_n19088__,
    new_new_n19089__, new_new_n19090__, new_new_n19091__, new_new_n19092__,
    new_new_n19093__, new_new_n19094__, new_new_n19095__, new_new_n19096__,
    new_new_n19097__, new_new_n19098__, new_new_n19099__, new_new_n19100__,
    new_new_n19101__, new_new_n19102__, new_new_n19103__, new_new_n19104__,
    new_new_n19105__, new_new_n19106__, new_new_n19107__, new_new_n19108__,
    new_new_n19109__, new_new_n19110__, new_new_n19111__, new_new_n19112__,
    new_new_n19113__, new_new_n19114__, new_new_n19115__, new_new_n19116__,
    new_new_n19117__, new_new_n19118__, new_new_n19119__, new_new_n19120__,
    new_new_n19121__, new_new_n19122__, new_new_n19123__, new_new_n19124__,
    new_new_n19125__, new_new_n19126__, new_new_n19127__, new_new_n19128__,
    new_new_n19129__, new_new_n19130__, new_new_n19131__, new_new_n19132__,
    new_new_n19133__, new_new_n19134__, new_new_n19135__, new_new_n19136__,
    new_new_n19137__, new_new_n19138__, new_new_n19139__, new_new_n19140__,
    new_new_n19141__, new_new_n19142__, new_new_n19143__, new_new_n19144__,
    new_new_n19145__, new_new_n19146__, new_new_n19147__, new_new_n19148__,
    new_new_n19149__, new_new_n19150__, new_new_n19151__, new_new_n19152__,
    new_new_n19154__, new_new_n19155__, new_new_n19156__, new_new_n19157__,
    new_new_n19158__, new_new_n19159__, new_new_n19160__, new_new_n19161__,
    new_new_n19162__, new_new_n19163__, new_new_n19164__, new_new_n19165__,
    new_new_n19166__, new_new_n19167__, new_new_n19168__, new_new_n19169__,
    new_new_n19170__, new_new_n19171__, new_new_n19172__, new_new_n19173__,
    new_new_n19174__, new_new_n19175__, new_new_n19176__, new_new_n19177__,
    new_new_n19178__, new_new_n19179__, new_new_n19180__, new_new_n19181__,
    new_new_n19182__, new_new_n19183__, new_new_n19184__, new_new_n19185__,
    new_new_n19186__, new_new_n19187__, new_new_n19188__, new_new_n19189__,
    new_new_n19190__, new_new_n19191__, new_new_n19192__, new_new_n19193__,
    new_new_n19194__, new_new_n19195__, new_new_n19196__, new_new_n19197__,
    new_new_n19198__, new_new_n19199__, new_new_n19200__, new_new_n19201__,
    new_new_n19202__, new_new_n19203__, new_new_n19204__, new_new_n19205__,
    new_new_n19206__, new_new_n19207__, new_new_n19208__, new_new_n19209__,
    new_new_n19210__, new_new_n19211__, new_new_n19212__, new_new_n19213__,
    new_new_n19214__, new_new_n19215__, new_new_n19216__, new_new_n19217__,
    new_new_n19218__, new_new_n19219__, new_new_n19220__, new_new_n19221__,
    new_new_n19222__, new_new_n19223__, new_new_n19224__, new_new_n19225__,
    new_new_n19226__, new_new_n19227__, new_new_n19228__, new_new_n19229__,
    new_new_n19230__, new_new_n19231__, new_new_n19232__, new_new_n19233__,
    new_new_n19234__, new_new_n19235__, new_new_n19236__, new_new_n19237__,
    new_new_n19239__, new_new_n19240__, new_new_n19241__, new_new_n19242__,
    new_new_n19243__, new_new_n19244__, new_new_n19245__, new_new_n19246__,
    new_new_n19247__, new_new_n19248__, new_new_n19249__, new_new_n19250__,
    new_new_n19251__, new_new_n19252__, new_new_n19253__, new_new_n19254__,
    new_new_n19255__, new_new_n19256__, new_new_n19257__, new_new_n19258__,
    new_new_n19259__, new_new_n19260__, new_new_n19261__, new_new_n19262__,
    new_new_n19263__, new_new_n19264__, new_new_n19265__, new_new_n19266__,
    new_new_n19267__, new_new_n19268__, new_new_n19269__, new_new_n19270__,
    new_new_n19271__, new_new_n19272__, new_new_n19273__, new_new_n19274__,
    new_new_n19275__, new_new_n19276__, new_new_n19277__, new_new_n19278__,
    new_new_n19279__, new_new_n19280__, new_new_n19281__, new_new_n19282__,
    new_new_n19283__, new_new_n19284__, new_new_n19285__, new_new_n19286__,
    new_new_n19287__, new_new_n19288__, new_new_n19289__, new_new_n19290__,
    new_new_n19291__, new_new_n19292__, new_new_n19293__, new_new_n19294__,
    new_new_n19295__, new_new_n19296__, new_new_n19297__, new_new_n19298__,
    new_new_n19299__, new_new_n19300__, new_new_n19301__, new_new_n19302__,
    new_new_n19303__, new_new_n19304__, new_new_n19305__, new_new_n19306__,
    new_new_n19307__, new_new_n19308__, new_new_n19309__, new_new_n19310__,
    new_new_n19311__, new_new_n19312__, new_new_n19313__, new_new_n19314__,
    new_new_n19315__, new_new_n19316__, new_new_n19317__, new_new_n19318__,
    new_new_n19319__, new_new_n19320__, new_new_n19321__, new_new_n19322__,
    new_new_n19323__, new_new_n19324__, new_new_n19325__, new_new_n19326__,
    new_new_n19327__, new_new_n19328__, new_new_n19329__, new_new_n19330__,
    new_new_n19331__, new_new_n19332__, new_new_n19333__, new_new_n19334__,
    new_new_n19335__, new_new_n19336__, new_new_n19337__, new_new_n19338__,
    new_new_n19339__, new_new_n19340__, new_new_n19341__, new_new_n19342__,
    new_new_n19343__, new_new_n19344__, new_new_n19345__, new_new_n19346__,
    new_new_n19348__, new_new_n19349__, new_new_n19350__, new_new_n19351__,
    new_new_n19352__, new_new_n19353__, new_new_n19354__, new_new_n19355__,
    new_new_n19356__, new_new_n19357__, new_new_n19358__, new_new_n19359__,
    new_new_n19360__, new_new_n19361__, new_new_n19362__, new_new_n19363__,
    new_new_n19364__, new_new_n19365__, new_new_n19366__, new_new_n19367__,
    new_new_n19368__, new_new_n19369__, new_new_n19370__, new_new_n19371__,
    new_new_n19372__, new_new_n19373__, new_new_n19374__, new_new_n19375__,
    new_new_n19376__, new_new_n19377__, new_new_n19378__, new_new_n19379__,
    new_new_n19380__, new_new_n19381__, new_new_n19382__, new_new_n19383__,
    new_new_n19384__, new_new_n19385__, new_new_n19386__, new_new_n19387__,
    new_new_n19388__, new_new_n19389__, new_new_n19390__, new_new_n19391__,
    new_new_n19392__, new_new_n19393__, new_new_n19394__, new_new_n19395__,
    new_new_n19396__, new_new_n19397__, new_new_n19398__, new_new_n19399__,
    new_new_n19400__, new_new_n19401__, new_new_n19402__, new_new_n19403__,
    new_new_n19404__, new_new_n19405__, new_new_n19406__, new_new_n19407__,
    new_new_n19408__, new_new_n19409__, new_new_n19410__, new_new_n19411__,
    new_new_n19412__, new_new_n19413__, new_new_n19414__, new_new_n19415__,
    new_new_n19416__, new_new_n19417__, new_new_n19418__, new_new_n19419__,
    new_new_n19420__, new_new_n19421__, new_new_n19422__, new_new_n19423__,
    new_new_n19424__, new_new_n19425__, new_new_n19426__, new_new_n19427__,
    new_new_n19428__, new_new_n19430__, new_new_n19431__, new_new_n19432__,
    new_new_n19433__, new_new_n19434__, new_new_n19435__, new_new_n19436__,
    new_new_n19437__, new_new_n19438__, new_new_n19439__, new_new_n19440__,
    new_new_n19441__, new_new_n19442__, new_new_n19443__, new_new_n19444__,
    new_new_n19445__, new_new_n19446__, new_new_n19447__, new_new_n19448__,
    new_new_n19449__, new_new_n19450__, new_new_n19451__, new_new_n19452__,
    new_new_n19453__, new_new_n19454__, new_new_n19455__, new_new_n19456__,
    new_new_n19457__, new_new_n19458__, new_new_n19459__, new_new_n19460__,
    new_new_n19461__, new_new_n19462__, new_new_n19463__, new_new_n19464__,
    new_new_n19465__, new_new_n19466__, new_new_n19467__, new_new_n19468__,
    new_new_n19469__, new_new_n19470__, new_new_n19471__, new_new_n19472__,
    new_new_n19473__, new_new_n19474__, new_new_n19475__, new_new_n19476__,
    new_new_n19477__, new_new_n19478__, new_new_n19479__, new_new_n19480__,
    new_new_n19481__, new_new_n19482__, new_new_n19483__, new_new_n19484__,
    new_new_n19485__, new_new_n19486__, new_new_n19487__, new_new_n19488__,
    new_new_n19489__, new_new_n19490__, new_new_n19491__, new_new_n19492__,
    new_new_n19493__, new_new_n19494__, new_new_n19495__, new_new_n19496__,
    new_new_n19497__, new_new_n19498__, new_new_n19499__, new_new_n19500__,
    new_new_n19501__, new_new_n19502__, new_new_n19503__, new_new_n19504__,
    new_new_n19505__, new_new_n19506__, new_new_n19507__, new_new_n19508__,
    new_new_n19509__, new_new_n19510__, new_new_n19511__, new_new_n19512__,
    new_new_n19513__, new_new_n19514__, new_new_n19515__, new_new_n19516__,
    new_new_n19517__, new_new_n19518__, new_new_n19519__, new_new_n19520__,
    new_new_n19522__, new_new_n19523__, new_new_n19524__, new_new_n19525__,
    new_new_n19526__, new_new_n19527__, new_new_n19528__, new_new_n19529__,
    new_new_n19530__, new_new_n19531__, new_new_n19532__, new_new_n19533__,
    new_new_n19534__, new_new_n19535__, new_new_n19536__, new_new_n19537__,
    new_new_n19538__, new_new_n19539__, new_new_n19540__, new_new_n19541__,
    new_new_n19542__, new_new_n19543__, new_new_n19544__, new_new_n19545__,
    new_new_n19546__, new_new_n19547__, new_new_n19548__, new_new_n19549__,
    new_new_n19550__, new_new_n19551__, new_new_n19552__, new_new_n19553__,
    new_new_n19554__, new_new_n19555__, new_new_n19556__, new_new_n19557__,
    new_new_n19558__, new_new_n19559__, new_new_n19560__, new_new_n19561__,
    new_new_n19562__, new_new_n19563__, new_new_n19564__, new_new_n19565__,
    new_new_n19566__, new_new_n19567__, new_new_n19568__, new_new_n19569__,
    new_new_n19570__, new_new_n19571__, new_new_n19572__, new_new_n19573__,
    new_new_n19574__, new_new_n19575__, new_new_n19576__, new_new_n19577__,
    new_new_n19578__, new_new_n19579__, new_new_n19580__, new_new_n19581__,
    new_new_n19582__, new_new_n19583__, new_new_n19584__, new_new_n19585__,
    new_new_n19586__, new_new_n19587__, new_new_n19588__, new_new_n19589__,
    new_new_n19590__, new_new_n19591__, new_new_n19592__, new_new_n19593__,
    new_new_n19595__, new_new_n19596__, new_new_n19597__, new_new_n19598__,
    new_new_n19599__, new_new_n19600__, new_new_n19601__, new_new_n19602__,
    new_new_n19603__, new_new_n19604__, new_new_n19605__, new_new_n19606__,
    new_new_n19607__, new_new_n19608__, new_new_n19609__, new_new_n19610__,
    new_new_n19611__, new_new_n19612__, new_new_n19613__, new_new_n19614__,
    new_new_n19615__, new_new_n19616__, new_new_n19617__, new_new_n19618__,
    new_new_n19619__, new_new_n19620__, new_new_n19621__, new_new_n19622__,
    new_new_n19623__, new_new_n19624__, new_new_n19625__, new_new_n19626__,
    new_new_n19627__, new_new_n19628__, new_new_n19629__, new_new_n19630__,
    new_new_n19631__, new_new_n19632__, new_new_n19633__, new_new_n19634__,
    new_new_n19635__, new_new_n19636__, new_new_n19637__, new_new_n19638__,
    new_new_n19639__, new_new_n19640__, new_new_n19641__, new_new_n19642__,
    new_new_n19643__, new_new_n19644__, new_new_n19645__, new_new_n19646__,
    new_new_n19647__, new_new_n19648__, new_new_n19649__, new_new_n19650__,
    new_new_n19651__, new_new_n19652__, new_new_n19653__, new_new_n19654__,
    new_new_n19655__, new_new_n19656__, new_new_n19657__, new_new_n19658__,
    new_new_n19659__, new_new_n19660__, new_new_n19661__, new_new_n19662__,
    new_new_n19663__, new_new_n19664__, new_new_n19665__, new_new_n19666__,
    new_new_n19667__, new_new_n19668__, new_new_n19669__, new_new_n19670__,
    new_new_n19671__, new_new_n19672__, new_new_n19673__, new_new_n19675__,
    new_new_n19676__, new_new_n19677__, new_new_n19678__, new_new_n19679__,
    new_new_n19680__, new_new_n19681__, new_new_n19682__, new_new_n19683__,
    new_new_n19684__, new_new_n19685__, new_new_n19686__, new_new_n19687__,
    new_new_n19688__, new_new_n19689__, new_new_n19690__, new_new_n19691__,
    new_new_n19692__, new_new_n19693__, new_new_n19694__, new_new_n19695__,
    new_new_n19696__, new_new_n19697__, new_new_n19698__, new_new_n19699__,
    new_new_n19700__, new_new_n19701__, new_new_n19702__, new_new_n19703__,
    new_new_n19704__, new_new_n19705__, new_new_n19706__, new_new_n19707__,
    new_new_n19708__, new_new_n19709__, new_new_n19710__, new_new_n19711__,
    new_new_n19712__, new_new_n19713__, new_new_n19714__, new_new_n19715__,
    new_new_n19716__, new_new_n19717__, new_new_n19718__, new_new_n19719__,
    new_new_n19720__, new_new_n19721__, new_new_n19722__, new_new_n19723__,
    new_new_n19724__, new_new_n19725__, new_new_n19726__, new_new_n19727__,
    new_new_n19728__, new_new_n19729__, new_new_n19730__, new_new_n19731__,
    new_new_n19732__, new_new_n19733__, new_new_n19734__, new_new_n19735__,
    new_new_n19736__, new_new_n19737__, new_new_n19738__, new_new_n19739__,
    new_new_n19740__, new_new_n19741__, new_new_n19742__, new_new_n19743__,
    new_new_n19744__, new_new_n19745__, new_new_n19746__, new_new_n19747__,
    new_new_n19748__, new_new_n19749__, new_new_n19750__, new_new_n19751__,
    new_new_n19752__, new_new_n19753__, new_new_n19754__, new_new_n19755__,
    new_new_n19756__, new_new_n19757__, new_new_n19758__, new_new_n19759__,
    new_new_n19760__, new_new_n19761__, new_new_n19762__, new_new_n19763__,
    new_new_n19765__, new_new_n19766__, new_new_n19767__, new_new_n19768__,
    new_new_n19769__, new_new_n19770__, new_new_n19771__, new_new_n19772__,
    new_new_n19773__, new_new_n19774__, new_new_n19775__, new_new_n19776__,
    new_new_n19777__, new_new_n19778__, new_new_n19779__, new_new_n19780__,
    new_new_n19781__, new_new_n19782__, new_new_n19783__, new_new_n19784__,
    new_new_n19785__, new_new_n19786__, new_new_n19787__, new_new_n19788__,
    new_new_n19789__, new_new_n19790__, new_new_n19791__, new_new_n19792__,
    new_new_n19793__, new_new_n19794__, new_new_n19795__, new_new_n19796__,
    new_new_n19797__, new_new_n19798__, new_new_n19799__, new_new_n19800__,
    new_new_n19801__, new_new_n19802__, new_new_n19803__, new_new_n19804__,
    new_new_n19805__, new_new_n19806__, new_new_n19807__, new_new_n19808__,
    new_new_n19809__, new_new_n19810__, new_new_n19811__, new_new_n19812__,
    new_new_n19813__, new_new_n19814__, new_new_n19815__, new_new_n19816__,
    new_new_n19817__, new_new_n19818__, new_new_n19819__, new_new_n19820__,
    new_new_n19821__, new_new_n19822__, new_new_n19823__, new_new_n19824__,
    new_new_n19825__, new_new_n19826__, new_new_n19827__, new_new_n19828__,
    new_new_n19830__, new_new_n19831__, new_new_n19832__, new_new_n19833__,
    new_new_n19834__, new_new_n19835__, new_new_n19836__, new_new_n19837__,
    new_new_n19838__, new_new_n19839__, new_new_n19840__, new_new_n19841__,
    new_new_n19842__, new_new_n19843__, new_new_n19844__, new_new_n19845__,
    new_new_n19846__, new_new_n19847__, new_new_n19848__, new_new_n19849__,
    new_new_n19850__, new_new_n19851__, new_new_n19852__, new_new_n19853__,
    new_new_n19854__, new_new_n19855__, new_new_n19856__, new_new_n19857__,
    new_new_n19858__, new_new_n19859__, new_new_n19860__, new_new_n19861__,
    new_new_n19862__, new_new_n19863__, new_new_n19864__, new_new_n19865__,
    new_new_n19866__, new_new_n19867__, new_new_n19868__, new_new_n19869__,
    new_new_n19870__, new_new_n19871__, new_new_n19872__, new_new_n19873__,
    new_new_n19874__, new_new_n19875__, new_new_n19876__, new_new_n19877__,
    new_new_n19878__, new_new_n19879__, new_new_n19880__, new_new_n19881__,
    new_new_n19882__, new_new_n19883__, new_new_n19884__, new_new_n19885__,
    new_new_n19886__, new_new_n19887__, new_new_n19888__, new_new_n19889__,
    new_new_n19890__, new_new_n19891__, new_new_n19892__, new_new_n19893__,
    new_new_n19894__, new_new_n19895__, new_new_n19896__, new_new_n19897__,
    new_new_n19898__, new_new_n19900__, new_new_n19901__, new_new_n19902__,
    new_new_n19903__, new_new_n19904__, new_new_n19905__, new_new_n19906__,
    new_new_n19907__, new_new_n19908__, new_new_n19909__, new_new_n19910__,
    new_new_n19911__, new_new_n19912__, new_new_n19913__, new_new_n19914__,
    new_new_n19915__, new_new_n19916__, new_new_n19917__, new_new_n19918__,
    new_new_n19919__, new_new_n19920__, new_new_n19921__, new_new_n19922__,
    new_new_n19923__, new_new_n19924__, new_new_n19925__, new_new_n19926__,
    new_new_n19927__, new_new_n19928__, new_new_n19929__, new_new_n19930__,
    new_new_n19931__, new_new_n19932__, new_new_n19933__, new_new_n19934__,
    new_new_n19935__, new_new_n19936__, new_new_n19937__, new_new_n19938__,
    new_new_n19939__, new_new_n19940__, new_new_n19941__, new_new_n19942__,
    new_new_n19943__, new_new_n19944__, new_new_n19945__, new_new_n19946__,
    new_new_n19947__, new_new_n19948__, new_new_n19949__, new_new_n19950__,
    new_new_n19951__, new_new_n19952__, new_new_n19953__, new_new_n19955__,
    new_new_n19956__, new_new_n19957__, new_new_n19958__, new_new_n19959__,
    new_new_n19960__, new_new_n19961__, new_new_n19962__, new_new_n19963__,
    new_new_n19964__, new_new_n19965__, new_new_n19966__, new_new_n19967__,
    new_new_n19968__, new_new_n19969__, new_new_n19970__, new_new_n19971__,
    new_new_n19972__, new_new_n19973__, new_new_n19974__, new_new_n19975__,
    new_new_n19976__, new_new_n19977__, new_new_n19978__, new_new_n19979__,
    new_new_n19980__, new_new_n19981__, new_new_n19982__, new_new_n19983__,
    new_new_n19984__, new_new_n19985__, new_new_n19986__, new_new_n19987__,
    new_new_n19988__, new_new_n19989__, new_new_n19990__, new_new_n19991__,
    new_new_n19992__, new_new_n19993__, new_new_n19994__, new_new_n19995__,
    new_new_n19996__, new_new_n19997__, new_new_n19998__, new_new_n19999__,
    new_new_n20000__, new_new_n20001__, new_new_n20002__, new_new_n20003__,
    new_new_n20004__, new_new_n20005__, new_new_n20006__, new_new_n20007__,
    new_new_n20008__, new_new_n20009__, new_new_n20010__, new_new_n20011__,
    new_new_n20012__, new_new_n20013__, new_new_n20014__, new_new_n20015__,
    new_new_n20016__, new_new_n20018__, new_new_n20019__, new_new_n20020__,
    new_new_n20021__, new_new_n20022__, new_new_n20023__, new_new_n20024__,
    new_new_n20025__, new_new_n20026__, new_new_n20027__, new_new_n20028__,
    new_new_n20029__, new_new_n20030__, new_new_n20031__, new_new_n20032__,
    new_new_n20033__, new_new_n20034__, new_new_n20035__, new_new_n20036__,
    new_new_n20037__, new_new_n20038__, new_new_n20039__, new_new_n20040__,
    new_new_n20041__, new_new_n20042__, new_new_n20043__, new_new_n20044__,
    new_new_n20045__, new_new_n20046__, new_new_n20047__, new_new_n20048__,
    new_new_n20049__, new_new_n20050__, new_new_n20051__, new_new_n20052__,
    new_new_n20053__, new_new_n20054__, new_new_n20055__, new_new_n20056__,
    new_new_n20057__, new_new_n20058__, new_new_n20059__, new_new_n20060__,
    new_new_n20061__, new_new_n20062__, new_new_n20063__, new_new_n20064__,
    new_new_n20066__, new_new_n20067__, new_new_n20068__, new_new_n20069__,
    new_new_n20070__, new_new_n20071__, new_new_n20072__, new_new_n20073__,
    new_new_n20074__, new_new_n20075__, new_new_n20076__, new_new_n20077__,
    new_new_n20078__, new_new_n20079__, new_new_n20080__, new_new_n20081__,
    new_new_n20082__, new_new_n20083__, new_new_n20084__, new_new_n20085__,
    new_new_n20086__, new_new_n20087__, new_new_n20088__, new_new_n20089__,
    new_new_n20090__, new_new_n20091__, new_new_n20092__, new_new_n20093__,
    new_new_n20094__, new_new_n20095__, new_new_n20096__, new_new_n20097__,
    new_new_n20098__, new_new_n20099__, new_new_n20100__, new_new_n20101__,
    new_new_n20102__, new_new_n20104__, new_new_n20105__, new_new_n20106__,
    new_new_n20107__, new_new_n20108__, new_new_n20109__, new_new_n20110__,
    new_new_n20111__, new_new_n20112__, new_new_n20113__, new_new_n20114__,
    new_new_n20115__, new_new_n20116__, new_new_n20117__, new_new_n20118__,
    new_new_n20119__, new_new_n20120__, new_new_n20121__, new_new_n20122__,
    new_new_n20123__, new_new_n20124__, new_new_n20125__, new_new_n20126__,
    new_new_n20127__, new_new_n20128__, new_new_n20129__, new_new_n20130__,
    new_new_n20131__, new_new_n20132__, new_new_n20133__, new_new_n20134__,
    new_new_n20135__, new_new_n20136__, new_new_n20137__, new_new_n20138__,
    new_new_n20139__, new_new_n20140__, new_new_n20141__, new_new_n20142__,
    new_new_n20143__, new_new_n20144__, new_new_n20145__, new_new_n20146__,
    new_new_n20147__, new_new_n20148__, new_new_n20149__, new_new_n20150__,
    new_new_n20151__, new_new_n20152__, new_new_n20153__, new_new_n20154__,
    new_new_n20155__, new_new_n20156__, new_new_n20157__, new_new_n20159__,
    new_new_n20160__, new_new_n20161__, new_new_n20162__, new_new_n20163__,
    new_new_n20164__, new_new_n20165__, new_new_n20166__, new_new_n20167__,
    new_new_n20168__, new_new_n20169__, new_new_n20170__, new_new_n20171__,
    new_new_n20172__, new_new_n20173__, new_new_n20174__, new_new_n20175__,
    new_new_n20176__, new_new_n20177__, new_new_n20178__, new_new_n20179__,
    new_new_n20180__, new_new_n20181__, new_new_n20182__, new_new_n20183__,
    new_new_n20184__, new_new_n20185__, new_new_n20186__, new_new_n20187__,
    new_new_n20188__, new_new_n20189__, new_new_n20190__, new_new_n20191__,
    new_new_n20192__, new_new_n20194__, new_new_n20195__, new_new_n20196__,
    new_new_n20197__, new_new_n20198__, new_new_n20199__, new_new_n20200__,
    new_new_n20201__, new_new_n20202__, new_new_n20203__, new_new_n20204__,
    new_new_n20205__, new_new_n20206__, new_new_n20207__, new_new_n20208__,
    new_new_n20209__, new_new_n20210__, new_new_n20211__, new_new_n20212__,
    new_new_n20213__, new_new_n20215__, new_new_n20216__, new_new_n20217__,
    new_new_n20218__, new_new_n20219__, new_new_n20220__, new_new_n20221__;
  assign po002 = ~pi00 & pi01;
  assign new_new_n195__ = ~pi01 & pi02;
  assign new_new_n196__ = pi01 & ~pi02;
  assign new_new_n197__ = ~new_new_n195__ & ~new_new_n196__;
  assign po003 = pi00 & ~new_new_n197__;
  assign new_new_n199__ = pi02 & pi03;
  assign new_new_n200__ = ~pi02 & ~pi03;
  assign new_new_n201__ = ~new_new_n199__ & ~new_new_n200__;
  assign new_new_n202__ = pi00 & new_new_n201__;
  assign new_new_n203__ = ~pi00 & ~pi01;
  assign new_new_n204__ = pi02 & new_new_n203__;
  assign po004 = new_new_n202__ | new_new_n204__;
  assign new_new_n206__ = pi00 & pi04;
  assign new_new_n207__ = pi01 & new_new_n201__;
  assign new_new_n208__ = pi00 & pi03;
  assign new_new_n209__ = pi02 & new_new_n208__;
  assign new_new_n210__ = ~new_new_n207__ & ~new_new_n209__;
  assign new_new_n211__ = new_new_n206__ & ~new_new_n210__;
  assign new_new_n212__ = ~new_new_n206__ & new_new_n210__;
  assign po005 = ~new_new_n211__ & ~new_new_n212__;
  assign new_new_n214__ = ~pi03 & pi04;
  assign new_new_n215__ = pi03 & ~pi04;
  assign new_new_n216__ = ~new_new_n214__ & ~new_new_n215__;
  assign new_new_n217__ = ~pi00 & ~new_new_n216__;
  assign new_new_n218__ = ~pi02 & new_new_n214__;
  assign new_new_n219__ = ~new_new_n215__ & ~new_new_n218__;
  assign new_new_n220__ = ~pi05 & ~new_new_n219__;
  assign new_new_n221__ = ~new_new_n217__ & ~new_new_n220__;
  assign new_new_n222__ = pi01 & ~new_new_n221__;
  assign new_new_n223__ = pi01 & pi04;
  assign new_new_n224__ = ~pi03 & new_new_n223__;
  assign new_new_n225__ = pi00 & ~pi01;
  assign new_new_n226__ = ~pi04 & new_new_n225__;
  assign new_new_n227__ = ~new_new_n224__ & ~new_new_n226__;
  assign new_new_n228__ = pi02 & ~new_new_n227__;
  assign new_new_n229__ = pi00 & ~pi03;
  assign new_new_n230__ = ~new_new_n223__ & new_new_n229__;
  assign new_new_n231__ = ~new_new_n228__ & ~new_new_n230__;
  assign new_new_n232__ = pi05 & ~new_new_n231__;
  assign new_new_n233__ = ~pi02 & ~pi04;
  assign new_new_n234__ = ~new_new_n206__ & ~new_new_n233__;
  assign new_new_n235__ = ~pi05 & ~new_new_n234__;
  assign new_new_n236__ = ~pi02 & new_new_n203__;
  assign new_new_n237__ = ~new_new_n235__ & ~new_new_n236__;
  assign new_new_n238__ = pi03 & ~new_new_n237__;
  assign new_new_n239__ = ~new_new_n222__ & ~new_new_n238__;
  assign po006 = new_new_n232__ | ~new_new_n239__;
  assign new_new_n241__ = pi02 & ~new_new_n216__;
  assign new_new_n242__ = pi01 & pi05;
  assign new_new_n243__ = pi00 & pi06;
  assign new_new_n244__ = new_new_n242__ & new_new_n243__;
  assign new_new_n245__ = ~new_new_n242__ & ~new_new_n243__;
  assign new_new_n246__ = ~new_new_n244__ & ~new_new_n245__;
  assign new_new_n247__ = new_new_n241__ & ~new_new_n246__;
  assign new_new_n248__ = ~new_new_n241__ & new_new_n246__;
  assign new_new_n249__ = ~new_new_n247__ & ~new_new_n248__;
  assign new_new_n250__ = ~pi03 & ~pi05;
  assign new_new_n251__ = pi00 & new_new_n223__;
  assign new_new_n252__ = ~new_new_n250__ & new_new_n251__;
  assign new_new_n253__ = ~new_new_n249__ & new_new_n252__;
  assign new_new_n254__ = new_new_n249__ & ~new_new_n252__;
  assign new_new_n255__ = ~new_new_n253__ & ~new_new_n254__;
  assign new_new_n256__ = pi03 & pi05;
  assign new_new_n257__ = ~pi04 & new_new_n195__;
  assign new_new_n258__ = pi00 & new_new_n256__;
  assign new_new_n259__ = ~new_new_n257__ & new_new_n258__;
  assign new_new_n260__ = pi00 & pi02;
  assign new_new_n261__ = ~pi05 & new_new_n260__;
  assign new_new_n262__ = ~pi03 & ~new_new_n261__;
  assign new_new_n263__ = ~new_new_n208__ & new_new_n223__;
  assign new_new_n264__ = ~new_new_n262__ & new_new_n263__;
  assign new_new_n265__ = ~new_new_n259__ & ~new_new_n264__;
  assign new_new_n266__ = new_new_n255__ & new_new_n265__;
  assign new_new_n267__ = ~new_new_n255__ & ~new_new_n265__;
  assign po007 = new_new_n266__ | new_new_n267__;
  assign new_new_n269__ = pi03 & pi04;
  assign new_new_n270__ = pi02 & pi05;
  assign new_new_n271__ = pi00 & pi07;
  assign new_new_n272__ = ~new_new_n270__ & ~new_new_n271__;
  assign new_new_n273__ = new_new_n270__ & new_new_n271__;
  assign new_new_n274__ = ~new_new_n272__ & ~new_new_n273__;
  assign new_new_n275__ = new_new_n269__ & ~new_new_n274__;
  assign new_new_n276__ = ~new_new_n269__ & new_new_n274__;
  assign new_new_n277__ = ~new_new_n275__ & ~new_new_n276__;
  assign new_new_n278__ = pi04 & ~new_new_n243__;
  assign new_new_n279__ = pi03 & ~new_new_n245__;
  assign new_new_n280__ = ~new_new_n278__ & new_new_n279__;
  assign new_new_n281__ = ~pi03 & ~new_new_n243__;
  assign new_new_n282__ = pi04 & ~new_new_n242__;
  assign new_new_n283__ = ~new_new_n281__ & new_new_n282__;
  assign new_new_n284__ = ~new_new_n280__ & ~new_new_n283__;
  assign new_new_n285__ = pi02 & ~new_new_n284__;
  assign new_new_n286__ = pi02 & pi04;
  assign new_new_n287__ = new_new_n244__ & ~new_new_n286__;
  assign new_new_n288__ = ~new_new_n285__ & ~new_new_n287__;
  assign new_new_n289__ = pi06 & new_new_n288__;
  assign new_new_n290__ = pi01 & pi06;
  assign new_new_n291__ = ~new_new_n288__ & ~new_new_n290__;
  assign new_new_n292__ = ~pi05 & ~new_new_n291__;
  assign new_new_n293__ = ~new_new_n289__ & new_new_n292__;
  assign new_new_n294__ = ~pi02 & ~new_new_n289__;
  assign new_new_n295__ = pi05 & pi06;
  assign new_new_n296__ = pi02 & new_new_n295__;
  assign new_new_n297__ = pi01 & ~new_new_n296__;
  assign new_new_n298__ = new_new_n288__ & ~new_new_n297__;
  assign new_new_n299__ = pi04 & ~new_new_n298__;
  assign new_new_n300__ = ~new_new_n294__ & new_new_n299__;
  assign new_new_n301__ = ~new_new_n293__ & new_new_n300__;
  assign new_new_n302__ = new_new_n288__ & new_new_n290__;
  assign new_new_n303__ = ~pi04 & ~new_new_n291__;
  assign new_new_n304__ = ~new_new_n302__ & new_new_n303__;
  assign new_new_n305__ = ~new_new_n301__ & ~new_new_n304__;
  assign new_new_n306__ = new_new_n277__ & ~new_new_n305__;
  assign new_new_n307__ = ~new_new_n277__ & new_new_n305__;
  assign new_new_n308__ = ~new_new_n306__ & ~new_new_n307__;
  assign new_new_n309__ = ~new_new_n254__ & ~new_new_n265__;
  assign new_new_n310__ = ~new_new_n253__ & ~new_new_n309__;
  assign new_new_n311__ = new_new_n308__ & new_new_n310__;
  assign new_new_n312__ = ~new_new_n308__ & ~new_new_n310__;
  assign po008 = new_new_n311__ | new_new_n312__;
  assign new_new_n314__ = ~new_new_n306__ & ~new_new_n310__;
  assign new_new_n315__ = ~new_new_n307__ & ~new_new_n314__;
  assign new_new_n316__ = pi01 & ~pi06;
  assign new_new_n317__ = new_new_n288__ & ~new_new_n316__;
  assign new_new_n318__ = new_new_n286__ & ~new_new_n317__;
  assign new_new_n319__ = ~new_new_n292__ & new_new_n318__;
  assign new_new_n320__ = ~pi04 & new_new_n290__;
  assign new_new_n321__ = ~new_new_n288__ & new_new_n320__;
  assign new_new_n322__ = ~new_new_n319__ & ~new_new_n321__;
  assign new_new_n323__ = new_new_n315__ & new_new_n322__;
  assign new_new_n324__ = ~new_new_n315__ & ~new_new_n322__;
  assign new_new_n325__ = ~new_new_n323__ & ~new_new_n324__;
  assign new_new_n326__ = ~new_new_n269__ & ~new_new_n273__;
  assign new_new_n327__ = ~new_new_n272__ & ~new_new_n326__;
  assign new_new_n328__ = pi01 & pi07;
  assign new_new_n329__ = ~new_new_n256__ & new_new_n328__;
  assign new_new_n330__ = new_new_n256__ & ~new_new_n328__;
  assign new_new_n331__ = ~new_new_n329__ & ~new_new_n330__;
  assign new_new_n332__ = ~new_new_n327__ & new_new_n331__;
  assign new_new_n333__ = new_new_n327__ & ~new_new_n331__;
  assign new_new_n334__ = ~new_new_n332__ & ~new_new_n333__;
  assign new_new_n335__ = new_new_n325__ & ~new_new_n334__;
  assign new_new_n336__ = ~new_new_n325__ & ~new_new_n333__;
  assign new_new_n337__ = ~new_new_n335__ & ~new_new_n336__;
  assign new_new_n338__ = new_new_n323__ & new_new_n332__;
  assign new_new_n339__ = ~new_new_n337__ & ~new_new_n338__;
  assign new_new_n340__ = pi00 & pi08;
  assign new_new_n341__ = pi02 & new_new_n223__;
  assign new_new_n342__ = ~pi02 & ~new_new_n223__;
  assign new_new_n343__ = pi06 & ~new_new_n342__;
  assign new_new_n344__ = ~new_new_n341__ & new_new_n343__;
  assign new_new_n345__ = new_new_n340__ & ~new_new_n344__;
  assign new_new_n346__ = ~new_new_n340__ & new_new_n344__;
  assign new_new_n347__ = ~new_new_n345__ & ~new_new_n346__;
  assign new_new_n348__ = ~new_new_n339__ & ~new_new_n347__;
  assign new_new_n349__ = new_new_n324__ & ~new_new_n327__;
  assign new_new_n350__ = ~new_new_n325__ & new_new_n334__;
  assign new_new_n351__ = ~new_new_n335__ & ~new_new_n349__;
  assign new_new_n352__ = ~new_new_n350__ & new_new_n351__;
  assign new_new_n353__ = new_new_n347__ & ~new_new_n352__;
  assign po009 = new_new_n348__ | new_new_n353__;
  assign new_new_n355__ = ~new_new_n323__ & ~new_new_n347__;
  assign new_new_n356__ = ~new_new_n324__ & ~new_new_n355__;
  assign new_new_n357__ = new_new_n333__ & ~new_new_n356__;
  assign new_new_n358__ = new_new_n324__ & ~new_new_n347__;
  assign new_new_n359__ = new_new_n323__ & new_new_n347__;
  assign new_new_n360__ = ~new_new_n327__ & new_new_n359__;
  assign new_new_n361__ = new_new_n327__ & ~new_new_n359__;
  assign new_new_n362__ = new_new_n331__ & ~new_new_n355__;
  assign new_new_n363__ = ~new_new_n361__ & new_new_n362__;
  assign new_new_n364__ = ~new_new_n358__ & ~new_new_n360__;
  assign new_new_n365__ = ~new_new_n357__ & new_new_n364__;
  assign new_new_n366__ = ~new_new_n363__ & new_new_n365__;
  assign new_new_n367__ = ~new_new_n340__ & ~new_new_n341__;
  assign new_new_n368__ = new_new_n343__ & ~new_new_n367__;
  assign new_new_n369__ = pi04 & pi05;
  assign new_new_n370__ = pi03 & pi06;
  assign new_new_n371__ = pi02 & pi07;
  assign new_new_n372__ = ~new_new_n370__ & ~new_new_n371__;
  assign new_new_n373__ = new_new_n370__ & new_new_n371__;
  assign new_new_n374__ = ~new_new_n372__ & ~new_new_n373__;
  assign new_new_n375__ = new_new_n369__ & ~new_new_n374__;
  assign new_new_n376__ = ~new_new_n369__ & new_new_n374__;
  assign new_new_n377__ = ~new_new_n375__ & ~new_new_n376__;
  assign new_new_n378__ = pi00 & pi09;
  assign new_new_n379__ = pi05 & pi08;
  assign new_new_n380__ = ~new_new_n378__ & ~new_new_n379__;
  assign new_new_n381__ = pi03 & pi07;
  assign new_new_n382__ = pi01 & ~pi08;
  assign new_new_n383__ = new_new_n378__ & ~new_new_n382__;
  assign new_new_n384__ = ~new_new_n380__ & new_new_n381__;
  assign new_new_n385__ = ~new_new_n383__ & new_new_n384__;
  assign new_new_n386__ = new_new_n242__ & new_new_n381__;
  assign new_new_n387__ = pi01 & pi08;
  assign new_new_n388__ = ~new_new_n378__ & new_new_n387__;
  assign new_new_n389__ = new_new_n378__ & ~new_new_n387__;
  assign new_new_n390__ = ~new_new_n388__ & ~new_new_n389__;
  assign new_new_n391__ = pi05 & ~new_new_n390__;
  assign new_new_n392__ = ~pi05 & new_new_n390__;
  assign new_new_n393__ = ~new_new_n386__ & ~new_new_n391__;
  assign new_new_n394__ = ~new_new_n392__ & new_new_n393__;
  assign new_new_n395__ = ~new_new_n385__ & ~new_new_n394__;
  assign new_new_n396__ = ~new_new_n377__ & ~new_new_n395__;
  assign new_new_n397__ = new_new_n377__ & new_new_n395__;
  assign new_new_n398__ = ~new_new_n396__ & ~new_new_n397__;
  assign new_new_n399__ = new_new_n368__ & new_new_n398__;
  assign new_new_n400__ = ~new_new_n368__ & ~new_new_n398__;
  assign new_new_n401__ = ~new_new_n399__ & ~new_new_n400__;
  assign new_new_n402__ = ~new_new_n366__ & new_new_n401__;
  assign new_new_n403__ = ~new_new_n323__ & ~new_new_n331__;
  assign new_new_n404__ = ~new_new_n327__ & new_new_n347__;
  assign new_new_n405__ = new_new_n403__ & new_new_n404__;
  assign new_new_n406__ = new_new_n327__ & ~new_new_n347__;
  assign new_new_n407__ = ~new_new_n324__ & new_new_n406__;
  assign new_new_n408__ = ~new_new_n403__ & new_new_n407__;
  assign new_new_n409__ = new_new_n324__ & ~new_new_n331__;
  assign new_new_n410__ = new_new_n323__ & new_new_n331__;
  assign new_new_n411__ = ~new_new_n404__ & ~new_new_n406__;
  assign new_new_n412__ = ~new_new_n409__ & new_new_n411__;
  assign new_new_n413__ = ~new_new_n410__ & new_new_n412__;
  assign new_new_n414__ = ~new_new_n405__ & ~new_new_n408__;
  assign new_new_n415__ = ~new_new_n413__ & new_new_n414__;
  assign new_new_n416__ = ~new_new_n401__ & ~new_new_n415__;
  assign po010 = new_new_n402__ | new_new_n416__;
  assign new_new_n418__ = ~new_new_n333__ & new_new_n347__;
  assign new_new_n419__ = ~new_new_n315__ & ~new_new_n418__;
  assign new_new_n420__ = ~new_new_n333__ & ~new_new_n401__;
  assign new_new_n421__ = ~new_new_n332__ & new_new_n401__;
  assign new_new_n422__ = new_new_n347__ & ~new_new_n421__;
  assign new_new_n423__ = ~new_new_n420__ & ~new_new_n422__;
  assign new_new_n424__ = ~new_new_n419__ & ~new_new_n423__;
  assign new_new_n425__ = ~new_new_n322__ & ~new_new_n424__;
  assign new_new_n426__ = ~new_new_n315__ & new_new_n423__;
  assign new_new_n427__ = ~new_new_n418__ & new_new_n421__;
  assign new_new_n428__ = ~new_new_n426__ & ~new_new_n427__;
  assign new_new_n429__ = ~new_new_n425__ & new_new_n428__;
  assign new_new_n430__ = new_new_n368__ & ~new_new_n397__;
  assign new_new_n431__ = ~new_new_n396__ & ~new_new_n430__;
  assign new_new_n432__ = ~new_new_n429__ & ~new_new_n431__;
  assign new_new_n433__ = new_new_n429__ & new_new_n431__;
  assign new_new_n434__ = ~new_new_n432__ & ~new_new_n433__;
  assign new_new_n435__ = pi04 & pi06;
  assign new_new_n436__ = ~new_new_n369__ & ~new_new_n373__;
  assign new_new_n437__ = ~new_new_n372__ & ~new_new_n436__;
  assign new_new_n438__ = new_new_n435__ & new_new_n437__;
  assign new_new_n439__ = ~new_new_n435__ & ~new_new_n437__;
  assign new_new_n440__ = ~new_new_n438__ & ~new_new_n439__;
  assign new_new_n441__ = ~pi09 & ~new_new_n379__;
  assign new_new_n442__ = pi05 & pi09;
  assign new_new_n443__ = pi08 & new_new_n442__;
  assign new_new_n444__ = pi01 & ~new_new_n441__;
  assign new_new_n445__ = ~new_new_n443__ & new_new_n444__;
  assign new_new_n446__ = new_new_n440__ & ~new_new_n445__;
  assign new_new_n447__ = ~new_new_n440__ & new_new_n445__;
  assign new_new_n448__ = ~new_new_n446__ & ~new_new_n447__;
  assign new_new_n449__ = ~new_new_n378__ & ~new_new_n382__;
  assign new_new_n450__ = new_new_n381__ & ~new_new_n449__;
  assign new_new_n451__ = ~new_new_n389__ & ~new_new_n450__;
  assign new_new_n452__ = pi05 & ~new_new_n451__;
  assign new_new_n453__ = ~pi05 & new_new_n378__;
  assign new_new_n454__ = new_new_n387__ & new_new_n453__;
  assign new_new_n455__ = ~new_new_n452__ & ~new_new_n454__;
  assign new_new_n456__ = new_new_n448__ & new_new_n455__;
  assign new_new_n457__ = ~new_new_n448__ & ~new_new_n455__;
  assign new_new_n458__ = ~new_new_n456__ & ~new_new_n457__;
  assign new_new_n459__ = pi02 & pi08;
  assign new_new_n460__ = pi00 & pi10;
  assign new_new_n461__ = ~new_new_n459__ & ~new_new_n460__;
  assign new_new_n462__ = new_new_n459__ & new_new_n460__;
  assign new_new_n463__ = ~new_new_n461__ & ~new_new_n462__;
  assign new_new_n464__ = new_new_n381__ & ~new_new_n463__;
  assign new_new_n465__ = ~new_new_n381__ & new_new_n463__;
  assign new_new_n466__ = ~new_new_n464__ & ~new_new_n465__;
  assign new_new_n467__ = new_new_n458__ & ~new_new_n466__;
  assign new_new_n468__ = ~new_new_n458__ & new_new_n466__;
  assign new_new_n469__ = ~new_new_n467__ & ~new_new_n468__;
  assign new_new_n470__ = new_new_n434__ & new_new_n469__;
  assign new_new_n471__ = ~new_new_n434__ & ~new_new_n469__;
  assign po011 = ~new_new_n470__ & ~new_new_n471__;
  assign new_new_n473__ = ~new_new_n381__ & ~new_new_n462__;
  assign new_new_n474__ = ~new_new_n461__ & ~new_new_n473__;
  assign new_new_n475__ = pi03 & pi08;
  assign new_new_n476__ = pi06 & new_new_n223__;
  assign new_new_n477__ = ~pi02 & ~new_new_n476__;
  assign new_new_n478__ = pi09 & ~new_new_n477__;
  assign new_new_n479__ = pi06 & new_new_n341__;
  assign new_new_n480__ = new_new_n478__ & ~new_new_n479__;
  assign new_new_n481__ = new_new_n475__ & ~new_new_n480__;
  assign new_new_n482__ = ~new_new_n475__ & new_new_n480__;
  assign new_new_n483__ = ~new_new_n481__ & ~new_new_n482__;
  assign new_new_n484__ = new_new_n474__ & ~new_new_n483__;
  assign new_new_n485__ = ~new_new_n474__ & new_new_n483__;
  assign new_new_n486__ = ~new_new_n484__ & ~new_new_n485__;
  assign new_new_n487__ = ~new_new_n379__ & ~new_new_n437__;
  assign new_new_n488__ = pi09 & ~new_new_n435__;
  assign new_new_n489__ = ~new_new_n487__ & new_new_n488__;
  assign new_new_n490__ = ~pi09 & new_new_n435__;
  assign new_new_n491__ = ~new_new_n437__ & ~new_new_n490__;
  assign new_new_n492__ = new_new_n379__ & ~new_new_n491__;
  assign new_new_n493__ = ~new_new_n489__ & ~new_new_n492__;
  assign new_new_n494__ = pi01 & ~new_new_n493__;
  assign new_new_n495__ = pi01 & pi09;
  assign new_new_n496__ = new_new_n438__ & ~new_new_n495__;
  assign new_new_n497__ = ~new_new_n494__ & ~new_new_n496__;
  assign new_new_n498__ = pi01 & pi10;
  assign new_new_n499__ = new_new_n497__ & ~new_new_n498__;
  assign new_new_n500__ = ~new_new_n497__ & new_new_n498__;
  assign new_new_n501__ = ~new_new_n499__ & ~new_new_n500__;
  assign new_new_n502__ = new_new_n486__ & ~new_new_n501__;
  assign new_new_n503__ = ~new_new_n486__ & new_new_n501__;
  assign new_new_n504__ = ~new_new_n502__ & ~new_new_n503__;
  assign new_new_n505__ = pi04 & pi07;
  assign new_new_n506__ = pi00 & pi11;
  assign new_new_n507__ = ~new_new_n505__ & ~new_new_n506__;
  assign new_new_n508__ = new_new_n505__ & new_new_n506__;
  assign new_new_n509__ = ~new_new_n507__ & ~new_new_n508__;
  assign new_new_n510__ = new_new_n295__ & ~new_new_n509__;
  assign new_new_n511__ = ~new_new_n295__ & new_new_n509__;
  assign new_new_n512__ = ~new_new_n510__ & ~new_new_n511__;
  assign new_new_n513__ = pi06 & ~new_new_n512__;
  assign new_new_n514__ = ~pi06 & ~new_new_n509__;
  assign new_new_n515__ = ~new_new_n513__ & ~new_new_n514__;
  assign new_new_n516__ = new_new_n504__ & new_new_n515__;
  assign new_new_n517__ = ~new_new_n504__ & ~new_new_n515__;
  assign new_new_n518__ = ~new_new_n516__ & ~new_new_n517__;
  assign new_new_n519__ = ~new_new_n456__ & ~new_new_n466__;
  assign new_new_n520__ = ~new_new_n457__ & ~new_new_n519__;
  assign new_new_n521__ = ~new_new_n432__ & new_new_n520__;
  assign new_new_n522__ = ~new_new_n433__ & ~new_new_n520__;
  assign new_new_n523__ = ~new_new_n521__ & ~new_new_n522__;
  assign new_new_n524__ = new_new_n456__ & new_new_n466__;
  assign new_new_n525__ = new_new_n457__ & ~new_new_n466__;
  assign new_new_n526__ = ~new_new_n524__ & ~new_new_n525__;
  assign new_new_n527__ = new_new_n434__ & new_new_n526__;
  assign new_new_n528__ = ~new_new_n523__ & ~new_new_n527__;
  assign new_new_n529__ = new_new_n518__ & ~new_new_n528__;
  assign new_new_n530__ = new_new_n432__ & new_new_n457__;
  assign new_new_n531__ = new_new_n432__ & ~new_new_n448__;
  assign new_new_n532__ = ~new_new_n432__ & new_new_n448__;
  assign new_new_n533__ = ~new_new_n433__ & ~new_new_n455__;
  assign new_new_n534__ = ~new_new_n532__ & new_new_n533__;
  assign new_new_n535__ = ~new_new_n531__ & ~new_new_n534__;
  assign new_new_n536__ = ~new_new_n466__ & ~new_new_n535__;
  assign new_new_n537__ = new_new_n433__ & ~new_new_n457__;
  assign new_new_n538__ = new_new_n455__ & new_new_n532__;
  assign new_new_n539__ = ~new_new_n537__ & ~new_new_n538__;
  assign new_new_n540__ = new_new_n466__ & ~new_new_n539__;
  assign new_new_n541__ = new_new_n433__ & new_new_n456__;
  assign new_new_n542__ = ~new_new_n530__ & ~new_new_n541__;
  assign new_new_n543__ = ~new_new_n536__ & new_new_n542__;
  assign new_new_n544__ = ~new_new_n540__ & new_new_n543__;
  assign new_new_n545__ = ~new_new_n518__ & ~new_new_n544__;
  assign po012 = new_new_n529__ | new_new_n545__;
  assign new_new_n547__ = ~new_new_n518__ & ~new_new_n521__;
  assign new_new_n548__ = new_new_n432__ & ~new_new_n520__;
  assign new_new_n549__ = new_new_n518__ & ~new_new_n525__;
  assign new_new_n550__ = ~new_new_n524__ & ~new_new_n549__;
  assign new_new_n551__ = ~new_new_n433__ & new_new_n550__;
  assign new_new_n552__ = ~new_new_n548__ & ~new_new_n551__;
  assign new_new_n553__ = ~new_new_n547__ & new_new_n552__;
  assign new_new_n554__ = pi06 & ~new_new_n498__;
  assign new_new_n555__ = pi10 & new_new_n316__;
  assign new_new_n556__ = ~new_new_n554__ & ~new_new_n555__;
  assign new_new_n557__ = ~new_new_n485__ & ~new_new_n556__;
  assign new_new_n558__ = ~new_new_n484__ & ~new_new_n557__;
  assign new_new_n559__ = pi04 & pi08;
  assign new_new_n560__ = pi05 & pi07;
  assign new_new_n561__ = pi01 & pi11;
  assign new_new_n562__ = ~new_new_n560__ & ~new_new_n561__;
  assign new_new_n563__ = new_new_n560__ & new_new_n561__;
  assign new_new_n564__ = ~new_new_n562__ & ~new_new_n563__;
  assign new_new_n565__ = new_new_n559__ & new_new_n564__;
  assign new_new_n566__ = ~new_new_n559__ & ~new_new_n564__;
  assign new_new_n567__ = ~new_new_n565__ & ~new_new_n566__;
  assign new_new_n568__ = pi10 & new_new_n290__;
  assign new_new_n569__ = ~new_new_n567__ & new_new_n568__;
  assign new_new_n570__ = new_new_n567__ & ~new_new_n568__;
  assign new_new_n571__ = ~new_new_n569__ & ~new_new_n570__;
  assign new_new_n572__ = ~new_new_n558__ & ~new_new_n571__;
  assign new_new_n573__ = new_new_n558__ & new_new_n571__;
  assign new_new_n574__ = ~new_new_n572__ & ~new_new_n573__;
  assign new_new_n575__ = ~new_new_n295__ & ~new_new_n508__;
  assign new_new_n576__ = ~new_new_n507__ & ~new_new_n575__;
  assign new_new_n577__ = pi03 & pi09;
  assign new_new_n578__ = pi02 & pi10;
  assign new_new_n579__ = pi00 & pi12;
  assign new_new_n580__ = ~new_new_n578__ & ~new_new_n579__;
  assign new_new_n581__ = new_new_n578__ & new_new_n579__;
  assign new_new_n582__ = ~new_new_n580__ & ~new_new_n581__;
  assign new_new_n583__ = new_new_n577__ & ~new_new_n582__;
  assign new_new_n584__ = ~new_new_n577__ & new_new_n582__;
  assign new_new_n585__ = ~new_new_n583__ & ~new_new_n584__;
  assign new_new_n586__ = new_new_n576__ & ~new_new_n585__;
  assign new_new_n587__ = ~new_new_n576__ & new_new_n585__;
  assign new_new_n588__ = ~new_new_n586__ & ~new_new_n587__;
  assign new_new_n589__ = ~new_new_n475__ & ~new_new_n479__;
  assign new_new_n590__ = new_new_n478__ & ~new_new_n589__;
  assign new_new_n591__ = new_new_n588__ & ~new_new_n590__;
  assign new_new_n592__ = ~new_new_n588__ & new_new_n590__;
  assign new_new_n593__ = ~new_new_n591__ & ~new_new_n592__;
  assign new_new_n594__ = new_new_n574__ & new_new_n593__;
  assign new_new_n595__ = ~new_new_n574__ & ~new_new_n593__;
  assign new_new_n596__ = ~new_new_n594__ & ~new_new_n595__;
  assign new_new_n597__ = ~new_new_n553__ & ~new_new_n596__;
  assign new_new_n598__ = new_new_n553__ & new_new_n596__;
  assign new_new_n599__ = ~new_new_n597__ & ~new_new_n598__;
  assign new_new_n600__ = ~new_new_n497__ & ~new_new_n512__;
  assign new_new_n601__ = new_new_n497__ & new_new_n512__;
  assign new_new_n602__ = ~pi06 & new_new_n498__;
  assign new_new_n603__ = ~new_new_n554__ & ~new_new_n602__;
  assign new_new_n604__ = ~new_new_n486__ & ~new_new_n603__;
  assign new_new_n605__ = new_new_n486__ & new_new_n603__;
  assign new_new_n606__ = ~new_new_n604__ & ~new_new_n605__;
  assign new_new_n607__ = ~new_new_n601__ & ~new_new_n606__;
  assign new_new_n608__ = ~new_new_n600__ & ~new_new_n607__;
  assign new_new_n609__ = new_new_n599__ & ~new_new_n608__;
  assign new_new_n610__ = ~new_new_n599__ & new_new_n608__;
  assign po013 = ~new_new_n609__ & ~new_new_n610__;
  assign new_new_n612__ = pi05 & pi11;
  assign new_new_n613__ = pi01 & ~pi12;
  assign new_new_n614__ = ~new_new_n577__ & ~new_new_n581__;
  assign new_new_n615__ = ~new_new_n580__ & ~new_new_n614__;
  assign new_new_n616__ = ~new_new_n613__ & ~new_new_n615__;
  assign new_new_n617__ = new_new_n612__ & ~new_new_n616__;
  assign new_new_n618__ = pi07 & pi12;
  assign new_new_n619__ = new_new_n615__ & ~new_new_n618__;
  assign new_new_n620__ = new_new_n617__ & ~new_new_n619__;
  assign new_new_n621__ = pi01 & pi12;
  assign new_new_n622__ = new_new_n615__ & ~new_new_n621__;
  assign new_new_n623__ = ~new_new_n615__ & new_new_n621__;
  assign new_new_n624__ = ~new_new_n622__ & ~new_new_n623__;
  assign new_new_n625__ = pi07 & new_new_n624__;
  assign new_new_n626__ = ~pi07 & ~new_new_n624__;
  assign new_new_n627__ = ~new_new_n563__ & ~new_new_n625__;
  assign new_new_n628__ = ~new_new_n626__ & new_new_n627__;
  assign new_new_n629__ = ~new_new_n620__ & ~new_new_n628__;
  assign new_new_n630__ = ~new_new_n586__ & ~new_new_n590__;
  assign new_new_n631__ = ~new_new_n587__ & ~new_new_n630__;
  assign new_new_n632__ = new_new_n573__ & new_new_n631__;
  assign new_new_n633__ = new_new_n587__ & ~new_new_n590__;
  assign new_new_n634__ = new_new_n586__ & new_new_n590__;
  assign new_new_n635__ = ~new_new_n633__ & ~new_new_n634__;
  assign new_new_n636__ = new_new_n574__ & new_new_n635__;
  assign new_new_n637__ = new_new_n572__ & ~new_new_n631__;
  assign new_new_n638__ = ~new_new_n632__ & ~new_new_n637__;
  assign new_new_n639__ = ~new_new_n636__ & new_new_n638__;
  assign new_new_n640__ = new_new_n629__ & ~new_new_n639__;
  assign new_new_n641__ = new_new_n572__ & new_new_n590__;
  assign new_new_n642__ = new_new_n576__ & new_new_n641__;
  assign new_new_n643__ = ~new_new_n576__ & ~new_new_n641__;
  assign new_new_n644__ = ~new_new_n573__ & new_new_n590__;
  assign new_new_n645__ = ~new_new_n572__ & ~new_new_n644__;
  assign new_new_n646__ = ~new_new_n585__ & ~new_new_n643__;
  assign new_new_n647__ = ~new_new_n645__ & new_new_n646__;
  assign new_new_n648__ = new_new_n573__ & ~new_new_n590__;
  assign new_new_n649__ = new_new_n576__ & ~new_new_n648__;
  assign new_new_n650__ = new_new_n585__ & new_new_n645__;
  assign new_new_n651__ = ~new_new_n649__ & new_new_n650__;
  assign new_new_n652__ = ~new_new_n576__ & new_new_n648__;
  assign new_new_n653__ = ~new_new_n642__ & ~new_new_n652__;
  assign new_new_n654__ = ~new_new_n647__ & new_new_n653__;
  assign new_new_n655__ = ~new_new_n651__ & new_new_n654__;
  assign new_new_n656__ = ~new_new_n629__ & ~new_new_n655__;
  assign new_new_n657__ = ~new_new_n640__ & ~new_new_n656__;
  assign new_new_n658__ = ~new_new_n565__ & ~new_new_n568__;
  assign new_new_n659__ = ~new_new_n566__ & ~new_new_n658__;
  assign new_new_n660__ = pi06 & pi07;
  assign new_new_n661__ = pi02 & pi11;
  assign new_new_n662__ = ~new_new_n379__ & ~new_new_n661__;
  assign new_new_n663__ = new_new_n379__ & new_new_n661__;
  assign new_new_n664__ = ~new_new_n662__ & ~new_new_n663__;
  assign new_new_n665__ = new_new_n660__ & ~new_new_n664__;
  assign new_new_n666__ = ~new_new_n660__ & new_new_n664__;
  assign new_new_n667__ = ~new_new_n665__ & ~new_new_n666__;
  assign new_new_n668__ = ~new_new_n659__ & new_new_n667__;
  assign new_new_n669__ = new_new_n659__ & ~new_new_n667__;
  assign new_new_n670__ = ~new_new_n668__ & ~new_new_n669__;
  assign new_new_n671__ = pi04 & pi09;
  assign new_new_n672__ = pi03 & pi10;
  assign new_new_n673__ = pi00 & pi13;
  assign new_new_n674__ = ~new_new_n672__ & ~new_new_n673__;
  assign new_new_n675__ = new_new_n672__ & new_new_n673__;
  assign new_new_n676__ = ~new_new_n674__ & ~new_new_n675__;
  assign new_new_n677__ = new_new_n671__ & ~new_new_n676__;
  assign new_new_n678__ = ~new_new_n671__ & new_new_n676__;
  assign new_new_n679__ = ~new_new_n677__ & ~new_new_n678__;
  assign new_new_n680__ = new_new_n670__ & new_new_n679__;
  assign new_new_n681__ = ~new_new_n670__ & ~new_new_n679__;
  assign new_new_n682__ = ~new_new_n680__ & ~new_new_n681__;
  assign new_new_n683__ = new_new_n657__ & ~new_new_n682__;
  assign new_new_n684__ = ~new_new_n657__ & new_new_n682__;
  assign new_new_n685__ = ~new_new_n683__ & ~new_new_n684__;
  assign new_new_n686__ = ~new_new_n598__ & ~new_new_n608__;
  assign new_new_n687__ = ~new_new_n597__ & ~new_new_n686__;
  assign new_new_n688__ = new_new_n685__ & new_new_n687__;
  assign new_new_n689__ = ~new_new_n685__ & ~new_new_n687__;
  assign po014 = new_new_n688__ | new_new_n689__;
  assign new_new_n691__ = pi07 & new_new_n621__;
  assign new_new_n692__ = pi04 & pi10;
  assign new_new_n693__ = ~new_new_n442__ & ~new_new_n692__;
  assign new_new_n694__ = new_new_n442__ & new_new_n692__;
  assign new_new_n695__ = ~new_new_n693__ & ~new_new_n694__;
  assign new_new_n696__ = new_new_n691__ & ~new_new_n695__;
  assign new_new_n697__ = ~new_new_n691__ & new_new_n695__;
  assign new_new_n698__ = ~new_new_n696__ & ~new_new_n697__;
  assign new_new_n699__ = ~new_new_n617__ & ~new_new_n622__;
  assign new_new_n700__ = pi07 & ~new_new_n699__;
  assign new_new_n701__ = ~pi07 & new_new_n621__;
  assign new_new_n702__ = new_new_n615__ & new_new_n701__;
  assign new_new_n703__ = ~new_new_n700__ & ~new_new_n702__;
  assign new_new_n704__ = new_new_n698__ & new_new_n703__;
  assign new_new_n705__ = ~new_new_n698__ & ~new_new_n703__;
  assign new_new_n706__ = ~new_new_n704__ & ~new_new_n705__;
  assign new_new_n707__ = pi03 & pi11;
  assign new_new_n708__ = pi02 & pi12;
  assign new_new_n709__ = pi00 & pi14;
  assign new_new_n710__ = ~new_new_n708__ & ~new_new_n709__;
  assign new_new_n711__ = new_new_n708__ & new_new_n709__;
  assign new_new_n712__ = ~new_new_n710__ & ~new_new_n711__;
  assign new_new_n713__ = new_new_n707__ & ~new_new_n712__;
  assign new_new_n714__ = ~new_new_n707__ & new_new_n712__;
  assign new_new_n715__ = ~new_new_n713__ & ~new_new_n714__;
  assign new_new_n716__ = new_new_n706__ & ~new_new_n715__;
  assign new_new_n717__ = ~new_new_n706__ & new_new_n715__;
  assign new_new_n718__ = ~new_new_n716__ & ~new_new_n717__;
  assign new_new_n719__ = ~new_new_n668__ & ~new_new_n679__;
  assign new_new_n720__ = ~new_new_n669__ & ~new_new_n719__;
  assign new_new_n721__ = new_new_n718__ & ~new_new_n720__;
  assign new_new_n722__ = ~new_new_n718__ & new_new_n720__;
  assign new_new_n723__ = ~new_new_n721__ & ~new_new_n722__;
  assign new_new_n724__ = ~new_new_n684__ & ~new_new_n687__;
  assign new_new_n725__ = ~new_new_n683__ & ~new_new_n724__;
  assign new_new_n726__ = ~new_new_n572__ & ~new_new_n629__;
  assign new_new_n727__ = new_new_n631__ & ~new_new_n726__;
  assign new_new_n728__ = new_new_n629__ & ~new_new_n633__;
  assign new_new_n729__ = ~new_new_n634__ & ~new_new_n728__;
  assign new_new_n730__ = ~new_new_n573__ & ~new_new_n729__;
  assign new_new_n731__ = new_new_n572__ & new_new_n629__;
  assign new_new_n732__ = ~new_new_n727__ & ~new_new_n731__;
  assign new_new_n733__ = ~new_new_n730__ & new_new_n732__;
  assign new_new_n734__ = new_new_n725__ & new_new_n733__;
  assign new_new_n735__ = ~new_new_n725__ & ~new_new_n733__;
  assign new_new_n736__ = ~new_new_n734__ & ~new_new_n735__;
  assign new_new_n737__ = pi01 & pi13;
  assign new_new_n738__ = pi06 & pi08;
  assign new_new_n739__ = new_new_n737__ & ~new_new_n738__;
  assign new_new_n740__ = ~new_new_n737__ & new_new_n738__;
  assign new_new_n741__ = ~new_new_n739__ & ~new_new_n740__;
  assign new_new_n742__ = ~new_new_n671__ & ~new_new_n675__;
  assign new_new_n743__ = ~new_new_n674__ & ~new_new_n742__;
  assign new_new_n744__ = ~new_new_n660__ & ~new_new_n663__;
  assign new_new_n745__ = ~new_new_n662__ & ~new_new_n744__;
  assign new_new_n746__ = new_new_n743__ & new_new_n745__;
  assign new_new_n747__ = ~new_new_n743__ & ~new_new_n745__;
  assign new_new_n748__ = ~new_new_n746__ & ~new_new_n747__;
  assign new_new_n749__ = new_new_n741__ & new_new_n748__;
  assign new_new_n750__ = ~new_new_n741__ & ~new_new_n748__;
  assign new_new_n751__ = ~new_new_n749__ & ~new_new_n750__;
  assign new_new_n752__ = new_new_n736__ & ~new_new_n751__;
  assign new_new_n753__ = ~new_new_n736__ & new_new_n751__;
  assign new_new_n754__ = ~new_new_n752__ & ~new_new_n753__;
  assign new_new_n755__ = new_new_n723__ & new_new_n754__;
  assign new_new_n756__ = ~new_new_n723__ & ~new_new_n754__;
  assign po015 = ~new_new_n755__ & ~new_new_n756__;
  assign new_new_n758__ = ~new_new_n704__ & ~new_new_n715__;
  assign new_new_n759__ = ~new_new_n705__ & ~new_new_n758__;
  assign new_new_n760__ = ~new_new_n691__ & ~new_new_n694__;
  assign new_new_n761__ = ~new_new_n693__ & ~new_new_n760__;
  assign new_new_n762__ = pi05 & pi10;
  assign new_new_n763__ = pi03 & pi12;
  assign new_new_n764__ = pi00 & pi15;
  assign new_new_n765__ = ~new_new_n763__ & ~new_new_n764__;
  assign new_new_n766__ = new_new_n763__ & new_new_n764__;
  assign new_new_n767__ = ~new_new_n765__ & ~new_new_n766__;
  assign new_new_n768__ = new_new_n762__ & ~new_new_n767__;
  assign new_new_n769__ = ~new_new_n762__ & new_new_n767__;
  assign new_new_n770__ = ~new_new_n768__ & ~new_new_n769__;
  assign new_new_n771__ = ~new_new_n761__ & new_new_n770__;
  assign new_new_n772__ = new_new_n761__ & ~new_new_n770__;
  assign new_new_n773__ = ~new_new_n771__ & ~new_new_n772__;
  assign new_new_n774__ = ~new_new_n707__ & ~new_new_n711__;
  assign new_new_n775__ = ~new_new_n710__ & ~new_new_n774__;
  assign new_new_n776__ = new_new_n773__ & ~new_new_n775__;
  assign new_new_n777__ = ~new_new_n773__ & new_new_n775__;
  assign new_new_n778__ = ~new_new_n776__ & ~new_new_n777__;
  assign new_new_n779__ = ~new_new_n759__ & ~new_new_n778__;
  assign new_new_n780__ = new_new_n759__ & new_new_n778__;
  assign new_new_n781__ = ~new_new_n779__ & ~new_new_n780__;
  assign new_new_n782__ = new_new_n741__ & ~new_new_n746__;
  assign new_new_n783__ = ~new_new_n747__ & ~new_new_n782__;
  assign new_new_n784__ = pi06 & pi13;
  assign new_new_n785__ = pi01 & new_new_n784__;
  assign new_new_n786__ = pi08 & ~new_new_n785__;
  assign new_new_n787__ = pi04 & pi11;
  assign new_new_n788__ = pi01 & pi14;
  assign new_new_n789__ = new_new_n787__ & ~new_new_n788__;
  assign new_new_n790__ = ~new_new_n787__ & new_new_n788__;
  assign new_new_n791__ = ~new_new_n789__ & ~new_new_n790__;
  assign new_new_n792__ = new_new_n786__ & new_new_n791__;
  assign new_new_n793__ = ~new_new_n786__ & ~new_new_n791__;
  assign new_new_n794__ = ~new_new_n792__ & ~new_new_n793__;
  assign new_new_n795__ = ~new_new_n783__ & new_new_n794__;
  assign new_new_n796__ = new_new_n783__ & ~new_new_n794__;
  assign new_new_n797__ = ~new_new_n795__ & ~new_new_n796__;
  assign new_new_n798__ = pi07 & pi08;
  assign new_new_n799__ = pi06 & pi09;
  assign new_new_n800__ = pi02 & pi13;
  assign new_new_n801__ = ~new_new_n799__ & ~new_new_n800__;
  assign new_new_n802__ = new_new_n799__ & new_new_n800__;
  assign new_new_n803__ = ~new_new_n801__ & ~new_new_n802__;
  assign new_new_n804__ = new_new_n798__ & ~new_new_n803__;
  assign new_new_n805__ = ~new_new_n798__ & new_new_n803__;
  assign new_new_n806__ = ~new_new_n804__ & ~new_new_n805__;
  assign new_new_n807__ = new_new_n797__ & new_new_n806__;
  assign new_new_n808__ = ~new_new_n797__ & ~new_new_n806__;
  assign new_new_n809__ = ~new_new_n807__ & ~new_new_n808__;
  assign new_new_n810__ = new_new_n781__ & ~new_new_n809__;
  assign new_new_n811__ = ~new_new_n781__ & new_new_n809__;
  assign new_new_n812__ = ~new_new_n810__ & ~new_new_n811__;
  assign new_new_n813__ = new_new_n722__ & new_new_n751__;
  assign new_new_n814__ = new_new_n721__ & ~new_new_n751__;
  assign new_new_n815__ = ~new_new_n813__ & ~new_new_n814__;
  assign new_new_n816__ = new_new_n736__ & new_new_n815__;
  assign new_new_n817__ = ~new_new_n722__ & ~new_new_n751__;
  assign new_new_n818__ = ~new_new_n721__ & ~new_new_n817__;
  assign new_new_n819__ = new_new_n734__ & ~new_new_n818__;
  assign new_new_n820__ = new_new_n735__ & new_new_n818__;
  assign new_new_n821__ = ~new_new_n812__ & ~new_new_n819__;
  assign new_new_n822__ = ~new_new_n820__ & new_new_n821__;
  assign new_new_n823__ = ~new_new_n816__ & new_new_n822__;
  assign new_new_n824__ = ~new_new_n720__ & ~new_new_n733__;
  assign new_new_n825__ = ~new_new_n725__ & new_new_n824__;
  assign new_new_n826__ = new_new_n718__ & new_new_n825__;
  assign new_new_n827__ = ~new_new_n720__ & ~new_new_n734__;
  assign new_new_n828__ = ~new_new_n735__ & ~new_new_n827__;
  assign new_new_n829__ = new_new_n718__ & ~new_new_n828__;
  assign new_new_n830__ = ~new_new_n825__ & ~new_new_n829__;
  assign new_new_n831__ = ~new_new_n751__ & ~new_new_n830__;
  assign new_new_n832__ = ~new_new_n718__ & new_new_n828__;
  assign new_new_n833__ = new_new_n720__ & new_new_n733__;
  assign new_new_n834__ = new_new_n725__ & new_new_n833__;
  assign new_new_n835__ = ~new_new_n832__ & ~new_new_n834__;
  assign new_new_n836__ = new_new_n751__ & ~new_new_n835__;
  assign new_new_n837__ = ~new_new_n718__ & new_new_n725__;
  assign new_new_n838__ = new_new_n833__ & new_new_n837__;
  assign new_new_n839__ = new_new_n812__ & ~new_new_n826__;
  assign new_new_n840__ = ~new_new_n838__ & new_new_n839__;
  assign new_new_n841__ = ~new_new_n831__ & new_new_n840__;
  assign new_new_n842__ = ~new_new_n836__ & new_new_n841__;
  assign po016 = ~new_new_n823__ & ~new_new_n842__;
  assign new_new_n844__ = ~new_new_n795__ & ~new_new_n806__;
  assign new_new_n845__ = ~new_new_n796__ & ~new_new_n844__;
  assign new_new_n846__ = ~new_new_n779__ & new_new_n809__;
  assign new_new_n847__ = ~new_new_n780__ & ~new_new_n846__;
  assign new_new_n848__ = ~new_new_n762__ & ~new_new_n766__;
  assign new_new_n849__ = ~new_new_n765__ & ~new_new_n848__;
  assign new_new_n850__ = pi14 & ~new_new_n787__;
  assign new_new_n851__ = new_new_n785__ & ~new_new_n850__;
  assign new_new_n852__ = ~new_new_n789__ & ~new_new_n851__;
  assign new_new_n853__ = pi08 & ~new_new_n852__;
  assign new_new_n854__ = ~pi08 & new_new_n787__;
  assign new_new_n855__ = new_new_n788__ & new_new_n854__;
  assign new_new_n856__ = ~new_new_n853__ & ~new_new_n855__;
  assign new_new_n857__ = ~new_new_n849__ & new_new_n856__;
  assign new_new_n858__ = new_new_n849__ & ~new_new_n856__;
  assign new_new_n859__ = ~new_new_n857__ & ~new_new_n858__;
  assign new_new_n860__ = pi06 & pi10;
  assign new_new_n861__ = pi00 & pi16;
  assign new_new_n862__ = ~new_new_n612__ & ~new_new_n861__;
  assign new_new_n863__ = new_new_n612__ & new_new_n861__;
  assign new_new_n864__ = ~new_new_n862__ & ~new_new_n863__;
  assign new_new_n865__ = new_new_n860__ & ~new_new_n864__;
  assign new_new_n866__ = ~new_new_n860__ & new_new_n864__;
  assign new_new_n867__ = ~new_new_n865__ & ~new_new_n866__;
  assign new_new_n868__ = new_new_n859__ & new_new_n867__;
  assign new_new_n869__ = ~new_new_n859__ & ~new_new_n867__;
  assign new_new_n870__ = ~new_new_n868__ & ~new_new_n869__;
  assign new_new_n871__ = ~new_new_n847__ & new_new_n870__;
  assign new_new_n872__ = new_new_n847__ & ~new_new_n870__;
  assign new_new_n873__ = ~new_new_n871__ & ~new_new_n872__;
  assign new_new_n874__ = pi04 & pi12;
  assign new_new_n875__ = pi03 & pi13;
  assign new_new_n876__ = pi02 & pi14;
  assign new_new_n877__ = ~new_new_n875__ & ~new_new_n876__;
  assign new_new_n878__ = new_new_n875__ & new_new_n876__;
  assign new_new_n879__ = ~new_new_n877__ & ~new_new_n878__;
  assign new_new_n880__ = new_new_n874__ & ~new_new_n879__;
  assign new_new_n881__ = ~new_new_n874__ & new_new_n879__;
  assign new_new_n882__ = ~new_new_n880__ & ~new_new_n881__;
  assign new_new_n883__ = ~new_new_n798__ & ~new_new_n802__;
  assign new_new_n884__ = ~new_new_n801__ & ~new_new_n883__;
  assign new_new_n885__ = pi07 & pi09;
  assign new_new_n886__ = pi08 & pi14;
  assign new_new_n887__ = ~pi15 & ~new_new_n886__;
  assign new_new_n888__ = pi08 & pi15;
  assign new_new_n889__ = pi14 & new_new_n888__;
  assign new_new_n890__ = pi01 & ~new_new_n887__;
  assign new_new_n891__ = ~new_new_n889__ & new_new_n890__;
  assign new_new_n892__ = new_new_n885__ & ~new_new_n891__;
  assign new_new_n893__ = ~new_new_n885__ & new_new_n891__;
  assign new_new_n894__ = ~new_new_n892__ & ~new_new_n893__;
  assign new_new_n895__ = new_new_n884__ & new_new_n894__;
  assign new_new_n896__ = ~new_new_n884__ & ~new_new_n894__;
  assign new_new_n897__ = ~new_new_n895__ & ~new_new_n896__;
  assign new_new_n898__ = ~new_new_n882__ & ~new_new_n897__;
  assign new_new_n899__ = new_new_n882__ & new_new_n897__;
  assign new_new_n900__ = ~new_new_n898__ & ~new_new_n899__;
  assign new_new_n901__ = ~new_new_n772__ & ~new_new_n775__;
  assign new_new_n902__ = ~new_new_n771__ & ~new_new_n901__;
  assign new_new_n903__ = new_new_n900__ & new_new_n902__;
  assign new_new_n904__ = ~new_new_n900__ & ~new_new_n902__;
  assign new_new_n905__ = ~new_new_n903__ & ~new_new_n904__;
  assign new_new_n906__ = new_new_n751__ & ~new_new_n824__;
  assign new_new_n907__ = ~new_new_n833__ & ~new_new_n906__;
  assign new_new_n908__ = new_new_n812__ & new_new_n907__;
  assign new_new_n909__ = new_new_n837__ & ~new_new_n908__;
  assign new_new_n910__ = new_new_n718__ & ~new_new_n725__;
  assign new_new_n911__ = ~new_new_n751__ & new_new_n824__;
  assign new_new_n912__ = ~new_new_n812__ & ~new_new_n911__;
  assign new_new_n913__ = new_new_n751__ & new_new_n833__;
  assign new_new_n914__ = ~new_new_n912__ & ~new_new_n913__;
  assign new_new_n915__ = ~new_new_n910__ & ~new_new_n914__;
  assign new_new_n916__ = ~new_new_n812__ & ~new_new_n907__;
  assign new_new_n917__ = ~new_new_n909__ & ~new_new_n916__;
  assign new_new_n918__ = ~new_new_n915__ & new_new_n917__;
  assign new_new_n919__ = new_new_n905__ & new_new_n918__;
  assign new_new_n920__ = ~new_new_n905__ & ~new_new_n918__;
  assign new_new_n921__ = ~new_new_n919__ & ~new_new_n920__;
  assign new_new_n922__ = new_new_n873__ & ~new_new_n921__;
  assign new_new_n923__ = ~new_new_n873__ & new_new_n921__;
  assign new_new_n924__ = ~new_new_n922__ & ~new_new_n923__;
  assign new_new_n925__ = new_new_n845__ & new_new_n924__;
  assign new_new_n926__ = ~new_new_n845__ & ~new_new_n924__;
  assign po017 = ~new_new_n925__ & ~new_new_n926__;
  assign new_new_n928__ = ~new_new_n845__ & ~new_new_n871__;
  assign new_new_n929__ = ~new_new_n872__ & ~new_new_n928__;
  assign new_new_n930__ = ~new_new_n920__ & ~new_new_n929__;
  assign new_new_n931__ = ~new_new_n919__ & new_new_n929__;
  assign new_new_n932__ = ~new_new_n930__ & ~new_new_n931__;
  assign new_new_n933__ = ~new_new_n898__ & ~new_new_n902__;
  assign new_new_n934__ = ~new_new_n899__ & ~new_new_n933__;
  assign new_new_n935__ = ~new_new_n874__ & ~new_new_n878__;
  assign new_new_n936__ = ~new_new_n877__ & ~new_new_n935__;
  assign new_new_n937__ = ~new_new_n860__ & ~new_new_n863__;
  assign new_new_n938__ = ~new_new_n862__ & ~new_new_n937__;
  assign new_new_n939__ = new_new_n936__ & new_new_n938__;
  assign new_new_n940__ = pi01 & pi16;
  assign new_new_n941__ = pi09 & new_new_n940__;
  assign new_new_n942__ = ~new_new_n936__ & ~new_new_n938__;
  assign new_new_n943__ = ~pi09 & ~new_new_n940__;
  assign new_new_n944__ = ~new_new_n941__ & ~new_new_n943__;
  assign new_new_n945__ = ~new_new_n942__ & new_new_n944__;
  assign new_new_n946__ = ~new_new_n939__ & new_new_n945__;
  assign new_new_n947__ = pi09 & pi16;
  assign new_new_n948__ = pi01 & new_new_n947__;
  assign new_new_n949__ = ~new_new_n943__ & ~new_new_n948__;
  assign new_new_n950__ = ~new_new_n939__ & ~new_new_n942__;
  assign new_new_n951__ = ~new_new_n949__ & ~new_new_n950__;
  assign new_new_n952__ = ~new_new_n946__ & ~new_new_n951__;
  assign new_new_n953__ = ~new_new_n884__ & ~new_new_n886__;
  assign new_new_n954__ = pi15 & ~new_new_n885__;
  assign new_new_n955__ = ~new_new_n953__ & new_new_n954__;
  assign new_new_n956__ = ~pi15 & new_new_n885__;
  assign new_new_n957__ = ~new_new_n884__ & ~new_new_n956__;
  assign new_new_n958__ = new_new_n886__ & ~new_new_n957__;
  assign new_new_n959__ = ~new_new_n955__ & ~new_new_n958__;
  assign new_new_n960__ = pi01 & ~new_new_n959__;
  assign new_new_n961__ = pi01 & pi15;
  assign new_new_n962__ = new_new_n885__ & ~new_new_n961__;
  assign new_new_n963__ = new_new_n884__ & new_new_n962__;
  assign new_new_n964__ = ~new_new_n960__ & ~new_new_n963__;
  assign new_new_n965__ = ~new_new_n952__ & new_new_n964__;
  assign new_new_n966__ = new_new_n952__ & ~new_new_n964__;
  assign new_new_n967__ = ~new_new_n965__ & ~new_new_n966__;
  assign new_new_n968__ = ~new_new_n857__ & ~new_new_n867__;
  assign new_new_n969__ = ~new_new_n858__ & ~new_new_n968__;
  assign new_new_n970__ = new_new_n967__ & new_new_n969__;
  assign new_new_n971__ = ~new_new_n967__ & ~new_new_n969__;
  assign new_new_n972__ = ~new_new_n970__ & ~new_new_n971__;
  assign new_new_n973__ = ~new_new_n934__ & new_new_n972__;
  assign new_new_n974__ = new_new_n934__ & ~new_new_n972__;
  assign new_new_n975__ = ~new_new_n973__ & ~new_new_n974__;
  assign new_new_n976__ = pi05 & pi12;
  assign new_new_n977__ = pi00 & pi17;
  assign new_new_n978__ = ~new_new_n976__ & ~new_new_n977__;
  assign new_new_n979__ = new_new_n976__ & new_new_n977__;
  assign new_new_n980__ = ~new_new_n978__ & ~new_new_n979__;
  assign new_new_n981__ = pi07 & pi15;
  assign new_new_n982__ = new_new_n495__ & new_new_n981__;
  assign new_new_n983__ = ~new_new_n980__ & new_new_n982__;
  assign new_new_n984__ = new_new_n980__ & ~new_new_n982__;
  assign new_new_n985__ = ~new_new_n983__ & ~new_new_n984__;
  assign new_new_n986__ = pi06 & pi11;
  assign new_new_n987__ = pi04 & pi13;
  assign new_new_n988__ = pi02 & pi15;
  assign new_new_n989__ = ~new_new_n987__ & ~new_new_n988__;
  assign new_new_n990__ = new_new_n987__ & new_new_n988__;
  assign new_new_n991__ = ~new_new_n989__ & ~new_new_n990__;
  assign new_new_n992__ = new_new_n986__ & ~new_new_n991__;
  assign new_new_n993__ = ~new_new_n986__ & new_new_n991__;
  assign new_new_n994__ = ~new_new_n992__ & ~new_new_n993__;
  assign new_new_n995__ = new_new_n985__ & new_new_n994__;
  assign new_new_n996__ = ~new_new_n985__ & ~new_new_n994__;
  assign new_new_n997__ = ~new_new_n995__ & ~new_new_n996__;
  assign new_new_n998__ = pi08 & pi09;
  assign new_new_n999__ = pi03 & pi14;
  assign new_new_n1000__ = pi07 & pi10;
  assign new_new_n1001__ = ~new_new_n999__ & ~new_new_n1000__;
  assign new_new_n1002__ = new_new_n999__ & new_new_n1000__;
  assign new_new_n1003__ = ~new_new_n1001__ & ~new_new_n1002__;
  assign new_new_n1004__ = new_new_n998__ & ~new_new_n1003__;
  assign new_new_n1005__ = ~new_new_n998__ & new_new_n1003__;
  assign new_new_n1006__ = ~new_new_n1004__ & ~new_new_n1005__;
  assign new_new_n1007__ = ~new_new_n997__ & new_new_n1006__;
  assign new_new_n1008__ = new_new_n997__ & ~new_new_n1006__;
  assign new_new_n1009__ = ~new_new_n1007__ & ~new_new_n1008__;
  assign new_new_n1010__ = new_new_n975__ & new_new_n1009__;
  assign new_new_n1011__ = ~new_new_n975__ & ~new_new_n1009__;
  assign new_new_n1012__ = ~new_new_n1010__ & ~new_new_n1011__;
  assign new_new_n1013__ = new_new_n845__ & new_new_n871__;
  assign new_new_n1014__ = ~new_new_n845__ & new_new_n872__;
  assign new_new_n1015__ = ~new_new_n1013__ & ~new_new_n1014__;
  assign new_new_n1016__ = new_new_n921__ & new_new_n1015__;
  assign new_new_n1017__ = ~new_new_n932__ & ~new_new_n1012__;
  assign new_new_n1018__ = ~new_new_n1016__ & new_new_n1017__;
  assign new_new_n1019__ = new_new_n871__ & new_new_n920__;
  assign new_new_n1020__ = new_new_n847__ & new_new_n919__;
  assign new_new_n1021__ = ~new_new_n870__ & new_new_n1020__;
  assign new_new_n1022__ = ~new_new_n847__ & ~new_new_n919__;
  assign new_new_n1023__ = new_new_n870__ & new_new_n1022__;
  assign new_new_n1024__ = ~new_new_n872__ & new_new_n920__;
  assign new_new_n1025__ = new_new_n845__ & ~new_new_n1024__;
  assign new_new_n1026__ = ~new_new_n1023__ & new_new_n1025__;
  assign new_new_n1027__ = ~new_new_n870__ & ~new_new_n920__;
  assign new_new_n1028__ = ~new_new_n1022__ & new_new_n1027__;
  assign new_new_n1029__ = ~new_new_n845__ & ~new_new_n1020__;
  assign new_new_n1030__ = ~new_new_n1028__ & new_new_n1029__;
  assign new_new_n1031__ = ~new_new_n1026__ & ~new_new_n1030__;
  assign new_new_n1032__ = new_new_n1012__ & ~new_new_n1019__;
  assign new_new_n1033__ = ~new_new_n1021__ & new_new_n1032__;
  assign new_new_n1034__ = ~new_new_n1031__ & new_new_n1033__;
  assign po018 = ~new_new_n1018__ & ~new_new_n1034__;
  assign new_new_n1036__ = ~new_new_n930__ & ~new_new_n1012__;
  assign new_new_n1037__ = new_new_n920__ & new_new_n929__;
  assign new_new_n1038__ = ~new_new_n1012__ & ~new_new_n1014__;
  assign new_new_n1039__ = ~new_new_n1013__ & ~new_new_n1038__;
  assign new_new_n1040__ = ~new_new_n919__ & ~new_new_n1039__;
  assign new_new_n1041__ = ~new_new_n1037__ & ~new_new_n1040__;
  assign new_new_n1042__ = ~new_new_n1036__ & new_new_n1041__;
  assign new_new_n1043__ = ~new_new_n974__ & ~new_new_n1009__;
  assign new_new_n1044__ = ~new_new_n973__ & ~new_new_n1043__;
  assign new_new_n1045__ = new_new_n1042__ & new_new_n1044__;
  assign new_new_n1046__ = ~new_new_n1042__ & ~new_new_n1044__;
  assign new_new_n1047__ = ~new_new_n1045__ & ~new_new_n1046__;
  assign new_new_n1048__ = ~new_new_n965__ & ~new_new_n969__;
  assign new_new_n1049__ = ~new_new_n966__ & ~new_new_n1048__;
  assign new_new_n1050__ = ~new_new_n986__ & ~new_new_n990__;
  assign new_new_n1051__ = ~new_new_n989__ & ~new_new_n1050__;
  assign new_new_n1052__ = ~new_new_n979__ & ~new_new_n982__;
  assign new_new_n1053__ = ~new_new_n978__ & ~new_new_n1052__;
  assign new_new_n1054__ = ~new_new_n1051__ & ~new_new_n1053__;
  assign new_new_n1055__ = new_new_n1051__ & new_new_n1053__;
  assign new_new_n1056__ = ~new_new_n1054__ & ~new_new_n1055__;
  assign new_new_n1057__ = ~new_new_n998__ & ~new_new_n1002__;
  assign new_new_n1058__ = ~new_new_n1001__ & ~new_new_n1057__;
  assign new_new_n1059__ = ~new_new_n1056__ & new_new_n1058__;
  assign new_new_n1060__ = ~new_new_n1055__ & ~new_new_n1058__;
  assign new_new_n1061__ = ~new_new_n1054__ & new_new_n1060__;
  assign new_new_n1062__ = ~new_new_n1059__ & ~new_new_n1061__;
  assign new_new_n1063__ = ~new_new_n939__ & ~new_new_n945__;
  assign new_new_n1064__ = ~new_new_n996__ & new_new_n1006__;
  assign new_new_n1065__ = ~new_new_n995__ & ~new_new_n1064__;
  assign new_new_n1066__ = ~new_new_n1063__ & new_new_n1065__;
  assign new_new_n1067__ = new_new_n1063__ & ~new_new_n1065__;
  assign new_new_n1068__ = ~new_new_n1066__ & ~new_new_n1067__;
  assign new_new_n1069__ = new_new_n1062__ & new_new_n1068__;
  assign new_new_n1070__ = ~new_new_n1062__ & ~new_new_n1068__;
  assign new_new_n1071__ = ~new_new_n1069__ & ~new_new_n1070__;
  assign new_new_n1072__ = new_new_n1049__ & new_new_n1071__;
  assign new_new_n1073__ = ~new_new_n1049__ & ~new_new_n1071__;
  assign new_new_n1074__ = ~new_new_n1072__ & ~new_new_n1073__;
  assign new_new_n1075__ = pi07 & pi11;
  assign new_new_n1076__ = pi05 & pi13;
  assign new_new_n1077__ = pi00 & pi18;
  assign new_new_n1078__ = ~new_new_n1076__ & ~new_new_n1077__;
  assign new_new_n1079__ = new_new_n1076__ & new_new_n1077__;
  assign new_new_n1080__ = ~new_new_n1078__ & ~new_new_n1079__;
  assign new_new_n1081__ = new_new_n1075__ & ~new_new_n1080__;
  assign new_new_n1082__ = ~new_new_n1075__ & new_new_n1080__;
  assign new_new_n1083__ = ~new_new_n1081__ & ~new_new_n1082__;
  assign new_new_n1084__ = pi06 & pi12;
  assign new_new_n1085__ = pi08 & pi10;
  assign new_new_n1086__ = pi01 & pi17;
  assign new_new_n1087__ = ~new_new_n1085__ & new_new_n1086__;
  assign new_new_n1088__ = new_new_n1085__ & ~new_new_n1086__;
  assign new_new_n1089__ = ~new_new_n1087__ & ~new_new_n1088__;
  assign new_new_n1090__ = ~new_new_n1084__ & new_new_n1089__;
  assign new_new_n1091__ = new_new_n1084__ & ~new_new_n1089__;
  assign new_new_n1092__ = ~new_new_n1090__ & ~new_new_n1091__;
  assign new_new_n1093__ = new_new_n941__ & ~new_new_n1092__;
  assign new_new_n1094__ = ~new_new_n941__ & new_new_n1092__;
  assign new_new_n1095__ = ~new_new_n1093__ & ~new_new_n1094__;
  assign new_new_n1096__ = ~new_new_n1083__ & ~new_new_n1095__;
  assign new_new_n1097__ = new_new_n1083__ & new_new_n1095__;
  assign new_new_n1098__ = ~new_new_n1096__ & ~new_new_n1097__;
  assign new_new_n1099__ = pi04 & pi14;
  assign new_new_n1100__ = pi03 & pi15;
  assign new_new_n1101__ = pi02 & pi16;
  assign new_new_n1102__ = ~new_new_n1100__ & ~new_new_n1101__;
  assign new_new_n1103__ = new_new_n1100__ & new_new_n1101__;
  assign new_new_n1104__ = ~new_new_n1102__ & ~new_new_n1103__;
  assign new_new_n1105__ = new_new_n1099__ & ~new_new_n1104__;
  assign new_new_n1106__ = ~new_new_n1099__ & new_new_n1104__;
  assign new_new_n1107__ = ~new_new_n1105__ & ~new_new_n1106__;
  assign new_new_n1108__ = ~new_new_n1098__ & new_new_n1107__;
  assign new_new_n1109__ = new_new_n1098__ & ~new_new_n1107__;
  assign new_new_n1110__ = ~new_new_n1108__ & ~new_new_n1109__;
  assign new_new_n1111__ = new_new_n1074__ & ~new_new_n1110__;
  assign new_new_n1112__ = ~new_new_n1074__ & new_new_n1110__;
  assign new_new_n1113__ = ~new_new_n1111__ & ~new_new_n1112__;
  assign new_new_n1114__ = new_new_n1047__ & new_new_n1113__;
  assign new_new_n1115__ = ~new_new_n1047__ & ~new_new_n1113__;
  assign po019 = new_new_n1114__ | new_new_n1115__;
  assign new_new_n1117__ = ~new_new_n1062__ & ~new_new_n1067__;
  assign new_new_n1118__ = ~new_new_n1066__ & ~new_new_n1117__;
  assign new_new_n1119__ = ~new_new_n1097__ & ~new_new_n1107__;
  assign new_new_n1120__ = ~new_new_n1096__ & ~new_new_n1119__;
  assign new_new_n1121__ = ~new_new_n1099__ & ~new_new_n1103__;
  assign new_new_n1122__ = ~new_new_n1102__ & ~new_new_n1121__;
  assign new_new_n1123__ = pi10 & pi18;
  assign new_new_n1124__ = ~new_new_n1122__ & ~new_new_n1123__;
  assign new_new_n1125__ = pi08 & pi17;
  assign new_new_n1126__ = pi01 & ~pi18;
  assign new_new_n1127__ = new_new_n1122__ & ~new_new_n1126__;
  assign new_new_n1128__ = ~new_new_n1124__ & new_new_n1125__;
  assign new_new_n1129__ = ~new_new_n1127__ & new_new_n1128__;
  assign new_new_n1130__ = new_new_n1085__ & new_new_n1086__;
  assign new_new_n1131__ = pi01 & pi18;
  assign new_new_n1132__ = ~new_new_n1122__ & new_new_n1131__;
  assign new_new_n1133__ = new_new_n1122__ & ~new_new_n1131__;
  assign new_new_n1134__ = ~new_new_n1132__ & ~new_new_n1133__;
  assign new_new_n1135__ = pi10 & ~new_new_n1134__;
  assign new_new_n1136__ = ~pi10 & new_new_n1134__;
  assign new_new_n1137__ = ~new_new_n1130__ & ~new_new_n1135__;
  assign new_new_n1138__ = ~new_new_n1136__ & new_new_n1137__;
  assign new_new_n1139__ = ~new_new_n1129__ & ~new_new_n1138__;
  assign new_new_n1140__ = ~new_new_n1120__ & ~new_new_n1139__;
  assign new_new_n1141__ = new_new_n1120__ & new_new_n1139__;
  assign new_new_n1142__ = ~new_new_n1140__ & ~new_new_n1141__;
  assign new_new_n1143__ = ~new_new_n1075__ & ~new_new_n1079__;
  assign new_new_n1144__ = ~new_new_n1078__ & ~new_new_n1143__;
  assign new_new_n1145__ = ~new_new_n941__ & ~new_new_n1091__;
  assign new_new_n1146__ = ~new_new_n1090__ & ~new_new_n1145__;
  assign new_new_n1147__ = ~new_new_n1144__ & ~new_new_n1146__;
  assign new_new_n1148__ = new_new_n1144__ & new_new_n1146__;
  assign new_new_n1149__ = ~new_new_n1147__ & ~new_new_n1148__;
  assign new_new_n1150__ = pi09 & pi10;
  assign new_new_n1151__ = pi03 & pi16;
  assign new_new_n1152__ = pi08 & pi11;
  assign new_new_n1153__ = ~new_new_n1151__ & ~new_new_n1152__;
  assign new_new_n1154__ = new_new_n1151__ & new_new_n1152__;
  assign new_new_n1155__ = ~new_new_n1153__ & ~new_new_n1154__;
  assign new_new_n1156__ = new_new_n1150__ & ~new_new_n1155__;
  assign new_new_n1157__ = ~new_new_n1150__ & new_new_n1155__;
  assign new_new_n1158__ = ~new_new_n1156__ & ~new_new_n1157__;
  assign new_new_n1159__ = new_new_n1149__ & ~new_new_n1158__;
  assign new_new_n1160__ = ~new_new_n1149__ & new_new_n1158__;
  assign new_new_n1161__ = ~new_new_n1159__ & ~new_new_n1160__;
  assign new_new_n1162__ = new_new_n1142__ & ~new_new_n1161__;
  assign new_new_n1163__ = ~new_new_n1142__ & new_new_n1161__;
  assign new_new_n1164__ = ~new_new_n1162__ & ~new_new_n1163__;
  assign new_new_n1165__ = new_new_n1118__ & new_new_n1164__;
  assign new_new_n1166__ = ~new_new_n1118__ & ~new_new_n1164__;
  assign new_new_n1167__ = ~new_new_n1165__ & ~new_new_n1166__;
  assign new_new_n1168__ = ~new_new_n1054__ & ~new_new_n1060__;
  assign new_new_n1169__ = pi04 & pi15;
  assign new_new_n1170__ = pi02 & pi17;
  assign new_new_n1171__ = pi00 & pi19;
  assign new_new_n1172__ = ~new_new_n1170__ & ~new_new_n1171__;
  assign new_new_n1173__ = new_new_n1170__ & new_new_n1171__;
  assign new_new_n1174__ = ~new_new_n1172__ & ~new_new_n1173__;
  assign new_new_n1175__ = new_new_n1169__ & ~new_new_n1174__;
  assign new_new_n1176__ = ~new_new_n1169__ & new_new_n1174__;
  assign new_new_n1177__ = ~new_new_n1175__ & ~new_new_n1176__;
  assign new_new_n1178__ = ~new_new_n1168__ & new_new_n1177__;
  assign new_new_n1179__ = new_new_n1168__ & ~new_new_n1177__;
  assign new_new_n1180__ = ~new_new_n1178__ & ~new_new_n1179__;
  assign new_new_n1181__ = pi05 & pi14;
  assign new_new_n1182__ = ~new_new_n784__ & ~new_new_n1181__;
  assign new_new_n1183__ = new_new_n784__ & new_new_n1181__;
  assign new_new_n1184__ = ~new_new_n1182__ & ~new_new_n1183__;
  assign new_new_n1185__ = new_new_n618__ & ~new_new_n1184__;
  assign new_new_n1186__ = ~new_new_n618__ & new_new_n1184__;
  assign new_new_n1187__ = ~new_new_n1185__ & ~new_new_n1186__;
  assign new_new_n1188__ = new_new_n1180__ & new_new_n1187__;
  assign new_new_n1189__ = ~new_new_n1180__ & ~new_new_n1187__;
  assign new_new_n1190__ = ~new_new_n1188__ & ~new_new_n1189__;
  assign new_new_n1191__ = new_new_n1167__ & ~new_new_n1190__;
  assign new_new_n1192__ = ~new_new_n1167__ & new_new_n1190__;
  assign new_new_n1193__ = ~new_new_n1191__ & ~new_new_n1192__;
  assign new_new_n1194__ = ~new_new_n1072__ & new_new_n1110__;
  assign new_new_n1195__ = ~new_new_n1073__ & ~new_new_n1194__;
  assign new_new_n1196__ = new_new_n1045__ & new_new_n1195__;
  assign new_new_n1197__ = new_new_n1072__ & ~new_new_n1110__;
  assign new_new_n1198__ = new_new_n1073__ & new_new_n1110__;
  assign new_new_n1199__ = ~new_new_n1197__ & ~new_new_n1198__;
  assign new_new_n1200__ = new_new_n1047__ & new_new_n1199__;
  assign new_new_n1201__ = new_new_n1046__ & ~new_new_n1195__;
  assign new_new_n1202__ = ~new_new_n1196__ & ~new_new_n1201__;
  assign new_new_n1203__ = ~new_new_n1200__ & new_new_n1202__;
  assign new_new_n1204__ = ~new_new_n1193__ & ~new_new_n1203__;
  assign new_new_n1205__ = new_new_n1045__ & ~new_new_n1071__;
  assign new_new_n1206__ = ~new_new_n1049__ & new_new_n1205__;
  assign new_new_n1207__ = ~new_new_n1045__ & new_new_n1071__;
  assign new_new_n1208__ = ~new_new_n1046__ & ~new_new_n1049__;
  assign new_new_n1209__ = ~new_new_n1207__ & new_new_n1208__;
  assign new_new_n1210__ = ~new_new_n1205__ & ~new_new_n1209__;
  assign new_new_n1211__ = new_new_n1110__ & ~new_new_n1210__;
  assign new_new_n1212__ = new_new_n1046__ & new_new_n1072__;
  assign new_new_n1213__ = new_new_n1046__ & ~new_new_n1073__;
  assign new_new_n1214__ = new_new_n1049__ & new_new_n1207__;
  assign new_new_n1215__ = ~new_new_n1213__ & ~new_new_n1214__;
  assign new_new_n1216__ = ~new_new_n1110__ & ~new_new_n1215__;
  assign new_new_n1217__ = ~new_new_n1206__ & ~new_new_n1212__;
  assign new_new_n1218__ = ~new_new_n1211__ & new_new_n1217__;
  assign new_new_n1219__ = ~new_new_n1216__ & new_new_n1218__;
  assign new_new_n1220__ = new_new_n1193__ & ~new_new_n1219__;
  assign po020 = new_new_n1204__ | new_new_n1220__;
  assign new_new_n1222__ = ~new_new_n1178__ & ~new_new_n1188__;
  assign new_new_n1223__ = pi01 & pi19;
  assign new_new_n1224__ = pi09 & pi11;
  assign new_new_n1225__ = new_new_n1223__ & ~new_new_n1224__;
  assign new_new_n1226__ = ~new_new_n1223__ & new_new_n1224__;
  assign new_new_n1227__ = ~new_new_n1225__ & ~new_new_n1226__;
  assign new_new_n1228__ = ~new_new_n1169__ & ~new_new_n1173__;
  assign new_new_n1229__ = ~new_new_n1172__ & ~new_new_n1228__;
  assign new_new_n1230__ = ~new_new_n1150__ & ~new_new_n1154__;
  assign new_new_n1231__ = ~new_new_n1153__ & ~new_new_n1230__;
  assign new_new_n1232__ = new_new_n1229__ & new_new_n1231__;
  assign new_new_n1233__ = ~new_new_n1229__ & ~new_new_n1231__;
  assign new_new_n1234__ = ~new_new_n1232__ & ~new_new_n1233__;
  assign new_new_n1235__ = new_new_n1227__ & new_new_n1234__;
  assign new_new_n1236__ = ~new_new_n1227__ & ~new_new_n1234__;
  assign new_new_n1237__ = ~new_new_n1235__ & ~new_new_n1236__;
  assign new_new_n1238__ = ~new_new_n1222__ & new_new_n1237__;
  assign new_new_n1239__ = new_new_n1222__ & ~new_new_n1237__;
  assign new_new_n1240__ = ~new_new_n1238__ & ~new_new_n1239__;
  assign new_new_n1241__ = ~new_new_n618__ & ~new_new_n1183__;
  assign new_new_n1242__ = ~new_new_n1182__ & ~new_new_n1241__;
  assign new_new_n1243__ = pi08 & pi12;
  assign new_new_n1244__ = pi06 & pi14;
  assign new_new_n1245__ = pi05 & pi15;
  assign new_new_n1246__ = ~new_new_n1244__ & ~new_new_n1245__;
  assign new_new_n1247__ = new_new_n1244__ & new_new_n1245__;
  assign new_new_n1248__ = ~new_new_n1246__ & ~new_new_n1247__;
  assign new_new_n1249__ = new_new_n1243__ & ~new_new_n1248__;
  assign new_new_n1250__ = ~new_new_n1243__ & new_new_n1248__;
  assign new_new_n1251__ = ~new_new_n1249__ & ~new_new_n1250__;
  assign new_new_n1252__ = pi18 & new_new_n498__;
  assign new_new_n1253__ = pi07 & pi13;
  assign new_new_n1254__ = pi00 & pi20;
  assign new_new_n1255__ = ~new_new_n1253__ & ~new_new_n1254__;
  assign new_new_n1256__ = new_new_n1253__ & new_new_n1254__;
  assign new_new_n1257__ = ~new_new_n1255__ & ~new_new_n1256__;
  assign new_new_n1258__ = new_new_n1252__ & ~new_new_n1257__;
  assign new_new_n1259__ = ~new_new_n1252__ & new_new_n1257__;
  assign new_new_n1260__ = ~new_new_n1258__ & ~new_new_n1259__;
  assign new_new_n1261__ = new_new_n1251__ & new_new_n1260__;
  assign new_new_n1262__ = ~new_new_n1251__ & ~new_new_n1260__;
  assign new_new_n1263__ = ~new_new_n1261__ & ~new_new_n1262__;
  assign new_new_n1264__ = new_new_n1242__ & ~new_new_n1263__;
  assign new_new_n1265__ = ~new_new_n1242__ & new_new_n1263__;
  assign new_new_n1266__ = ~new_new_n1264__ & ~new_new_n1265__;
  assign new_new_n1267__ = new_new_n1240__ & ~new_new_n1266__;
  assign new_new_n1268__ = ~new_new_n1240__ & new_new_n1266__;
  assign new_new_n1269__ = ~new_new_n1267__ & ~new_new_n1268__;
  assign new_new_n1270__ = new_new_n1193__ & ~new_new_n1195__;
  assign new_new_n1271__ = new_new_n1193__ & ~new_new_n1197__;
  assign new_new_n1272__ = ~new_new_n1198__ & ~new_new_n1271__;
  assign new_new_n1273__ = ~new_new_n1046__ & ~new_new_n1272__;
  assign new_new_n1274__ = ~new_new_n1193__ & new_new_n1195__;
  assign new_new_n1275__ = new_new_n1045__ & ~new_new_n1274__;
  assign new_new_n1276__ = ~new_new_n1270__ & ~new_new_n1273__;
  assign new_new_n1277__ = ~new_new_n1275__ & new_new_n1276__;
  assign new_new_n1278__ = ~new_new_n1269__ & new_new_n1277__;
  assign new_new_n1279__ = new_new_n1269__ & ~new_new_n1277__;
  assign new_new_n1280__ = ~new_new_n1278__ & ~new_new_n1279__;
  assign new_new_n1281__ = ~new_new_n1165__ & ~new_new_n1190__;
  assign new_new_n1282__ = ~new_new_n1166__ & ~new_new_n1281__;
  assign new_new_n1283__ = pi04 & pi16;
  assign new_new_n1284__ = pi03 & pi17;
  assign new_new_n1285__ = pi02 & pi18;
  assign new_new_n1286__ = ~new_new_n1284__ & ~new_new_n1285__;
  assign new_new_n1287__ = new_new_n1284__ & new_new_n1285__;
  assign new_new_n1288__ = ~new_new_n1286__ & ~new_new_n1287__;
  assign new_new_n1289__ = new_new_n1283__ & ~new_new_n1288__;
  assign new_new_n1290__ = ~new_new_n1283__ & new_new_n1288__;
  assign new_new_n1291__ = ~new_new_n1289__ & ~new_new_n1290__;
  assign new_new_n1292__ = ~new_new_n1122__ & ~new_new_n1126__;
  assign new_new_n1293__ = new_new_n1125__ & ~new_new_n1292__;
  assign new_new_n1294__ = ~new_new_n1133__ & ~new_new_n1293__;
  assign new_new_n1295__ = pi10 & ~new_new_n1294__;
  assign new_new_n1296__ = ~pi10 & new_new_n1131__;
  assign new_new_n1297__ = new_new_n1122__ & new_new_n1296__;
  assign new_new_n1298__ = ~new_new_n1295__ & ~new_new_n1297__;
  assign new_new_n1299__ = new_new_n1291__ & new_new_n1298__;
  assign new_new_n1300__ = ~new_new_n1291__ & ~new_new_n1298__;
  assign new_new_n1301__ = ~new_new_n1299__ & ~new_new_n1300__;
  assign new_new_n1302__ = ~new_new_n1148__ & new_new_n1158__;
  assign new_new_n1303__ = ~new_new_n1147__ & ~new_new_n1302__;
  assign new_new_n1304__ = new_new_n1301__ & new_new_n1303__;
  assign new_new_n1305__ = ~new_new_n1301__ & ~new_new_n1303__;
  assign new_new_n1306__ = ~new_new_n1304__ & ~new_new_n1305__;
  assign new_new_n1307__ = new_new_n1282__ & ~new_new_n1306__;
  assign new_new_n1308__ = ~new_new_n1282__ & new_new_n1306__;
  assign new_new_n1309__ = ~new_new_n1307__ & ~new_new_n1308__;
  assign new_new_n1310__ = ~new_new_n1141__ & new_new_n1161__;
  assign new_new_n1311__ = ~new_new_n1140__ & ~new_new_n1310__;
  assign new_new_n1312__ = new_new_n1309__ & ~new_new_n1311__;
  assign new_new_n1313__ = ~new_new_n1309__ & new_new_n1311__;
  assign new_new_n1314__ = ~new_new_n1312__ & ~new_new_n1313__;
  assign new_new_n1315__ = new_new_n1280__ & new_new_n1314__;
  assign new_new_n1316__ = ~new_new_n1280__ & ~new_new_n1314__;
  assign po021 = ~new_new_n1315__ & ~new_new_n1316__;
  assign new_new_n1318__ = new_new_n1242__ & ~new_new_n1261__;
  assign new_new_n1319__ = ~new_new_n1262__ & ~new_new_n1318__;
  assign new_new_n1320__ = pi09 & pi19;
  assign new_new_n1321__ = pi00 & pi21;
  assign new_new_n1322__ = pi01 & ~pi20;
  assign new_new_n1323__ = ~new_new_n1321__ & ~new_new_n1322__;
  assign new_new_n1324__ = new_new_n1320__ & ~new_new_n1323__;
  assign new_new_n1325__ = pi11 & pi20;
  assign new_new_n1326__ = new_new_n1321__ & ~new_new_n1325__;
  assign new_new_n1327__ = new_new_n1324__ & ~new_new_n1326__;
  assign new_new_n1328__ = new_new_n1223__ & new_new_n1224__;
  assign new_new_n1329__ = pi01 & pi20;
  assign new_new_n1330__ = new_new_n1321__ & ~new_new_n1329__;
  assign new_new_n1331__ = ~new_new_n1321__ & new_new_n1329__;
  assign new_new_n1332__ = ~new_new_n1330__ & ~new_new_n1331__;
  assign new_new_n1333__ = pi11 & new_new_n1332__;
  assign new_new_n1334__ = ~pi11 & ~new_new_n1332__;
  assign new_new_n1335__ = ~new_new_n1328__ & ~new_new_n1333__;
  assign new_new_n1336__ = ~new_new_n1334__ & new_new_n1335__;
  assign new_new_n1337__ = ~new_new_n1327__ & ~new_new_n1336__;
  assign new_new_n1338__ = new_new_n1227__ & ~new_new_n1232__;
  assign new_new_n1339__ = ~new_new_n1233__ & ~new_new_n1338__;
  assign new_new_n1340__ = ~new_new_n1337__ & ~new_new_n1339__;
  assign new_new_n1341__ = new_new_n1337__ & new_new_n1339__;
  assign new_new_n1342__ = ~new_new_n1340__ & ~new_new_n1341__;
  assign new_new_n1343__ = new_new_n1319__ & new_new_n1342__;
  assign new_new_n1344__ = ~new_new_n1319__ & ~new_new_n1342__;
  assign new_new_n1345__ = ~new_new_n1343__ & ~new_new_n1344__;
  assign new_new_n1346__ = ~new_new_n1239__ & new_new_n1266__;
  assign new_new_n1347__ = ~new_new_n1238__ & ~new_new_n1346__;
  assign new_new_n1348__ = ~new_new_n1299__ & new_new_n1303__;
  assign new_new_n1349__ = ~new_new_n1300__ & ~new_new_n1348__;
  assign new_new_n1350__ = ~new_new_n1283__ & ~new_new_n1287__;
  assign new_new_n1351__ = ~new_new_n1286__ & ~new_new_n1350__;
  assign new_new_n1352__ = ~new_new_n1243__ & ~new_new_n1247__;
  assign new_new_n1353__ = ~new_new_n1246__ & ~new_new_n1352__;
  assign new_new_n1354__ = ~new_new_n1252__ & ~new_new_n1256__;
  assign new_new_n1355__ = ~new_new_n1255__ & ~new_new_n1354__;
  assign new_new_n1356__ = new_new_n1353__ & new_new_n1355__;
  assign new_new_n1357__ = ~new_new_n1353__ & ~new_new_n1355__;
  assign new_new_n1358__ = ~new_new_n1356__ & ~new_new_n1357__;
  assign new_new_n1359__ = new_new_n1351__ & ~new_new_n1358__;
  assign new_new_n1360__ = ~new_new_n1351__ & new_new_n1358__;
  assign new_new_n1361__ = ~new_new_n1359__ & ~new_new_n1360__;
  assign new_new_n1362__ = new_new_n1349__ & new_new_n1361__;
  assign new_new_n1363__ = ~new_new_n1349__ & ~new_new_n1361__;
  assign new_new_n1364__ = ~new_new_n1362__ & ~new_new_n1363__;
  assign new_new_n1365__ = pi05 & pi16;
  assign new_new_n1366__ = pi02 & pi19;
  assign new_new_n1367__ = pi03 & pi18;
  assign new_new_n1368__ = ~new_new_n1366__ & ~new_new_n1367__;
  assign new_new_n1369__ = new_new_n1366__ & new_new_n1367__;
  assign new_new_n1370__ = ~new_new_n1368__ & ~new_new_n1369__;
  assign new_new_n1371__ = new_new_n1365__ & ~new_new_n1370__;
  assign new_new_n1372__ = ~new_new_n1365__ & new_new_n1370__;
  assign new_new_n1373__ = ~new_new_n1371__ & ~new_new_n1372__;
  assign new_new_n1374__ = pi08 & pi13;
  assign new_new_n1375__ = pi07 & pi14;
  assign new_new_n1376__ = pi06 & pi15;
  assign new_new_n1377__ = ~new_new_n1375__ & ~new_new_n1376__;
  assign new_new_n1378__ = new_new_n1375__ & new_new_n1376__;
  assign new_new_n1379__ = ~new_new_n1377__ & ~new_new_n1378__;
  assign new_new_n1380__ = new_new_n1374__ & ~new_new_n1379__;
  assign new_new_n1381__ = ~new_new_n1374__ & new_new_n1379__;
  assign new_new_n1382__ = ~new_new_n1380__ & ~new_new_n1381__;
  assign new_new_n1383__ = new_new_n1373__ & new_new_n1382__;
  assign new_new_n1384__ = ~new_new_n1373__ & ~new_new_n1382__;
  assign new_new_n1385__ = ~new_new_n1383__ & ~new_new_n1384__;
  assign new_new_n1386__ = pi10 & pi11;
  assign new_new_n1387__ = pi09 & pi12;
  assign new_new_n1388__ = pi04 & pi17;
  assign new_new_n1389__ = ~new_new_n1387__ & ~new_new_n1388__;
  assign new_new_n1390__ = new_new_n1387__ & new_new_n1388__;
  assign new_new_n1391__ = ~new_new_n1389__ & ~new_new_n1390__;
  assign new_new_n1392__ = new_new_n1386__ & ~new_new_n1391__;
  assign new_new_n1393__ = ~new_new_n1386__ & new_new_n1391__;
  assign new_new_n1394__ = ~new_new_n1392__ & ~new_new_n1393__;
  assign new_new_n1395__ = ~new_new_n1385__ & new_new_n1394__;
  assign new_new_n1396__ = new_new_n1385__ & ~new_new_n1394__;
  assign new_new_n1397__ = ~new_new_n1395__ & ~new_new_n1396__;
  assign new_new_n1398__ = new_new_n1364__ & new_new_n1397__;
  assign new_new_n1399__ = ~new_new_n1364__ & ~new_new_n1397__;
  assign new_new_n1400__ = ~new_new_n1398__ & ~new_new_n1399__;
  assign new_new_n1401__ = ~new_new_n1347__ & ~new_new_n1400__;
  assign new_new_n1402__ = new_new_n1347__ & new_new_n1400__;
  assign new_new_n1403__ = ~new_new_n1401__ & ~new_new_n1402__;
  assign new_new_n1404__ = new_new_n1345__ & ~new_new_n1403__;
  assign new_new_n1405__ = ~new_new_n1345__ & new_new_n1403__;
  assign new_new_n1406__ = ~new_new_n1404__ & ~new_new_n1405__;
  assign new_new_n1407__ = ~new_new_n1308__ & new_new_n1311__;
  assign new_new_n1408__ = ~new_new_n1307__ & ~new_new_n1407__;
  assign new_new_n1409__ = ~new_new_n1279__ & ~new_new_n1408__;
  assign new_new_n1410__ = ~new_new_n1278__ & new_new_n1408__;
  assign new_new_n1411__ = ~new_new_n1409__ & ~new_new_n1410__;
  assign new_new_n1412__ = new_new_n1308__ & ~new_new_n1311__;
  assign new_new_n1413__ = new_new_n1307__ & new_new_n1311__;
  assign new_new_n1414__ = ~new_new_n1412__ & ~new_new_n1413__;
  assign new_new_n1415__ = new_new_n1280__ & new_new_n1414__;
  assign new_new_n1416__ = ~new_new_n1411__ & ~new_new_n1415__;
  assign new_new_n1417__ = ~new_new_n1406__ & ~new_new_n1416__;
  assign new_new_n1418__ = new_new_n1278__ & new_new_n1307__;
  assign new_new_n1419__ = new_new_n1278__ & new_new_n1282__;
  assign new_new_n1420__ = ~new_new_n1278__ & ~new_new_n1282__;
  assign new_new_n1421__ = ~new_new_n1279__ & ~new_new_n1306__;
  assign new_new_n1422__ = ~new_new_n1420__ & new_new_n1421__;
  assign new_new_n1423__ = ~new_new_n1419__ & ~new_new_n1422__;
  assign new_new_n1424__ = new_new_n1311__ & ~new_new_n1423__;
  assign new_new_n1425__ = new_new_n1279__ & ~new_new_n1307__;
  assign new_new_n1426__ = new_new_n1306__ & new_new_n1420__;
  assign new_new_n1427__ = ~new_new_n1425__ & ~new_new_n1426__;
  assign new_new_n1428__ = ~new_new_n1311__ & ~new_new_n1427__;
  assign new_new_n1429__ = new_new_n1279__ & new_new_n1308__;
  assign new_new_n1430__ = ~new_new_n1418__ & ~new_new_n1429__;
  assign new_new_n1431__ = ~new_new_n1424__ & new_new_n1430__;
  assign new_new_n1432__ = ~new_new_n1428__ & new_new_n1431__;
  assign new_new_n1433__ = new_new_n1406__ & ~new_new_n1432__;
  assign po022 = new_new_n1417__ | new_new_n1433__;
  assign new_new_n1435__ = new_new_n1345__ & ~new_new_n1402__;
  assign new_new_n1436__ = ~new_new_n1401__ & ~new_new_n1435__;
  assign new_new_n1437__ = new_new_n1406__ & ~new_new_n1409__;
  assign new_new_n1438__ = new_new_n1279__ & new_new_n1408__;
  assign new_new_n1439__ = ~new_new_n1406__ & ~new_new_n1412__;
  assign new_new_n1440__ = ~new_new_n1413__ & ~new_new_n1439__;
  assign new_new_n1441__ = ~new_new_n1278__ & new_new_n1440__;
  assign new_new_n1442__ = ~new_new_n1438__ & ~new_new_n1441__;
  assign new_new_n1443__ = ~new_new_n1437__ & new_new_n1442__;
  assign new_new_n1444__ = new_new_n1436__ & ~new_new_n1443__;
  assign new_new_n1445__ = ~new_new_n1436__ & new_new_n1443__;
  assign new_new_n1446__ = ~new_new_n1444__ & ~new_new_n1445__;
  assign new_new_n1447__ = ~new_new_n1363__ & ~new_new_n1397__;
  assign new_new_n1448__ = ~new_new_n1362__ & ~new_new_n1447__;
  assign new_new_n1449__ = pi10 & pi12;
  assign new_new_n1450__ = ~new_new_n1386__ & ~new_new_n1390__;
  assign new_new_n1451__ = ~new_new_n1389__ & ~new_new_n1450__;
  assign new_new_n1452__ = new_new_n1449__ & new_new_n1451__;
  assign new_new_n1453__ = ~new_new_n1449__ & ~new_new_n1451__;
  assign new_new_n1454__ = ~new_new_n1452__ & ~new_new_n1453__;
  assign new_new_n1455__ = ~pi21 & ~new_new_n1325__;
  assign new_new_n1456__ = pi11 & pi21;
  assign new_new_n1457__ = pi20 & new_new_n1456__;
  assign new_new_n1458__ = pi01 & ~new_new_n1455__;
  assign new_new_n1459__ = ~new_new_n1457__ & new_new_n1458__;
  assign new_new_n1460__ = new_new_n1454__ & ~new_new_n1459__;
  assign new_new_n1461__ = ~new_new_n1454__ & new_new_n1459__;
  assign new_new_n1462__ = ~new_new_n1460__ & ~new_new_n1461__;
  assign new_new_n1463__ = ~new_new_n1351__ & ~new_new_n1356__;
  assign new_new_n1464__ = ~new_new_n1357__ & ~new_new_n1463__;
  assign new_new_n1465__ = ~new_new_n1462__ & new_new_n1464__;
  assign new_new_n1466__ = new_new_n1462__ & ~new_new_n1464__;
  assign new_new_n1467__ = ~new_new_n1465__ & ~new_new_n1466__;
  assign new_new_n1468__ = ~new_new_n1384__ & new_new_n1394__;
  assign new_new_n1469__ = ~new_new_n1383__ & ~new_new_n1468__;
  assign new_new_n1470__ = new_new_n1467__ & ~new_new_n1469__;
  assign new_new_n1471__ = ~new_new_n1467__ & new_new_n1469__;
  assign new_new_n1472__ = ~new_new_n1470__ & ~new_new_n1471__;
  assign new_new_n1473__ = ~new_new_n1340__ & ~new_new_n1343__;
  assign new_new_n1474__ = pi00 & pi22;
  assign new_new_n1475__ = ~new_new_n981__ & ~new_new_n1474__;
  assign new_new_n1476__ = new_new_n981__ & new_new_n1474__;
  assign new_new_n1477__ = ~new_new_n1475__ & ~new_new_n1476__;
  assign new_new_n1478__ = new_new_n886__ & ~new_new_n1477__;
  assign new_new_n1479__ = ~new_new_n886__ & new_new_n1477__;
  assign new_new_n1480__ = ~new_new_n1478__ & ~new_new_n1479__;
  assign new_new_n1481__ = pi05 & pi17;
  assign new_new_n1482__ = pi03 & pi19;
  assign new_new_n1483__ = pi04 & pi18;
  assign new_new_n1484__ = ~new_new_n1482__ & ~new_new_n1483__;
  assign new_new_n1485__ = new_new_n1482__ & new_new_n1483__;
  assign new_new_n1486__ = ~new_new_n1484__ & ~new_new_n1485__;
  assign new_new_n1487__ = new_new_n1481__ & ~new_new_n1486__;
  assign new_new_n1488__ = ~new_new_n1481__ & new_new_n1486__;
  assign new_new_n1489__ = ~new_new_n1487__ & ~new_new_n1488__;
  assign new_new_n1490__ = new_new_n1480__ & new_new_n1489__;
  assign new_new_n1491__ = ~new_new_n1480__ & ~new_new_n1489__;
  assign new_new_n1492__ = ~new_new_n1490__ & ~new_new_n1491__;
  assign new_new_n1493__ = pi09 & pi13;
  assign new_new_n1494__ = pi06 & pi16;
  assign new_new_n1495__ = pi02 & pi20;
  assign new_new_n1496__ = ~new_new_n1494__ & ~new_new_n1495__;
  assign new_new_n1497__ = new_new_n1494__ & new_new_n1495__;
  assign new_new_n1498__ = ~new_new_n1496__ & ~new_new_n1497__;
  assign new_new_n1499__ = new_new_n1493__ & ~new_new_n1498__;
  assign new_new_n1500__ = ~new_new_n1493__ & new_new_n1498__;
  assign new_new_n1501__ = ~new_new_n1499__ & ~new_new_n1500__;
  assign new_new_n1502__ = new_new_n1492__ & ~new_new_n1501__;
  assign new_new_n1503__ = ~new_new_n1492__ & new_new_n1501__;
  assign new_new_n1504__ = ~new_new_n1502__ & ~new_new_n1503__;
  assign new_new_n1505__ = new_new_n1473__ & new_new_n1504__;
  assign new_new_n1506__ = ~new_new_n1473__ & ~new_new_n1504__;
  assign new_new_n1507__ = ~new_new_n1505__ & ~new_new_n1506__;
  assign new_new_n1508__ = ~new_new_n1324__ & ~new_new_n1330__;
  assign new_new_n1509__ = pi11 & ~new_new_n1508__;
  assign new_new_n1510__ = ~pi11 & new_new_n1321__;
  assign new_new_n1511__ = new_new_n1329__ & new_new_n1510__;
  assign new_new_n1512__ = ~new_new_n1509__ & ~new_new_n1511__;
  assign new_new_n1513__ = ~new_new_n1365__ & ~new_new_n1369__;
  assign new_new_n1514__ = ~new_new_n1368__ & ~new_new_n1513__;
  assign new_new_n1515__ = new_new_n1512__ & ~new_new_n1514__;
  assign new_new_n1516__ = ~new_new_n1512__ & new_new_n1514__;
  assign new_new_n1517__ = ~new_new_n1515__ & ~new_new_n1516__;
  assign new_new_n1518__ = ~new_new_n1374__ & ~new_new_n1378__;
  assign new_new_n1519__ = ~new_new_n1377__ & ~new_new_n1518__;
  assign new_new_n1520__ = new_new_n1517__ & new_new_n1519__;
  assign new_new_n1521__ = ~new_new_n1517__ & ~new_new_n1519__;
  assign new_new_n1522__ = ~new_new_n1520__ & ~new_new_n1521__;
  assign new_new_n1523__ = new_new_n1507__ & ~new_new_n1522__;
  assign new_new_n1524__ = ~new_new_n1507__ & new_new_n1522__;
  assign new_new_n1525__ = ~new_new_n1523__ & ~new_new_n1524__;
  assign new_new_n1526__ = new_new_n1472__ & new_new_n1525__;
  assign new_new_n1527__ = ~new_new_n1472__ & ~new_new_n1525__;
  assign new_new_n1528__ = ~new_new_n1526__ & ~new_new_n1527__;
  assign new_new_n1529__ = ~new_new_n1448__ & new_new_n1528__;
  assign new_new_n1530__ = new_new_n1448__ & ~new_new_n1528__;
  assign new_new_n1531__ = ~new_new_n1529__ & ~new_new_n1530__;
  assign new_new_n1532__ = new_new_n1446__ & new_new_n1531__;
  assign new_new_n1533__ = ~new_new_n1446__ & ~new_new_n1531__;
  assign po023 = new_new_n1532__ | new_new_n1533__;
  assign new_new_n1535__ = pi01 & pi22;
  assign new_new_n1536__ = ~pi12 & ~new_new_n1535__;
  assign new_new_n1537__ = pi22 & new_new_n621__;
  assign new_new_n1538__ = ~new_new_n1536__ & ~new_new_n1537__;
  assign new_new_n1539__ = ~new_new_n1481__ & ~new_new_n1485__;
  assign new_new_n1540__ = ~new_new_n1484__ & ~new_new_n1539__;
  assign new_new_n1541__ = ~new_new_n1493__ & ~new_new_n1497__;
  assign new_new_n1542__ = ~new_new_n1496__ & ~new_new_n1541__;
  assign new_new_n1543__ = ~new_new_n1540__ & ~new_new_n1542__;
  assign new_new_n1544__ = new_new_n1540__ & new_new_n1542__;
  assign new_new_n1545__ = ~new_new_n1543__ & ~new_new_n1544__;
  assign new_new_n1546__ = ~new_new_n1538__ & new_new_n1545__;
  assign new_new_n1547__ = pi12 & new_new_n1535__;
  assign new_new_n1548__ = ~new_new_n1536__ & ~new_new_n1547__;
  assign new_new_n1549__ = ~new_new_n1545__ & new_new_n1548__;
  assign new_new_n1550__ = ~new_new_n1546__ & ~new_new_n1549__;
  assign new_new_n1551__ = ~new_new_n1491__ & new_new_n1501__;
  assign new_new_n1552__ = ~new_new_n1490__ & ~new_new_n1551__;
  assign new_new_n1553__ = new_new_n1550__ & ~new_new_n1552__;
  assign new_new_n1554__ = ~new_new_n1550__ & new_new_n1552__;
  assign new_new_n1555__ = ~new_new_n1553__ & ~new_new_n1554__;
  assign new_new_n1556__ = ~new_new_n1516__ & ~new_new_n1519__;
  assign new_new_n1557__ = ~new_new_n1515__ & ~new_new_n1556__;
  assign new_new_n1558__ = new_new_n1555__ & ~new_new_n1557__;
  assign new_new_n1559__ = ~new_new_n1555__ & new_new_n1557__;
  assign new_new_n1560__ = ~new_new_n1558__ & ~new_new_n1559__;
  assign new_new_n1561__ = ~new_new_n1506__ & new_new_n1522__;
  assign new_new_n1562__ = ~new_new_n1505__ & ~new_new_n1561__;
  assign new_new_n1563__ = ~new_new_n1465__ & ~new_new_n1469__;
  assign new_new_n1564__ = ~new_new_n1466__ & ~new_new_n1563__;
  assign new_new_n1565__ = pi10 & pi13;
  assign new_new_n1566__ = pi04 & pi19;
  assign new_new_n1567__ = ~new_new_n1325__ & ~new_new_n1451__;
  assign new_new_n1568__ = pi21 & ~new_new_n1449__;
  assign new_new_n1569__ = ~new_new_n1567__ & new_new_n1568__;
  assign new_new_n1570__ = ~pi21 & new_new_n1449__;
  assign new_new_n1571__ = ~new_new_n1451__ & ~new_new_n1570__;
  assign new_new_n1572__ = new_new_n1325__ & ~new_new_n1571__;
  assign new_new_n1573__ = ~new_new_n1569__ & ~new_new_n1572__;
  assign new_new_n1574__ = pi01 & ~new_new_n1573__;
  assign new_new_n1575__ = pi01 & pi21;
  assign new_new_n1576__ = new_new_n1452__ & ~new_new_n1575__;
  assign new_new_n1577__ = ~new_new_n1574__ & ~new_new_n1576__;
  assign new_new_n1578__ = pi11 & pi12;
  assign new_new_n1579__ = pi06 & pi17;
  assign new_new_n1580__ = pi05 & pi18;
  assign new_new_n1581__ = pi03 & pi20;
  assign new_new_n1582__ = ~new_new_n1580__ & ~new_new_n1581__;
  assign new_new_n1583__ = new_new_n1580__ & new_new_n1581__;
  assign new_new_n1584__ = ~new_new_n1582__ & ~new_new_n1583__;
  assign new_new_n1585__ = new_new_n1579__ & ~new_new_n1584__;
  assign new_new_n1586__ = ~new_new_n1579__ & new_new_n1584__;
  assign new_new_n1587__ = ~new_new_n1585__ & ~new_new_n1586__;
  assign new_new_n1588__ = new_new_n1578__ & ~new_new_n1587__;
  assign new_new_n1589__ = ~new_new_n1578__ & new_new_n1587__;
  assign new_new_n1590__ = ~new_new_n1588__ & ~new_new_n1589__;
  assign new_new_n1591__ = new_new_n1577__ & new_new_n1590__;
  assign new_new_n1592__ = ~new_new_n1577__ & ~new_new_n1590__;
  assign new_new_n1593__ = ~new_new_n1591__ & ~new_new_n1592__;
  assign new_new_n1594__ = new_new_n1566__ & ~new_new_n1593__;
  assign new_new_n1595__ = ~new_new_n1566__ & new_new_n1593__;
  assign new_new_n1596__ = ~new_new_n1594__ & ~new_new_n1595__;
  assign new_new_n1597__ = new_new_n1565__ & new_new_n1596__;
  assign new_new_n1598__ = ~new_new_n1565__ & ~new_new_n1596__;
  assign new_new_n1599__ = ~new_new_n1597__ & ~new_new_n1598__;
  assign new_new_n1600__ = new_new_n1564__ & new_new_n1599__;
  assign new_new_n1601__ = ~new_new_n1564__ & ~new_new_n1599__;
  assign new_new_n1602__ = ~new_new_n1600__ & ~new_new_n1601__;
  assign new_new_n1603__ = pi09 & pi14;
  assign new_new_n1604__ = pi07 & pi16;
  assign new_new_n1605__ = ~new_new_n888__ & ~new_new_n1604__;
  assign new_new_n1606__ = new_new_n888__ & new_new_n1604__;
  assign new_new_n1607__ = ~new_new_n1605__ & ~new_new_n1606__;
  assign new_new_n1608__ = new_new_n1603__ & ~new_new_n1607__;
  assign new_new_n1609__ = ~new_new_n1603__ & new_new_n1607__;
  assign new_new_n1610__ = ~new_new_n1608__ & ~new_new_n1609__;
  assign new_new_n1611__ = pi00 & pi23;
  assign new_new_n1612__ = pi12 & new_new_n498__;
  assign new_new_n1613__ = ~pi02 & ~new_new_n1612__;
  assign new_new_n1614__ = pi21 & ~new_new_n1613__;
  assign new_new_n1615__ = new_new_n498__ & new_new_n708__;
  assign new_new_n1616__ = new_new_n1614__ & ~new_new_n1615__;
  assign new_new_n1617__ = new_new_n1611__ & ~new_new_n1616__;
  assign new_new_n1618__ = ~new_new_n1611__ & new_new_n1616__;
  assign new_new_n1619__ = ~new_new_n1617__ & ~new_new_n1618__;
  assign new_new_n1620__ = new_new_n1610__ & new_new_n1619__;
  assign new_new_n1621__ = ~new_new_n1610__ & ~new_new_n1619__;
  assign new_new_n1622__ = ~new_new_n1620__ & ~new_new_n1621__;
  assign new_new_n1623__ = ~new_new_n886__ & ~new_new_n1476__;
  assign new_new_n1624__ = ~new_new_n1475__ & ~new_new_n1623__;
  assign new_new_n1625__ = new_new_n1622__ & new_new_n1624__;
  assign new_new_n1626__ = ~new_new_n1622__ & ~new_new_n1624__;
  assign new_new_n1627__ = ~new_new_n1625__ & ~new_new_n1626__;
  assign new_new_n1628__ = new_new_n1602__ & ~new_new_n1627__;
  assign new_new_n1629__ = ~new_new_n1602__ & new_new_n1627__;
  assign new_new_n1630__ = ~new_new_n1628__ & ~new_new_n1629__;
  assign new_new_n1631__ = new_new_n1562__ & new_new_n1630__;
  assign new_new_n1632__ = ~new_new_n1562__ & ~new_new_n1630__;
  assign new_new_n1633__ = ~new_new_n1631__ & ~new_new_n1632__;
  assign new_new_n1634__ = ~new_new_n1448__ & ~new_new_n1527__;
  assign new_new_n1635__ = ~new_new_n1526__ & ~new_new_n1634__;
  assign new_new_n1636__ = ~new_new_n1445__ & ~new_new_n1531__;
  assign new_new_n1637__ = ~new_new_n1444__ & ~new_new_n1636__;
  assign new_new_n1638__ = new_new_n1635__ & ~new_new_n1637__;
  assign new_new_n1639__ = ~new_new_n1635__ & new_new_n1637__;
  assign new_new_n1640__ = ~new_new_n1638__ & ~new_new_n1639__;
  assign new_new_n1641__ = new_new_n1633__ & ~new_new_n1640__;
  assign new_new_n1642__ = ~new_new_n1633__ & new_new_n1640__;
  assign new_new_n1643__ = ~new_new_n1641__ & ~new_new_n1642__;
  assign new_new_n1644__ = new_new_n1560__ & new_new_n1643__;
  assign new_new_n1645__ = ~new_new_n1560__ & ~new_new_n1643__;
  assign po024 = ~new_new_n1644__ & ~new_new_n1645__;
  assign new_new_n1647__ = ~new_new_n1601__ & new_new_n1627__;
  assign new_new_n1648__ = ~new_new_n1600__ & ~new_new_n1647__;
  assign new_new_n1649__ = ~new_new_n1603__ & ~new_new_n1606__;
  assign new_new_n1650__ = ~new_new_n1605__ & ~new_new_n1649__;
  assign new_new_n1651__ = ~new_new_n1579__ & ~new_new_n1583__;
  assign new_new_n1652__ = ~new_new_n1582__ & ~new_new_n1651__;
  assign new_new_n1653__ = ~new_new_n1650__ & ~new_new_n1652__;
  assign new_new_n1654__ = new_new_n1650__ & new_new_n1652__;
  assign new_new_n1655__ = ~new_new_n1653__ & ~new_new_n1654__;
  assign new_new_n1656__ = ~new_new_n1565__ & ~new_new_n1578__;
  assign new_new_n1657__ = new_new_n1565__ & new_new_n1578__;
  assign new_new_n1658__ = ~new_new_n1566__ & ~new_new_n1657__;
  assign new_new_n1659__ = ~new_new_n1656__ & ~new_new_n1658__;
  assign new_new_n1660__ = ~new_new_n1655__ & new_new_n1659__;
  assign new_new_n1661__ = new_new_n1655__ & ~new_new_n1659__;
  assign new_new_n1662__ = ~new_new_n1660__ & ~new_new_n1661__;
  assign new_new_n1663__ = new_new_n1577__ & new_new_n1587__;
  assign new_new_n1664__ = ~new_new_n1577__ & ~new_new_n1587__;
  assign new_new_n1665__ = ~new_new_n1656__ & ~new_new_n1657__;
  assign new_new_n1666__ = new_new_n1566__ & ~new_new_n1665__;
  assign new_new_n1667__ = ~new_new_n1566__ & new_new_n1665__;
  assign new_new_n1668__ = ~new_new_n1666__ & ~new_new_n1667__;
  assign new_new_n1669__ = ~new_new_n1664__ & new_new_n1668__;
  assign new_new_n1670__ = ~new_new_n1663__ & ~new_new_n1669__;
  assign new_new_n1671__ = ~new_new_n1662__ & new_new_n1670__;
  assign new_new_n1672__ = new_new_n1662__ & ~new_new_n1670__;
  assign new_new_n1673__ = ~new_new_n1671__ & ~new_new_n1672__;
  assign new_new_n1674__ = ~new_new_n1621__ & ~new_new_n1624__;
  assign new_new_n1675__ = ~new_new_n1620__ & ~new_new_n1674__;
  assign new_new_n1676__ = new_new_n1673__ & ~new_new_n1675__;
  assign new_new_n1677__ = ~new_new_n1673__ & new_new_n1675__;
  assign new_new_n1678__ = ~new_new_n1676__ & ~new_new_n1677__;
  assign new_new_n1679__ = new_new_n1648__ & new_new_n1678__;
  assign new_new_n1680__ = ~new_new_n1648__ & ~new_new_n1678__;
  assign new_new_n1681__ = ~new_new_n1679__ & ~new_new_n1680__;
  assign new_new_n1682__ = ~new_new_n1611__ & ~new_new_n1615__;
  assign new_new_n1683__ = new_new_n1614__ & ~new_new_n1682__;
  assign new_new_n1684__ = pi10 & pi14;
  assign new_new_n1685__ = pi08 & pi16;
  assign new_new_n1686__ = pi09 & pi15;
  assign new_new_n1687__ = ~new_new_n1685__ & ~new_new_n1686__;
  assign new_new_n1688__ = new_new_n1685__ & new_new_n1686__;
  assign new_new_n1689__ = ~new_new_n1687__ & ~new_new_n1688__;
  assign new_new_n1690__ = new_new_n1684__ & ~new_new_n1689__;
  assign new_new_n1691__ = ~new_new_n1684__ & new_new_n1689__;
  assign new_new_n1692__ = ~new_new_n1690__ & ~new_new_n1691__;
  assign new_new_n1693__ = new_new_n1683__ & ~new_new_n1692__;
  assign new_new_n1694__ = ~new_new_n1683__ & new_new_n1692__;
  assign new_new_n1695__ = ~new_new_n1693__ & ~new_new_n1694__;
  assign new_new_n1696__ = pi05 & pi19;
  assign new_new_n1697__ = pi04 & pi20;
  assign new_new_n1698__ = pi03 & pi21;
  assign new_new_n1699__ = ~new_new_n1697__ & ~new_new_n1698__;
  assign new_new_n1700__ = new_new_n1697__ & new_new_n1698__;
  assign new_new_n1701__ = ~new_new_n1699__ & ~new_new_n1700__;
  assign new_new_n1702__ = new_new_n1696__ & ~new_new_n1701__;
  assign new_new_n1703__ = ~new_new_n1696__ & new_new_n1701__;
  assign new_new_n1704__ = ~new_new_n1702__ & ~new_new_n1703__;
  assign new_new_n1705__ = new_new_n1695__ & ~new_new_n1704__;
  assign new_new_n1706__ = ~new_new_n1695__ & new_new_n1704__;
  assign new_new_n1707__ = ~new_new_n1705__ & ~new_new_n1706__;
  assign new_new_n1708__ = ~new_new_n1554__ & ~new_new_n1557__;
  assign new_new_n1709__ = ~new_new_n1553__ & ~new_new_n1708__;
  assign new_new_n1710__ = ~new_new_n1707__ & ~new_new_n1709__;
  assign new_new_n1711__ = new_new_n1707__ & new_new_n1709__;
  assign new_new_n1712__ = ~new_new_n1710__ & ~new_new_n1711__;
  assign new_new_n1713__ = ~new_new_n1538__ & ~new_new_n1544__;
  assign new_new_n1714__ = ~new_new_n1543__ & ~new_new_n1713__;
  assign new_new_n1715__ = pi07 & pi17;
  assign new_new_n1716__ = pi06 & pi18;
  assign new_new_n1717__ = pi02 & pi22;
  assign new_new_n1718__ = ~new_new_n1716__ & ~new_new_n1717__;
  assign new_new_n1719__ = new_new_n1716__ & new_new_n1717__;
  assign new_new_n1720__ = ~new_new_n1718__ & ~new_new_n1719__;
  assign new_new_n1721__ = new_new_n1715__ & ~new_new_n1720__;
  assign new_new_n1722__ = ~new_new_n1715__ & new_new_n1720__;
  assign new_new_n1723__ = ~new_new_n1721__ & ~new_new_n1722__;
  assign new_new_n1724__ = new_new_n1714__ & ~new_new_n1723__;
  assign new_new_n1725__ = ~new_new_n1714__ & new_new_n1723__;
  assign new_new_n1726__ = ~new_new_n1724__ & ~new_new_n1725__;
  assign new_new_n1727__ = pi00 & pi24;
  assign new_new_n1728__ = pi11 & pi13;
  assign new_new_n1729__ = pi01 & pi23;
  assign new_new_n1730__ = ~new_new_n1728__ & ~new_new_n1729__;
  assign new_new_n1731__ = new_new_n1728__ & new_new_n1729__;
  assign new_new_n1732__ = ~new_new_n1730__ & ~new_new_n1731__;
  assign new_new_n1733__ = ~new_new_n1727__ & ~new_new_n1732__;
  assign new_new_n1734__ = new_new_n1727__ & new_new_n1732__;
  assign new_new_n1735__ = ~new_new_n1733__ & ~new_new_n1734__;
  assign new_new_n1736__ = ~new_new_n1547__ & new_new_n1735__;
  assign new_new_n1737__ = new_new_n1537__ & ~new_new_n1735__;
  assign new_new_n1738__ = ~new_new_n1736__ & ~new_new_n1737__;
  assign new_new_n1739__ = ~new_new_n1726__ & new_new_n1738__;
  assign new_new_n1740__ = new_new_n1726__ & ~new_new_n1738__;
  assign new_new_n1741__ = ~new_new_n1739__ & ~new_new_n1740__;
  assign new_new_n1742__ = new_new_n1712__ & new_new_n1741__;
  assign new_new_n1743__ = ~new_new_n1712__ & ~new_new_n1741__;
  assign new_new_n1744__ = ~new_new_n1742__ & ~new_new_n1743__;
  assign new_new_n1745__ = new_new_n1681__ & ~new_new_n1744__;
  assign new_new_n1746__ = ~new_new_n1681__ & new_new_n1744__;
  assign new_new_n1747__ = ~new_new_n1745__ & ~new_new_n1746__;
  assign new_new_n1748__ = ~new_new_n1560__ & ~new_new_n1631__;
  assign new_new_n1749__ = ~new_new_n1632__ & ~new_new_n1748__;
  assign new_new_n1750__ = ~new_new_n1638__ & new_new_n1749__;
  assign new_new_n1751__ = ~new_new_n1639__ & ~new_new_n1749__;
  assign new_new_n1752__ = ~new_new_n1750__ & ~new_new_n1751__;
  assign new_new_n1753__ = ~new_new_n1560__ & new_new_n1632__;
  assign new_new_n1754__ = new_new_n1560__ & new_new_n1631__;
  assign new_new_n1755__ = ~new_new_n1753__ & ~new_new_n1754__;
  assign new_new_n1756__ = new_new_n1640__ & new_new_n1755__;
  assign new_new_n1757__ = new_new_n1747__ & ~new_new_n1752__;
  assign new_new_n1758__ = ~new_new_n1756__ & new_new_n1757__;
  assign new_new_n1759__ = ~new_new_n1630__ & new_new_n1638__;
  assign new_new_n1760__ = ~new_new_n1562__ & new_new_n1759__;
  assign new_new_n1761__ = new_new_n1630__ & ~new_new_n1638__;
  assign new_new_n1762__ = ~new_new_n1562__ & ~new_new_n1639__;
  assign new_new_n1763__ = ~new_new_n1761__ & new_new_n1762__;
  assign new_new_n1764__ = ~new_new_n1759__ & ~new_new_n1763__;
  assign new_new_n1765__ = ~new_new_n1560__ & ~new_new_n1764__;
  assign new_new_n1766__ = new_new_n1631__ & new_new_n1639__;
  assign new_new_n1767__ = ~new_new_n1632__ & new_new_n1639__;
  assign new_new_n1768__ = new_new_n1562__ & new_new_n1761__;
  assign new_new_n1769__ = ~new_new_n1767__ & ~new_new_n1768__;
  assign new_new_n1770__ = new_new_n1560__ & ~new_new_n1769__;
  assign new_new_n1771__ = ~new_new_n1747__ & ~new_new_n1766__;
  assign new_new_n1772__ = ~new_new_n1760__ & new_new_n1771__;
  assign new_new_n1773__ = ~new_new_n1765__ & new_new_n1772__;
  assign new_new_n1774__ = ~new_new_n1770__ & new_new_n1773__;
  assign po025 = ~new_new_n1758__ & ~new_new_n1774__;
  assign new_new_n1776__ = ~new_new_n1747__ & ~new_new_n1750__;
  assign new_new_n1777__ = new_new_n1638__ & ~new_new_n1749__;
  assign new_new_n1778__ = new_new_n1747__ & ~new_new_n1753__;
  assign new_new_n1779__ = ~new_new_n1754__ & ~new_new_n1778__;
  assign new_new_n1780__ = ~new_new_n1639__ & new_new_n1779__;
  assign new_new_n1781__ = ~new_new_n1777__ & ~new_new_n1780__;
  assign new_new_n1782__ = ~new_new_n1776__ & new_new_n1781__;
  assign new_new_n1783__ = ~new_new_n1680__ & ~new_new_n1744__;
  assign new_new_n1784__ = ~new_new_n1679__ & ~new_new_n1783__;
  assign new_new_n1785__ = new_new_n1782__ & ~new_new_n1784__;
  assign new_new_n1786__ = ~new_new_n1782__ & new_new_n1784__;
  assign new_new_n1787__ = ~new_new_n1785__ & ~new_new_n1786__;
  assign new_new_n1788__ = ~new_new_n1671__ & ~new_new_n1675__;
  assign new_new_n1789__ = ~new_new_n1672__ & ~new_new_n1788__;
  assign new_new_n1790__ = pi06 & pi19;
  assign new_new_n1791__ = pi04 & pi21;
  assign new_new_n1792__ = pi03 & pi22;
  assign new_new_n1793__ = ~new_new_n1791__ & ~new_new_n1792__;
  assign new_new_n1794__ = new_new_n1791__ & new_new_n1792__;
  assign new_new_n1795__ = ~new_new_n1793__ & ~new_new_n1794__;
  assign new_new_n1796__ = new_new_n1790__ & ~new_new_n1795__;
  assign new_new_n1797__ = ~new_new_n1790__ & new_new_n1795__;
  assign new_new_n1798__ = ~new_new_n1796__ & ~new_new_n1797__;
  assign new_new_n1799__ = pi07 & pi18;
  assign new_new_n1800__ = ~new_new_n1125__ & ~new_new_n1799__;
  assign new_new_n1801__ = new_new_n1125__ & new_new_n1799__;
  assign new_new_n1802__ = ~new_new_n1800__ & ~new_new_n1801__;
  assign new_new_n1803__ = new_new_n947__ & ~new_new_n1802__;
  assign new_new_n1804__ = ~new_new_n947__ & new_new_n1802__;
  assign new_new_n1805__ = ~new_new_n1803__ & ~new_new_n1804__;
  assign new_new_n1806__ = new_new_n1798__ & new_new_n1805__;
  assign new_new_n1807__ = ~new_new_n1798__ & ~new_new_n1805__;
  assign new_new_n1808__ = ~new_new_n1806__ & ~new_new_n1807__;
  assign new_new_n1809__ = pi10 & pi15;
  assign new_new_n1810__ = pi02 & pi23;
  assign new_new_n1811__ = pi00 & pi25;
  assign new_new_n1812__ = ~new_new_n1810__ & ~new_new_n1811__;
  assign new_new_n1813__ = new_new_n1810__ & new_new_n1811__;
  assign new_new_n1814__ = ~new_new_n1812__ & ~new_new_n1813__;
  assign new_new_n1815__ = new_new_n1809__ & ~new_new_n1814__;
  assign new_new_n1816__ = ~new_new_n1809__ & new_new_n1814__;
  assign new_new_n1817__ = ~new_new_n1815__ & ~new_new_n1816__;
  assign new_new_n1818__ = ~new_new_n1808__ & new_new_n1817__;
  assign new_new_n1819__ = new_new_n1808__ & ~new_new_n1817__;
  assign new_new_n1820__ = ~new_new_n1818__ & ~new_new_n1819__;
  assign new_new_n1821__ = new_new_n1789__ & new_new_n1820__;
  assign new_new_n1822__ = ~new_new_n1789__ & ~new_new_n1820__;
  assign new_new_n1823__ = ~new_new_n1821__ & ~new_new_n1822__;
  assign new_new_n1824__ = pi12 & pi13;
  assign new_new_n1825__ = pi05 & pi20;
  assign new_new_n1826__ = pi11 & pi14;
  assign new_new_n1827__ = ~new_new_n1825__ & ~new_new_n1826__;
  assign new_new_n1828__ = new_new_n1825__ & new_new_n1826__;
  assign new_new_n1829__ = ~new_new_n1827__ & ~new_new_n1828__;
  assign new_new_n1830__ = new_new_n1824__ & ~new_new_n1829__;
  assign new_new_n1831__ = ~new_new_n1824__ & new_new_n1829__;
  assign new_new_n1832__ = ~new_new_n1830__ & ~new_new_n1831__;
  assign new_new_n1833__ = ~new_new_n1654__ & ~new_new_n1659__;
  assign new_new_n1834__ = ~new_new_n1653__ & ~new_new_n1833__;
  assign new_new_n1835__ = pi11 & pi23;
  assign new_new_n1836__ = ~new_new_n1696__ & ~new_new_n1700__;
  assign new_new_n1837__ = ~new_new_n1699__ & ~new_new_n1836__;
  assign new_new_n1838__ = pi01 & ~pi24;
  assign new_new_n1839__ = ~new_new_n1837__ & ~new_new_n1838__;
  assign new_new_n1840__ = new_new_n1835__ & ~new_new_n1839__;
  assign new_new_n1841__ = pi13 & pi24;
  assign new_new_n1842__ = new_new_n1837__ & ~new_new_n1841__;
  assign new_new_n1843__ = new_new_n1840__ & ~new_new_n1842__;
  assign new_new_n1844__ = pi01 & pi24;
  assign new_new_n1845__ = new_new_n1837__ & ~new_new_n1844__;
  assign new_new_n1846__ = ~new_new_n1837__ & new_new_n1844__;
  assign new_new_n1847__ = ~new_new_n1845__ & ~new_new_n1846__;
  assign new_new_n1848__ = pi13 & new_new_n1847__;
  assign new_new_n1849__ = ~pi13 & ~new_new_n1847__;
  assign new_new_n1850__ = ~new_new_n1731__ & ~new_new_n1848__;
  assign new_new_n1851__ = ~new_new_n1849__ & new_new_n1850__;
  assign new_new_n1852__ = ~new_new_n1843__ & ~new_new_n1851__;
  assign new_new_n1853__ = new_new_n1834__ & new_new_n1852__;
  assign new_new_n1854__ = ~new_new_n1834__ & ~new_new_n1852__;
  assign new_new_n1855__ = new_new_n1832__ & ~new_new_n1853__;
  assign new_new_n1856__ = ~new_new_n1854__ & ~new_new_n1855__;
  assign new_new_n1857__ = ~new_new_n1853__ & new_new_n1856__;
  assign new_new_n1858__ = ~new_new_n1832__ & ~new_new_n1857__;
  assign new_new_n1859__ = ~new_new_n1854__ & new_new_n1855__;
  assign new_new_n1860__ = ~new_new_n1858__ & ~new_new_n1859__;
  assign new_new_n1861__ = new_new_n1823__ & ~new_new_n1860__;
  assign new_new_n1862__ = ~new_new_n1823__ & new_new_n1860__;
  assign new_new_n1863__ = ~new_new_n1861__ & ~new_new_n1862__;
  assign new_new_n1864__ = ~new_new_n1715__ & ~new_new_n1719__;
  assign new_new_n1865__ = ~new_new_n1718__ & ~new_new_n1864__;
  assign new_new_n1866__ = ~new_new_n1537__ & ~new_new_n1734__;
  assign new_new_n1867__ = ~new_new_n1733__ & ~new_new_n1866__;
  assign new_new_n1868__ = ~new_new_n1865__ & ~new_new_n1867__;
  assign new_new_n1869__ = new_new_n1865__ & new_new_n1867__;
  assign new_new_n1870__ = ~new_new_n1868__ & ~new_new_n1869__;
  assign new_new_n1871__ = ~new_new_n1684__ & ~new_new_n1688__;
  assign new_new_n1872__ = ~new_new_n1687__ & ~new_new_n1871__;
  assign new_new_n1873__ = ~new_new_n1870__ & new_new_n1872__;
  assign new_new_n1874__ = new_new_n1870__ & ~new_new_n1872__;
  assign new_new_n1875__ = ~new_new_n1873__ & ~new_new_n1874__;
  assign new_new_n1876__ = ~new_new_n1725__ & ~new_new_n1738__;
  assign new_new_n1877__ = ~new_new_n1724__ & ~new_new_n1876__;
  assign new_new_n1878__ = ~new_new_n1694__ & ~new_new_n1704__;
  assign new_new_n1879__ = ~new_new_n1693__ & ~new_new_n1878__;
  assign new_new_n1880__ = new_new_n1877__ & new_new_n1879__;
  assign new_new_n1881__ = ~new_new_n1877__ & ~new_new_n1879__;
  assign new_new_n1882__ = ~new_new_n1880__ & ~new_new_n1881__;
  assign new_new_n1883__ = new_new_n1875__ & new_new_n1882__;
  assign new_new_n1884__ = ~new_new_n1875__ & ~new_new_n1882__;
  assign new_new_n1885__ = ~new_new_n1883__ & ~new_new_n1884__;
  assign new_new_n1886__ = ~new_new_n1863__ & new_new_n1885__;
  assign new_new_n1887__ = new_new_n1863__ & ~new_new_n1885__;
  assign new_new_n1888__ = ~new_new_n1886__ & ~new_new_n1887__;
  assign new_new_n1889__ = ~new_new_n1711__ & ~new_new_n1741__;
  assign new_new_n1890__ = ~new_new_n1710__ & ~new_new_n1889__;
  assign new_new_n1891__ = new_new_n1888__ & ~new_new_n1890__;
  assign new_new_n1892__ = ~new_new_n1888__ & new_new_n1890__;
  assign new_new_n1893__ = ~new_new_n1891__ & ~new_new_n1892__;
  assign new_new_n1894__ = new_new_n1787__ & new_new_n1893__;
  assign new_new_n1895__ = ~new_new_n1787__ & ~new_new_n1893__;
  assign po026 = new_new_n1894__ | new_new_n1895__;
  assign new_new_n1897__ = ~new_new_n1806__ & ~new_new_n1817__;
  assign new_new_n1898__ = ~new_new_n1807__ & ~new_new_n1897__;
  assign new_new_n1899__ = ~new_new_n1824__ & ~new_new_n1828__;
  assign new_new_n1900__ = ~new_new_n1827__ & ~new_new_n1899__;
  assign new_new_n1901__ = ~new_new_n1790__ & ~new_new_n1794__;
  assign new_new_n1902__ = ~new_new_n1793__ & ~new_new_n1901__;
  assign new_new_n1903__ = ~new_new_n1900__ & ~new_new_n1902__;
  assign new_new_n1904__ = new_new_n1900__ & new_new_n1902__;
  assign new_new_n1905__ = ~new_new_n1903__ & ~new_new_n1904__;
  assign new_new_n1906__ = pi12 & pi14;
  assign new_new_n1907__ = pi01 & pi25;
  assign new_new_n1908__ = ~new_new_n1906__ & new_new_n1907__;
  assign new_new_n1909__ = new_new_n1906__ & ~new_new_n1907__;
  assign new_new_n1910__ = ~new_new_n1908__ & ~new_new_n1909__;
  assign new_new_n1911__ = new_new_n1905__ & new_new_n1910__;
  assign new_new_n1912__ = ~new_new_n1905__ & ~new_new_n1910__;
  assign new_new_n1913__ = ~new_new_n1911__ & ~new_new_n1912__;
  assign new_new_n1914__ = ~new_new_n1898__ & ~new_new_n1913__;
  assign new_new_n1915__ = new_new_n1898__ & new_new_n1913__;
  assign new_new_n1916__ = ~new_new_n1914__ & ~new_new_n1915__;
  assign new_new_n1917__ = ~new_new_n1856__ & ~new_new_n1916__;
  assign new_new_n1918__ = new_new_n1856__ & new_new_n1916__;
  assign new_new_n1919__ = ~new_new_n1917__ & ~new_new_n1918__;
  assign new_new_n1920__ = ~new_new_n1821__ & new_new_n1860__;
  assign new_new_n1921__ = ~new_new_n1822__ & ~new_new_n1920__;
  assign new_new_n1922__ = ~new_new_n1869__ & ~new_new_n1872__;
  assign new_new_n1923__ = ~new_new_n1868__ & ~new_new_n1922__;
  assign new_new_n1924__ = pi08 & pi18;
  assign new_new_n1925__ = pi24 & new_new_n737__;
  assign new_new_n1926__ = ~new_new_n947__ & ~new_new_n1801__;
  assign new_new_n1927__ = ~new_new_n1800__ & ~new_new_n1926__;
  assign new_new_n1928__ = new_new_n1925__ & ~new_new_n1927__;
  assign new_new_n1929__ = ~new_new_n1925__ & new_new_n1927__;
  assign new_new_n1930__ = ~new_new_n1928__ & ~new_new_n1929__;
  assign new_new_n1931__ = new_new_n1924__ & ~new_new_n1930__;
  assign new_new_n1932__ = ~new_new_n1924__ & new_new_n1930__;
  assign new_new_n1933__ = ~new_new_n1931__ & ~new_new_n1932__;
  assign new_new_n1934__ = pi00 & pi26;
  assign new_new_n1935__ = ~new_new_n1809__ & ~new_new_n1813__;
  assign new_new_n1936__ = ~new_new_n1812__ & ~new_new_n1935__;
  assign new_new_n1937__ = new_new_n1934__ & ~new_new_n1936__;
  assign new_new_n1938__ = ~new_new_n1934__ & new_new_n1936__;
  assign new_new_n1939__ = ~new_new_n1937__ & ~new_new_n1938__;
  assign new_new_n1940__ = new_new_n1933__ & new_new_n1939__;
  assign new_new_n1941__ = ~new_new_n1933__ & ~new_new_n1939__;
  assign new_new_n1942__ = ~new_new_n1940__ & ~new_new_n1941__;
  assign new_new_n1943__ = ~new_new_n1840__ & ~new_new_n1845__;
  assign new_new_n1944__ = pi13 & ~new_new_n1943__;
  assign new_new_n1945__ = ~pi13 & new_new_n1844__;
  assign new_new_n1946__ = new_new_n1837__ & new_new_n1945__;
  assign new_new_n1947__ = ~new_new_n1944__ & ~new_new_n1946__;
  assign new_new_n1948__ = new_new_n1942__ & new_new_n1947__;
  assign new_new_n1949__ = ~new_new_n1942__ & ~new_new_n1947__;
  assign new_new_n1950__ = ~new_new_n1948__ & ~new_new_n1949__;
  assign new_new_n1951__ = new_new_n1923__ & ~new_new_n1950__;
  assign new_new_n1952__ = ~new_new_n1923__ & new_new_n1950__;
  assign new_new_n1953__ = ~new_new_n1951__ & ~new_new_n1952__;
  assign new_new_n1954__ = ~new_new_n1875__ & ~new_new_n1880__;
  assign new_new_n1955__ = ~new_new_n1881__ & ~new_new_n1954__;
  assign new_new_n1956__ = ~new_new_n1953__ & ~new_new_n1955__;
  assign new_new_n1957__ = new_new_n1953__ & new_new_n1955__;
  assign new_new_n1958__ = ~new_new_n1956__ & ~new_new_n1957__;
  assign new_new_n1959__ = pi11 & pi15;
  assign new_new_n1960__ = pi09 & pi17;
  assign new_new_n1961__ = pi10 & pi16;
  assign new_new_n1962__ = ~new_new_n1960__ & ~new_new_n1961__;
  assign new_new_n1963__ = new_new_n1960__ & new_new_n1961__;
  assign new_new_n1964__ = ~new_new_n1962__ & ~new_new_n1963__;
  assign new_new_n1965__ = new_new_n1959__ & ~new_new_n1964__;
  assign new_new_n1966__ = ~new_new_n1959__ & new_new_n1964__;
  assign new_new_n1967__ = ~new_new_n1965__ & ~new_new_n1966__;
  assign new_new_n1968__ = pi06 & pi20;
  assign new_new_n1969__ = pi04 & pi22;
  assign new_new_n1970__ = pi05 & pi21;
  assign new_new_n1971__ = ~new_new_n1969__ & ~new_new_n1970__;
  assign new_new_n1972__ = new_new_n1969__ & new_new_n1970__;
  assign new_new_n1973__ = ~new_new_n1971__ & ~new_new_n1972__;
  assign new_new_n1974__ = new_new_n1968__ & ~new_new_n1973__;
  assign new_new_n1975__ = ~new_new_n1968__ & new_new_n1973__;
  assign new_new_n1976__ = ~new_new_n1974__ & ~new_new_n1975__;
  assign new_new_n1977__ = new_new_n1967__ & new_new_n1976__;
  assign new_new_n1978__ = ~new_new_n1967__ & ~new_new_n1976__;
  assign new_new_n1979__ = ~new_new_n1977__ & ~new_new_n1978__;
  assign new_new_n1980__ = pi07 & pi19;
  assign new_new_n1981__ = pi03 & pi23;
  assign new_new_n1982__ = pi02 & pi24;
  assign new_new_n1983__ = ~new_new_n1981__ & ~new_new_n1982__;
  assign new_new_n1984__ = new_new_n1981__ & new_new_n1982__;
  assign new_new_n1985__ = ~new_new_n1983__ & ~new_new_n1984__;
  assign new_new_n1986__ = new_new_n1980__ & ~new_new_n1985__;
  assign new_new_n1987__ = ~new_new_n1980__ & new_new_n1985__;
  assign new_new_n1988__ = ~new_new_n1986__ & ~new_new_n1987__;
  assign new_new_n1989__ = new_new_n1979__ & ~new_new_n1988__;
  assign new_new_n1990__ = ~new_new_n1979__ & new_new_n1988__;
  assign new_new_n1991__ = ~new_new_n1989__ & ~new_new_n1990__;
  assign new_new_n1992__ = new_new_n1958__ & ~new_new_n1991__;
  assign new_new_n1993__ = ~new_new_n1958__ & new_new_n1991__;
  assign new_new_n1994__ = ~new_new_n1992__ & ~new_new_n1993__;
  assign new_new_n1995__ = new_new_n1921__ & ~new_new_n1994__;
  assign new_new_n1996__ = ~new_new_n1921__ & new_new_n1994__;
  assign new_new_n1997__ = ~new_new_n1995__ & ~new_new_n1996__;
  assign new_new_n1998__ = new_new_n1919__ & ~new_new_n1997__;
  assign new_new_n1999__ = ~new_new_n1919__ & new_new_n1997__;
  assign new_new_n2000__ = ~new_new_n1998__ & ~new_new_n1999__;
  assign new_new_n2001__ = new_new_n1887__ & new_new_n1890__;
  assign new_new_n2002__ = new_new_n1886__ & ~new_new_n1890__;
  assign new_new_n2003__ = ~new_new_n2001__ & ~new_new_n2002__;
  assign new_new_n2004__ = new_new_n1787__ & new_new_n2003__;
  assign new_new_n2005__ = ~new_new_n1887__ & ~new_new_n1890__;
  assign new_new_n2006__ = ~new_new_n1886__ & ~new_new_n2005__;
  assign new_new_n2007__ = new_new_n1786__ & ~new_new_n2006__;
  assign new_new_n2008__ = new_new_n1785__ & new_new_n2006__;
  assign new_new_n2009__ = ~new_new_n2007__ & ~new_new_n2008__;
  assign new_new_n2010__ = ~new_new_n2004__ & new_new_n2009__;
  assign new_new_n2011__ = new_new_n2000__ & ~new_new_n2010__;
  assign new_new_n2012__ = new_new_n1782__ & new_new_n1885__;
  assign new_new_n2013__ = ~new_new_n1782__ & ~new_new_n1885__;
  assign new_new_n2014__ = ~new_new_n1784__ & ~new_new_n2013__;
  assign new_new_n2015__ = ~new_new_n2012__ & ~new_new_n2014__;
  assign new_new_n2016__ = new_new_n1863__ & new_new_n2015__;
  assign new_new_n2017__ = new_new_n1786__ & ~new_new_n1885__;
  assign new_new_n2018__ = ~new_new_n2016__ & ~new_new_n2017__;
  assign new_new_n2019__ = new_new_n1890__ & ~new_new_n2018__;
  assign new_new_n2020__ = ~new_new_n1863__ & ~new_new_n2015__;
  assign new_new_n2021__ = new_new_n1785__ & new_new_n1885__;
  assign new_new_n2022__ = ~new_new_n2020__ & ~new_new_n2021__;
  assign new_new_n2023__ = ~new_new_n1890__ & ~new_new_n2022__;
  assign new_new_n2024__ = new_new_n1784__ & new_new_n1863__;
  assign new_new_n2025__ = ~new_new_n2012__ & ~new_new_n2024__;
  assign new_new_n2026__ = ~new_new_n1784__ & ~new_new_n1863__;
  assign new_new_n2027__ = ~new_new_n2013__ & ~new_new_n2026__;
  assign new_new_n2028__ = ~new_new_n2025__ & ~new_new_n2027__;
  assign new_new_n2029__ = ~new_new_n2019__ & ~new_new_n2028__;
  assign new_new_n2030__ = ~new_new_n2023__ & new_new_n2029__;
  assign new_new_n2031__ = ~new_new_n2000__ & ~new_new_n2030__;
  assign po027 = new_new_n2011__ | new_new_n2031__;
  assign new_new_n2033__ = ~new_new_n1956__ & ~new_new_n1991__;
  assign new_new_n2034__ = ~new_new_n1957__ & ~new_new_n2033__;
  assign new_new_n2035__ = new_new_n1923__ & ~new_new_n1948__;
  assign new_new_n2036__ = ~new_new_n1949__ & ~new_new_n2035__;
  assign new_new_n2037__ = ~new_new_n1980__ & ~new_new_n1984__;
  assign new_new_n2038__ = ~new_new_n1983__ & ~new_new_n2037__;
  assign new_new_n2039__ = ~new_new_n1959__ & ~new_new_n1963__;
  assign new_new_n2040__ = ~new_new_n1962__ & ~new_new_n2039__;
  assign new_new_n2041__ = ~new_new_n1968__ & ~new_new_n1972__;
  assign new_new_n2042__ = ~new_new_n1971__ & ~new_new_n2041__;
  assign new_new_n2043__ = new_new_n2040__ & new_new_n2042__;
  assign new_new_n2044__ = ~new_new_n2040__ & ~new_new_n2042__;
  assign new_new_n2045__ = ~new_new_n2043__ & ~new_new_n2044__;
  assign new_new_n2046__ = new_new_n2038__ & ~new_new_n2045__;
  assign new_new_n2047__ = ~new_new_n2038__ & new_new_n2045__;
  assign new_new_n2048__ = ~new_new_n2046__ & ~new_new_n2047__;
  assign new_new_n2049__ = ~new_new_n2036__ & ~new_new_n2048__;
  assign new_new_n2050__ = new_new_n2036__ & new_new_n2048__;
  assign new_new_n2051__ = ~new_new_n2049__ & ~new_new_n2050__;
  assign new_new_n2052__ = pi13 & pi14;
  assign new_new_n2053__ = pi05 & pi22;
  assign new_new_n2054__ = pi12 & pi15;
  assign new_new_n2055__ = ~new_new_n2053__ & ~new_new_n2054__;
  assign new_new_n2056__ = new_new_n2053__ & new_new_n2054__;
  assign new_new_n2057__ = ~new_new_n2055__ & ~new_new_n2056__;
  assign new_new_n2058__ = new_new_n2052__ & ~new_new_n2057__;
  assign new_new_n2059__ = ~new_new_n2052__ & new_new_n2057__;
  assign new_new_n2060__ = ~new_new_n2058__ & ~new_new_n2059__;
  assign new_new_n2061__ = pi12 & pi25;
  assign new_new_n2062__ = pi01 & new_new_n2061__;
  assign new_new_n2063__ = pi14 & ~new_new_n2062__;
  assign new_new_n2064__ = pi00 & pi27;
  assign new_new_n2065__ = pi01 & pi26;
  assign new_new_n2066__ = new_new_n2064__ & ~new_new_n2065__;
  assign new_new_n2067__ = ~new_new_n2064__ & new_new_n2065__;
  assign new_new_n2068__ = ~new_new_n2066__ & ~new_new_n2067__;
  assign new_new_n2069__ = new_new_n2063__ & new_new_n2068__;
  assign new_new_n2070__ = ~new_new_n2063__ & ~new_new_n2068__;
  assign new_new_n2071__ = ~new_new_n2069__ & ~new_new_n2070__;
  assign new_new_n2072__ = ~new_new_n2060__ & ~new_new_n2071__;
  assign new_new_n2073__ = new_new_n2060__ & new_new_n2071__;
  assign new_new_n2074__ = ~new_new_n2072__ & ~new_new_n2073__;
  assign new_new_n2075__ = pi06 & pi21;
  assign new_new_n2076__ = pi03 & pi24;
  assign new_new_n2077__ = pi04 & pi23;
  assign new_new_n2078__ = ~new_new_n2076__ & ~new_new_n2077__;
  assign new_new_n2079__ = new_new_n2076__ & new_new_n2077__;
  assign new_new_n2080__ = ~new_new_n2078__ & ~new_new_n2079__;
  assign new_new_n2081__ = new_new_n2075__ & ~new_new_n2080__;
  assign new_new_n2082__ = ~new_new_n2075__ & new_new_n2080__;
  assign new_new_n2083__ = ~new_new_n2081__ & ~new_new_n2082__;
  assign new_new_n2084__ = new_new_n2074__ & ~new_new_n2083__;
  assign new_new_n2085__ = ~new_new_n2074__ & new_new_n2083__;
  assign new_new_n2086__ = ~new_new_n2084__ & ~new_new_n2085__;
  assign new_new_n2087__ = new_new_n2051__ & ~new_new_n2086__;
  assign new_new_n2088__ = ~new_new_n2051__ & new_new_n2086__;
  assign new_new_n2089__ = ~new_new_n2087__ & ~new_new_n2088__;
  assign new_new_n2090__ = new_new_n2034__ & ~new_new_n2089__;
  assign new_new_n2091__ = ~new_new_n2034__ & new_new_n2089__;
  assign new_new_n2092__ = ~new_new_n2090__ & ~new_new_n2091__;
  assign new_new_n2093__ = ~new_new_n1914__ & ~new_new_n1918__;
  assign new_new_n2094__ = ~new_new_n1977__ & ~new_new_n1988__;
  assign new_new_n2095__ = ~new_new_n1978__ & ~new_new_n2094__;
  assign new_new_n2096__ = ~new_new_n1927__ & ~new_new_n1936__;
  assign new_new_n2097__ = new_new_n1927__ & new_new_n1936__;
  assign new_new_n2098__ = new_new_n1924__ & new_new_n1925__;
  assign new_new_n2099__ = ~new_new_n1924__ & ~new_new_n1925__;
  assign new_new_n2100__ = ~new_new_n2098__ & ~new_new_n2099__;
  assign new_new_n2101__ = new_new_n1934__ & ~new_new_n2100__;
  assign new_new_n2102__ = ~new_new_n1934__ & new_new_n2100__;
  assign new_new_n2103__ = ~new_new_n2097__ & ~new_new_n2101__;
  assign new_new_n2104__ = ~new_new_n2102__ & new_new_n2103__;
  assign new_new_n2105__ = ~new_new_n2096__ & ~new_new_n2104__;
  assign new_new_n2106__ = ~new_new_n1903__ & ~new_new_n1910__;
  assign new_new_n2107__ = ~new_new_n1904__ & ~new_new_n2106__;
  assign new_new_n2108__ = ~new_new_n2105__ & new_new_n2107__;
  assign new_new_n2109__ = new_new_n2105__ & ~new_new_n2107__;
  assign new_new_n2110__ = ~new_new_n2108__ & ~new_new_n2109__;
  assign new_new_n2111__ = new_new_n2095__ & new_new_n2110__;
  assign new_new_n2112__ = ~new_new_n2095__ & ~new_new_n2110__;
  assign new_new_n2113__ = ~new_new_n2111__ & ~new_new_n2112__;
  assign new_new_n2114__ = new_new_n2093__ & new_new_n2113__;
  assign new_new_n2115__ = ~new_new_n2093__ & ~new_new_n2113__;
  assign new_new_n2116__ = ~new_new_n2114__ & ~new_new_n2115__;
  assign new_new_n2117__ = pi11 & pi16;
  assign new_new_n2118__ = pi07 & pi20;
  assign new_new_n2119__ = pi02 & pi25;
  assign new_new_n2120__ = ~new_new_n2118__ & ~new_new_n2119__;
  assign new_new_n2121__ = new_new_n2118__ & new_new_n2119__;
  assign new_new_n2122__ = ~new_new_n2120__ & ~new_new_n2121__;
  assign new_new_n2123__ = new_new_n2117__ & ~new_new_n2122__;
  assign new_new_n2124__ = ~new_new_n2117__ & new_new_n2122__;
  assign new_new_n2125__ = ~new_new_n2123__ & ~new_new_n2124__;
  assign new_new_n2126__ = pi10 & pi17;
  assign new_new_n2127__ = pi09 & pi18;
  assign new_new_n2128__ = pi08 & pi19;
  assign new_new_n2129__ = ~new_new_n2127__ & ~new_new_n2128__;
  assign new_new_n2130__ = new_new_n2127__ & new_new_n2128__;
  assign new_new_n2131__ = ~new_new_n2129__ & ~new_new_n2130__;
  assign new_new_n2132__ = new_new_n2126__ & ~new_new_n2131__;
  assign new_new_n2133__ = ~new_new_n2126__ & new_new_n2131__;
  assign new_new_n2134__ = ~new_new_n2132__ & ~new_new_n2133__;
  assign new_new_n2135__ = new_new_n2125__ & new_new_n2134__;
  assign new_new_n2136__ = ~new_new_n2125__ & ~new_new_n2134__;
  assign new_new_n2137__ = ~new_new_n2135__ & ~new_new_n2136__;
  assign new_new_n2138__ = ~new_new_n1934__ & ~new_new_n2098__;
  assign new_new_n2139__ = ~new_new_n2099__ & ~new_new_n2138__;
  assign new_new_n2140__ = new_new_n2137__ & new_new_n2139__;
  assign new_new_n2141__ = ~new_new_n2137__ & ~new_new_n2139__;
  assign new_new_n2142__ = ~new_new_n2140__ & ~new_new_n2141__;
  assign new_new_n2143__ = new_new_n2116__ & ~new_new_n2142__;
  assign new_new_n2144__ = ~new_new_n2116__ & new_new_n2142__;
  assign new_new_n2145__ = ~new_new_n2143__ & ~new_new_n2144__;
  assign new_new_n2146__ = new_new_n2092__ & new_new_n2145__;
  assign new_new_n2147__ = ~new_new_n2092__ & ~new_new_n2145__;
  assign new_new_n2148__ = ~new_new_n2146__ & ~new_new_n2147__;
  assign new_new_n2149__ = ~new_new_n1890__ & ~new_new_n2024__;
  assign new_new_n2150__ = new_new_n2000__ & ~new_new_n2013__;
  assign new_new_n2151__ = ~new_new_n2026__ & ~new_new_n2149__;
  assign new_new_n2152__ = ~new_new_n2150__ & new_new_n2151__;
  assign new_new_n2153__ = ~new_new_n1890__ & new_new_n2026__;
  assign new_new_n2154__ = ~new_new_n2000__ & ~new_new_n2153__;
  assign new_new_n2155__ = new_new_n1890__ & new_new_n2024__;
  assign new_new_n2156__ = ~new_new_n2154__ & ~new_new_n2155__;
  assign new_new_n2157__ = ~new_new_n2012__ & ~new_new_n2156__;
  assign new_new_n2158__ = ~new_new_n2000__ & new_new_n2013__;
  assign new_new_n2159__ = ~new_new_n2157__ & ~new_new_n2158__;
  assign new_new_n2160__ = ~new_new_n2152__ & new_new_n2159__;
  assign new_new_n2161__ = ~new_new_n2148__ & ~new_new_n2160__;
  assign new_new_n2162__ = new_new_n2148__ & new_new_n2160__;
  assign new_new_n2163__ = ~new_new_n2161__ & ~new_new_n2162__;
  assign new_new_n2164__ = new_new_n1919__ & ~new_new_n1996__;
  assign new_new_n2165__ = ~new_new_n1995__ & ~new_new_n2164__;
  assign new_new_n2166__ = new_new_n2163__ & ~new_new_n2165__;
  assign new_new_n2167__ = ~new_new_n2163__ & new_new_n2165__;
  assign po028 = ~new_new_n2166__ & ~new_new_n2167__;
  assign new_new_n2169__ = ~new_new_n2089__ & ~new_new_n2113__;
  assign new_new_n2170__ = new_new_n2034__ & ~new_new_n2093__;
  assign new_new_n2171__ = new_new_n2169__ & new_new_n2170__;
  assign new_new_n2172__ = ~new_new_n2095__ & ~new_new_n2108__;
  assign new_new_n2173__ = ~new_new_n2109__ & ~new_new_n2172__;
  assign new_new_n2174__ = pi02 & pi26;
  assign new_new_n2175__ = ~new_new_n1320__ & ~new_new_n2174__;
  assign new_new_n2176__ = new_new_n1320__ & new_new_n2174__;
  assign new_new_n2177__ = ~new_new_n2175__ & ~new_new_n2176__;
  assign new_new_n2178__ = new_new_n1123__ & ~new_new_n2177__;
  assign new_new_n2179__ = ~new_new_n1123__ & new_new_n2177__;
  assign new_new_n2180__ = ~new_new_n2178__ & ~new_new_n2179__;
  assign new_new_n2181__ = pi12 & pi16;
  assign new_new_n2182__ = pi11 & pi17;
  assign new_new_n2183__ = pi00 & pi28;
  assign new_new_n2184__ = ~new_new_n2182__ & ~new_new_n2183__;
  assign new_new_n2185__ = new_new_n2182__ & new_new_n2183__;
  assign new_new_n2186__ = ~new_new_n2184__ & ~new_new_n2185__;
  assign new_new_n2187__ = new_new_n2181__ & ~new_new_n2186__;
  assign new_new_n2188__ = ~new_new_n2181__ & new_new_n2186__;
  assign new_new_n2189__ = ~new_new_n2187__ & ~new_new_n2188__;
  assign new_new_n2190__ = ~new_new_n2180__ & ~new_new_n2189__;
  assign new_new_n2191__ = new_new_n2180__ & new_new_n2189__;
  assign new_new_n2192__ = ~new_new_n2190__ & ~new_new_n2191__;
  assign new_new_n2193__ = ~new_new_n2038__ & ~new_new_n2043__;
  assign new_new_n2194__ = ~new_new_n2044__ & ~new_new_n2193__;
  assign new_new_n2195__ = new_new_n2192__ & ~new_new_n2194__;
  assign new_new_n2196__ = ~new_new_n2192__ & new_new_n2194__;
  assign new_new_n2197__ = ~new_new_n2195__ & ~new_new_n2196__;
  assign new_new_n2198__ = new_new_n2173__ & new_new_n2197__;
  assign new_new_n2199__ = ~new_new_n2173__ & ~new_new_n2197__;
  assign new_new_n2200__ = ~new_new_n2198__ & ~new_new_n2199__;
  assign new_new_n2201__ = ~new_new_n2126__ & ~new_new_n2130__;
  assign new_new_n2202__ = ~new_new_n2129__ & ~new_new_n2201__;
  assign new_new_n2203__ = ~new_new_n2117__ & ~new_new_n2121__;
  assign new_new_n2204__ = ~new_new_n2120__ & ~new_new_n2203__;
  assign new_new_n2205__ = ~new_new_n2075__ & ~new_new_n2079__;
  assign new_new_n2206__ = ~new_new_n2078__ & ~new_new_n2205__;
  assign new_new_n2207__ = ~new_new_n2204__ & ~new_new_n2206__;
  assign new_new_n2208__ = new_new_n2204__ & new_new_n2206__;
  assign new_new_n2209__ = ~new_new_n2207__ & ~new_new_n2208__;
  assign new_new_n2210__ = new_new_n2202__ & ~new_new_n2209__;
  assign new_new_n2211__ = ~new_new_n2202__ & new_new_n2209__;
  assign new_new_n2212__ = ~new_new_n2210__ & ~new_new_n2211__;
  assign new_new_n2213__ = new_new_n2200__ & new_new_n2212__;
  assign new_new_n2214__ = ~new_new_n2200__ & ~new_new_n2212__;
  assign new_new_n2215__ = ~new_new_n2213__ & ~new_new_n2214__;
  assign new_new_n2216__ = new_new_n2091__ & new_new_n2113__;
  assign new_new_n2217__ = ~new_new_n2091__ & ~new_new_n2113__;
  assign new_new_n2218__ = ~new_new_n2090__ & ~new_new_n2217__;
  assign new_new_n2219__ = new_new_n2093__ & new_new_n2218__;
  assign new_new_n2220__ = ~new_new_n2142__ & ~new_new_n2216__;
  assign new_new_n2221__ = ~new_new_n2219__ & new_new_n2220__;
  assign new_new_n2222__ = new_new_n2090__ & ~new_new_n2113__;
  assign new_new_n2223__ = ~new_new_n2093__ & ~new_new_n2218__;
  assign new_new_n2224__ = new_new_n2142__ & ~new_new_n2222__;
  assign new_new_n2225__ = ~new_new_n2223__ & new_new_n2224__;
  assign new_new_n2226__ = ~new_new_n2221__ & ~new_new_n2225__;
  assign new_new_n2227__ = new_new_n2089__ & new_new_n2113__;
  assign new_new_n2228__ = ~new_new_n2034__ & new_new_n2093__;
  assign new_new_n2229__ = new_new_n2227__ & new_new_n2228__;
  assign new_new_n2230__ = ~new_new_n2171__ & new_new_n2215__;
  assign new_new_n2231__ = ~new_new_n2229__ & new_new_n2230__;
  assign new_new_n2232__ = ~new_new_n2226__ & new_new_n2231__;
  assign new_new_n2233__ = ~new_new_n2114__ & new_new_n2142__;
  assign new_new_n2234__ = ~new_new_n2115__ & ~new_new_n2233__;
  assign new_new_n2235__ = new_new_n2090__ & new_new_n2234__;
  assign new_new_n2236__ = new_new_n2115__ & new_new_n2142__;
  assign new_new_n2237__ = new_new_n2114__ & ~new_new_n2142__;
  assign new_new_n2238__ = ~new_new_n2236__ & ~new_new_n2237__;
  assign new_new_n2239__ = new_new_n2092__ & new_new_n2238__;
  assign new_new_n2240__ = new_new_n2091__ & ~new_new_n2234__;
  assign new_new_n2241__ = ~new_new_n2215__ & ~new_new_n2235__;
  assign new_new_n2242__ = ~new_new_n2240__ & new_new_n2241__;
  assign new_new_n2243__ = ~new_new_n2239__ & new_new_n2242__;
  assign new_new_n2244__ = ~new_new_n2232__ & ~new_new_n2243__;
  assign new_new_n2245__ = ~new_new_n2162__ & ~new_new_n2165__;
  assign new_new_n2246__ = ~new_new_n2161__ & ~new_new_n2245__;
  assign new_new_n2247__ = new_new_n2244__ & new_new_n2246__;
  assign new_new_n2248__ = ~new_new_n2244__ & ~new_new_n2246__;
  assign new_new_n2249__ = ~new_new_n2247__ & ~new_new_n2248__;
  assign new_new_n2250__ = ~new_new_n2049__ & ~new_new_n2086__;
  assign new_new_n2251__ = ~new_new_n2050__ & ~new_new_n2250__;
  assign new_new_n2252__ = pi07 & pi21;
  assign new_new_n2253__ = pi06 & pi22;
  assign new_new_n2254__ = pi05 & pi23;
  assign new_new_n2255__ = ~new_new_n2253__ & ~new_new_n2254__;
  assign new_new_n2256__ = new_new_n2253__ & new_new_n2254__;
  assign new_new_n2257__ = ~new_new_n2255__ & ~new_new_n2256__;
  assign new_new_n2258__ = new_new_n2252__ & ~new_new_n2257__;
  assign new_new_n2259__ = ~new_new_n2252__ & new_new_n2257__;
  assign new_new_n2260__ = ~new_new_n2258__ & ~new_new_n2259__;
  assign new_new_n2261__ = pi26 & ~new_new_n2064__;
  assign new_new_n2262__ = new_new_n2062__ & ~new_new_n2261__;
  assign new_new_n2263__ = ~new_new_n2066__ & ~new_new_n2262__;
  assign new_new_n2264__ = pi14 & ~new_new_n2263__;
  assign new_new_n2265__ = ~pi14 & new_new_n2064__;
  assign new_new_n2266__ = new_new_n2065__ & new_new_n2265__;
  assign new_new_n2267__ = ~new_new_n2264__ & ~new_new_n2266__;
  assign new_new_n2268__ = new_new_n2260__ & new_new_n2267__;
  assign new_new_n2269__ = ~new_new_n2260__ & ~new_new_n2267__;
  assign new_new_n2270__ = ~new_new_n2268__ & ~new_new_n2269__;
  assign new_new_n2271__ = pi08 & pi20;
  assign new_new_n2272__ = pi04 & pi24;
  assign new_new_n2273__ = pi03 & pi25;
  assign new_new_n2274__ = ~new_new_n2272__ & ~new_new_n2273__;
  assign new_new_n2275__ = new_new_n2272__ & new_new_n2273__;
  assign new_new_n2276__ = ~new_new_n2274__ & ~new_new_n2275__;
  assign new_new_n2277__ = new_new_n2271__ & ~new_new_n2276__;
  assign new_new_n2278__ = ~new_new_n2271__ & new_new_n2276__;
  assign new_new_n2279__ = ~new_new_n2277__ & ~new_new_n2278__;
  assign new_new_n2280__ = new_new_n2270__ & ~new_new_n2279__;
  assign new_new_n2281__ = ~new_new_n2270__ & new_new_n2279__;
  assign new_new_n2282__ = ~new_new_n2280__ & ~new_new_n2281__;
  assign new_new_n2283__ = ~new_new_n2251__ & ~new_new_n2282__;
  assign new_new_n2284__ = new_new_n2251__ & new_new_n2282__;
  assign new_new_n2285__ = ~new_new_n2073__ & ~new_new_n2083__;
  assign new_new_n2286__ = ~new_new_n2072__ & ~new_new_n2285__;
  assign new_new_n2287__ = ~new_new_n2136__ & ~new_new_n2139__;
  assign new_new_n2288__ = ~new_new_n2135__ & ~new_new_n2287__;
  assign new_new_n2289__ = new_new_n2286__ & ~new_new_n2288__;
  assign new_new_n2290__ = ~new_new_n2286__ & new_new_n2288__;
  assign new_new_n2291__ = ~new_new_n2289__ & ~new_new_n2290__;
  assign new_new_n2292__ = ~pi01 & pi27;
  assign new_new_n2293__ = pi14 & new_new_n2065__;
  assign new_new_n2294__ = ~new_new_n2292__ & ~new_new_n2293__;
  assign new_new_n2295__ = pi13 & pi15;
  assign new_new_n2296__ = pi27 & ~new_new_n2295__;
  assign new_new_n2297__ = ~pi27 & new_new_n2295__;
  assign new_new_n2298__ = ~new_new_n2296__ & ~new_new_n2297__;
  assign new_new_n2299__ = ~new_new_n2052__ & ~new_new_n2056__;
  assign new_new_n2300__ = ~new_new_n2055__ & ~new_new_n2299__;
  assign new_new_n2301__ = new_new_n2298__ & ~new_new_n2300__;
  assign new_new_n2302__ = ~new_new_n2298__ & new_new_n2300__;
  assign new_new_n2303__ = ~new_new_n2301__ & ~new_new_n2302__;
  assign new_new_n2304__ = new_new_n2294__ & new_new_n2303__;
  assign new_new_n2305__ = ~new_new_n2294__ & ~new_new_n2303__;
  assign new_new_n2306__ = ~new_new_n2304__ & ~new_new_n2305__;
  assign new_new_n2307__ = new_new_n2291__ & new_new_n2306__;
  assign new_new_n2308__ = ~new_new_n2291__ & ~new_new_n2306__;
  assign new_new_n2309__ = ~new_new_n2307__ & ~new_new_n2308__;
  assign new_new_n2310__ = ~new_new_n2283__ & ~new_new_n2309__;
  assign new_new_n2311__ = ~new_new_n2284__ & ~new_new_n2310__;
  assign new_new_n2312__ = ~new_new_n2283__ & new_new_n2311__;
  assign new_new_n2313__ = ~new_new_n2284__ & new_new_n2310__;
  assign new_new_n2314__ = ~new_new_n2309__ & ~new_new_n2313__;
  assign new_new_n2315__ = ~new_new_n2312__ & ~new_new_n2314__;
  assign new_new_n2316__ = new_new_n2249__ & ~new_new_n2315__;
  assign new_new_n2317__ = ~new_new_n2249__ & new_new_n2315__;
  assign po029 = ~new_new_n2316__ & ~new_new_n2317__;
  assign new_new_n2319__ = ~new_new_n2198__ & ~new_new_n2212__;
  assign new_new_n2320__ = ~new_new_n2199__ & ~new_new_n2319__;
  assign new_new_n2321__ = ~new_new_n2290__ & new_new_n2306__;
  assign new_new_n2322__ = ~new_new_n2289__ & ~new_new_n2321__;
  assign new_new_n2323__ = new_new_n2320__ & ~new_new_n2322__;
  assign new_new_n2324__ = ~new_new_n2320__ & new_new_n2322__;
  assign new_new_n2325__ = ~new_new_n2323__ & ~new_new_n2324__;
  assign new_new_n2326__ = ~new_new_n2191__ & new_new_n2194__;
  assign new_new_n2327__ = ~new_new_n2190__ & ~new_new_n2326__;
  assign new_new_n2328__ = ~new_new_n2268__ & ~new_new_n2279__;
  assign new_new_n2329__ = ~new_new_n2269__ & ~new_new_n2328__;
  assign new_new_n2330__ = ~new_new_n1123__ & ~new_new_n2176__;
  assign new_new_n2331__ = ~new_new_n2175__ & ~new_new_n2330__;
  assign new_new_n2332__ = ~new_new_n2181__ & ~new_new_n2185__;
  assign new_new_n2333__ = ~new_new_n2184__ & ~new_new_n2332__;
  assign new_new_n2334__ = pi00 & pi29;
  assign new_new_n2335__ = pi15 & new_new_n737__;
  assign new_new_n2336__ = ~pi02 & ~new_new_n2335__;
  assign new_new_n2337__ = pi27 & ~new_new_n2336__;
  assign new_new_n2338__ = new_new_n737__ & new_new_n988__;
  assign new_new_n2339__ = new_new_n2337__ & ~new_new_n2338__;
  assign new_new_n2340__ = new_new_n2334__ & ~new_new_n2339__;
  assign new_new_n2341__ = ~new_new_n2334__ & new_new_n2339__;
  assign new_new_n2342__ = ~new_new_n2340__ & ~new_new_n2341__;
  assign new_new_n2343__ = ~new_new_n2333__ & new_new_n2342__;
  assign new_new_n2344__ = new_new_n2333__ & ~new_new_n2342__;
  assign new_new_n2345__ = ~new_new_n2343__ & ~new_new_n2344__;
  assign new_new_n2346__ = ~new_new_n2331__ & ~new_new_n2345__;
  assign new_new_n2347__ = new_new_n2331__ & new_new_n2345__;
  assign new_new_n2348__ = ~new_new_n2346__ & ~new_new_n2347__;
  assign new_new_n2349__ = new_new_n2329__ & ~new_new_n2348__;
  assign new_new_n2350__ = ~new_new_n2329__ & new_new_n2348__;
  assign new_new_n2351__ = ~new_new_n2349__ & ~new_new_n2350__;
  assign new_new_n2352__ = new_new_n2327__ & ~new_new_n2351__;
  assign new_new_n2353__ = ~new_new_n2327__ & new_new_n2351__;
  assign new_new_n2354__ = ~new_new_n2352__ & ~new_new_n2353__;
  assign new_new_n2355__ = new_new_n2325__ & ~new_new_n2354__;
  assign new_new_n2356__ = ~new_new_n2325__ & new_new_n2354__;
  assign new_new_n2357__ = ~new_new_n2355__ & ~new_new_n2356__;
  assign new_new_n2358__ = ~new_new_n2247__ & ~new_new_n2315__;
  assign new_new_n2359__ = ~new_new_n2248__ & ~new_new_n2358__;
  assign new_new_n2360__ = ~new_new_n2357__ & ~new_new_n2359__;
  assign new_new_n2361__ = new_new_n2357__ & new_new_n2359__;
  assign new_new_n2362__ = ~new_new_n2360__ & ~new_new_n2361__;
  assign new_new_n2363__ = ~new_new_n2271__ & ~new_new_n2275__;
  assign new_new_n2364__ = ~new_new_n2274__ & ~new_new_n2363__;
  assign new_new_n2365__ = ~new_new_n2252__ & ~new_new_n2256__;
  assign new_new_n2366__ = ~new_new_n2255__ & ~new_new_n2365__;
  assign new_new_n2367__ = new_new_n2364__ & new_new_n2366__;
  assign new_new_n2368__ = ~new_new_n2364__ & ~new_new_n2366__;
  assign new_new_n2369__ = ~new_new_n2367__ & ~new_new_n2368__;
  assign new_new_n2370__ = pi01 & pi28;
  assign new_new_n2371__ = ~pi15 & ~new_new_n2370__;
  assign new_new_n2372__ = pi15 & new_new_n2370__;
  assign new_new_n2373__ = ~new_new_n2371__ & ~new_new_n2372__;
  assign new_new_n2374__ = new_new_n2369__ & ~new_new_n2373__;
  assign new_new_n2375__ = ~new_new_n2369__ & new_new_n2373__;
  assign new_new_n2376__ = ~new_new_n2374__ & ~new_new_n2375__;
  assign new_new_n2377__ = ~new_new_n2202__ & ~new_new_n2208__;
  assign new_new_n2378__ = ~new_new_n2207__ & ~new_new_n2377__;
  assign new_new_n2379__ = pi14 & pi26;
  assign new_new_n2380__ = ~new_new_n2301__ & new_new_n2379__;
  assign new_new_n2381__ = new_new_n2296__ & new_new_n2300__;
  assign new_new_n2382__ = ~new_new_n2380__ & ~new_new_n2381__;
  assign new_new_n2383__ = pi01 & ~new_new_n2382__;
  assign new_new_n2384__ = pi01 & pi27;
  assign new_new_n2385__ = new_new_n2295__ & ~new_new_n2384__;
  assign new_new_n2386__ = new_new_n2300__ & new_new_n2385__;
  assign new_new_n2387__ = ~new_new_n2383__ & ~new_new_n2386__;
  assign new_new_n2388__ = ~new_new_n2378__ & new_new_n2387__;
  assign new_new_n2389__ = new_new_n2378__ & ~new_new_n2387__;
  assign new_new_n2390__ = ~new_new_n2388__ & ~new_new_n2389__;
  assign new_new_n2391__ = pi14 & pi15;
  assign new_new_n2392__ = pi06 & pi23;
  assign new_new_n2393__ = pi13 & pi16;
  assign new_new_n2394__ = new_new_n2392__ & ~new_new_n2393__;
  assign new_new_n2395__ = ~new_new_n2392__ & new_new_n2393__;
  assign new_new_n2396__ = ~new_new_n2394__ & ~new_new_n2395__;
  assign new_new_n2397__ = new_new_n2391__ & new_new_n2396__;
  assign new_new_n2398__ = ~new_new_n2391__ & ~new_new_n2396__;
  assign new_new_n2399__ = ~new_new_n2397__ & ~new_new_n2398__;
  assign new_new_n2400__ = ~new_new_n2390__ & new_new_n2399__;
  assign new_new_n2401__ = new_new_n2390__ & ~new_new_n2399__;
  assign new_new_n2402__ = ~new_new_n2400__ & ~new_new_n2401__;
  assign new_new_n2403__ = ~new_new_n2376__ & new_new_n2402__;
  assign new_new_n2404__ = new_new_n2376__ & ~new_new_n2402__;
  assign new_new_n2405__ = ~new_new_n2403__ & ~new_new_n2404__;
  assign new_new_n2406__ = pi07 & pi22;
  assign new_new_n2407__ = pi04 & pi25;
  assign new_new_n2408__ = pi05 & pi24;
  assign new_new_n2409__ = ~new_new_n2407__ & ~new_new_n2408__;
  assign new_new_n2410__ = new_new_n2407__ & new_new_n2408__;
  assign new_new_n2411__ = ~new_new_n2409__ & ~new_new_n2410__;
  assign new_new_n2412__ = new_new_n2406__ & ~new_new_n2411__;
  assign new_new_n2413__ = ~new_new_n2406__ & new_new_n2411__;
  assign new_new_n2414__ = ~new_new_n2412__ & ~new_new_n2413__;
  assign new_new_n2415__ = pi11 & pi18;
  assign new_new_n2416__ = pi10 & pi19;
  assign new_new_n2417__ = pi09 & pi20;
  assign new_new_n2418__ = ~new_new_n2416__ & ~new_new_n2417__;
  assign new_new_n2419__ = new_new_n2416__ & new_new_n2417__;
  assign new_new_n2420__ = ~new_new_n2418__ & ~new_new_n2419__;
  assign new_new_n2421__ = new_new_n2415__ & ~new_new_n2420__;
  assign new_new_n2422__ = ~new_new_n2415__ & new_new_n2420__;
  assign new_new_n2423__ = ~new_new_n2421__ & ~new_new_n2422__;
  assign new_new_n2424__ = new_new_n2414__ & new_new_n2423__;
  assign new_new_n2425__ = ~new_new_n2414__ & ~new_new_n2423__;
  assign new_new_n2426__ = ~new_new_n2424__ & ~new_new_n2425__;
  assign new_new_n2427__ = pi12 & pi17;
  assign new_new_n2428__ = pi08 & pi21;
  assign new_new_n2429__ = pi03 & pi26;
  assign new_new_n2430__ = ~new_new_n2428__ & ~new_new_n2429__;
  assign new_new_n2431__ = new_new_n2428__ & new_new_n2429__;
  assign new_new_n2432__ = ~new_new_n2430__ & ~new_new_n2431__;
  assign new_new_n2433__ = new_new_n2427__ & ~new_new_n2432__;
  assign new_new_n2434__ = ~new_new_n2427__ & new_new_n2432__;
  assign new_new_n2435__ = ~new_new_n2433__ & ~new_new_n2434__;
  assign new_new_n2436__ = new_new_n2426__ & ~new_new_n2435__;
  assign new_new_n2437__ = ~new_new_n2426__ & new_new_n2435__;
  assign new_new_n2438__ = ~new_new_n2436__ & ~new_new_n2437__;
  assign new_new_n2439__ = new_new_n2405__ & ~new_new_n2438__;
  assign new_new_n2440__ = ~new_new_n2405__ & new_new_n2438__;
  assign new_new_n2441__ = ~new_new_n2439__ & ~new_new_n2440__;
  assign new_new_n2442__ = ~new_new_n2142__ & ~new_new_n2169__;
  assign new_new_n2443__ = ~new_new_n2170__ & new_new_n2215__;
  assign new_new_n2444__ = ~new_new_n2227__ & ~new_new_n2442__;
  assign new_new_n2445__ = ~new_new_n2443__ & new_new_n2444__;
  assign new_new_n2446__ = new_new_n2170__ & ~new_new_n2215__;
  assign new_new_n2447__ = ~new_new_n2169__ & new_new_n2215__;
  assign new_new_n2448__ = ~new_new_n2215__ & ~new_new_n2227__;
  assign new_new_n2449__ = ~new_new_n2142__ & ~new_new_n2448__;
  assign new_new_n2450__ = ~new_new_n2228__ & ~new_new_n2447__;
  assign new_new_n2451__ = ~new_new_n2449__ & new_new_n2450__;
  assign new_new_n2452__ = ~new_new_n2445__ & ~new_new_n2446__;
  assign new_new_n2453__ = ~new_new_n2451__ & new_new_n2452__;
  assign new_new_n2454__ = ~new_new_n2441__ & ~new_new_n2453__;
  assign new_new_n2455__ = new_new_n2441__ & new_new_n2453__;
  assign new_new_n2456__ = ~new_new_n2454__ & ~new_new_n2455__;
  assign new_new_n2457__ = new_new_n2311__ & ~new_new_n2456__;
  assign new_new_n2458__ = ~new_new_n2311__ & new_new_n2456__;
  assign new_new_n2459__ = ~new_new_n2457__ & ~new_new_n2458__;
  assign new_new_n2460__ = new_new_n2362__ & new_new_n2459__;
  assign new_new_n2461__ = ~new_new_n2362__ & ~new_new_n2459__;
  assign po030 = ~new_new_n2460__ & ~new_new_n2461__;
  assign new_new_n2463__ = ~new_new_n2311__ & ~new_new_n2455__;
  assign new_new_n2464__ = ~new_new_n2454__ & ~new_new_n2463__;
  assign new_new_n2465__ = new_new_n2360__ & new_new_n2464__;
  assign new_new_n2466__ = ~new_new_n2311__ & new_new_n2454__;
  assign new_new_n2467__ = new_new_n2311__ & new_new_n2455__;
  assign new_new_n2468__ = ~new_new_n2466__ & ~new_new_n2467__;
  assign new_new_n2469__ = new_new_n2362__ & new_new_n2468__;
  assign new_new_n2470__ = pi00 & pi30;
  assign new_new_n2471__ = pi14 & pi16;
  assign new_new_n2472__ = pi01 & pi29;
  assign new_new_n2473__ = ~new_new_n2471__ & new_new_n2472__;
  assign new_new_n2474__ = new_new_n2471__ & ~new_new_n2472__;
  assign new_new_n2475__ = ~new_new_n2473__ & ~new_new_n2474__;
  assign new_new_n2476__ = new_new_n2372__ & ~new_new_n2475__;
  assign new_new_n2477__ = ~new_new_n2372__ & new_new_n2475__;
  assign new_new_n2478__ = ~new_new_n2476__ & ~new_new_n2477__;
  assign new_new_n2479__ = new_new_n2470__ & new_new_n2478__;
  assign new_new_n2480__ = ~new_new_n2470__ & ~new_new_n2478__;
  assign new_new_n2481__ = ~new_new_n2479__ & ~new_new_n2480__;
  assign new_new_n2482__ = ~new_new_n2368__ & new_new_n2373__;
  assign new_new_n2483__ = ~new_new_n2367__ & ~new_new_n2482__;
  assign new_new_n2484__ = ~new_new_n2481__ & new_new_n2483__;
  assign new_new_n2485__ = new_new_n2331__ & ~new_new_n2343__;
  assign new_new_n2486__ = new_new_n2481__ & ~new_new_n2483__;
  assign new_new_n2487__ = ~new_new_n2344__ & ~new_new_n2486__;
  assign new_new_n2488__ = ~new_new_n2485__ & new_new_n2487__;
  assign new_new_n2489__ = ~new_new_n2484__ & new_new_n2488__;
  assign new_new_n2490__ = new_new_n2333__ & new_new_n2486__;
  assign new_new_n2491__ = new_new_n2331__ & new_new_n2484__;
  assign new_new_n2492__ = ~new_new_n2490__ & ~new_new_n2491__;
  assign new_new_n2493__ = ~new_new_n2348__ & ~new_new_n2492__;
  assign new_new_n2494__ = new_new_n2333__ & new_new_n2484__;
  assign new_new_n2495__ = new_new_n2331__ & new_new_n2486__;
  assign new_new_n2496__ = ~new_new_n2494__ & ~new_new_n2495__;
  assign new_new_n2497__ = ~new_new_n2342__ & ~new_new_n2496__;
  assign new_new_n2498__ = ~new_new_n2489__ & ~new_new_n2497__;
  assign new_new_n2499__ = ~new_new_n2493__ & new_new_n2498__;
  assign new_new_n2500__ = ~new_new_n2424__ & ~new_new_n2435__;
  assign new_new_n2501__ = ~new_new_n2425__ & ~new_new_n2500__;
  assign new_new_n2502__ = ~new_new_n2427__ & ~new_new_n2431__;
  assign new_new_n2503__ = ~new_new_n2430__ & ~new_new_n2502__;
  assign new_new_n2504__ = ~new_new_n2334__ & ~new_new_n2338__;
  assign new_new_n2505__ = new_new_n2337__ & ~new_new_n2504__;
  assign new_new_n2506__ = ~new_new_n2415__ & ~new_new_n2419__;
  assign new_new_n2507__ = ~new_new_n2418__ & ~new_new_n2506__;
  assign new_new_n2508__ = ~new_new_n2505__ & ~new_new_n2507__;
  assign new_new_n2509__ = new_new_n2505__ & new_new_n2507__;
  assign new_new_n2510__ = ~new_new_n2508__ & ~new_new_n2509__;
  assign new_new_n2511__ = ~new_new_n2503__ & new_new_n2510__;
  assign new_new_n2512__ = new_new_n2503__ & ~new_new_n2510__;
  assign new_new_n2513__ = ~new_new_n2511__ & ~new_new_n2512__;
  assign new_new_n2514__ = ~new_new_n2406__ & ~new_new_n2410__;
  assign new_new_n2515__ = ~new_new_n2409__ & ~new_new_n2514__;
  assign new_new_n2516__ = pi13 & pi17;
  assign new_new_n2517__ = pi09 & pi21;
  assign new_new_n2518__ = pi02 & pi28;
  assign new_new_n2519__ = ~new_new_n2517__ & ~new_new_n2518__;
  assign new_new_n2520__ = new_new_n2517__ & new_new_n2518__;
  assign new_new_n2521__ = ~new_new_n2519__ & ~new_new_n2520__;
  assign new_new_n2522__ = new_new_n2516__ & ~new_new_n2521__;
  assign new_new_n2523__ = ~new_new_n2516__ & new_new_n2521__;
  assign new_new_n2524__ = ~new_new_n2522__ & ~new_new_n2523__;
  assign new_new_n2525__ = ~new_new_n2515__ & new_new_n2524__;
  assign new_new_n2526__ = new_new_n2515__ & ~new_new_n2524__;
  assign new_new_n2527__ = ~new_new_n2525__ & ~new_new_n2526__;
  assign new_new_n2528__ = ~new_new_n2392__ & ~new_new_n2393__;
  assign new_new_n2529__ = new_new_n2392__ & new_new_n2393__;
  assign new_new_n2530__ = ~new_new_n2391__ & ~new_new_n2529__;
  assign new_new_n2531__ = ~new_new_n2528__ & ~new_new_n2530__;
  assign new_new_n2532__ = new_new_n2527__ & ~new_new_n2531__;
  assign new_new_n2533__ = ~new_new_n2527__ & new_new_n2531__;
  assign new_new_n2534__ = ~new_new_n2532__ & ~new_new_n2533__;
  assign new_new_n2535__ = ~new_new_n2513__ & ~new_new_n2534__;
  assign new_new_n2536__ = new_new_n2513__ & new_new_n2534__;
  assign new_new_n2537__ = ~new_new_n2535__ & ~new_new_n2536__;
  assign new_new_n2538__ = new_new_n2501__ & ~new_new_n2537__;
  assign new_new_n2539__ = ~new_new_n2501__ & new_new_n2537__;
  assign new_new_n2540__ = ~new_new_n2538__ & ~new_new_n2539__;
  assign new_new_n2541__ = ~new_new_n2499__ & new_new_n2540__;
  assign new_new_n2542__ = new_new_n2499__ & ~new_new_n2540__;
  assign new_new_n2543__ = ~new_new_n2541__ & ~new_new_n2542__;
  assign new_new_n2544__ = ~new_new_n2403__ & ~new_new_n2438__;
  assign new_new_n2545__ = ~new_new_n2404__ & ~new_new_n2544__;
  assign new_new_n2546__ = new_new_n2543__ & ~new_new_n2545__;
  assign new_new_n2547__ = ~new_new_n2543__ & new_new_n2545__;
  assign new_new_n2548__ = ~new_new_n2546__ & ~new_new_n2547__;
  assign new_new_n2549__ = ~new_new_n2323__ & new_new_n2354__;
  assign new_new_n2550__ = ~new_new_n2324__ & ~new_new_n2549__;
  assign new_new_n2551__ = new_new_n2548__ & new_new_n2550__;
  assign new_new_n2552__ = ~new_new_n2548__ & ~new_new_n2550__;
  assign new_new_n2553__ = ~new_new_n2551__ & ~new_new_n2552__;
  assign new_new_n2554__ = ~new_new_n2388__ & ~new_new_n2399__;
  assign new_new_n2555__ = ~new_new_n2389__ & ~new_new_n2554__;
  assign new_new_n2556__ = new_new_n2327__ & ~new_new_n2350__;
  assign new_new_n2557__ = ~new_new_n2349__ & ~new_new_n2556__;
  assign new_new_n2558__ = new_new_n2555__ & ~new_new_n2557__;
  assign new_new_n2559__ = ~new_new_n2555__ & new_new_n2557__;
  assign new_new_n2560__ = ~new_new_n2558__ & ~new_new_n2559__;
  assign new_new_n2561__ = pi07 & pi23;
  assign new_new_n2562__ = pi05 & pi25;
  assign new_new_n2563__ = pi06 & pi24;
  assign new_new_n2564__ = ~new_new_n2562__ & ~new_new_n2563__;
  assign new_new_n2565__ = new_new_n2562__ & new_new_n2563__;
  assign new_new_n2566__ = ~new_new_n2564__ & ~new_new_n2565__;
  assign new_new_n2567__ = new_new_n2561__ & ~new_new_n2566__;
  assign new_new_n2568__ = ~new_new_n2561__ & new_new_n2566__;
  assign new_new_n2569__ = ~new_new_n2567__ & ~new_new_n2568__;
  assign new_new_n2570__ = pi08 & pi22;
  assign new_new_n2571__ = pi04 & pi26;
  assign new_new_n2572__ = pi03 & pi27;
  assign new_new_n2573__ = ~new_new_n2571__ & ~new_new_n2572__;
  assign new_new_n2574__ = new_new_n2571__ & new_new_n2572__;
  assign new_new_n2575__ = ~new_new_n2573__ & ~new_new_n2574__;
  assign new_new_n2576__ = new_new_n2570__ & ~new_new_n2575__;
  assign new_new_n2577__ = ~new_new_n2570__ & new_new_n2575__;
  assign new_new_n2578__ = ~new_new_n2576__ & ~new_new_n2577__;
  assign new_new_n2579__ = new_new_n2569__ & new_new_n2578__;
  assign new_new_n2580__ = ~new_new_n2569__ & ~new_new_n2578__;
  assign new_new_n2581__ = ~new_new_n2579__ & ~new_new_n2580__;
  assign new_new_n2582__ = pi12 & pi18;
  assign new_new_n2583__ = pi11 & pi19;
  assign new_new_n2584__ = pi10 & pi20;
  assign new_new_n2585__ = ~new_new_n2583__ & ~new_new_n2584__;
  assign new_new_n2586__ = new_new_n2583__ & new_new_n2584__;
  assign new_new_n2587__ = ~new_new_n2585__ & ~new_new_n2586__;
  assign new_new_n2588__ = new_new_n2582__ & ~new_new_n2587__;
  assign new_new_n2589__ = ~new_new_n2582__ & new_new_n2587__;
  assign new_new_n2590__ = ~new_new_n2588__ & ~new_new_n2589__;
  assign new_new_n2591__ = ~new_new_n2581__ & new_new_n2590__;
  assign new_new_n2592__ = new_new_n2581__ & ~new_new_n2590__;
  assign new_new_n2593__ = ~new_new_n2591__ & ~new_new_n2592__;
  assign new_new_n2594__ = new_new_n2560__ & new_new_n2593__;
  assign new_new_n2595__ = ~new_new_n2560__ & ~new_new_n2593__;
  assign new_new_n2596__ = ~new_new_n2594__ & ~new_new_n2595__;
  assign new_new_n2597__ = ~new_new_n2553__ & new_new_n2596__;
  assign new_new_n2598__ = new_new_n2553__ & ~new_new_n2596__;
  assign new_new_n2599__ = ~new_new_n2597__ & ~new_new_n2598__;
  assign new_new_n2600__ = new_new_n2361__ & ~new_new_n2464__;
  assign new_new_n2601__ = ~new_new_n2465__ & new_new_n2599__;
  assign new_new_n2602__ = ~new_new_n2600__ & new_new_n2601__;
  assign new_new_n2603__ = ~new_new_n2469__ & new_new_n2602__;
  assign new_new_n2604__ = ~new_new_n2360__ & new_new_n2453__;
  assign new_new_n2605__ = new_new_n2441__ & new_new_n2604__;
  assign new_new_n2606__ = new_new_n2361__ & ~new_new_n2454__;
  assign new_new_n2607__ = new_new_n2311__ & ~new_new_n2606__;
  assign new_new_n2608__ = ~new_new_n2605__ & new_new_n2607__;
  assign new_new_n2609__ = new_new_n2360__ & ~new_new_n2453__;
  assign new_new_n2610__ = ~new_new_n2361__ & ~new_new_n2441__;
  assign new_new_n2611__ = ~new_new_n2604__ & new_new_n2610__;
  assign new_new_n2612__ = ~new_new_n2311__ & ~new_new_n2609__;
  assign new_new_n2613__ = ~new_new_n2611__ & new_new_n2612__;
  assign new_new_n2614__ = ~new_new_n2608__ & ~new_new_n2613__;
  assign new_new_n2615__ = ~new_new_n2441__ & new_new_n2609__;
  assign new_new_n2616__ = new_new_n2361__ & new_new_n2455__;
  assign new_new_n2617__ = ~new_new_n2599__ & ~new_new_n2616__;
  assign new_new_n2618__ = ~new_new_n2615__ & new_new_n2617__;
  assign new_new_n2619__ = ~new_new_n2614__ & new_new_n2618__;
  assign po031 = ~new_new_n2603__ & ~new_new_n2619__;
  assign new_new_n2621__ = ~new_new_n2466__ & new_new_n2599__;
  assign new_new_n2622__ = ~new_new_n2467__ & ~new_new_n2621__;
  assign new_new_n2623__ = ~new_new_n2361__ & new_new_n2622__;
  assign new_new_n2624__ = new_new_n2464__ & new_new_n2599__;
  assign new_new_n2625__ = ~new_new_n2464__ & ~new_new_n2599__;
  assign new_new_n2626__ = ~new_new_n2360__ & ~new_new_n2625__;
  assign new_new_n2627__ = ~new_new_n2624__ & ~new_new_n2626__;
  assign new_new_n2628__ = ~new_new_n2623__ & ~new_new_n2627__;
  assign new_new_n2629__ = ~new_new_n2558__ & new_new_n2593__;
  assign new_new_n2630__ = ~new_new_n2559__ & ~new_new_n2629__;
  assign new_new_n2631__ = ~new_new_n2582__ & ~new_new_n2586__;
  assign new_new_n2632__ = ~new_new_n2585__ & ~new_new_n2631__;
  assign new_new_n2633__ = ~new_new_n2570__ & ~new_new_n2574__;
  assign new_new_n2634__ = ~new_new_n2573__ & ~new_new_n2633__;
  assign new_new_n2635__ = new_new_n2632__ & new_new_n2634__;
  assign new_new_n2636__ = ~new_new_n2632__ & ~new_new_n2634__;
  assign new_new_n2637__ = ~new_new_n2635__ & ~new_new_n2636__;
  assign new_new_n2638__ = ~new_new_n2516__ & ~new_new_n2520__;
  assign new_new_n2639__ = ~new_new_n2519__ & ~new_new_n2638__;
  assign new_new_n2640__ = ~new_new_n2637__ & new_new_n2639__;
  assign new_new_n2641__ = ~new_new_n2635__ & ~new_new_n2639__;
  assign new_new_n2642__ = ~new_new_n2636__ & new_new_n2641__;
  assign new_new_n2643__ = ~new_new_n2640__ & ~new_new_n2642__;
  assign new_new_n2644__ = ~new_new_n2484__ & ~new_new_n2488__;
  assign new_new_n2645__ = ~new_new_n2579__ & ~new_new_n2590__;
  assign new_new_n2646__ = ~new_new_n2580__ & ~new_new_n2645__;
  assign new_new_n2647__ = new_new_n2644__ & ~new_new_n2646__;
  assign new_new_n2648__ = ~new_new_n2644__ & new_new_n2646__;
  assign new_new_n2649__ = ~new_new_n2647__ & ~new_new_n2648__;
  assign new_new_n2650__ = new_new_n2643__ & new_new_n2649__;
  assign new_new_n2651__ = ~new_new_n2643__ & ~new_new_n2649__;
  assign new_new_n2652__ = ~new_new_n2650__ & ~new_new_n2651__;
  assign new_new_n2653__ = ~new_new_n2541__ & ~new_new_n2545__;
  assign new_new_n2654__ = ~new_new_n2542__ & ~new_new_n2653__;
  assign new_new_n2655__ = ~new_new_n2501__ & ~new_new_n2536__;
  assign new_new_n2656__ = ~new_new_n2535__ & ~new_new_n2655__;
  assign new_new_n2657__ = pi10 & pi21;
  assign new_new_n2658__ = pi09 & pi22;
  assign new_new_n2659__ = pi00 & pi31;
  assign new_new_n2660__ = ~new_new_n2658__ & ~new_new_n2659__;
  assign new_new_n2661__ = new_new_n2658__ & new_new_n2659__;
  assign new_new_n2662__ = ~new_new_n2660__ & ~new_new_n2661__;
  assign new_new_n2663__ = new_new_n2657__ & ~new_new_n2662__;
  assign new_new_n2664__ = ~new_new_n2657__ & new_new_n2662__;
  assign new_new_n2665__ = ~new_new_n2663__ & ~new_new_n2664__;
  assign new_new_n2666__ = pi13 & pi18;
  assign new_new_n2667__ = pi12 & pi19;
  assign new_new_n2668__ = ~new_new_n1325__ & ~new_new_n2667__;
  assign new_new_n2669__ = new_new_n1325__ & new_new_n2667__;
  assign new_new_n2670__ = ~new_new_n2668__ & ~new_new_n2669__;
  assign new_new_n2671__ = new_new_n2666__ & ~new_new_n2670__;
  assign new_new_n2672__ = ~new_new_n2666__ & new_new_n2670__;
  assign new_new_n2673__ = ~new_new_n2671__ & ~new_new_n2672__;
  assign new_new_n2674__ = new_new_n2665__ & new_new_n2673__;
  assign new_new_n2675__ = ~new_new_n2665__ & ~new_new_n2673__;
  assign new_new_n2676__ = ~new_new_n2674__ & ~new_new_n2675__;
  assign new_new_n2677__ = ~new_new_n2470__ & ~new_new_n2476__;
  assign new_new_n2678__ = ~new_new_n2477__ & ~new_new_n2677__;
  assign new_new_n2679__ = new_new_n2676__ & ~new_new_n2678__;
  assign new_new_n2680__ = ~new_new_n2676__ & new_new_n2678__;
  assign new_new_n2681__ = ~new_new_n2679__ & ~new_new_n2680__;
  assign new_new_n2682__ = new_new_n2656__ & new_new_n2681__;
  assign new_new_n2683__ = ~new_new_n2656__ & ~new_new_n2681__;
  assign new_new_n2684__ = ~new_new_n2682__ & ~new_new_n2683__;
  assign new_new_n2685__ = pi15 & pi16;
  assign new_new_n2686__ = pi06 & pi25;
  assign new_new_n2687__ = pi14 & pi17;
  assign new_new_n2688__ = ~new_new_n2686__ & ~new_new_n2687__;
  assign new_new_n2689__ = new_new_n2686__ & new_new_n2687__;
  assign new_new_n2690__ = ~new_new_n2688__ & ~new_new_n2689__;
  assign new_new_n2691__ = new_new_n2685__ & ~new_new_n2690__;
  assign new_new_n2692__ = ~new_new_n2685__ & new_new_n2690__;
  assign new_new_n2693__ = ~new_new_n2691__ & ~new_new_n2692__;
  assign new_new_n2694__ = pi04 & pi27;
  assign new_new_n2695__ = pi03 & pi28;
  assign new_new_n2696__ = pi02 & pi29;
  assign new_new_n2697__ = ~new_new_n2695__ & ~new_new_n2696__;
  assign new_new_n2698__ = new_new_n2695__ & new_new_n2696__;
  assign new_new_n2699__ = ~new_new_n2697__ & ~new_new_n2698__;
  assign new_new_n2700__ = new_new_n2694__ & ~new_new_n2699__;
  assign new_new_n2701__ = ~new_new_n2694__ & new_new_n2699__;
  assign new_new_n2702__ = ~new_new_n2700__ & ~new_new_n2701__;
  assign new_new_n2703__ = ~new_new_n2693__ & ~new_new_n2702__;
  assign new_new_n2704__ = new_new_n2693__ & new_new_n2702__;
  assign new_new_n2705__ = ~new_new_n2703__ & ~new_new_n2704__;
  assign new_new_n2706__ = pi08 & pi23;
  assign new_new_n2707__ = pi07 & pi24;
  assign new_new_n2708__ = pi05 & pi26;
  assign new_new_n2709__ = ~new_new_n2707__ & ~new_new_n2708__;
  assign new_new_n2710__ = new_new_n2707__ & new_new_n2708__;
  assign new_new_n2711__ = ~new_new_n2709__ & ~new_new_n2710__;
  assign new_new_n2712__ = new_new_n2706__ & ~new_new_n2711__;
  assign new_new_n2713__ = ~new_new_n2706__ & new_new_n2711__;
  assign new_new_n2714__ = ~new_new_n2712__ & ~new_new_n2713__;
  assign new_new_n2715__ = ~new_new_n2705__ & new_new_n2714__;
  assign new_new_n2716__ = new_new_n2705__ & ~new_new_n2714__;
  assign new_new_n2717__ = ~new_new_n2715__ & ~new_new_n2716__;
  assign new_new_n2718__ = new_new_n2684__ & new_new_n2717__;
  assign new_new_n2719__ = ~new_new_n2684__ & ~new_new_n2717__;
  assign new_new_n2720__ = ~new_new_n2718__ & ~new_new_n2719__;
  assign new_new_n2721__ = new_new_n2654__ & new_new_n2720__;
  assign new_new_n2722__ = ~new_new_n2654__ & ~new_new_n2720__;
  assign new_new_n2723__ = ~new_new_n2721__ & ~new_new_n2722__;
  assign new_new_n2724__ = ~new_new_n2525__ & new_new_n2531__;
  assign new_new_n2725__ = ~new_new_n2526__ & ~new_new_n2724__;
  assign new_new_n2726__ = ~new_new_n2561__ & ~new_new_n2565__;
  assign new_new_n2727__ = ~new_new_n2564__ & ~new_new_n2726__;
  assign new_new_n2728__ = pi16 & pi30;
  assign new_new_n2729__ = ~new_new_n2727__ & ~new_new_n2728__;
  assign new_new_n2730__ = pi14 & pi29;
  assign new_new_n2731__ = pi01 & ~pi30;
  assign new_new_n2732__ = new_new_n2727__ & ~new_new_n2731__;
  assign new_new_n2733__ = ~new_new_n2729__ & new_new_n2730__;
  assign new_new_n2734__ = ~new_new_n2732__ & new_new_n2733__;
  assign new_new_n2735__ = new_new_n2471__ & new_new_n2472__;
  assign new_new_n2736__ = pi01 & pi30;
  assign new_new_n2737__ = ~new_new_n2727__ & new_new_n2736__;
  assign new_new_n2738__ = new_new_n2727__ & ~new_new_n2736__;
  assign new_new_n2739__ = ~new_new_n2737__ & ~new_new_n2738__;
  assign new_new_n2740__ = pi16 & ~new_new_n2739__;
  assign new_new_n2741__ = ~pi16 & new_new_n2739__;
  assign new_new_n2742__ = ~new_new_n2735__ & ~new_new_n2740__;
  assign new_new_n2743__ = ~new_new_n2741__ & new_new_n2742__;
  assign new_new_n2744__ = ~new_new_n2734__ & ~new_new_n2743__;
  assign new_new_n2745__ = ~new_new_n2725__ & ~new_new_n2744__;
  assign new_new_n2746__ = new_new_n2725__ & new_new_n2744__;
  assign new_new_n2747__ = ~new_new_n2745__ & ~new_new_n2746__;
  assign new_new_n2748__ = ~new_new_n2503__ & ~new_new_n2509__;
  assign new_new_n2749__ = ~new_new_n2508__ & ~new_new_n2748__;
  assign new_new_n2750__ = new_new_n2747__ & ~new_new_n2749__;
  assign new_new_n2751__ = ~new_new_n2747__ & new_new_n2749__;
  assign new_new_n2752__ = ~new_new_n2750__ & ~new_new_n2751__;
  assign new_new_n2753__ = new_new_n2723__ & ~new_new_n2752__;
  assign new_new_n2754__ = ~new_new_n2723__ & new_new_n2752__;
  assign new_new_n2755__ = ~new_new_n2753__ & ~new_new_n2754__;
  assign new_new_n2756__ = new_new_n2652__ & ~new_new_n2755__;
  assign new_new_n2757__ = ~new_new_n2652__ & new_new_n2755__;
  assign new_new_n2758__ = ~new_new_n2756__ & ~new_new_n2757__;
  assign new_new_n2759__ = new_new_n2630__ & new_new_n2758__;
  assign new_new_n2760__ = ~new_new_n2630__ & ~new_new_n2758__;
  assign new_new_n2761__ = ~new_new_n2759__ & ~new_new_n2760__;
  assign new_new_n2762__ = new_new_n2628__ & new_new_n2761__;
  assign new_new_n2763__ = ~new_new_n2628__ & ~new_new_n2761__;
  assign new_new_n2764__ = ~new_new_n2762__ & ~new_new_n2763__;
  assign new_new_n2765__ = ~new_new_n2551__ & new_new_n2596__;
  assign new_new_n2766__ = ~new_new_n2552__ & ~new_new_n2765__;
  assign new_new_n2767__ = new_new_n2764__ & ~new_new_n2766__;
  assign new_new_n2768__ = ~new_new_n2764__ & new_new_n2766__;
  assign po032 = ~new_new_n2767__ & ~new_new_n2768__;
  assign new_new_n2770__ = ~new_new_n2762__ & ~new_new_n2766__;
  assign new_new_n2771__ = ~new_new_n2763__ & ~new_new_n2770__;
  assign new_new_n2772__ = new_new_n2630__ & new_new_n2652__;
  assign new_new_n2773__ = ~new_new_n2630__ & ~new_new_n2652__;
  assign new_new_n2774__ = ~new_new_n2772__ & ~new_new_n2773__;
  assign new_new_n2775__ = new_new_n2752__ & ~new_new_n2774__;
  assign new_new_n2776__ = ~new_new_n2752__ & new_new_n2774__;
  assign new_new_n2777__ = ~new_new_n2722__ & ~new_new_n2775__;
  assign new_new_n2778__ = ~new_new_n2776__ & new_new_n2777__;
  assign new_new_n2779__ = ~new_new_n2721__ & ~new_new_n2778__;
  assign new_new_n2780__ = ~new_new_n2771__ & ~new_new_n2779__;
  assign new_new_n2781__ = new_new_n2771__ & new_new_n2779__;
  assign new_new_n2782__ = ~new_new_n2780__ & ~new_new_n2781__;
  assign new_new_n2783__ = ~new_new_n2636__ & ~new_new_n2641__;
  assign new_new_n2784__ = ~new_new_n2704__ & ~new_new_n2714__;
  assign new_new_n2785__ = ~new_new_n2703__ & ~new_new_n2784__;
  assign new_new_n2786__ = ~new_new_n2675__ & ~new_new_n2678__;
  assign new_new_n2787__ = ~new_new_n2674__ & ~new_new_n2786__;
  assign new_new_n2788__ = ~new_new_n2785__ & new_new_n2787__;
  assign new_new_n2789__ = new_new_n2785__ & ~new_new_n2787__;
  assign new_new_n2790__ = ~new_new_n2788__ & ~new_new_n2789__;
  assign new_new_n2791__ = new_new_n2783__ & new_new_n2790__;
  assign new_new_n2792__ = ~new_new_n2783__ & ~new_new_n2790__;
  assign new_new_n2793__ = ~new_new_n2791__ & ~new_new_n2792__;
  assign new_new_n2794__ = ~new_new_n2745__ & ~new_new_n2749__;
  assign new_new_n2795__ = ~new_new_n2746__ & ~new_new_n2794__;
  assign new_new_n2796__ = ~new_new_n2685__ & ~new_new_n2689__;
  assign new_new_n2797__ = ~new_new_n2688__ & ~new_new_n2796__;
  assign new_new_n2798__ = ~new_new_n2706__ & ~new_new_n2710__;
  assign new_new_n2799__ = ~new_new_n2709__ & ~new_new_n2798__;
  assign new_new_n2800__ = ~new_new_n2797__ & ~new_new_n2799__;
  assign new_new_n2801__ = new_new_n2797__ & new_new_n2799__;
  assign new_new_n2802__ = ~new_new_n2800__ & ~new_new_n2801__;
  assign new_new_n2803__ = pi01 & pi31;
  assign new_new_n2804__ = pi15 & pi17;
  assign new_new_n2805__ = new_new_n2803__ & ~new_new_n2804__;
  assign new_new_n2806__ = ~new_new_n2803__ & new_new_n2804__;
  assign new_new_n2807__ = ~new_new_n2805__ & ~new_new_n2806__;
  assign new_new_n2808__ = new_new_n2802__ & new_new_n2807__;
  assign new_new_n2809__ = ~new_new_n2802__ & ~new_new_n2807__;
  assign new_new_n2810__ = ~new_new_n2808__ & ~new_new_n2809__;
  assign new_new_n2811__ = new_new_n2795__ & ~new_new_n2810__;
  assign new_new_n2812__ = ~new_new_n2795__ & new_new_n2810__;
  assign new_new_n2813__ = ~new_new_n2811__ & ~new_new_n2812__;
  assign new_new_n2814__ = ~new_new_n2666__ & ~new_new_n2669__;
  assign new_new_n2815__ = ~new_new_n2668__ & ~new_new_n2814__;
  assign new_new_n2816__ = ~new_new_n2657__ & ~new_new_n2661__;
  assign new_new_n2817__ = ~new_new_n2660__ & ~new_new_n2816__;
  assign new_new_n2818__ = ~new_new_n2694__ & ~new_new_n2698__;
  assign new_new_n2819__ = ~new_new_n2697__ & ~new_new_n2818__;
  assign new_new_n2820__ = ~new_new_n2817__ & ~new_new_n2819__;
  assign new_new_n2821__ = new_new_n2817__ & new_new_n2819__;
  assign new_new_n2822__ = ~new_new_n2820__ & ~new_new_n2821__;
  assign new_new_n2823__ = new_new_n2815__ & ~new_new_n2822__;
  assign new_new_n2824__ = ~new_new_n2815__ & new_new_n2822__;
  assign new_new_n2825__ = ~new_new_n2823__ & ~new_new_n2824__;
  assign new_new_n2826__ = new_new_n2813__ & new_new_n2825__;
  assign new_new_n2827__ = ~new_new_n2813__ & ~new_new_n2825__;
  assign new_new_n2828__ = ~new_new_n2826__ & ~new_new_n2827__;
  assign new_new_n2829__ = new_new_n2793__ & ~new_new_n2828__;
  assign new_new_n2830__ = ~new_new_n2793__ & new_new_n2828__;
  assign new_new_n2831__ = ~new_new_n2829__ & ~new_new_n2830__;
  assign new_new_n2832__ = ~new_new_n2683__ & ~new_new_n2717__;
  assign new_new_n2833__ = ~new_new_n2682__ & ~new_new_n2832__;
  assign new_new_n2834__ = new_new_n2831__ & new_new_n2833__;
  assign new_new_n2835__ = ~new_new_n2831__ & ~new_new_n2833__;
  assign new_new_n2836__ = ~new_new_n2834__ & ~new_new_n2835__;
  assign new_new_n2837__ = ~new_new_n2643__ & ~new_new_n2648__;
  assign new_new_n2838__ = ~new_new_n2647__ & ~new_new_n2837__;
  assign new_new_n2839__ = pi14 & pi18;
  assign new_new_n2840__ = pi03 & pi29;
  assign new_new_n2841__ = pi10 & pi22;
  assign new_new_n2842__ = ~new_new_n2840__ & ~new_new_n2841__;
  assign new_new_n2843__ = new_new_n2840__ & new_new_n2841__;
  assign new_new_n2844__ = ~new_new_n2842__ & ~new_new_n2843__;
  assign new_new_n2845__ = new_new_n2839__ & ~new_new_n2844__;
  assign new_new_n2846__ = ~new_new_n2839__ & new_new_n2844__;
  assign new_new_n2847__ = ~new_new_n2845__ & ~new_new_n2846__;
  assign new_new_n2848__ = pi00 & pi32;
  assign new_new_n2849__ = pi02 & new_new_n940__;
  assign new_new_n2850__ = ~pi02 & ~new_new_n940__;
  assign new_new_n2851__ = pi30 & ~new_new_n2850__;
  assign new_new_n2852__ = ~new_new_n2849__ & new_new_n2851__;
  assign new_new_n2853__ = new_new_n2848__ & ~new_new_n2852__;
  assign new_new_n2854__ = ~new_new_n2848__ & new_new_n2852__;
  assign new_new_n2855__ = ~new_new_n2853__ & ~new_new_n2854__;
  assign new_new_n2856__ = new_new_n2847__ & new_new_n2855__;
  assign new_new_n2857__ = ~new_new_n2847__ & ~new_new_n2855__;
  assign new_new_n2858__ = ~new_new_n2856__ & ~new_new_n2857__;
  assign new_new_n2859__ = pi13 & pi19;
  assign new_new_n2860__ = pi12 & pi20;
  assign new_new_n2861__ = ~new_new_n1456__ & ~new_new_n2860__;
  assign new_new_n2862__ = new_new_n1456__ & new_new_n2860__;
  assign new_new_n2863__ = ~new_new_n2861__ & ~new_new_n2862__;
  assign new_new_n2864__ = new_new_n2859__ & ~new_new_n2863__;
  assign new_new_n2865__ = ~new_new_n2859__ & new_new_n2863__;
  assign new_new_n2866__ = ~new_new_n2864__ & ~new_new_n2865__;
  assign new_new_n2867__ = ~new_new_n2858__ & new_new_n2866__;
  assign new_new_n2868__ = new_new_n2858__ & ~new_new_n2866__;
  assign new_new_n2869__ = ~new_new_n2867__ & ~new_new_n2868__;
  assign new_new_n2870__ = ~new_new_n2838__ & new_new_n2869__;
  assign new_new_n2871__ = new_new_n2838__ & ~new_new_n2869__;
  assign new_new_n2872__ = ~new_new_n2870__ & ~new_new_n2871__;
  assign new_new_n2873__ = pi08 & pi24;
  assign new_new_n2874__ = pi07 & pi25;
  assign new_new_n2875__ = pi06 & pi26;
  assign new_new_n2876__ = ~new_new_n2874__ & ~new_new_n2875__;
  assign new_new_n2877__ = new_new_n2874__ & new_new_n2875__;
  assign new_new_n2878__ = ~new_new_n2876__ & ~new_new_n2877__;
  assign new_new_n2879__ = new_new_n2873__ & ~new_new_n2878__;
  assign new_new_n2880__ = ~new_new_n2873__ & new_new_n2878__;
  assign new_new_n2881__ = ~new_new_n2879__ & ~new_new_n2880__;
  assign new_new_n2882__ = ~new_new_n2727__ & ~new_new_n2731__;
  assign new_new_n2883__ = new_new_n2730__ & ~new_new_n2882__;
  assign new_new_n2884__ = ~new_new_n2738__ & ~new_new_n2883__;
  assign new_new_n2885__ = pi16 & ~new_new_n2884__;
  assign new_new_n2886__ = ~pi16 & new_new_n2736__;
  assign new_new_n2887__ = new_new_n2727__ & new_new_n2886__;
  assign new_new_n2888__ = ~new_new_n2885__ & ~new_new_n2887__;
  assign new_new_n2889__ = ~new_new_n2881__ & ~new_new_n2888__;
  assign new_new_n2890__ = new_new_n2881__ & new_new_n2888__;
  assign new_new_n2891__ = ~new_new_n2889__ & ~new_new_n2890__;
  assign new_new_n2892__ = pi09 & pi23;
  assign new_new_n2893__ = pi05 & pi27;
  assign new_new_n2894__ = pi04 & pi28;
  assign new_new_n2895__ = ~new_new_n2893__ & ~new_new_n2894__;
  assign new_new_n2896__ = new_new_n2893__ & new_new_n2894__;
  assign new_new_n2897__ = ~new_new_n2895__ & ~new_new_n2896__;
  assign new_new_n2898__ = new_new_n2892__ & ~new_new_n2897__;
  assign new_new_n2899__ = ~new_new_n2892__ & new_new_n2897__;
  assign new_new_n2900__ = ~new_new_n2898__ & ~new_new_n2899__;
  assign new_new_n2901__ = new_new_n2891__ & ~new_new_n2900__;
  assign new_new_n2902__ = ~new_new_n2891__ & new_new_n2900__;
  assign new_new_n2903__ = ~new_new_n2901__ & ~new_new_n2902__;
  assign new_new_n2904__ = new_new_n2872__ & ~new_new_n2903__;
  assign new_new_n2905__ = ~new_new_n2872__ & new_new_n2903__;
  assign new_new_n2906__ = ~new_new_n2904__ & ~new_new_n2905__;
  assign new_new_n2907__ = ~new_new_n2836__ & new_new_n2906__;
  assign new_new_n2908__ = new_new_n2836__ & ~new_new_n2906__;
  assign new_new_n2909__ = ~new_new_n2907__ & ~new_new_n2908__;
  assign new_new_n2910__ = ~new_new_n2752__ & ~new_new_n2772__;
  assign new_new_n2911__ = ~new_new_n2773__ & ~new_new_n2910__;
  assign new_new_n2912__ = new_new_n2909__ & ~new_new_n2911__;
  assign new_new_n2913__ = ~new_new_n2909__ & new_new_n2911__;
  assign new_new_n2914__ = ~new_new_n2912__ & ~new_new_n2913__;
  assign new_new_n2915__ = new_new_n2782__ & new_new_n2914__;
  assign new_new_n2916__ = ~new_new_n2782__ & ~new_new_n2914__;
  assign po033 = ~new_new_n2915__ & ~new_new_n2916__;
  assign new_new_n2918__ = ~new_new_n2815__ & ~new_new_n2821__;
  assign new_new_n2919__ = ~new_new_n2820__ & ~new_new_n2918__;
  assign new_new_n2920__ = ~new_new_n2890__ & ~new_new_n2900__;
  assign new_new_n2921__ = ~new_new_n2889__ & ~new_new_n2920__;
  assign new_new_n2922__ = ~new_new_n2856__ & ~new_new_n2866__;
  assign new_new_n2923__ = ~new_new_n2857__ & ~new_new_n2922__;
  assign new_new_n2924__ = new_new_n2921__ & new_new_n2923__;
  assign new_new_n2925__ = ~new_new_n2921__ & ~new_new_n2923__;
  assign new_new_n2926__ = ~new_new_n2924__ & ~new_new_n2925__;
  assign new_new_n2927__ = ~new_new_n2919__ & new_new_n2926__;
  assign new_new_n2928__ = new_new_n2919__ & ~new_new_n2926__;
  assign new_new_n2929__ = ~new_new_n2927__ & ~new_new_n2928__;
  assign new_new_n2930__ = ~new_new_n2870__ & ~new_new_n2903__;
  assign new_new_n2931__ = ~new_new_n2871__ & ~new_new_n2930__;
  assign new_new_n2932__ = pi08 & pi25;
  assign new_new_n2933__ = pi05 & pi28;
  assign new_new_n2934__ = pi06 & pi27;
  assign new_new_n2935__ = ~new_new_n2933__ & ~new_new_n2934__;
  assign new_new_n2936__ = new_new_n2933__ & new_new_n2934__;
  assign new_new_n2937__ = ~new_new_n2935__ & ~new_new_n2936__;
  assign new_new_n2938__ = new_new_n2932__ & ~new_new_n2937__;
  assign new_new_n2939__ = ~new_new_n2932__ & new_new_n2937__;
  assign new_new_n2940__ = ~new_new_n2938__ & ~new_new_n2939__;
  assign new_new_n2941__ = pi16 & pi17;
  assign new_new_n2942__ = pi07 & pi26;
  assign new_new_n2943__ = pi15 & pi18;
  assign new_new_n2944__ = ~new_new_n2942__ & ~new_new_n2943__;
  assign new_new_n2945__ = new_new_n2942__ & new_new_n2943__;
  assign new_new_n2946__ = ~new_new_n2944__ & ~new_new_n2945__;
  assign new_new_n2947__ = new_new_n2941__ & ~new_new_n2946__;
  assign new_new_n2948__ = ~new_new_n2941__ & new_new_n2946__;
  assign new_new_n2949__ = ~new_new_n2947__ & ~new_new_n2948__;
  assign new_new_n2950__ = new_new_n2940__ & new_new_n2949__;
  assign new_new_n2951__ = ~new_new_n2940__ & ~new_new_n2949__;
  assign new_new_n2952__ = ~new_new_n2950__ & ~new_new_n2951__;
  assign new_new_n2953__ = pi09 & pi24;
  assign new_new_n2954__ = pi04 & pi29;
  assign new_new_n2955__ = pi03 & pi30;
  assign new_new_n2956__ = ~new_new_n2954__ & ~new_new_n2955__;
  assign new_new_n2957__ = new_new_n2954__ & new_new_n2955__;
  assign new_new_n2958__ = ~new_new_n2956__ & ~new_new_n2957__;
  assign new_new_n2959__ = new_new_n2953__ & ~new_new_n2958__;
  assign new_new_n2960__ = ~new_new_n2953__ & new_new_n2958__;
  assign new_new_n2961__ = ~new_new_n2959__ & ~new_new_n2960__;
  assign new_new_n2962__ = new_new_n2952__ & ~new_new_n2961__;
  assign new_new_n2963__ = ~new_new_n2952__ & new_new_n2961__;
  assign new_new_n2964__ = ~new_new_n2962__ & ~new_new_n2963__;
  assign new_new_n2965__ = ~new_new_n2848__ & ~new_new_n2849__;
  assign new_new_n2966__ = new_new_n2851__ & ~new_new_n2965__;
  assign new_new_n2967__ = ~new_new_n2859__ & ~new_new_n2862__;
  assign new_new_n2968__ = ~new_new_n2861__ & ~new_new_n2967__;
  assign new_new_n2969__ = ~new_new_n2839__ & ~new_new_n2843__;
  assign new_new_n2970__ = ~new_new_n2842__ & ~new_new_n2969__;
  assign new_new_n2971__ = ~new_new_n2968__ & ~new_new_n2970__;
  assign new_new_n2972__ = new_new_n2968__ & new_new_n2970__;
  assign new_new_n2973__ = ~new_new_n2971__ & ~new_new_n2972__;
  assign new_new_n2974__ = new_new_n2966__ & ~new_new_n2973__;
  assign new_new_n2975__ = ~new_new_n2966__ & new_new_n2973__;
  assign new_new_n2976__ = ~new_new_n2974__ & ~new_new_n2975__;
  assign new_new_n2977__ = ~new_new_n2964__ & new_new_n2976__;
  assign new_new_n2978__ = new_new_n2964__ & ~new_new_n2976__;
  assign new_new_n2979__ = ~new_new_n2977__ & ~new_new_n2978__;
  assign new_new_n2980__ = ~new_new_n2873__ & ~new_new_n2877__;
  assign new_new_n2981__ = ~new_new_n2876__ & ~new_new_n2980__;
  assign new_new_n2982__ = ~new_new_n2892__ & ~new_new_n2896__;
  assign new_new_n2983__ = ~new_new_n2895__ & ~new_new_n2982__;
  assign new_new_n2984__ = pi11 & pi22;
  assign new_new_n2985__ = pi02 & pi31;
  assign new_new_n2986__ = pi00 & pi33;
  assign new_new_n2987__ = ~new_new_n2985__ & ~new_new_n2986__;
  assign new_new_n2988__ = new_new_n2985__ & new_new_n2986__;
  assign new_new_n2989__ = ~new_new_n2987__ & ~new_new_n2988__;
  assign new_new_n2990__ = new_new_n2984__ & ~new_new_n2989__;
  assign new_new_n2991__ = ~new_new_n2984__ & new_new_n2989__;
  assign new_new_n2992__ = ~new_new_n2990__ & ~new_new_n2991__;
  assign new_new_n2993__ = ~new_new_n2983__ & new_new_n2992__;
  assign new_new_n2994__ = new_new_n2983__ & ~new_new_n2992__;
  assign new_new_n2995__ = ~new_new_n2993__ & ~new_new_n2994__;
  assign new_new_n2996__ = new_new_n2981__ & new_new_n2995__;
  assign new_new_n2997__ = ~new_new_n2981__ & ~new_new_n2995__;
  assign new_new_n2998__ = ~new_new_n2996__ & ~new_new_n2997__;
  assign new_new_n2999__ = new_new_n2979__ & new_new_n2998__;
  assign new_new_n3000__ = ~new_new_n2979__ & ~new_new_n2998__;
  assign new_new_n3001__ = ~new_new_n2999__ & ~new_new_n3000__;
  assign new_new_n3002__ = new_new_n2931__ & new_new_n3001__;
  assign new_new_n3003__ = ~new_new_n2931__ & ~new_new_n3001__;
  assign new_new_n3004__ = ~new_new_n3002__ & ~new_new_n3003__;
  assign new_new_n3005__ = new_new_n2929__ & new_new_n3004__;
  assign new_new_n3006__ = ~new_new_n2929__ & ~new_new_n3004__;
  assign new_new_n3007__ = ~new_new_n3005__ & ~new_new_n3006__;
  assign new_new_n3008__ = ~new_new_n2829__ & ~new_new_n2833__;
  assign new_new_n3009__ = ~new_new_n2830__ & ~new_new_n3008__;
  assign new_new_n3010__ = new_new_n3007__ & ~new_new_n3009__;
  assign new_new_n3011__ = ~new_new_n3007__ & new_new_n3009__;
  assign new_new_n3012__ = ~new_new_n3010__ & ~new_new_n3011__;
  assign new_new_n3013__ = ~new_new_n2812__ & ~new_new_n2825__;
  assign new_new_n3014__ = ~new_new_n2811__ & ~new_new_n3013__;
  assign new_new_n3015__ = pi10 & pi23;
  assign new_new_n3016__ = pi15 & pi31;
  assign new_new_n3017__ = ~pi32 & ~new_new_n3016__;
  assign new_new_n3018__ = pi17 & ~new_new_n3016__;
  assign new_new_n3019__ = pi32 & ~new_new_n3018__;
  assign new_new_n3020__ = pi01 & ~new_new_n3017__;
  assign new_new_n3021__ = ~new_new_n3019__ & new_new_n3020__;
  assign new_new_n3022__ = pi17 & ~new_new_n3021__;
  assign new_new_n3023__ = pi01 & new_new_n3019__;
  assign new_new_n3024__ = ~new_new_n3022__ & ~new_new_n3023__;
  assign new_new_n3025__ = new_new_n3015__ & ~new_new_n3024__;
  assign new_new_n3026__ = ~new_new_n3015__ & new_new_n3024__;
  assign new_new_n3027__ = ~new_new_n3025__ & ~new_new_n3026__;
  assign new_new_n3028__ = ~new_new_n2800__ & ~new_new_n2807__;
  assign new_new_n3029__ = ~new_new_n2801__ & ~new_new_n3028__;
  assign new_new_n3030__ = ~new_new_n3027__ & new_new_n3029__;
  assign new_new_n3031__ = new_new_n3027__ & ~new_new_n3029__;
  assign new_new_n3032__ = ~new_new_n3030__ & ~new_new_n3031__;
  assign new_new_n3033__ = pi14 & pi19;
  assign new_new_n3034__ = pi12 & pi21;
  assign new_new_n3035__ = pi13 & pi20;
  assign new_new_n3036__ = ~new_new_n3034__ & ~new_new_n3035__;
  assign new_new_n3037__ = new_new_n3034__ & new_new_n3035__;
  assign new_new_n3038__ = ~new_new_n3036__ & ~new_new_n3037__;
  assign new_new_n3039__ = new_new_n3033__ & ~new_new_n3038__;
  assign new_new_n3040__ = ~new_new_n3033__ & new_new_n3038__;
  assign new_new_n3041__ = ~new_new_n3039__ & ~new_new_n3040__;
  assign new_new_n3042__ = new_new_n3032__ & ~new_new_n3041__;
  assign new_new_n3043__ = ~new_new_n3032__ & new_new_n3041__;
  assign new_new_n3044__ = ~new_new_n3042__ & ~new_new_n3043__;
  assign new_new_n3045__ = ~new_new_n3014__ & new_new_n3044__;
  assign new_new_n3046__ = new_new_n3014__ & ~new_new_n3044__;
  assign new_new_n3047__ = ~new_new_n3045__ & ~new_new_n3046__;
  assign new_new_n3048__ = new_new_n2783__ & ~new_new_n2789__;
  assign new_new_n3049__ = ~new_new_n2788__ & ~new_new_n3048__;
  assign new_new_n3050__ = new_new_n3047__ & new_new_n3049__;
  assign new_new_n3051__ = ~new_new_n3047__ & ~new_new_n3049__;
  assign new_new_n3052__ = ~new_new_n3050__ & ~new_new_n3051__;
  assign new_new_n3053__ = new_new_n3012__ & ~new_new_n3052__;
  assign new_new_n3054__ = ~new_new_n3012__ & new_new_n3052__;
  assign new_new_n3055__ = ~new_new_n3053__ & ~new_new_n3054__;
  assign new_new_n3056__ = ~new_new_n2907__ & ~new_new_n2911__;
  assign new_new_n3057__ = ~new_new_n2908__ & ~new_new_n3056__;
  assign new_new_n3058__ = new_new_n2780__ & new_new_n3057__;
  assign new_new_n3059__ = new_new_n2907__ & new_new_n2911__;
  assign new_new_n3060__ = new_new_n2908__ & ~new_new_n2911__;
  assign new_new_n3061__ = ~new_new_n3059__ & ~new_new_n3060__;
  assign new_new_n3062__ = new_new_n2782__ & new_new_n3061__;
  assign new_new_n3063__ = new_new_n2781__ & ~new_new_n3057__;
  assign new_new_n3064__ = ~new_new_n3058__ & ~new_new_n3063__;
  assign new_new_n3065__ = ~new_new_n3062__ & new_new_n3064__;
  assign new_new_n3066__ = ~new_new_n3055__ & ~new_new_n3065__;
  assign new_new_n3067__ = new_new_n2780__ & new_new_n2908__;
  assign new_new_n3068__ = new_new_n2780__ & ~new_new_n2906__;
  assign new_new_n3069__ = ~new_new_n2780__ & new_new_n2906__;
  assign new_new_n3070__ = ~new_new_n2781__ & new_new_n2836__;
  assign new_new_n3071__ = ~new_new_n3069__ & new_new_n3070__;
  assign new_new_n3072__ = ~new_new_n3068__ & ~new_new_n3071__;
  assign new_new_n3073__ = ~new_new_n2911__ & ~new_new_n3072__;
  assign new_new_n3074__ = new_new_n2781__ & ~new_new_n2908__;
  assign new_new_n3075__ = ~new_new_n2836__ & new_new_n3069__;
  assign new_new_n3076__ = ~new_new_n3074__ & ~new_new_n3075__;
  assign new_new_n3077__ = new_new_n2911__ & ~new_new_n3076__;
  assign new_new_n3078__ = new_new_n2781__ & new_new_n2907__;
  assign new_new_n3079__ = ~new_new_n3067__ & ~new_new_n3078__;
  assign new_new_n3080__ = ~new_new_n3073__ & new_new_n3079__;
  assign new_new_n3081__ = ~new_new_n3077__ & new_new_n3080__;
  assign new_new_n3082__ = new_new_n3055__ & ~new_new_n3081__;
  assign po034 = new_new_n3066__ | new_new_n3082__;
  assign new_new_n3084__ = ~new_new_n3011__ & new_new_n3052__;
  assign new_new_n3085__ = ~new_new_n3010__ & ~new_new_n3084__;
  assign new_new_n3086__ = new_new_n3055__ & ~new_new_n3057__;
  assign new_new_n3087__ = ~new_new_n3055__ & new_new_n3057__;
  assign new_new_n3088__ = new_new_n2780__ & ~new_new_n3087__;
  assign new_new_n3089__ = ~new_new_n3055__ & ~new_new_n3060__;
  assign new_new_n3090__ = ~new_new_n3059__ & ~new_new_n3089__;
  assign new_new_n3091__ = ~new_new_n2781__ & new_new_n3090__;
  assign new_new_n3092__ = ~new_new_n3086__ & ~new_new_n3088__;
  assign new_new_n3093__ = ~new_new_n3091__ & new_new_n3092__;
  assign new_new_n3094__ = ~new_new_n3085__ & new_new_n3093__;
  assign new_new_n3095__ = new_new_n3085__ & ~new_new_n3093__;
  assign new_new_n3096__ = ~new_new_n3094__ & ~new_new_n3095__;
  assign new_new_n3097__ = new_new_n2929__ & ~new_new_n3002__;
  assign new_new_n3098__ = ~new_new_n3003__ & ~new_new_n3097__;
  assign new_new_n3099__ = ~new_new_n2924__ & ~new_new_n2927__;
  assign new_new_n3100__ = ~new_new_n2966__ & ~new_new_n2972__;
  assign new_new_n3101__ = ~new_new_n2971__ & ~new_new_n3100__;
  assign new_new_n3102__ = pi04 & pi30;
  assign new_new_n3103__ = pi03 & pi31;
  assign new_new_n3104__ = pi00 & pi34;
  assign new_new_n3105__ = ~new_new_n3103__ & ~new_new_n3104__;
  assign new_new_n3106__ = new_new_n3103__ & new_new_n3104__;
  assign new_new_n3107__ = ~new_new_n3105__ & ~new_new_n3106__;
  assign new_new_n3108__ = new_new_n3102__ & ~new_new_n3107__;
  assign new_new_n3109__ = ~new_new_n3102__ & new_new_n3107__;
  assign new_new_n3110__ = ~new_new_n3108__ & ~new_new_n3109__;
  assign new_new_n3111__ = ~new_new_n3101__ & new_new_n3110__;
  assign new_new_n3112__ = new_new_n3101__ & ~new_new_n3110__;
  assign new_new_n3113__ = ~new_new_n3111__ & ~new_new_n3112__;
  assign new_new_n3114__ = ~new_new_n2981__ & ~new_new_n2994__;
  assign new_new_n3115__ = ~new_new_n2993__ & ~new_new_n3114__;
  assign new_new_n3116__ = new_new_n3113__ & new_new_n3115__;
  assign new_new_n3117__ = ~new_new_n3113__ & ~new_new_n3115__;
  assign new_new_n3118__ = ~new_new_n3116__ & ~new_new_n3117__;
  assign new_new_n3119__ = ~new_new_n3099__ & ~new_new_n3118__;
  assign new_new_n3120__ = new_new_n3099__ & new_new_n3118__;
  assign new_new_n3121__ = ~new_new_n3119__ & ~new_new_n3120__;
  assign new_new_n3122__ = ~new_new_n2978__ & ~new_new_n2998__;
  assign new_new_n3123__ = ~new_new_n2977__ & ~new_new_n3122__;
  assign new_new_n3124__ = new_new_n3121__ & ~new_new_n3123__;
  assign new_new_n3125__ = ~new_new_n3121__ & new_new_n3123__;
  assign new_new_n3126__ = ~new_new_n3124__ & ~new_new_n3125__;
  assign new_new_n3127__ = new_new_n3098__ & ~new_new_n3126__;
  assign new_new_n3128__ = ~new_new_n3098__ & new_new_n3126__;
  assign new_new_n3129__ = ~new_new_n3127__ & ~new_new_n3128__;
  assign new_new_n3130__ = ~new_new_n3045__ & new_new_n3049__;
  assign new_new_n3131__ = ~new_new_n3046__ & ~new_new_n3130__;
  assign new_new_n3132__ = pi10 & pi24;
  assign new_new_n3133__ = pi09 & pi25;
  assign new_new_n3134__ = pi05 & pi29;
  assign new_new_n3135__ = ~new_new_n3133__ & ~new_new_n3134__;
  assign new_new_n3136__ = new_new_n3133__ & new_new_n3134__;
  assign new_new_n3137__ = ~new_new_n3135__ & ~new_new_n3136__;
  assign new_new_n3138__ = new_new_n3132__ & ~new_new_n3137__;
  assign new_new_n3139__ = ~new_new_n3132__ & new_new_n3137__;
  assign new_new_n3140__ = ~new_new_n3138__ & ~new_new_n3139__;
  assign new_new_n3141__ = pi08 & pi26;
  assign new_new_n3142__ = pi06 & pi28;
  assign new_new_n3143__ = pi07 & pi27;
  assign new_new_n3144__ = ~new_new_n3142__ & ~new_new_n3143__;
  assign new_new_n3145__ = new_new_n3142__ & new_new_n3143__;
  assign new_new_n3146__ = ~new_new_n3144__ & ~new_new_n3145__;
  assign new_new_n3147__ = new_new_n3141__ & ~new_new_n3146__;
  assign new_new_n3148__ = ~new_new_n3141__ & new_new_n3146__;
  assign new_new_n3149__ = ~new_new_n3147__ & ~new_new_n3148__;
  assign new_new_n3150__ = new_new_n3140__ & new_new_n3149__;
  assign new_new_n3151__ = ~new_new_n3140__ & ~new_new_n3149__;
  assign new_new_n3152__ = ~new_new_n3150__ & ~new_new_n3151__;
  assign new_new_n3153__ = pi15 & pi19;
  assign new_new_n3154__ = pi13 & pi21;
  assign new_new_n3155__ = pi14 & pi20;
  assign new_new_n3156__ = ~new_new_n3154__ & ~new_new_n3155__;
  assign new_new_n3157__ = new_new_n3154__ & new_new_n3155__;
  assign new_new_n3158__ = ~new_new_n3156__ & ~new_new_n3157__;
  assign new_new_n3159__ = new_new_n3153__ & ~new_new_n3158__;
  assign new_new_n3160__ = ~new_new_n3153__ & new_new_n3158__;
  assign new_new_n3161__ = ~new_new_n3159__ & ~new_new_n3160__;
  assign new_new_n3162__ = ~new_new_n3152__ & new_new_n3161__;
  assign new_new_n3163__ = new_new_n3152__ & ~new_new_n3161__;
  assign new_new_n3164__ = ~new_new_n3162__ & ~new_new_n3163__;
  assign new_new_n3165__ = pi12 & pi22;
  assign new_new_n3166__ = pi02 & pi32;
  assign new_new_n3167__ = ~new_new_n1835__ & ~new_new_n3166__;
  assign new_new_n3168__ = new_new_n1835__ & new_new_n3166__;
  assign new_new_n3169__ = ~new_new_n3167__ & ~new_new_n3168__;
  assign new_new_n3170__ = new_new_n3165__ & ~new_new_n3169__;
  assign new_new_n3171__ = ~new_new_n3165__ & new_new_n3169__;
  assign new_new_n3172__ = ~new_new_n3170__ & ~new_new_n3171__;
  assign new_new_n3173__ = pi01 & pi32;
  assign new_new_n3174__ = ~new_new_n3016__ & new_new_n3173__;
  assign new_new_n3175__ = new_new_n3015__ & ~new_new_n3174__;
  assign new_new_n3176__ = pi01 & ~pi32;
  assign new_new_n3177__ = new_new_n3016__ & new_new_n3176__;
  assign new_new_n3178__ = ~new_new_n3175__ & ~new_new_n3177__;
  assign new_new_n3179__ = pi17 & ~new_new_n3178__;
  assign new_new_n3180__ = ~pi17 & new_new_n3015__;
  assign new_new_n3181__ = new_new_n3173__ & new_new_n3180__;
  assign new_new_n3182__ = ~new_new_n3179__ & ~new_new_n3181__;
  assign new_new_n3183__ = new_new_n3172__ & new_new_n3182__;
  assign new_new_n3184__ = ~new_new_n3172__ & ~new_new_n3182__;
  assign new_new_n3185__ = ~new_new_n3183__ & ~new_new_n3184__;
  assign new_new_n3186__ = ~new_new_n3033__ & ~new_new_n3037__;
  assign new_new_n3187__ = ~new_new_n3036__ & ~new_new_n3186__;
  assign new_new_n3188__ = new_new_n3185__ & new_new_n3187__;
  assign new_new_n3189__ = ~new_new_n3185__ & ~new_new_n3187__;
  assign new_new_n3190__ = ~new_new_n3188__ & ~new_new_n3189__;
  assign new_new_n3191__ = new_new_n3164__ & new_new_n3190__;
  assign new_new_n3192__ = ~new_new_n3164__ & ~new_new_n3190__;
  assign new_new_n3193__ = ~new_new_n3191__ & ~new_new_n3192__;
  assign new_new_n3194__ = ~new_new_n3030__ & ~new_new_n3041__;
  assign new_new_n3195__ = ~new_new_n3031__ & ~new_new_n3194__;
  assign new_new_n3196__ = ~new_new_n3193__ & new_new_n3195__;
  assign new_new_n3197__ = new_new_n3193__ & ~new_new_n3195__;
  assign new_new_n3198__ = ~new_new_n3196__ & ~new_new_n3197__;
  assign new_new_n3199__ = ~new_new_n2950__ & ~new_new_n2961__;
  assign new_new_n3200__ = ~new_new_n2951__ & ~new_new_n3199__;
  assign new_new_n3201__ = pi16 & pi18;
  assign new_new_n3202__ = ~new_new_n2941__ & ~new_new_n2945__;
  assign new_new_n3203__ = ~new_new_n2944__ & ~new_new_n3202__;
  assign new_new_n3204__ = new_new_n3201__ & new_new_n3203__;
  assign new_new_n3205__ = ~new_new_n3201__ & ~new_new_n3203__;
  assign new_new_n3206__ = ~new_new_n3204__ & ~new_new_n3205__;
  assign new_new_n3207__ = pi17 & pi32;
  assign new_new_n3208__ = ~pi33 & ~new_new_n3207__;
  assign new_new_n3209__ = pi33 & new_new_n3207__;
  assign new_new_n3210__ = pi01 & ~new_new_n3208__;
  assign new_new_n3211__ = ~new_new_n3209__ & new_new_n3210__;
  assign new_new_n3212__ = ~new_new_n3206__ & new_new_n3211__;
  assign new_new_n3213__ = new_new_n3206__ & ~new_new_n3211__;
  assign new_new_n3214__ = ~new_new_n3212__ & ~new_new_n3213__;
  assign new_new_n3215__ = new_new_n3200__ & new_new_n3214__;
  assign new_new_n3216__ = ~new_new_n3200__ & ~new_new_n3214__;
  assign new_new_n3217__ = ~new_new_n3215__ & ~new_new_n3216__;
  assign new_new_n3218__ = ~new_new_n2953__ & ~new_new_n2957__;
  assign new_new_n3219__ = ~new_new_n2956__ & ~new_new_n3218__;
  assign new_new_n3220__ = ~new_new_n2932__ & ~new_new_n2936__;
  assign new_new_n3221__ = ~new_new_n2935__ & ~new_new_n3220__;
  assign new_new_n3222__ = ~new_new_n2984__ & ~new_new_n2988__;
  assign new_new_n3223__ = ~new_new_n2987__ & ~new_new_n3222__;
  assign new_new_n3224__ = ~new_new_n3221__ & ~new_new_n3223__;
  assign new_new_n3225__ = new_new_n3221__ & new_new_n3223__;
  assign new_new_n3226__ = ~new_new_n3224__ & ~new_new_n3225__;
  assign new_new_n3227__ = new_new_n3219__ & ~new_new_n3226__;
  assign new_new_n3228__ = ~new_new_n3219__ & new_new_n3226__;
  assign new_new_n3229__ = ~new_new_n3227__ & ~new_new_n3228__;
  assign new_new_n3230__ = new_new_n3217__ & new_new_n3229__;
  assign new_new_n3231__ = ~new_new_n3217__ & ~new_new_n3229__;
  assign new_new_n3232__ = ~new_new_n3230__ & ~new_new_n3231__;
  assign new_new_n3233__ = ~new_new_n3198__ & new_new_n3232__;
  assign new_new_n3234__ = new_new_n3198__ & ~new_new_n3232__;
  assign new_new_n3235__ = ~new_new_n3233__ & ~new_new_n3234__;
  assign new_new_n3236__ = new_new_n3131__ & new_new_n3235__;
  assign new_new_n3237__ = ~new_new_n3131__ & ~new_new_n3235__;
  assign new_new_n3238__ = ~new_new_n3236__ & ~new_new_n3237__;
  assign new_new_n3239__ = new_new_n3129__ & ~new_new_n3238__;
  assign new_new_n3240__ = ~new_new_n3129__ & new_new_n3238__;
  assign new_new_n3241__ = ~new_new_n3239__ & ~new_new_n3240__;
  assign new_new_n3242__ = new_new_n3096__ & new_new_n3241__;
  assign new_new_n3243__ = ~new_new_n3096__ & ~new_new_n3241__;
  assign po035 = new_new_n3242__ | new_new_n3243__;
  assign new_new_n3245__ = new_new_n3095__ & new_new_n3098__;
  assign new_new_n3246__ = new_new_n3093__ & ~new_new_n3098__;
  assign new_new_n3247__ = ~new_new_n3093__ & new_new_n3098__;
  assign new_new_n3248__ = ~new_new_n3085__ & ~new_new_n3247__;
  assign new_new_n3249__ = ~new_new_n3246__ & ~new_new_n3248__;
  assign new_new_n3250__ = ~new_new_n3126__ & new_new_n3249__;
  assign new_new_n3251__ = new_new_n3238__ & ~new_new_n3245__;
  assign new_new_n3252__ = ~new_new_n3250__ & new_new_n3251__;
  assign new_new_n3253__ = new_new_n3094__ & ~new_new_n3098__;
  assign new_new_n3254__ = new_new_n3126__ & ~new_new_n3249__;
  assign new_new_n3255__ = ~new_new_n3238__ & ~new_new_n3253__;
  assign new_new_n3256__ = ~new_new_n3254__ & new_new_n3255__;
  assign new_new_n3257__ = ~new_new_n3252__ & ~new_new_n3256__;
  assign new_new_n3258__ = new_new_n3085__ & ~new_new_n3126__;
  assign new_new_n3259__ = ~new_new_n3246__ & ~new_new_n3258__;
  assign new_new_n3260__ = ~new_new_n3085__ & new_new_n3126__;
  assign new_new_n3261__ = ~new_new_n3247__ & ~new_new_n3260__;
  assign new_new_n3262__ = ~new_new_n3259__ & ~new_new_n3261__;
  assign new_new_n3263__ = ~new_new_n3112__ & ~new_new_n3115__;
  assign new_new_n3264__ = ~new_new_n3111__ & ~new_new_n3263__;
  assign new_new_n3265__ = pi15 & pi20;
  assign new_new_n3266__ = pi14 & pi21;
  assign new_new_n3267__ = pi13 & pi22;
  assign new_new_n3268__ = ~new_new_n3266__ & ~new_new_n3267__;
  assign new_new_n3269__ = new_new_n3266__ & new_new_n3267__;
  assign new_new_n3270__ = ~new_new_n3268__ & ~new_new_n3269__;
  assign new_new_n3271__ = new_new_n3265__ & ~new_new_n3270__;
  assign new_new_n3272__ = ~new_new_n3265__ & new_new_n3270__;
  assign new_new_n3273__ = ~new_new_n3271__ & ~new_new_n3272__;
  assign new_new_n3274__ = pi00 & pi35;
  assign new_new_n3275__ = pi18 & new_new_n940__;
  assign new_new_n3276__ = ~pi02 & ~new_new_n3275__;
  assign new_new_n3277__ = pi33 & ~new_new_n3276__;
  assign new_new_n3278__ = new_new_n940__ & new_new_n1285__;
  assign new_new_n3279__ = new_new_n3277__ & ~new_new_n3278__;
  assign new_new_n3280__ = new_new_n3274__ & ~new_new_n3279__;
  assign new_new_n3281__ = ~new_new_n3274__ & new_new_n3279__;
  assign new_new_n3282__ = ~new_new_n3280__ & ~new_new_n3281__;
  assign new_new_n3283__ = new_new_n3273__ & new_new_n3282__;
  assign new_new_n3284__ = ~new_new_n3273__ & ~new_new_n3282__;
  assign new_new_n3285__ = ~new_new_n3283__ & ~new_new_n3284__;
  assign new_new_n3286__ = pi12 & pi23;
  assign new_new_n3287__ = pi11 & pi24;
  assign new_new_n3288__ = pi03 & pi32;
  assign new_new_n3289__ = ~new_new_n3287__ & ~new_new_n3288__;
  assign new_new_n3290__ = new_new_n3287__ & new_new_n3288__;
  assign new_new_n3291__ = ~new_new_n3289__ & ~new_new_n3290__;
  assign new_new_n3292__ = new_new_n3286__ & ~new_new_n3291__;
  assign new_new_n3293__ = ~new_new_n3286__ & new_new_n3291__;
  assign new_new_n3294__ = ~new_new_n3292__ & ~new_new_n3293__;
  assign new_new_n3295__ = new_new_n3285__ & ~new_new_n3294__;
  assign new_new_n3296__ = ~new_new_n3285__ & new_new_n3294__;
  assign new_new_n3297__ = ~new_new_n3295__ & ~new_new_n3296__;
  assign new_new_n3298__ = ~new_new_n3264__ & ~new_new_n3297__;
  assign new_new_n3299__ = new_new_n3264__ & new_new_n3297__;
  assign new_new_n3300__ = ~new_new_n3298__ & ~new_new_n3299__;
  assign new_new_n3301__ = pi17 & pi18;
  assign new_new_n3302__ = pi07 & pi28;
  assign new_new_n3303__ = pi16 & pi19;
  assign new_new_n3304__ = ~new_new_n3302__ & ~new_new_n3303__;
  assign new_new_n3305__ = new_new_n3302__ & new_new_n3303__;
  assign new_new_n3306__ = ~new_new_n3304__ & ~new_new_n3305__;
  assign new_new_n3307__ = new_new_n3301__ & ~new_new_n3306__;
  assign new_new_n3308__ = ~new_new_n3301__ & new_new_n3306__;
  assign new_new_n3309__ = ~new_new_n3307__ & ~new_new_n3308__;
  assign new_new_n3310__ = pi10 & pi25;
  assign new_new_n3311__ = pi09 & pi26;
  assign new_new_n3312__ = pi04 & pi31;
  assign new_new_n3313__ = ~new_new_n3311__ & ~new_new_n3312__;
  assign new_new_n3314__ = new_new_n3311__ & new_new_n3312__;
  assign new_new_n3315__ = ~new_new_n3313__ & ~new_new_n3314__;
  assign new_new_n3316__ = new_new_n3310__ & ~new_new_n3315__;
  assign new_new_n3317__ = ~new_new_n3310__ & new_new_n3315__;
  assign new_new_n3318__ = ~new_new_n3316__ & ~new_new_n3317__;
  assign new_new_n3319__ = new_new_n3309__ & new_new_n3318__;
  assign new_new_n3320__ = ~new_new_n3309__ & ~new_new_n3318__;
  assign new_new_n3321__ = ~new_new_n3319__ & ~new_new_n3320__;
  assign new_new_n3322__ = pi08 & pi27;
  assign new_new_n3323__ = pi06 & pi29;
  assign new_new_n3324__ = pi05 & pi30;
  assign new_new_n3325__ = ~new_new_n3323__ & ~new_new_n3324__;
  assign new_new_n3326__ = new_new_n3323__ & new_new_n3324__;
  assign new_new_n3327__ = ~new_new_n3325__ & ~new_new_n3326__;
  assign new_new_n3328__ = new_new_n3322__ & ~new_new_n3327__;
  assign new_new_n3329__ = ~new_new_n3322__ & new_new_n3327__;
  assign new_new_n3330__ = ~new_new_n3328__ & ~new_new_n3329__;
  assign new_new_n3331__ = new_new_n3321__ & ~new_new_n3330__;
  assign new_new_n3332__ = ~new_new_n3321__ & new_new_n3330__;
  assign new_new_n3333__ = ~new_new_n3331__ & ~new_new_n3332__;
  assign new_new_n3334__ = new_new_n3300__ & new_new_n3333__;
  assign new_new_n3335__ = ~new_new_n3300__ & ~new_new_n3333__;
  assign new_new_n3336__ = ~new_new_n3334__ & ~new_new_n3335__;
  assign new_new_n3337__ = ~new_new_n3150__ & ~new_new_n3161__;
  assign new_new_n3338__ = ~new_new_n3151__ & ~new_new_n3337__;
  assign new_new_n3339__ = ~new_new_n3141__ & ~new_new_n3145__;
  assign new_new_n3340__ = ~new_new_n3144__ & ~new_new_n3339__;
  assign new_new_n3341__ = ~new_new_n3132__ & ~new_new_n3136__;
  assign new_new_n3342__ = ~new_new_n3135__ & ~new_new_n3341__;
  assign new_new_n3343__ = ~new_new_n3340__ & ~new_new_n3342__;
  assign new_new_n3344__ = new_new_n3340__ & new_new_n3342__;
  assign new_new_n3345__ = pi18 & pi34;
  assign new_new_n3346__ = pi01 & new_new_n3345__;
  assign new_new_n3347__ = pi01 & pi34;
  assign new_new_n3348__ = ~pi18 & ~new_new_n3347__;
  assign new_new_n3349__ = ~new_new_n3346__ & ~new_new_n3348__;
  assign new_new_n3350__ = ~new_new_n3344__ & ~new_new_n3349__;
  assign new_new_n3351__ = ~new_new_n3343__ & new_new_n3350__;
  assign new_new_n3352__ = ~new_new_n3343__ & ~new_new_n3350__;
  assign new_new_n3353__ = ~new_new_n3344__ & new_new_n3352__;
  assign new_new_n3354__ = pi18 & new_new_n3347__;
  assign new_new_n3355__ = ~new_new_n3348__ & ~new_new_n3354__;
  assign new_new_n3356__ = ~new_new_n3353__ & new_new_n3355__;
  assign new_new_n3357__ = ~new_new_n3351__ & ~new_new_n3356__;
  assign new_new_n3358__ = new_new_n3338__ & new_new_n3357__;
  assign new_new_n3359__ = ~new_new_n3338__ & ~new_new_n3357__;
  assign new_new_n3360__ = ~new_new_n3358__ & ~new_new_n3359__;
  assign new_new_n3361__ = ~new_new_n3102__ & ~new_new_n3106__;
  assign new_new_n3362__ = ~new_new_n3105__ & ~new_new_n3361__;
  assign new_new_n3363__ = ~new_new_n3165__ & ~new_new_n3168__;
  assign new_new_n3364__ = ~new_new_n3167__ & ~new_new_n3363__;
  assign new_new_n3365__ = new_new_n3362__ & new_new_n3364__;
  assign new_new_n3366__ = ~new_new_n3362__ & ~new_new_n3364__;
  assign new_new_n3367__ = ~new_new_n3153__ & ~new_new_n3157__;
  assign new_new_n3368__ = ~new_new_n3156__ & ~new_new_n3367__;
  assign new_new_n3369__ = ~new_new_n3365__ & ~new_new_n3368__;
  assign new_new_n3370__ = ~new_new_n3366__ & ~new_new_n3369__;
  assign new_new_n3371__ = ~new_new_n3365__ & new_new_n3370__;
  assign new_new_n3372__ = ~new_new_n3366__ & new_new_n3369__;
  assign new_new_n3373__ = ~new_new_n3368__ & ~new_new_n3372__;
  assign new_new_n3374__ = ~new_new_n3371__ & ~new_new_n3373__;
  assign new_new_n3375__ = new_new_n3360__ & ~new_new_n3374__;
  assign new_new_n3376__ = ~new_new_n3360__ & new_new_n3374__;
  assign new_new_n3377__ = ~new_new_n3375__ & ~new_new_n3376__;
  assign new_new_n3378__ = ~new_new_n3336__ & new_new_n3377__;
  assign new_new_n3379__ = new_new_n3336__ & ~new_new_n3377__;
  assign new_new_n3380__ = ~new_new_n3378__ & ~new_new_n3379__;
  assign new_new_n3381__ = ~new_new_n3120__ & ~new_new_n3123__;
  assign new_new_n3382__ = ~new_new_n3119__ & ~new_new_n3381__;
  assign new_new_n3383__ = new_new_n3380__ & ~new_new_n3382__;
  assign new_new_n3384__ = ~new_new_n3380__ & new_new_n3382__;
  assign new_new_n3385__ = ~new_new_n3383__ & ~new_new_n3384__;
  assign new_new_n3386__ = new_new_n3131__ & ~new_new_n3233__;
  assign new_new_n3387__ = ~new_new_n3234__ & ~new_new_n3386__;
  assign new_new_n3388__ = new_new_n3385__ & new_new_n3387__;
  assign new_new_n3389__ = ~new_new_n3385__ & ~new_new_n3387__;
  assign new_new_n3390__ = ~new_new_n3388__ & ~new_new_n3389__;
  assign new_new_n3391__ = ~new_new_n3191__ & ~new_new_n3197__;
  assign new_new_n3392__ = ~new_new_n3183__ & new_new_n3187__;
  assign new_new_n3393__ = ~new_new_n3184__ & ~new_new_n3392__;
  assign new_new_n3394__ = ~new_new_n3219__ & ~new_new_n3225__;
  assign new_new_n3395__ = ~new_new_n3224__ & ~new_new_n3394__;
  assign new_new_n3396__ = ~new_new_n3203__ & ~new_new_n3207__;
  assign new_new_n3397__ = pi33 & ~new_new_n3201__;
  assign new_new_n3398__ = ~new_new_n3396__ & new_new_n3397__;
  assign new_new_n3399__ = ~pi33 & new_new_n3201__;
  assign new_new_n3400__ = ~new_new_n3203__ & ~new_new_n3399__;
  assign new_new_n3401__ = new_new_n3207__ & ~new_new_n3400__;
  assign new_new_n3402__ = ~new_new_n3398__ & ~new_new_n3401__;
  assign new_new_n3403__ = pi01 & ~new_new_n3402__;
  assign new_new_n3404__ = pi01 & pi33;
  assign new_new_n3405__ = new_new_n3204__ & ~new_new_n3404__;
  assign new_new_n3406__ = ~new_new_n3403__ & ~new_new_n3405__;
  assign new_new_n3407__ = new_new_n3395__ & ~new_new_n3406__;
  assign new_new_n3408__ = ~new_new_n3395__ & new_new_n3406__;
  assign new_new_n3409__ = ~new_new_n3407__ & ~new_new_n3408__;
  assign new_new_n3410__ = new_new_n3393__ & ~new_new_n3409__;
  assign new_new_n3411__ = ~new_new_n3393__ & new_new_n3409__;
  assign new_new_n3412__ = ~new_new_n3410__ & ~new_new_n3411__;
  assign new_new_n3413__ = new_new_n3391__ & ~new_new_n3412__;
  assign new_new_n3414__ = ~new_new_n3391__ & new_new_n3412__;
  assign new_new_n3415__ = ~new_new_n3413__ & ~new_new_n3414__;
  assign new_new_n3416__ = ~new_new_n3216__ & new_new_n3229__;
  assign new_new_n3417__ = ~new_new_n3215__ & ~new_new_n3416__;
  assign new_new_n3418__ = new_new_n3415__ & ~new_new_n3417__;
  assign new_new_n3419__ = ~new_new_n3415__ & new_new_n3417__;
  assign new_new_n3420__ = ~new_new_n3418__ & ~new_new_n3419__;
  assign new_new_n3421__ = new_new_n3390__ & ~new_new_n3420__;
  assign new_new_n3422__ = ~new_new_n3390__ & new_new_n3420__;
  assign new_new_n3423__ = ~new_new_n3421__ & ~new_new_n3422__;
  assign new_new_n3424__ = ~new_new_n3262__ & new_new_n3423__;
  assign new_new_n3425__ = ~new_new_n3257__ & new_new_n3424__;
  assign new_new_n3426__ = new_new_n3128__ & ~new_new_n3238__;
  assign new_new_n3427__ = new_new_n3127__ & new_new_n3238__;
  assign new_new_n3428__ = ~new_new_n3426__ & ~new_new_n3427__;
  assign new_new_n3429__ = new_new_n3096__ & new_new_n3428__;
  assign new_new_n3430__ = ~new_new_n3128__ & new_new_n3238__;
  assign new_new_n3431__ = ~new_new_n3127__ & ~new_new_n3430__;
  assign new_new_n3432__ = new_new_n3094__ & ~new_new_n3431__;
  assign new_new_n3433__ = new_new_n3095__ & new_new_n3431__;
  assign new_new_n3434__ = ~new_new_n3423__ & ~new_new_n3432__;
  assign new_new_n3435__ = ~new_new_n3433__ & new_new_n3434__;
  assign new_new_n3436__ = ~new_new_n3429__ & new_new_n3435__;
  assign po036 = ~new_new_n3425__ & ~new_new_n3436__;
  assign new_new_n3438__ = ~new_new_n3238__ & ~new_new_n3258__;
  assign new_new_n3439__ = ~new_new_n3260__ & ~new_new_n3438__;
  assign new_new_n3440__ = ~new_new_n3423__ & ~new_new_n3439__;
  assign new_new_n3441__ = new_new_n3247__ & ~new_new_n3440__;
  assign new_new_n3442__ = new_new_n3423__ & new_new_n3439__;
  assign new_new_n3443__ = ~new_new_n3258__ & ~new_new_n3423__;
  assign new_new_n3444__ = ~new_new_n3260__ & new_new_n3423__;
  assign new_new_n3445__ = ~new_new_n3238__ & ~new_new_n3444__;
  assign new_new_n3446__ = ~new_new_n3443__ & ~new_new_n3445__;
  assign new_new_n3447__ = ~new_new_n3246__ & new_new_n3446__;
  assign new_new_n3448__ = ~new_new_n3441__ & ~new_new_n3442__;
  assign new_new_n3449__ = ~new_new_n3447__ & new_new_n3448__;
  assign new_new_n3450__ = ~new_new_n3319__ & ~new_new_n3330__;
  assign new_new_n3451__ = ~new_new_n3320__ & ~new_new_n3450__;
  assign new_new_n3452__ = ~new_new_n3322__ & ~new_new_n3326__;
  assign new_new_n3453__ = ~new_new_n3325__ & ~new_new_n3452__;
  assign new_new_n3454__ = ~new_new_n3310__ & ~new_new_n3314__;
  assign new_new_n3455__ = ~new_new_n3313__ & ~new_new_n3454__;
  assign new_new_n3456__ = ~new_new_n3301__ & ~new_new_n3305__;
  assign new_new_n3457__ = ~new_new_n3304__ & ~new_new_n3456__;
  assign new_new_n3458__ = ~new_new_n3455__ & ~new_new_n3457__;
  assign new_new_n3459__ = new_new_n3455__ & new_new_n3457__;
  assign new_new_n3460__ = ~new_new_n3458__ & ~new_new_n3459__;
  assign new_new_n3461__ = new_new_n3453__ & ~new_new_n3460__;
  assign new_new_n3462__ = ~new_new_n3453__ & new_new_n3460__;
  assign new_new_n3463__ = ~new_new_n3461__ & ~new_new_n3462__;
  assign new_new_n3464__ = ~new_new_n3451__ & ~new_new_n3463__;
  assign new_new_n3465__ = new_new_n3451__ & new_new_n3463__;
  assign new_new_n3466__ = ~new_new_n3464__ & ~new_new_n3465__;
  assign new_new_n3467__ = ~new_new_n3286__ & ~new_new_n3290__;
  assign new_new_n3468__ = ~new_new_n3289__ & ~new_new_n3467__;
  assign new_new_n3469__ = ~new_new_n3274__ & ~new_new_n3278__;
  assign new_new_n3470__ = new_new_n3277__ & ~new_new_n3469__;
  assign new_new_n3471__ = ~new_new_n3265__ & ~new_new_n3269__;
  assign new_new_n3472__ = ~new_new_n3268__ & ~new_new_n3471__;
  assign new_new_n3473__ = new_new_n3470__ & new_new_n3472__;
  assign new_new_n3474__ = ~new_new_n3470__ & ~new_new_n3472__;
  assign new_new_n3475__ = ~new_new_n3473__ & ~new_new_n3474__;
  assign new_new_n3476__ = new_new_n3468__ & ~new_new_n3475__;
  assign new_new_n3477__ = ~new_new_n3468__ & new_new_n3475__;
  assign new_new_n3478__ = ~new_new_n3476__ & ~new_new_n3477__;
  assign new_new_n3479__ = new_new_n3466__ & new_new_n3478__;
  assign new_new_n3480__ = ~new_new_n3466__ & ~new_new_n3478__;
  assign new_new_n3481__ = ~new_new_n3479__ & ~new_new_n3480__;
  assign new_new_n3482__ = new_new_n3393__ & ~new_new_n3407__;
  assign new_new_n3483__ = ~new_new_n3408__ & ~new_new_n3482__;
  assign new_new_n3484__ = pi10 & pi26;
  assign new_new_n3485__ = pi09 & pi27;
  assign new_new_n3486__ = pi05 & pi31;
  assign new_new_n3487__ = ~new_new_n3485__ & ~new_new_n3486__;
  assign new_new_n3488__ = new_new_n3485__ & new_new_n3486__;
  assign new_new_n3489__ = ~new_new_n3487__ & ~new_new_n3488__;
  assign new_new_n3490__ = new_new_n3484__ & ~new_new_n3489__;
  assign new_new_n3491__ = ~new_new_n3484__ & new_new_n3489__;
  assign new_new_n3492__ = ~new_new_n3490__ & ~new_new_n3491__;
  assign new_new_n3493__ = pi13 & pi23;
  assign new_new_n3494__ = pi12 & pi24;
  assign new_new_n3495__ = pi02 & pi34;
  assign new_new_n3496__ = ~new_new_n3494__ & ~new_new_n3495__;
  assign new_new_n3497__ = new_new_n3494__ & new_new_n3495__;
  assign new_new_n3498__ = ~new_new_n3496__ & ~new_new_n3497__;
  assign new_new_n3499__ = new_new_n3493__ & ~new_new_n3498__;
  assign new_new_n3500__ = ~new_new_n3493__ & new_new_n3498__;
  assign new_new_n3501__ = ~new_new_n3499__ & ~new_new_n3500__;
  assign new_new_n3502__ = new_new_n3492__ & new_new_n3501__;
  assign new_new_n3503__ = ~new_new_n3492__ & ~new_new_n3501__;
  assign new_new_n3504__ = ~new_new_n3502__ & ~new_new_n3503__;
  assign new_new_n3505__ = pi08 & pi28;
  assign new_new_n3506__ = pi06 & pi30;
  assign new_new_n3507__ = pi07 & pi29;
  assign new_new_n3508__ = ~new_new_n3506__ & ~new_new_n3507__;
  assign new_new_n3509__ = new_new_n3506__ & new_new_n3507__;
  assign new_new_n3510__ = ~new_new_n3508__ & ~new_new_n3509__;
  assign new_new_n3511__ = new_new_n3505__ & ~new_new_n3510__;
  assign new_new_n3512__ = ~new_new_n3505__ & new_new_n3510__;
  assign new_new_n3513__ = ~new_new_n3511__ & ~new_new_n3512__;
  assign new_new_n3514__ = ~new_new_n3504__ & new_new_n3513__;
  assign new_new_n3515__ = new_new_n3504__ & ~new_new_n3513__;
  assign new_new_n3516__ = ~new_new_n3514__ & ~new_new_n3515__;
  assign new_new_n3517__ = new_new_n3483__ & new_new_n3516__;
  assign new_new_n3518__ = ~new_new_n3483__ & ~new_new_n3516__;
  assign new_new_n3519__ = ~new_new_n3517__ & ~new_new_n3518__;
  assign new_new_n3520__ = pi16 & pi20;
  assign new_new_n3521__ = pi14 & pi22;
  assign new_new_n3522__ = pi15 & pi21;
  assign new_new_n3523__ = ~new_new_n3521__ & ~new_new_n3522__;
  assign new_new_n3524__ = new_new_n3521__ & new_new_n3522__;
  assign new_new_n3525__ = ~new_new_n3523__ & ~new_new_n3524__;
  assign new_new_n3526__ = new_new_n3520__ & ~new_new_n3525__;
  assign new_new_n3527__ = ~new_new_n3520__ & new_new_n3525__;
  assign new_new_n3528__ = ~new_new_n3526__ & ~new_new_n3527__;
  assign new_new_n3529__ = pi00 & pi36;
  assign new_new_n3530__ = pi17 & pi19;
  assign new_new_n3531__ = pi01 & pi35;
  assign new_new_n3532__ = ~new_new_n3530__ & new_new_n3531__;
  assign new_new_n3533__ = new_new_n3530__ & ~new_new_n3531__;
  assign new_new_n3534__ = ~new_new_n3532__ & ~new_new_n3533__;
  assign new_new_n3535__ = ~new_new_n3529__ & new_new_n3534__;
  assign new_new_n3536__ = new_new_n3529__ & ~new_new_n3534__;
  assign new_new_n3537__ = ~new_new_n3535__ & ~new_new_n3536__;
  assign new_new_n3538__ = ~new_new_n3346__ & ~new_new_n3537__;
  assign new_new_n3539__ = new_new_n3354__ & new_new_n3537__;
  assign new_new_n3540__ = ~new_new_n3538__ & ~new_new_n3539__;
  assign new_new_n3541__ = ~new_new_n3528__ & new_new_n3540__;
  assign new_new_n3542__ = new_new_n3528__ & ~new_new_n3540__;
  assign new_new_n3543__ = ~new_new_n3541__ & ~new_new_n3542__;
  assign new_new_n3544__ = pi11 & pi25;
  assign new_new_n3545__ = pi04 & pi32;
  assign new_new_n3546__ = pi03 & pi33;
  assign new_new_n3547__ = ~new_new_n3545__ & ~new_new_n3546__;
  assign new_new_n3548__ = new_new_n3545__ & new_new_n3546__;
  assign new_new_n3549__ = ~new_new_n3547__ & ~new_new_n3548__;
  assign new_new_n3550__ = new_new_n3544__ & ~new_new_n3549__;
  assign new_new_n3551__ = ~new_new_n3544__ & new_new_n3549__;
  assign new_new_n3552__ = ~new_new_n3550__ & ~new_new_n3551__;
  assign new_new_n3553__ = ~new_new_n3543__ & new_new_n3552__;
  assign new_new_n3554__ = new_new_n3543__ & ~new_new_n3552__;
  assign new_new_n3555__ = ~new_new_n3553__ & ~new_new_n3554__;
  assign new_new_n3556__ = new_new_n3519__ & new_new_n3555__;
  assign new_new_n3557__ = ~new_new_n3519__ & ~new_new_n3555__;
  assign new_new_n3558__ = ~new_new_n3556__ & ~new_new_n3557__;
  assign new_new_n3559__ = new_new_n3481__ & ~new_new_n3558__;
  assign new_new_n3560__ = ~new_new_n3481__ & new_new_n3558__;
  assign new_new_n3561__ = ~new_new_n3559__ & ~new_new_n3560__;
  assign new_new_n3562__ = ~new_new_n3414__ & ~new_new_n3417__;
  assign new_new_n3563__ = ~new_new_n3413__ & ~new_new_n3562__;
  assign new_new_n3564__ = new_new_n3561__ & new_new_n3563__;
  assign new_new_n3565__ = ~new_new_n3561__ & ~new_new_n3563__;
  assign new_new_n3566__ = ~new_new_n3564__ & ~new_new_n3565__;
  assign new_new_n3567__ = ~new_new_n3449__ & new_new_n3566__;
  assign new_new_n3568__ = new_new_n3449__ & ~new_new_n3566__;
  assign new_new_n3569__ = ~new_new_n3567__ & ~new_new_n3568__;
  assign new_new_n3570__ = new_new_n3352__ & new_new_n3370__;
  assign new_new_n3571__ = ~new_new_n3352__ & ~new_new_n3370__;
  assign new_new_n3572__ = ~new_new_n3570__ & ~new_new_n3571__;
  assign new_new_n3573__ = ~new_new_n3283__ & ~new_new_n3294__;
  assign new_new_n3574__ = ~new_new_n3284__ & ~new_new_n3573__;
  assign new_new_n3575__ = ~new_new_n3572__ & new_new_n3574__;
  assign new_new_n3576__ = ~new_new_n3571__ & ~new_new_n3574__;
  assign new_new_n3577__ = ~new_new_n3570__ & new_new_n3576__;
  assign new_new_n3578__ = ~new_new_n3575__ & ~new_new_n3577__;
  assign new_new_n3579__ = ~new_new_n3359__ & ~new_new_n3374__;
  assign new_new_n3580__ = ~new_new_n3358__ & ~new_new_n3579__;
  assign new_new_n3581__ = new_new_n3578__ & new_new_n3580__;
  assign new_new_n3582__ = ~new_new_n3578__ & ~new_new_n3580__;
  assign new_new_n3583__ = ~new_new_n3581__ & ~new_new_n3582__;
  assign new_new_n3584__ = ~new_new_n3299__ & ~new_new_n3333__;
  assign new_new_n3585__ = ~new_new_n3298__ & ~new_new_n3584__;
  assign new_new_n3586__ = new_new_n3583__ & ~new_new_n3585__;
  assign new_new_n3587__ = ~new_new_n3583__ & new_new_n3585__;
  assign new_new_n3588__ = ~new_new_n3586__ & ~new_new_n3587__;
  assign new_new_n3589__ = ~new_new_n3388__ & ~new_new_n3420__;
  assign new_new_n3590__ = ~new_new_n3389__ & ~new_new_n3589__;
  assign new_new_n3591__ = ~new_new_n3588__ & ~new_new_n3590__;
  assign new_new_n3592__ = new_new_n3588__ & new_new_n3590__;
  assign new_new_n3593__ = ~new_new_n3591__ & ~new_new_n3592__;
  assign new_new_n3594__ = ~new_new_n3379__ & ~new_new_n3382__;
  assign new_new_n3595__ = ~new_new_n3378__ & ~new_new_n3594__;
  assign new_new_n3596__ = new_new_n3593__ & ~new_new_n3595__;
  assign new_new_n3597__ = ~new_new_n3593__ & new_new_n3595__;
  assign new_new_n3598__ = ~new_new_n3596__ & ~new_new_n3597__;
  assign new_new_n3599__ = new_new_n3569__ & new_new_n3598__;
  assign new_new_n3600__ = ~new_new_n3569__ & ~new_new_n3598__;
  assign po037 = new_new_n3599__ | new_new_n3600__;
  assign new_new_n3602__ = ~new_new_n3560__ & ~new_new_n3563__;
  assign new_new_n3603__ = ~new_new_n3559__ & ~new_new_n3602__;
  assign new_new_n3604__ = ~new_new_n3581__ & ~new_new_n3585__;
  assign new_new_n3605__ = ~new_new_n3582__ & ~new_new_n3604__;
  assign new_new_n3606__ = ~new_new_n3520__ & ~new_new_n3524__;
  assign new_new_n3607__ = ~new_new_n3523__ & ~new_new_n3606__;
  assign new_new_n3608__ = ~new_new_n3493__ & ~new_new_n3497__;
  assign new_new_n3609__ = ~new_new_n3496__ & ~new_new_n3608__;
  assign new_new_n3610__ = ~new_new_n3607__ & ~new_new_n3609__;
  assign new_new_n3611__ = new_new_n3607__ & new_new_n3609__;
  assign new_new_n3612__ = ~new_new_n3610__ & ~new_new_n3611__;
  assign new_new_n3613__ = ~new_new_n3544__ & ~new_new_n3548__;
  assign new_new_n3614__ = ~new_new_n3547__ & ~new_new_n3613__;
  assign new_new_n3615__ = ~new_new_n3612__ & new_new_n3614__;
  assign new_new_n3616__ = new_new_n3612__ & ~new_new_n3614__;
  assign new_new_n3617__ = ~new_new_n3615__ & ~new_new_n3616__;
  assign new_new_n3618__ = ~new_new_n3541__ & new_new_n3552__;
  assign new_new_n3619__ = ~new_new_n3542__ & ~new_new_n3618__;
  assign new_new_n3620__ = new_new_n3617__ & ~new_new_n3619__;
  assign new_new_n3621__ = ~new_new_n3617__ & new_new_n3619__;
  assign new_new_n3622__ = ~new_new_n3620__ & ~new_new_n3621__;
  assign new_new_n3623__ = ~new_new_n3484__ & ~new_new_n3488__;
  assign new_new_n3624__ = ~new_new_n3487__ & ~new_new_n3623__;
  assign new_new_n3625__ = new_new_n3346__ & ~new_new_n3535__;
  assign new_new_n3626__ = ~new_new_n3536__ & ~new_new_n3625__;
  assign new_new_n3627__ = ~new_new_n3624__ & new_new_n3626__;
  assign new_new_n3628__ = new_new_n3624__ & ~new_new_n3626__;
  assign new_new_n3629__ = ~new_new_n3627__ & ~new_new_n3628__;
  assign new_new_n3630__ = pi15 & pi22;
  assign new_new_n3631__ = pi14 & pi23;
  assign new_new_n3632__ = ~new_new_n1841__ & ~new_new_n3631__;
  assign new_new_n3633__ = new_new_n1841__ & new_new_n3631__;
  assign new_new_n3634__ = ~new_new_n3632__ & ~new_new_n3633__;
  assign new_new_n3635__ = new_new_n3630__ & ~new_new_n3634__;
  assign new_new_n3636__ = ~new_new_n3630__ & new_new_n3634__;
  assign new_new_n3637__ = ~new_new_n3635__ & ~new_new_n3636__;
  assign new_new_n3638__ = ~new_new_n3629__ & new_new_n3637__;
  assign new_new_n3639__ = new_new_n3629__ & ~new_new_n3637__;
  assign new_new_n3640__ = ~new_new_n3638__ & ~new_new_n3639__;
  assign new_new_n3641__ = new_new_n3622__ & new_new_n3640__;
  assign new_new_n3642__ = ~new_new_n3622__ & ~new_new_n3640__;
  assign new_new_n3643__ = ~new_new_n3641__ & ~new_new_n3642__;
  assign new_new_n3644__ = new_new_n3605__ & new_new_n3643__;
  assign new_new_n3645__ = ~new_new_n3605__ & ~new_new_n3643__;
  assign new_new_n3646__ = ~new_new_n3644__ & ~new_new_n3645__;
  assign new_new_n3647__ = ~new_new_n3570__ & ~new_new_n3576__;
  assign new_new_n3648__ = ~new_new_n3468__ & ~new_new_n3473__;
  assign new_new_n3649__ = ~new_new_n3474__ & ~new_new_n3648__;
  assign new_new_n3650__ = pi11 & pi26;
  assign new_new_n3651__ = pi10 & pi27;
  assign new_new_n3652__ = pi05 & pi32;
  assign new_new_n3653__ = ~new_new_n3651__ & ~new_new_n3652__;
  assign new_new_n3654__ = new_new_n3651__ & new_new_n3652__;
  assign new_new_n3655__ = ~new_new_n3653__ & ~new_new_n3654__;
  assign new_new_n3656__ = new_new_n3650__ & ~new_new_n3655__;
  assign new_new_n3657__ = ~new_new_n3650__ & new_new_n3655__;
  assign new_new_n3658__ = ~new_new_n3656__ & ~new_new_n3657__;
  assign new_new_n3659__ = pi18 & pi19;
  assign new_new_n3660__ = pi17 & pi20;
  assign new_new_n3661__ = pi08 & pi29;
  assign new_new_n3662__ = ~new_new_n3660__ & ~new_new_n3661__;
  assign new_new_n3663__ = new_new_n3660__ & new_new_n3661__;
  assign new_new_n3664__ = ~new_new_n3662__ & ~new_new_n3663__;
  assign new_new_n3665__ = new_new_n3659__ & ~new_new_n3664__;
  assign new_new_n3666__ = ~new_new_n3659__ & new_new_n3664__;
  assign new_new_n3667__ = ~new_new_n3665__ & ~new_new_n3666__;
  assign new_new_n3668__ = new_new_n3658__ & new_new_n3667__;
  assign new_new_n3669__ = ~new_new_n3658__ & ~new_new_n3667__;
  assign new_new_n3670__ = ~new_new_n3668__ & ~new_new_n3669__;
  assign new_new_n3671__ = new_new_n3649__ & ~new_new_n3670__;
  assign new_new_n3672__ = ~new_new_n3649__ & new_new_n3670__;
  assign new_new_n3673__ = ~new_new_n3671__ & ~new_new_n3672__;
  assign new_new_n3674__ = ~new_new_n3647__ & ~new_new_n3673__;
  assign new_new_n3675__ = new_new_n3647__ & new_new_n3673__;
  assign new_new_n3676__ = ~new_new_n3674__ & ~new_new_n3675__;
  assign new_new_n3677__ = pi16 & pi21;
  assign new_new_n3678__ = pi03 & pi34;
  assign new_new_n3679__ = pi02 & pi35;
  assign new_new_n3680__ = ~new_new_n3678__ & ~new_new_n3679__;
  assign new_new_n3681__ = new_new_n3678__ & new_new_n3679__;
  assign new_new_n3682__ = ~new_new_n3680__ & ~new_new_n3681__;
  assign new_new_n3683__ = new_new_n3677__ & ~new_new_n3682__;
  assign new_new_n3684__ = ~new_new_n3677__ & new_new_n3682__;
  assign new_new_n3685__ = ~new_new_n3683__ & ~new_new_n3684__;
  assign new_new_n3686__ = pi09 & pi28;
  assign new_new_n3687__ = pi07 & pi30;
  assign new_new_n3688__ = pi06 & pi31;
  assign new_new_n3689__ = ~new_new_n3687__ & ~new_new_n3688__;
  assign new_new_n3690__ = new_new_n3687__ & new_new_n3688__;
  assign new_new_n3691__ = ~new_new_n3689__ & ~new_new_n3690__;
  assign new_new_n3692__ = new_new_n3686__ & ~new_new_n3691__;
  assign new_new_n3693__ = ~new_new_n3686__ & new_new_n3691__;
  assign new_new_n3694__ = ~new_new_n3692__ & ~new_new_n3693__;
  assign new_new_n3695__ = new_new_n3685__ & new_new_n3694__;
  assign new_new_n3696__ = ~new_new_n3685__ & ~new_new_n3694__;
  assign new_new_n3697__ = ~new_new_n3695__ & ~new_new_n3696__;
  assign new_new_n3698__ = pi00 & pi37;
  assign new_new_n3699__ = pi04 & pi33;
  assign new_new_n3700__ = ~new_new_n2061__ & ~new_new_n3699__;
  assign new_new_n3701__ = new_new_n2061__ & new_new_n3699__;
  assign new_new_n3702__ = ~new_new_n3700__ & ~new_new_n3701__;
  assign new_new_n3703__ = new_new_n3698__ & ~new_new_n3702__;
  assign new_new_n3704__ = ~new_new_n3698__ & new_new_n3702__;
  assign new_new_n3705__ = ~new_new_n3703__ & ~new_new_n3704__;
  assign new_new_n3706__ = new_new_n3697__ & ~new_new_n3705__;
  assign new_new_n3707__ = ~new_new_n3697__ & new_new_n3705__;
  assign new_new_n3708__ = ~new_new_n3706__ & ~new_new_n3707__;
  assign new_new_n3709__ = new_new_n3676__ & ~new_new_n3708__;
  assign new_new_n3710__ = ~new_new_n3676__ & new_new_n3708__;
  assign new_new_n3711__ = ~new_new_n3709__ & ~new_new_n3710__;
  assign new_new_n3712__ = new_new_n3646__ & ~new_new_n3711__;
  assign new_new_n3713__ = ~new_new_n3646__ & new_new_n3711__;
  assign new_new_n3714__ = ~new_new_n3712__ & ~new_new_n3713__;
  assign new_new_n3715__ = new_new_n3603__ & new_new_n3714__;
  assign new_new_n3716__ = ~new_new_n3603__ & ~new_new_n3714__;
  assign new_new_n3717__ = ~new_new_n3715__ & ~new_new_n3716__;
  assign new_new_n3718__ = ~new_new_n3517__ & ~new_new_n3555__;
  assign new_new_n3719__ = ~new_new_n3518__ & ~new_new_n3718__;
  assign new_new_n3720__ = ~new_new_n3502__ & ~new_new_n3513__;
  assign new_new_n3721__ = ~new_new_n3503__ & ~new_new_n3720__;
  assign new_new_n3722__ = pi17 & pi35;
  assign new_new_n3723__ = ~new_new_n3505__ & ~new_new_n3509__;
  assign new_new_n3724__ = ~new_new_n3508__ & ~new_new_n3723__;
  assign new_new_n3725__ = pi01 & ~pi36;
  assign new_new_n3726__ = ~new_new_n3724__ & ~new_new_n3725__;
  assign new_new_n3727__ = new_new_n3722__ & ~new_new_n3726__;
  assign new_new_n3728__ = pi19 & pi36;
  assign new_new_n3729__ = new_new_n3724__ & ~new_new_n3728__;
  assign new_new_n3730__ = new_new_n3727__ & ~new_new_n3729__;
  assign new_new_n3731__ = new_new_n3530__ & new_new_n3531__;
  assign new_new_n3732__ = pi01 & pi36;
  assign new_new_n3733__ = new_new_n3724__ & ~new_new_n3732__;
  assign new_new_n3734__ = ~new_new_n3724__ & new_new_n3732__;
  assign new_new_n3735__ = ~new_new_n3733__ & ~new_new_n3734__;
  assign new_new_n3736__ = pi19 & new_new_n3735__;
  assign new_new_n3737__ = ~pi19 & ~new_new_n3735__;
  assign new_new_n3738__ = ~new_new_n3731__ & ~new_new_n3736__;
  assign new_new_n3739__ = ~new_new_n3737__ & new_new_n3738__;
  assign new_new_n3740__ = ~new_new_n3730__ & ~new_new_n3739__;
  assign new_new_n3741__ = new_new_n3721__ & ~new_new_n3740__;
  assign new_new_n3742__ = new_new_n3453__ & ~new_new_n3458__;
  assign new_new_n3743__ = ~new_new_n3721__ & new_new_n3740__;
  assign new_new_n3744__ = ~new_new_n3459__ & ~new_new_n3742__;
  assign new_new_n3745__ = ~new_new_n3743__ & new_new_n3744__;
  assign new_new_n3746__ = ~new_new_n3741__ & new_new_n3745__;
  assign new_new_n3747__ = new_new_n3455__ & new_new_n3743__;
  assign new_new_n3748__ = new_new_n3453__ & new_new_n3741__;
  assign new_new_n3749__ = ~new_new_n3747__ & ~new_new_n3748__;
  assign new_new_n3750__ = new_new_n3457__ & ~new_new_n3749__;
  assign new_new_n3751__ = new_new_n3455__ & new_new_n3741__;
  assign new_new_n3752__ = new_new_n3453__ & new_new_n3743__;
  assign new_new_n3753__ = ~new_new_n3751__ & ~new_new_n3752__;
  assign new_new_n3754__ = new_new_n3463__ & ~new_new_n3753__;
  assign new_new_n3755__ = ~new_new_n3746__ & ~new_new_n3750__;
  assign new_new_n3756__ = ~new_new_n3754__ & new_new_n3755__;
  assign new_new_n3757__ = ~new_new_n3719__ & new_new_n3756__;
  assign new_new_n3758__ = new_new_n3719__ & ~new_new_n3756__;
  assign new_new_n3759__ = ~new_new_n3757__ & ~new_new_n3758__;
  assign new_new_n3760__ = ~new_new_n3465__ & ~new_new_n3478__;
  assign new_new_n3761__ = ~new_new_n3464__ & ~new_new_n3760__;
  assign new_new_n3762__ = new_new_n3759__ & ~new_new_n3761__;
  assign new_new_n3763__ = ~new_new_n3759__ & new_new_n3761__;
  assign new_new_n3764__ = ~new_new_n3762__ & ~new_new_n3763__;
  assign new_new_n3765__ = new_new_n3717__ & ~new_new_n3764__;
  assign new_new_n3766__ = ~new_new_n3717__ & new_new_n3764__;
  assign new_new_n3767__ = ~new_new_n3765__ & ~new_new_n3766__;
  assign new_new_n3768__ = new_new_n3568__ & new_new_n3590__;
  assign new_new_n3769__ = new_new_n3449__ & new_new_n3590__;
  assign new_new_n3770__ = ~new_new_n3449__ & ~new_new_n3590__;
  assign new_new_n3771__ = ~new_new_n3566__ & ~new_new_n3770__;
  assign new_new_n3772__ = ~new_new_n3769__ & ~new_new_n3771__;
  assign new_new_n3773__ = new_new_n3588__ & ~new_new_n3772__;
  assign new_new_n3774__ = ~new_new_n3595__ & ~new_new_n3768__;
  assign new_new_n3775__ = ~new_new_n3773__ & new_new_n3774__;
  assign new_new_n3776__ = new_new_n3567__ & ~new_new_n3590__;
  assign new_new_n3777__ = ~new_new_n3588__ & new_new_n3772__;
  assign new_new_n3778__ = new_new_n3595__ & ~new_new_n3776__;
  assign new_new_n3779__ = ~new_new_n3777__ & new_new_n3778__;
  assign new_new_n3780__ = ~new_new_n3775__ & ~new_new_n3779__;
  assign new_new_n3781__ = ~new_new_n3568__ & ~new_new_n3770__;
  assign new_new_n3782__ = new_new_n3566__ & ~new_new_n3588__;
  assign new_new_n3783__ = ~new_new_n3592__ & ~new_new_n3782__;
  assign new_new_n3784__ = ~new_new_n3781__ & ~new_new_n3783__;
  assign new_new_n3785__ = ~new_new_n3767__ & ~new_new_n3784__;
  assign new_new_n3786__ = ~new_new_n3780__ & new_new_n3785__;
  assign new_new_n3787__ = new_new_n3592__ & ~new_new_n3595__;
  assign new_new_n3788__ = new_new_n3591__ & new_new_n3595__;
  assign new_new_n3789__ = ~new_new_n3787__ & ~new_new_n3788__;
  assign new_new_n3790__ = new_new_n3569__ & new_new_n3789__;
  assign new_new_n3791__ = ~new_new_n3592__ & new_new_n3595__;
  assign new_new_n3792__ = ~new_new_n3591__ & ~new_new_n3791__;
  assign new_new_n3793__ = new_new_n3568__ & ~new_new_n3792__;
  assign new_new_n3794__ = new_new_n3567__ & new_new_n3792__;
  assign new_new_n3795__ = new_new_n3767__ & ~new_new_n3793__;
  assign new_new_n3796__ = ~new_new_n3794__ & new_new_n3795__;
  assign new_new_n3797__ = ~new_new_n3790__ & new_new_n3796__;
  assign po038 = ~new_new_n3786__ & ~new_new_n3797__;
  assign new_new_n3799__ = ~new_new_n3757__ & ~new_new_n3761__;
  assign new_new_n3800__ = ~new_new_n3758__ & ~new_new_n3799__;
  assign new_new_n3801__ = ~new_new_n3695__ & ~new_new_n3705__;
  assign new_new_n3802__ = ~new_new_n3696__ & ~new_new_n3801__;
  assign new_new_n3803__ = pi18 & pi20;
  assign new_new_n3804__ = pi01 & pi37;
  assign new_new_n3805__ = ~new_new_n3803__ & new_new_n3804__;
  assign new_new_n3806__ = new_new_n3803__ & ~new_new_n3804__;
  assign new_new_n3807__ = ~new_new_n3805__ & ~new_new_n3806__;
  assign new_new_n3808__ = ~new_new_n3686__ & ~new_new_n3690__;
  assign new_new_n3809__ = ~new_new_n3689__ & ~new_new_n3808__;
  assign new_new_n3810__ = ~new_new_n3659__ & ~new_new_n3663__;
  assign new_new_n3811__ = ~new_new_n3662__ & ~new_new_n3810__;
  assign new_new_n3812__ = new_new_n3809__ & new_new_n3811__;
  assign new_new_n3813__ = ~new_new_n3809__ & ~new_new_n3811__;
  assign new_new_n3814__ = ~new_new_n3812__ & ~new_new_n3813__;
  assign new_new_n3815__ = new_new_n3807__ & new_new_n3814__;
  assign new_new_n3816__ = ~new_new_n3807__ & ~new_new_n3814__;
  assign new_new_n3817__ = ~new_new_n3815__ & ~new_new_n3816__;
  assign new_new_n3818__ = new_new_n3802__ & new_new_n3817__;
  assign new_new_n3819__ = ~new_new_n3802__ & ~new_new_n3817__;
  assign new_new_n3820__ = ~new_new_n3818__ & ~new_new_n3819__;
  assign new_new_n3821__ = ~new_new_n3628__ & new_new_n3637__;
  assign new_new_n3822__ = ~new_new_n3627__ & ~new_new_n3821__;
  assign new_new_n3823__ = new_new_n3820__ & ~new_new_n3822__;
  assign new_new_n3824__ = ~new_new_n3820__ & new_new_n3822__;
  assign new_new_n3825__ = ~new_new_n3823__ & ~new_new_n3824__;
  assign new_new_n3826__ = ~new_new_n3741__ & ~new_new_n3745__;
  assign new_new_n3827__ = ~new_new_n3611__ & ~new_new_n3614__;
  assign new_new_n3828__ = ~new_new_n3610__ & ~new_new_n3827__;
  assign new_new_n3829__ = pi12 & pi26;
  assign new_new_n3830__ = pi11 & pi27;
  assign new_new_n3831__ = pi04 & pi34;
  assign new_new_n3832__ = ~new_new_n3830__ & ~new_new_n3831__;
  assign new_new_n3833__ = new_new_n3830__ & new_new_n3831__;
  assign new_new_n3834__ = ~new_new_n3832__ & ~new_new_n3833__;
  assign new_new_n3835__ = new_new_n3829__ & ~new_new_n3834__;
  assign new_new_n3836__ = ~new_new_n3829__ & new_new_n3834__;
  assign new_new_n3837__ = ~new_new_n3835__ & ~new_new_n3836__;
  assign new_new_n3838__ = ~new_new_n3727__ & ~new_new_n3733__;
  assign new_new_n3839__ = pi19 & ~new_new_n3838__;
  assign new_new_n3840__ = ~pi19 & new_new_n3732__;
  assign new_new_n3841__ = new_new_n3724__ & new_new_n3840__;
  assign new_new_n3842__ = ~new_new_n3839__ & ~new_new_n3841__;
  assign new_new_n3843__ = ~new_new_n3837__ & ~new_new_n3842__;
  assign new_new_n3844__ = new_new_n3837__ & new_new_n3842__;
  assign new_new_n3845__ = ~new_new_n3843__ & ~new_new_n3844__;
  assign new_new_n3846__ = new_new_n3828__ & new_new_n3845__;
  assign new_new_n3847__ = ~new_new_n3828__ & ~new_new_n3845__;
  assign new_new_n3848__ = ~new_new_n3846__ & ~new_new_n3847__;
  assign new_new_n3849__ = ~new_new_n3826__ & ~new_new_n3848__;
  assign new_new_n3850__ = new_new_n3826__ & new_new_n3848__;
  assign new_new_n3851__ = ~new_new_n3849__ & ~new_new_n3850__;
  assign new_new_n3852__ = pi14 & pi24;
  assign new_new_n3853__ = pi03 & pi35;
  assign new_new_n3854__ = pi13 & pi25;
  assign new_new_n3855__ = ~new_new_n3853__ & ~new_new_n3854__;
  assign new_new_n3856__ = new_new_n3853__ & new_new_n3854__;
  assign new_new_n3857__ = ~new_new_n3855__ & ~new_new_n3856__;
  assign new_new_n3858__ = new_new_n3852__ & ~new_new_n3857__;
  assign new_new_n3859__ = ~new_new_n3852__ & new_new_n3857__;
  assign new_new_n3860__ = ~new_new_n3858__ & ~new_new_n3859__;
  assign new_new_n3861__ = ~new_new_n3650__ & ~new_new_n3654__;
  assign new_new_n3862__ = ~new_new_n3653__ & ~new_new_n3861__;
  assign new_new_n3863__ = pi00 & pi38;
  assign new_new_n3864__ = pi02 & new_new_n1223__;
  assign new_new_n3865__ = ~pi02 & ~new_new_n1223__;
  assign new_new_n3866__ = pi36 & ~new_new_n3865__;
  assign new_new_n3867__ = ~new_new_n3864__ & new_new_n3866__;
  assign new_new_n3868__ = new_new_n3863__ & ~new_new_n3867__;
  assign new_new_n3869__ = ~new_new_n3863__ & new_new_n3867__;
  assign new_new_n3870__ = ~new_new_n3868__ & ~new_new_n3869__;
  assign new_new_n3871__ = new_new_n3862__ & ~new_new_n3870__;
  assign new_new_n3872__ = ~new_new_n3862__ & new_new_n3870__;
  assign new_new_n3873__ = ~new_new_n3871__ & ~new_new_n3872__;
  assign new_new_n3874__ = new_new_n3860__ & new_new_n3873__;
  assign new_new_n3875__ = ~new_new_n3860__ & ~new_new_n3873__;
  assign new_new_n3876__ = ~new_new_n3874__ & ~new_new_n3875__;
  assign new_new_n3877__ = new_new_n3851__ & ~new_new_n3876__;
  assign new_new_n3878__ = ~new_new_n3851__ & new_new_n3876__;
  assign new_new_n3879__ = ~new_new_n3877__ & ~new_new_n3878__;
  assign new_new_n3880__ = new_new_n3825__ & ~new_new_n3879__;
  assign new_new_n3881__ = ~new_new_n3825__ & new_new_n3879__;
  assign new_new_n3882__ = ~new_new_n3880__ & ~new_new_n3881__;
  assign new_new_n3883__ = new_new_n3800__ & new_new_n3882__;
  assign new_new_n3884__ = ~new_new_n3800__ & ~new_new_n3882__;
  assign new_new_n3885__ = ~new_new_n3883__ & ~new_new_n3884__;
  assign new_new_n3886__ = ~new_new_n3621__ & ~new_new_n3640__;
  assign new_new_n3887__ = ~new_new_n3620__ & ~new_new_n3886__;
  assign new_new_n3888__ = new_new_n3649__ & ~new_new_n3668__;
  assign new_new_n3889__ = ~new_new_n3669__ & ~new_new_n3888__;
  assign new_new_n3890__ = pi17 & pi21;
  assign new_new_n3891__ = pi16 & pi22;
  assign new_new_n3892__ = pi15 & pi23;
  assign new_new_n3893__ = ~new_new_n3891__ & ~new_new_n3892__;
  assign new_new_n3894__ = new_new_n3891__ & new_new_n3892__;
  assign new_new_n3895__ = ~new_new_n3893__ & ~new_new_n3894__;
  assign new_new_n3896__ = new_new_n3890__ & ~new_new_n3895__;
  assign new_new_n3897__ = ~new_new_n3890__ & new_new_n3895__;
  assign new_new_n3898__ = ~new_new_n3896__ & ~new_new_n3897__;
  assign new_new_n3899__ = pi10 & pi28;
  assign new_new_n3900__ = pi06 & pi32;
  assign new_new_n3901__ = pi05 & pi33;
  assign new_new_n3902__ = ~new_new_n3900__ & ~new_new_n3901__;
  assign new_new_n3903__ = new_new_n3900__ & new_new_n3901__;
  assign new_new_n3904__ = ~new_new_n3902__ & ~new_new_n3903__;
  assign new_new_n3905__ = new_new_n3899__ & ~new_new_n3904__;
  assign new_new_n3906__ = ~new_new_n3899__ & new_new_n3904__;
  assign new_new_n3907__ = ~new_new_n3905__ & ~new_new_n3906__;
  assign new_new_n3908__ = new_new_n3898__ & new_new_n3907__;
  assign new_new_n3909__ = ~new_new_n3898__ & ~new_new_n3907__;
  assign new_new_n3910__ = ~new_new_n3908__ & ~new_new_n3909__;
  assign new_new_n3911__ = pi09 & pi29;
  assign new_new_n3912__ = pi07 & pi31;
  assign new_new_n3913__ = pi08 & pi30;
  assign new_new_n3914__ = ~new_new_n3912__ & ~new_new_n3913__;
  assign new_new_n3915__ = new_new_n3912__ & new_new_n3913__;
  assign new_new_n3916__ = ~new_new_n3914__ & ~new_new_n3915__;
  assign new_new_n3917__ = new_new_n3911__ & ~new_new_n3916__;
  assign new_new_n3918__ = ~new_new_n3911__ & new_new_n3916__;
  assign new_new_n3919__ = ~new_new_n3917__ & ~new_new_n3918__;
  assign new_new_n3920__ = ~new_new_n3910__ & new_new_n3919__;
  assign new_new_n3921__ = new_new_n3910__ & ~new_new_n3919__;
  assign new_new_n3922__ = ~new_new_n3920__ & ~new_new_n3921__;
  assign new_new_n3923__ = ~new_new_n3889__ & new_new_n3922__;
  assign new_new_n3924__ = new_new_n3889__ & ~new_new_n3922__;
  assign new_new_n3925__ = ~new_new_n3923__ & ~new_new_n3924__;
  assign new_new_n3926__ = ~new_new_n3630__ & ~new_new_n3633__;
  assign new_new_n3927__ = ~new_new_n3632__ & ~new_new_n3926__;
  assign new_new_n3928__ = ~new_new_n3677__ & ~new_new_n3681__;
  assign new_new_n3929__ = ~new_new_n3680__ & ~new_new_n3928__;
  assign new_new_n3930__ = ~new_new_n3927__ & ~new_new_n3929__;
  assign new_new_n3931__ = new_new_n3927__ & new_new_n3929__;
  assign new_new_n3932__ = ~new_new_n3930__ & ~new_new_n3931__;
  assign new_new_n3933__ = ~new_new_n3698__ & ~new_new_n3701__;
  assign new_new_n3934__ = ~new_new_n3700__ & ~new_new_n3933__;
  assign new_new_n3935__ = new_new_n3932__ & ~new_new_n3934__;
  assign new_new_n3936__ = ~new_new_n3932__ & new_new_n3934__;
  assign new_new_n3937__ = ~new_new_n3935__ & ~new_new_n3936__;
  assign new_new_n3938__ = new_new_n3925__ & new_new_n3937__;
  assign new_new_n3939__ = ~new_new_n3925__ & ~new_new_n3937__;
  assign new_new_n3940__ = ~new_new_n3938__ & ~new_new_n3939__;
  assign new_new_n3941__ = ~new_new_n3887__ & new_new_n3940__;
  assign new_new_n3942__ = new_new_n3887__ & ~new_new_n3940__;
  assign new_new_n3943__ = ~new_new_n3941__ & ~new_new_n3942__;
  assign new_new_n3944__ = ~new_new_n3675__ & new_new_n3708__;
  assign new_new_n3945__ = ~new_new_n3674__ & ~new_new_n3944__;
  assign new_new_n3946__ = new_new_n3943__ & new_new_n3945__;
  assign new_new_n3947__ = ~new_new_n3943__ & ~new_new_n3945__;
  assign new_new_n3948__ = ~new_new_n3946__ & ~new_new_n3947__;
  assign new_new_n3949__ = ~new_new_n3885__ & ~new_new_n3948__;
  assign new_new_n3950__ = new_new_n3885__ & new_new_n3948__;
  assign new_new_n3951__ = ~new_new_n3949__ & ~new_new_n3950__;
  assign new_new_n3952__ = ~new_new_n3566__ & new_new_n3588__;
  assign new_new_n3953__ = ~new_new_n3767__ & ~new_new_n3952__;
  assign new_new_n3954__ = new_new_n3767__ & ~new_new_n3782__;
  assign new_new_n3955__ = new_new_n3595__ & ~new_new_n3954__;
  assign new_new_n3956__ = ~new_new_n3769__ & new_new_n3955__;
  assign new_new_n3957__ = ~new_new_n3770__ & ~new_new_n3953__;
  assign new_new_n3958__ = ~new_new_n3956__ & new_new_n3957__;
  assign new_new_n3959__ = new_new_n3767__ & new_new_n3952__;
  assign new_new_n3960__ = ~new_new_n3767__ & ~new_new_n3769__;
  assign new_new_n3961__ = ~new_new_n3595__ & ~new_new_n3782__;
  assign new_new_n3962__ = ~new_new_n3960__ & new_new_n3961__;
  assign new_new_n3963__ = ~new_new_n3958__ & ~new_new_n3959__;
  assign new_new_n3964__ = ~new_new_n3962__ & new_new_n3963__;
  assign new_new_n3965__ = ~new_new_n3715__ & ~new_new_n3764__;
  assign new_new_n3966__ = ~new_new_n3716__ & ~new_new_n3965__;
  assign new_new_n3967__ = new_new_n3964__ & new_new_n3966__;
  assign new_new_n3968__ = ~new_new_n3964__ & ~new_new_n3966__;
  assign new_new_n3969__ = ~new_new_n3967__ & ~new_new_n3968__;
  assign new_new_n3970__ = new_new_n3951__ & ~new_new_n3969__;
  assign new_new_n3971__ = ~new_new_n3951__ & new_new_n3969__;
  assign new_new_n3972__ = ~new_new_n3970__ & ~new_new_n3971__;
  assign new_new_n3973__ = ~new_new_n3644__ & new_new_n3711__;
  assign new_new_n3974__ = ~new_new_n3645__ & ~new_new_n3973__;
  assign new_new_n3975__ = new_new_n3972__ & new_new_n3974__;
  assign new_new_n3976__ = ~new_new_n3972__ & ~new_new_n3974__;
  assign po039 = new_new_n3975__ | new_new_n3976__;
  assign new_new_n3978__ = new_new_n3885__ & ~new_new_n3964__;
  assign new_new_n3979__ = new_new_n3948__ & ~new_new_n3966__;
  assign new_new_n3980__ = new_new_n3978__ & new_new_n3979__;
  assign new_new_n3981__ = new_new_n3800__ & ~new_new_n3881__;
  assign new_new_n3982__ = ~new_new_n3880__ & ~new_new_n3981__;
  assign new_new_n3983__ = ~new_new_n3941__ & ~new_new_n3945__;
  assign new_new_n3984__ = ~new_new_n3942__ & ~new_new_n3983__;
  assign new_new_n3985__ = new_new_n3828__ & ~new_new_n3844__;
  assign new_new_n3986__ = ~new_new_n3843__ & ~new_new_n3985__;
  assign new_new_n3987__ = ~new_new_n3899__ & ~new_new_n3903__;
  assign new_new_n3988__ = ~new_new_n3902__ & ~new_new_n3987__;
  assign new_new_n3989__ = ~new_new_n3911__ & ~new_new_n3915__;
  assign new_new_n3990__ = ~new_new_n3914__ & ~new_new_n3989__;
  assign new_new_n3991__ = ~new_new_n3829__ & ~new_new_n3833__;
  assign new_new_n3992__ = ~new_new_n3832__ & ~new_new_n3991__;
  assign new_new_n3993__ = new_new_n3990__ & new_new_n3992__;
  assign new_new_n3994__ = ~new_new_n3990__ & ~new_new_n3992__;
  assign new_new_n3995__ = ~new_new_n3993__ & ~new_new_n3994__;
  assign new_new_n3996__ = new_new_n3988__ & ~new_new_n3995__;
  assign new_new_n3997__ = ~new_new_n3988__ & new_new_n3995__;
  assign new_new_n3998__ = ~new_new_n3996__ & ~new_new_n3997__;
  assign new_new_n3999__ = new_new_n3986__ & new_new_n3998__;
  assign new_new_n4000__ = ~new_new_n3986__ & ~new_new_n3998__;
  assign new_new_n4001__ = ~new_new_n3999__ & ~new_new_n4000__;
  assign new_new_n4002__ = pi19 & pi20;
  assign new_new_n4003__ = pi08 & pi31;
  assign new_new_n4004__ = pi18 & pi21;
  assign new_new_n4005__ = ~new_new_n4003__ & ~new_new_n4004__;
  assign new_new_n4006__ = new_new_n4003__ & new_new_n4004__;
  assign new_new_n4007__ = ~new_new_n4005__ & ~new_new_n4006__;
  assign new_new_n4008__ = new_new_n4002__ & ~new_new_n4007__;
  assign new_new_n4009__ = ~new_new_n4002__ & new_new_n4007__;
  assign new_new_n4010__ = ~new_new_n4008__ & ~new_new_n4009__;
  assign new_new_n4011__ = pi11 & pi28;
  assign new_new_n4012__ = pi10 & pi29;
  assign new_new_n4013__ = pi05 & pi34;
  assign new_new_n4014__ = ~new_new_n4012__ & ~new_new_n4013__;
  assign new_new_n4015__ = new_new_n4012__ & new_new_n4013__;
  assign new_new_n4016__ = ~new_new_n4014__ & ~new_new_n4015__;
  assign new_new_n4017__ = new_new_n4011__ & ~new_new_n4016__;
  assign new_new_n4018__ = ~new_new_n4011__ & new_new_n4016__;
  assign new_new_n4019__ = ~new_new_n4017__ & ~new_new_n4018__;
  assign new_new_n4020__ = new_new_n4010__ & new_new_n4019__;
  assign new_new_n4021__ = ~new_new_n4010__ & ~new_new_n4019__;
  assign new_new_n4022__ = ~new_new_n4020__ & ~new_new_n4021__;
  assign new_new_n4023__ = pi17 & pi22;
  assign new_new_n4024__ = pi12 & pi27;
  assign new_new_n4025__ = pi04 & pi35;
  assign new_new_n4026__ = ~new_new_n4024__ & ~new_new_n4025__;
  assign new_new_n4027__ = new_new_n4024__ & new_new_n4025__;
  assign new_new_n4028__ = ~new_new_n4026__ & ~new_new_n4027__;
  assign new_new_n4029__ = new_new_n4023__ & ~new_new_n4028__;
  assign new_new_n4030__ = ~new_new_n4023__ & new_new_n4028__;
  assign new_new_n4031__ = ~new_new_n4029__ & ~new_new_n4030__;
  assign new_new_n4032__ = ~new_new_n4022__ & new_new_n4031__;
  assign new_new_n4033__ = new_new_n4022__ & ~new_new_n4031__;
  assign new_new_n4034__ = ~new_new_n4032__ & ~new_new_n4033__;
  assign new_new_n4035__ = new_new_n4001__ & new_new_n4034__;
  assign new_new_n4036__ = ~new_new_n4001__ & ~new_new_n4034__;
  assign new_new_n4037__ = ~new_new_n4035__ & ~new_new_n4036__;
  assign new_new_n4038__ = ~new_new_n3984__ & new_new_n4037__;
  assign new_new_n4039__ = new_new_n3984__ & ~new_new_n4037__;
  assign new_new_n4040__ = ~new_new_n4038__ & ~new_new_n4039__;
  assign new_new_n4041__ = ~new_new_n3819__ & ~new_new_n3822__;
  assign new_new_n4042__ = ~new_new_n3818__ & ~new_new_n4041__;
  assign new_new_n4043__ = ~new_new_n3924__ & ~new_new_n3937__;
  assign new_new_n4044__ = ~new_new_n3923__ & ~new_new_n4043__;
  assign new_new_n4045__ = new_new_n4042__ & ~new_new_n4044__;
  assign new_new_n4046__ = ~new_new_n4042__ & new_new_n4044__;
  assign new_new_n4047__ = ~new_new_n4045__ & ~new_new_n4046__;
  assign new_new_n4048__ = pi09 & pi30;
  assign new_new_n4049__ = pi06 & pi33;
  assign new_new_n4050__ = pi07 & pi32;
  assign new_new_n4051__ = ~new_new_n4049__ & ~new_new_n4050__;
  assign new_new_n4052__ = new_new_n4049__ & new_new_n4050__;
  assign new_new_n4053__ = ~new_new_n4051__ & ~new_new_n4052__;
  assign new_new_n4054__ = new_new_n4048__ & ~new_new_n4053__;
  assign new_new_n4055__ = ~new_new_n4048__ & new_new_n4053__;
  assign new_new_n4056__ = ~new_new_n4054__ & ~new_new_n4055__;
  assign new_new_n4057__ = pi13 & pi26;
  assign new_new_n4058__ = pi03 & pi36;
  assign new_new_n4059__ = pi02 & pi37;
  assign new_new_n4060__ = ~new_new_n4058__ & ~new_new_n4059__;
  assign new_new_n4061__ = new_new_n4058__ & new_new_n4059__;
  assign new_new_n4062__ = ~new_new_n4060__ & ~new_new_n4061__;
  assign new_new_n4063__ = new_new_n4057__ & ~new_new_n4062__;
  assign new_new_n4064__ = ~new_new_n4057__ & new_new_n4062__;
  assign new_new_n4065__ = ~new_new_n4063__ & ~new_new_n4064__;
  assign new_new_n4066__ = new_new_n4056__ & new_new_n4065__;
  assign new_new_n4067__ = ~new_new_n4056__ & ~new_new_n4065__;
  assign new_new_n4068__ = ~new_new_n4066__ & ~new_new_n4067__;
  assign new_new_n4069__ = pi16 & pi23;
  assign new_new_n4070__ = pi14 & pi25;
  assign new_new_n4071__ = pi15 & pi24;
  assign new_new_n4072__ = ~new_new_n4070__ & ~new_new_n4071__;
  assign new_new_n4073__ = new_new_n4070__ & new_new_n4071__;
  assign new_new_n4074__ = ~new_new_n4072__ & ~new_new_n4073__;
  assign new_new_n4075__ = new_new_n4069__ & ~new_new_n4074__;
  assign new_new_n4076__ = ~new_new_n4069__ & new_new_n4074__;
  assign new_new_n4077__ = ~new_new_n4075__ & ~new_new_n4076__;
  assign new_new_n4078__ = new_new_n4068__ & ~new_new_n4077__;
  assign new_new_n4079__ = ~new_new_n4068__ & new_new_n4077__;
  assign new_new_n4080__ = ~new_new_n4078__ & ~new_new_n4079__;
  assign new_new_n4081__ = new_new_n4047__ & ~new_new_n4080__;
  assign new_new_n4082__ = ~new_new_n4047__ & new_new_n4080__;
  assign new_new_n4083__ = ~new_new_n4081__ & ~new_new_n4082__;
  assign new_new_n4084__ = new_new_n4040__ & ~new_new_n4083__;
  assign new_new_n4085__ = ~new_new_n4040__ & new_new_n4083__;
  assign new_new_n4086__ = ~new_new_n4084__ & ~new_new_n4085__;
  assign new_new_n4087__ = new_new_n3982__ & new_new_n4086__;
  assign new_new_n4088__ = ~new_new_n3982__ & ~new_new_n4086__;
  assign new_new_n4089__ = ~new_new_n4087__ & ~new_new_n4088__;
  assign new_new_n4090__ = new_new_n3807__ & ~new_new_n3812__;
  assign new_new_n4091__ = ~new_new_n3813__ & ~new_new_n4090__;
  assign new_new_n4092__ = pi00 & pi39;
  assign new_new_n4093__ = pi20 & pi38;
  assign new_new_n4094__ = ~new_new_n4092__ & ~new_new_n4093__;
  assign new_new_n4095__ = pi18 & pi37;
  assign new_new_n4096__ = pi01 & ~pi38;
  assign new_new_n4097__ = new_new_n4092__ & ~new_new_n4096__;
  assign new_new_n4098__ = ~new_new_n4094__ & new_new_n4095__;
  assign new_new_n4099__ = ~new_new_n4097__ & new_new_n4098__;
  assign new_new_n4100__ = new_new_n3803__ & new_new_n3804__;
  assign new_new_n4101__ = pi01 & pi38;
  assign new_new_n4102__ = ~new_new_n4092__ & new_new_n4101__;
  assign new_new_n4103__ = new_new_n4092__ & ~new_new_n4101__;
  assign new_new_n4104__ = ~new_new_n4102__ & ~new_new_n4103__;
  assign new_new_n4105__ = pi20 & ~new_new_n4104__;
  assign new_new_n4106__ = ~pi20 & new_new_n4104__;
  assign new_new_n4107__ = ~new_new_n4100__ & ~new_new_n4105__;
  assign new_new_n4108__ = ~new_new_n4106__ & new_new_n4107__;
  assign new_new_n4109__ = ~new_new_n4099__ & ~new_new_n4108__;
  assign new_new_n4110__ = ~new_new_n4091__ & new_new_n4109__;
  assign new_new_n4111__ = new_new_n4091__ & ~new_new_n4109__;
  assign new_new_n4112__ = ~new_new_n4110__ & ~new_new_n4111__;
  assign new_new_n4113__ = ~new_new_n3931__ & ~new_new_n3934__;
  assign new_new_n4114__ = ~new_new_n3930__ & ~new_new_n4113__;
  assign new_new_n4115__ = new_new_n4112__ & new_new_n4114__;
  assign new_new_n4116__ = ~new_new_n4112__ & ~new_new_n4114__;
  assign new_new_n4117__ = ~new_new_n4115__ & ~new_new_n4116__;
  assign new_new_n4118__ = ~new_new_n3850__ & new_new_n3876__;
  assign new_new_n4119__ = ~new_new_n3849__ & ~new_new_n4118__;
  assign new_new_n4120__ = ~new_new_n4117__ & ~new_new_n4119__;
  assign new_new_n4121__ = new_new_n4117__ & new_new_n4119__;
  assign new_new_n4122__ = ~new_new_n4120__ & ~new_new_n4121__;
  assign new_new_n4123__ = ~new_new_n3908__ & ~new_new_n3919__;
  assign new_new_n4124__ = ~new_new_n3909__ & ~new_new_n4123__;
  assign new_new_n4125__ = new_new_n3860__ & ~new_new_n3871__;
  assign new_new_n4126__ = ~new_new_n3872__ & ~new_new_n4125__;
  assign new_new_n4127__ = ~new_new_n3890__ & ~new_new_n3894__;
  assign new_new_n4128__ = ~new_new_n3893__ & ~new_new_n4127__;
  assign new_new_n4129__ = ~new_new_n3863__ & ~new_new_n3864__;
  assign new_new_n4130__ = new_new_n3866__ & ~new_new_n4129__;
  assign new_new_n4131__ = ~new_new_n3852__ & ~new_new_n3856__;
  assign new_new_n4132__ = ~new_new_n3855__ & ~new_new_n4131__;
  assign new_new_n4133__ = new_new_n4130__ & new_new_n4132__;
  assign new_new_n4134__ = ~new_new_n4130__ & ~new_new_n4132__;
  assign new_new_n4135__ = ~new_new_n4133__ & ~new_new_n4134__;
  assign new_new_n4136__ = new_new_n4128__ & ~new_new_n4135__;
  assign new_new_n4137__ = ~new_new_n4128__ & new_new_n4135__;
  assign new_new_n4138__ = ~new_new_n4136__ & ~new_new_n4137__;
  assign new_new_n4139__ = new_new_n4126__ & ~new_new_n4138__;
  assign new_new_n4140__ = ~new_new_n4126__ & new_new_n4138__;
  assign new_new_n4141__ = ~new_new_n4139__ & ~new_new_n4140__;
  assign new_new_n4142__ = new_new_n4124__ & ~new_new_n4141__;
  assign new_new_n4143__ = ~new_new_n4124__ & new_new_n4141__;
  assign new_new_n4144__ = ~new_new_n4142__ & ~new_new_n4143__;
  assign new_new_n4145__ = new_new_n4122__ & new_new_n4144__;
  assign new_new_n4146__ = ~new_new_n4122__ & ~new_new_n4144__;
  assign new_new_n4147__ = ~new_new_n4145__ & ~new_new_n4146__;
  assign new_new_n4148__ = new_new_n4089__ & ~new_new_n4147__;
  assign new_new_n4149__ = ~new_new_n4089__ & new_new_n4147__;
  assign new_new_n4150__ = ~new_new_n4148__ & ~new_new_n4149__;
  assign new_new_n4151__ = new_new_n3948__ & new_new_n3968__;
  assign new_new_n4152__ = ~new_new_n3948__ & ~new_new_n3968__;
  assign new_new_n4153__ = ~new_new_n3967__ & ~new_new_n4152__;
  assign new_new_n4154__ = new_new_n3885__ & new_new_n4153__;
  assign new_new_n4155__ = ~new_new_n3974__ & ~new_new_n4151__;
  assign new_new_n4156__ = ~new_new_n4154__ & new_new_n4155__;
  assign new_new_n4157__ = ~new_new_n3948__ & new_new_n3967__;
  assign new_new_n4158__ = ~new_new_n3885__ & ~new_new_n4153__;
  assign new_new_n4159__ = new_new_n3974__ & ~new_new_n4157__;
  assign new_new_n4160__ = ~new_new_n4158__ & new_new_n4159__;
  assign new_new_n4161__ = ~new_new_n4156__ & ~new_new_n4160__;
  assign new_new_n4162__ = ~new_new_n3948__ & new_new_n3966__;
  assign new_new_n4163__ = ~new_new_n3885__ & new_new_n3964__;
  assign new_new_n4164__ = new_new_n4162__ & new_new_n4163__;
  assign new_new_n4165__ = ~new_new_n3980__ & ~new_new_n4150__;
  assign new_new_n4166__ = ~new_new_n4164__ & new_new_n4165__;
  assign new_new_n4167__ = ~new_new_n4161__ & new_new_n4166__;
  assign new_new_n4168__ = ~new_new_n3950__ & new_new_n3974__;
  assign new_new_n4169__ = ~new_new_n3949__ & ~new_new_n4168__;
  assign new_new_n4170__ = new_new_n3967__ & new_new_n4169__;
  assign new_new_n4171__ = new_new_n3949__ & new_new_n3974__;
  assign new_new_n4172__ = new_new_n3950__ & ~new_new_n3974__;
  assign new_new_n4173__ = ~new_new_n4171__ & ~new_new_n4172__;
  assign new_new_n4174__ = new_new_n3969__ & new_new_n4173__;
  assign new_new_n4175__ = new_new_n3968__ & ~new_new_n4169__;
  assign new_new_n4176__ = new_new_n4150__ & ~new_new_n4170__;
  assign new_new_n4177__ = ~new_new_n4175__ & new_new_n4176__;
  assign new_new_n4178__ = ~new_new_n4174__ & new_new_n4177__;
  assign po040 = ~new_new_n4167__ & ~new_new_n4178__;
  assign new_new_n4180__ = new_new_n3974__ & ~new_new_n3979__;
  assign new_new_n4181__ = ~new_new_n4162__ & ~new_new_n4180__;
  assign new_new_n4182__ = ~new_new_n4150__ & ~new_new_n4181__;
  assign new_new_n4183__ = new_new_n3978__ & ~new_new_n4182__;
  assign new_new_n4184__ = new_new_n4150__ & new_new_n4181__;
  assign new_new_n4185__ = ~new_new_n3979__ & ~new_new_n4150__;
  assign new_new_n4186__ = new_new_n4150__ & ~new_new_n4162__;
  assign new_new_n4187__ = new_new_n3974__ & ~new_new_n4186__;
  assign new_new_n4188__ = ~new_new_n4185__ & ~new_new_n4187__;
  assign new_new_n4189__ = ~new_new_n4163__ & new_new_n4188__;
  assign new_new_n4190__ = ~new_new_n4183__ & ~new_new_n4184__;
  assign new_new_n4191__ = ~new_new_n4189__ & new_new_n4190__;
  assign new_new_n4192__ = ~new_new_n4038__ & new_new_n4083__;
  assign new_new_n4193__ = ~new_new_n4039__ & ~new_new_n4192__;
  assign new_new_n4194__ = ~new_new_n4191__ & ~new_new_n4193__;
  assign new_new_n4195__ = new_new_n4191__ & new_new_n4193__;
  assign new_new_n4196__ = ~new_new_n4194__ & ~new_new_n4195__;
  assign new_new_n4197__ = ~new_new_n4000__ & ~new_new_n4034__;
  assign new_new_n4198__ = ~new_new_n3999__ & ~new_new_n4197__;
  assign new_new_n4199__ = ~new_new_n4020__ & ~new_new_n4031__;
  assign new_new_n4200__ = ~new_new_n4021__ & ~new_new_n4199__;
  assign new_new_n4201__ = ~new_new_n4067__ & new_new_n4077__;
  assign new_new_n4202__ = ~new_new_n4066__ & ~new_new_n4201__;
  assign new_new_n4203__ = ~new_new_n4200__ & new_new_n4202__;
  assign new_new_n4204__ = new_new_n4200__ & ~new_new_n4202__;
  assign new_new_n4205__ = ~new_new_n4203__ & ~new_new_n4204__;
  assign new_new_n4206__ = ~new_new_n4011__ & ~new_new_n4015__;
  assign new_new_n4207__ = ~new_new_n4014__ & ~new_new_n4206__;
  assign new_new_n4208__ = ~new_new_n4057__ & ~new_new_n4061__;
  assign new_new_n4209__ = ~new_new_n4060__ & ~new_new_n4208__;
  assign new_new_n4210__ = ~new_new_n4023__ & ~new_new_n4027__;
  assign new_new_n4211__ = ~new_new_n4026__ & ~new_new_n4210__;
  assign new_new_n4212__ = new_new_n4209__ & new_new_n4211__;
  assign new_new_n4213__ = ~new_new_n4209__ & ~new_new_n4211__;
  assign new_new_n4214__ = ~new_new_n4207__ & ~new_new_n4212__;
  assign new_new_n4215__ = ~new_new_n4213__ & ~new_new_n4214__;
  assign new_new_n4216__ = ~new_new_n4212__ & new_new_n4215__;
  assign new_new_n4217__ = new_new_n4207__ & ~new_new_n4216__;
  assign new_new_n4218__ = ~new_new_n4213__ & new_new_n4214__;
  assign new_new_n4219__ = ~new_new_n4217__ & ~new_new_n4218__;
  assign new_new_n4220__ = new_new_n4205__ & ~new_new_n4219__;
  assign new_new_n4221__ = ~new_new_n4205__ & new_new_n4219__;
  assign new_new_n4222__ = ~new_new_n4220__ & ~new_new_n4221__;
  assign new_new_n4223__ = ~new_new_n4198__ & ~new_new_n4222__;
  assign new_new_n4224__ = new_new_n4198__ & new_new_n4222__;
  assign new_new_n4225__ = ~new_new_n4223__ & ~new_new_n4224__;
  assign new_new_n4226__ = ~new_new_n4046__ & new_new_n4080__;
  assign new_new_n4227__ = ~new_new_n4045__ & ~new_new_n4226__;
  assign new_new_n4228__ = new_new_n4225__ & ~new_new_n4227__;
  assign new_new_n4229__ = ~new_new_n4225__ & new_new_n4227__;
  assign new_new_n4230__ = ~new_new_n4228__ & ~new_new_n4229__;
  assign new_new_n4231__ = pi12 & pi28;
  assign new_new_n4232__ = pi05 & pi35;
  assign new_new_n4233__ = pi04 & pi36;
  assign new_new_n4234__ = ~new_new_n4232__ & ~new_new_n4233__;
  assign new_new_n4235__ = new_new_n4232__ & new_new_n4233__;
  assign new_new_n4236__ = ~new_new_n4234__ & ~new_new_n4235__;
  assign new_new_n4237__ = new_new_n4231__ & ~new_new_n4236__;
  assign new_new_n4238__ = ~new_new_n4231__ & new_new_n4236__;
  assign new_new_n4239__ = ~new_new_n4237__ & ~new_new_n4238__;
  assign new_new_n4240__ = pi09 & pi31;
  assign new_new_n4241__ = pi07 & pi33;
  assign new_new_n4242__ = pi08 & pi32;
  assign new_new_n4243__ = ~new_new_n4241__ & ~new_new_n4242__;
  assign new_new_n4244__ = new_new_n4241__ & new_new_n4242__;
  assign new_new_n4245__ = ~new_new_n4243__ & ~new_new_n4244__;
  assign new_new_n4246__ = new_new_n4240__ & ~new_new_n4245__;
  assign new_new_n4247__ = ~new_new_n4240__ & new_new_n4245__;
  assign new_new_n4248__ = ~new_new_n4246__ & ~new_new_n4247__;
  assign new_new_n4249__ = new_new_n4239__ & new_new_n4248__;
  assign new_new_n4250__ = ~new_new_n4239__ & ~new_new_n4248__;
  assign new_new_n4251__ = ~new_new_n4249__ & ~new_new_n4250__;
  assign new_new_n4252__ = pi18 & pi22;
  assign new_new_n4253__ = pi02 & pi38;
  assign new_new_n4254__ = pi00 & pi40;
  assign new_new_n4255__ = ~new_new_n4253__ & ~new_new_n4254__;
  assign new_new_n4256__ = new_new_n4253__ & new_new_n4254__;
  assign new_new_n4257__ = ~new_new_n4255__ & ~new_new_n4256__;
  assign new_new_n4258__ = new_new_n4252__ & ~new_new_n4257__;
  assign new_new_n4259__ = ~new_new_n4252__ & new_new_n4257__;
  assign new_new_n4260__ = ~new_new_n4258__ & ~new_new_n4259__;
  assign new_new_n4261__ = new_new_n4251__ & ~new_new_n4260__;
  assign new_new_n4262__ = ~new_new_n4251__ & new_new_n4260__;
  assign new_new_n4263__ = ~new_new_n4261__ & ~new_new_n4262__;
  assign new_new_n4264__ = ~new_new_n4110__ & new_new_n4114__;
  assign new_new_n4265__ = ~new_new_n4111__ & ~new_new_n4264__;
  assign new_new_n4266__ = new_new_n4263__ & ~new_new_n4265__;
  assign new_new_n4267__ = ~new_new_n4263__ & new_new_n4265__;
  assign new_new_n4268__ = ~new_new_n4266__ & ~new_new_n4267__;
  assign new_new_n4269__ = ~new_new_n4048__ & ~new_new_n4052__;
  assign new_new_n4270__ = ~new_new_n4051__ & ~new_new_n4269__;
  assign new_new_n4271__ = ~new_new_n4069__ & ~new_new_n4073__;
  assign new_new_n4272__ = ~new_new_n4072__ & ~new_new_n4271__;
  assign new_new_n4273__ = ~new_new_n4092__ & ~new_new_n4096__;
  assign new_new_n4274__ = new_new_n4095__ & ~new_new_n4273__;
  assign new_new_n4275__ = ~new_new_n4103__ & ~new_new_n4274__;
  assign new_new_n4276__ = pi20 & ~new_new_n4275__;
  assign new_new_n4277__ = ~pi20 & new_new_n4092__;
  assign new_new_n4278__ = new_new_n4101__ & new_new_n4277__;
  assign new_new_n4279__ = ~new_new_n4276__ & ~new_new_n4278__;
  assign new_new_n4280__ = new_new_n4272__ & ~new_new_n4279__;
  assign new_new_n4281__ = ~new_new_n4272__ & new_new_n4279__;
  assign new_new_n4282__ = ~new_new_n4280__ & ~new_new_n4281__;
  assign new_new_n4283__ = new_new_n4270__ & new_new_n4282__;
  assign new_new_n4284__ = ~new_new_n4270__ & ~new_new_n4282__;
  assign new_new_n4285__ = ~new_new_n4283__ & ~new_new_n4284__;
  assign new_new_n4286__ = new_new_n4268__ & ~new_new_n4285__;
  assign new_new_n4287__ = ~new_new_n4268__ & new_new_n4285__;
  assign new_new_n4288__ = ~new_new_n4286__ & ~new_new_n4287__;
  assign new_new_n4289__ = ~new_new_n4124__ & ~new_new_n4140__;
  assign new_new_n4290__ = ~new_new_n4139__ & ~new_new_n4289__;
  assign new_new_n4291__ = pi19 & pi21;
  assign new_new_n4292__ = ~new_new_n4002__ & ~new_new_n4006__;
  assign new_new_n4293__ = ~new_new_n4005__ & ~new_new_n4292__;
  assign new_new_n4294__ = new_new_n4291__ & new_new_n4293__;
  assign new_new_n4295__ = ~new_new_n4291__ & ~new_new_n4293__;
  assign new_new_n4296__ = ~new_new_n4294__ & ~new_new_n4295__;
  assign new_new_n4297__ = ~pi39 & ~new_new_n4093__;
  assign new_new_n4298__ = pi20 & pi39;
  assign new_new_n4299__ = pi38 & new_new_n4298__;
  assign new_new_n4300__ = pi01 & ~new_new_n4297__;
  assign new_new_n4301__ = ~new_new_n4299__ & new_new_n4300__;
  assign new_new_n4302__ = new_new_n4296__ & ~new_new_n4301__;
  assign new_new_n4303__ = ~new_new_n4296__ & new_new_n4301__;
  assign new_new_n4304__ = ~new_new_n4302__ & ~new_new_n4303__;
  assign new_new_n4305__ = ~new_new_n3988__ & ~new_new_n3993__;
  assign new_new_n4306__ = ~new_new_n3994__ & ~new_new_n4305__;
  assign new_new_n4307__ = new_new_n4304__ & ~new_new_n4306__;
  assign new_new_n4308__ = ~new_new_n4304__ & new_new_n4306__;
  assign new_new_n4309__ = ~new_new_n4307__ & ~new_new_n4308__;
  assign new_new_n4310__ = ~new_new_n4128__ & ~new_new_n4133__;
  assign new_new_n4311__ = ~new_new_n4134__ & ~new_new_n4310__;
  assign new_new_n4312__ = new_new_n4309__ & ~new_new_n4311__;
  assign new_new_n4313__ = ~new_new_n4309__ & new_new_n4311__;
  assign new_new_n4314__ = ~new_new_n4312__ & ~new_new_n4313__;
  assign new_new_n4315__ = ~new_new_n4290__ & ~new_new_n4314__;
  assign new_new_n4316__ = new_new_n4290__ & new_new_n4314__;
  assign new_new_n4317__ = ~new_new_n4315__ & ~new_new_n4316__;
  assign new_new_n4318__ = pi17 & pi23;
  assign new_new_n4319__ = pi15 & pi25;
  assign new_new_n4320__ = pi16 & pi24;
  assign new_new_n4321__ = ~new_new_n4319__ & ~new_new_n4320__;
  assign new_new_n4322__ = new_new_n4319__ & new_new_n4320__;
  assign new_new_n4323__ = ~new_new_n4321__ & ~new_new_n4322__;
  assign new_new_n4324__ = new_new_n4318__ & ~new_new_n4323__;
  assign new_new_n4325__ = ~new_new_n4318__ & new_new_n4323__;
  assign new_new_n4326__ = ~new_new_n4324__ & ~new_new_n4325__;
  assign new_new_n4327__ = pi11 & pi29;
  assign new_new_n4328__ = pi10 & pi30;
  assign new_new_n4329__ = pi06 & pi34;
  assign new_new_n4330__ = ~new_new_n4328__ & ~new_new_n4329__;
  assign new_new_n4331__ = new_new_n4328__ & new_new_n4329__;
  assign new_new_n4332__ = ~new_new_n4330__ & ~new_new_n4331__;
  assign new_new_n4333__ = new_new_n4327__ & ~new_new_n4332__;
  assign new_new_n4334__ = ~new_new_n4327__ & new_new_n4332__;
  assign new_new_n4335__ = ~new_new_n4333__ & ~new_new_n4334__;
  assign new_new_n4336__ = new_new_n4326__ & new_new_n4335__;
  assign new_new_n4337__ = ~new_new_n4326__ & ~new_new_n4335__;
  assign new_new_n4338__ = ~new_new_n4336__ & ~new_new_n4337__;
  assign new_new_n4339__ = pi13 & pi27;
  assign new_new_n4340__ = pi03 & pi37;
  assign new_new_n4341__ = ~new_new_n4339__ & ~new_new_n4340__;
  assign new_new_n4342__ = new_new_n4339__ & new_new_n4340__;
  assign new_new_n4343__ = ~new_new_n4341__ & ~new_new_n4342__;
  assign new_new_n4344__ = new_new_n2379__ & ~new_new_n4343__;
  assign new_new_n4345__ = ~new_new_n2379__ & new_new_n4343__;
  assign new_new_n4346__ = ~new_new_n4344__ & ~new_new_n4345__;
  assign new_new_n4347__ = new_new_n4338__ & ~new_new_n4346__;
  assign new_new_n4348__ = ~new_new_n4338__ & new_new_n4346__;
  assign new_new_n4349__ = ~new_new_n4347__ & ~new_new_n4348__;
  assign new_new_n4350__ = new_new_n4317__ & ~new_new_n4349__;
  assign new_new_n4351__ = ~new_new_n4317__ & new_new_n4349__;
  assign new_new_n4352__ = ~new_new_n4350__ & ~new_new_n4351__;
  assign new_new_n4353__ = ~new_new_n4288__ & ~new_new_n4352__;
  assign new_new_n4354__ = new_new_n4288__ & new_new_n4352__;
  assign new_new_n4355__ = ~new_new_n4353__ & ~new_new_n4354__;
  assign new_new_n4356__ = ~new_new_n4121__ & ~new_new_n4144__;
  assign new_new_n4357__ = ~new_new_n4120__ & ~new_new_n4356__;
  assign new_new_n4358__ = new_new_n4355__ & ~new_new_n4357__;
  assign new_new_n4359__ = ~new_new_n4355__ & new_new_n4357__;
  assign new_new_n4360__ = ~new_new_n4358__ & ~new_new_n4359__;
  assign new_new_n4361__ = ~new_new_n4230__ & new_new_n4360__;
  assign new_new_n4362__ = new_new_n4230__ & ~new_new_n4360__;
  assign new_new_n4363__ = ~new_new_n4361__ & ~new_new_n4362__;
  assign new_new_n4364__ = ~new_new_n4088__ & new_new_n4147__;
  assign new_new_n4365__ = ~new_new_n4087__ & ~new_new_n4364__;
  assign new_new_n4366__ = new_new_n4363__ & ~new_new_n4365__;
  assign new_new_n4367__ = ~new_new_n4363__ & new_new_n4365__;
  assign new_new_n4368__ = ~new_new_n4366__ & ~new_new_n4367__;
  assign new_new_n4369__ = new_new_n4196__ & new_new_n4368__;
  assign new_new_n4370__ = ~new_new_n4196__ & ~new_new_n4368__;
  assign po041 = ~new_new_n4369__ & ~new_new_n4370__;
  assign new_new_n4372__ = ~new_new_n4361__ & ~new_new_n4365__;
  assign new_new_n4373__ = ~new_new_n4354__ & new_new_n4357__;
  assign new_new_n4374__ = ~new_new_n4353__ & ~new_new_n4373__;
  assign new_new_n4375__ = ~new_new_n4223__ & ~new_new_n4227__;
  assign new_new_n4376__ = ~new_new_n4224__ & ~new_new_n4375__;
  assign new_new_n4377__ = ~new_new_n4336__ & ~new_new_n4346__;
  assign new_new_n4378__ = ~new_new_n4337__ & ~new_new_n4377__;
  assign new_new_n4379__ = ~new_new_n4270__ & ~new_new_n4280__;
  assign new_new_n4380__ = ~new_new_n4281__ & ~new_new_n4379__;
  assign new_new_n4381__ = ~new_new_n4215__ & ~new_new_n4380__;
  assign new_new_n4382__ = new_new_n4215__ & new_new_n4380__;
  assign new_new_n4383__ = ~new_new_n4381__ & ~new_new_n4382__;
  assign new_new_n4384__ = new_new_n4378__ & ~new_new_n4383__;
  assign new_new_n4385__ = ~new_new_n4378__ & new_new_n4383__;
  assign new_new_n4386__ = ~new_new_n4384__ & ~new_new_n4385__;
  assign new_new_n4387__ = ~new_new_n4203__ & new_new_n4219__;
  assign new_new_n4388__ = ~new_new_n4204__ & ~new_new_n4387__;
  assign new_new_n4389__ = ~new_new_n4386__ & ~new_new_n4388__;
  assign new_new_n4390__ = new_new_n4386__ & new_new_n4388__;
  assign new_new_n4391__ = ~new_new_n4389__ & ~new_new_n4390__;
  assign new_new_n4392__ = pi15 & pi26;
  assign new_new_n4393__ = pi13 & pi28;
  assign new_new_n4394__ = pi03 & pi38;
  assign new_new_n4395__ = ~new_new_n4393__ & ~new_new_n4394__;
  assign new_new_n4396__ = new_new_n4393__ & new_new_n4394__;
  assign new_new_n4397__ = ~new_new_n4395__ & ~new_new_n4396__;
  assign new_new_n4398__ = new_new_n4392__ & ~new_new_n4397__;
  assign new_new_n4399__ = ~new_new_n4392__ & new_new_n4397__;
  assign new_new_n4400__ = ~new_new_n4398__ & ~new_new_n4399__;
  assign new_new_n4401__ = pi00 & pi41;
  assign new_new_n4402__ = pi21 & new_new_n1223__;
  assign new_new_n4403__ = ~pi02 & ~new_new_n4402__;
  assign new_new_n4404__ = pi39 & ~new_new_n4403__;
  assign new_new_n4405__ = pi21 & new_new_n3864__;
  assign new_new_n4406__ = new_new_n4404__ & ~new_new_n4405__;
  assign new_new_n4407__ = new_new_n4401__ & ~new_new_n4406__;
  assign new_new_n4408__ = ~new_new_n4401__ & new_new_n4406__;
  assign new_new_n4409__ = ~new_new_n4407__ & ~new_new_n4408__;
  assign new_new_n4410__ = new_new_n4400__ & new_new_n4409__;
  assign new_new_n4411__ = ~new_new_n4400__ & ~new_new_n4409__;
  assign new_new_n4412__ = ~new_new_n4410__ & ~new_new_n4411__;
  assign new_new_n4413__ = ~new_new_n4231__ & ~new_new_n4235__;
  assign new_new_n4414__ = ~new_new_n4234__ & ~new_new_n4413__;
  assign new_new_n4415__ = new_new_n4412__ & ~new_new_n4414__;
  assign new_new_n4416__ = ~new_new_n4412__ & new_new_n4414__;
  assign new_new_n4417__ = ~new_new_n4415__ & ~new_new_n4416__;
  assign new_new_n4418__ = new_new_n4391__ & ~new_new_n4417__;
  assign new_new_n4419__ = ~new_new_n4391__ & new_new_n4417__;
  assign new_new_n4420__ = ~new_new_n4418__ & ~new_new_n4419__;
  assign new_new_n4421__ = ~new_new_n4376__ & new_new_n4420__;
  assign new_new_n4422__ = new_new_n4376__ & ~new_new_n4420__;
  assign new_new_n4423__ = ~new_new_n4421__ & ~new_new_n4422__;
  assign new_new_n4424__ = ~new_new_n4308__ & ~new_new_n4311__;
  assign new_new_n4425__ = ~new_new_n4307__ & ~new_new_n4424__;
  assign new_new_n4426__ = ~new_new_n4093__ & ~new_new_n4293__;
  assign new_new_n4427__ = pi39 & ~new_new_n4291__;
  assign new_new_n4428__ = ~new_new_n4426__ & new_new_n4427__;
  assign new_new_n4429__ = ~pi39 & new_new_n4291__;
  assign new_new_n4430__ = ~new_new_n4293__ & ~new_new_n4429__;
  assign new_new_n4431__ = new_new_n4093__ & ~new_new_n4430__;
  assign new_new_n4432__ = ~new_new_n4428__ & ~new_new_n4431__;
  assign new_new_n4433__ = pi01 & ~new_new_n4432__;
  assign new_new_n4434__ = pi01 & pi39;
  assign new_new_n4435__ = new_new_n4294__ & ~new_new_n4434__;
  assign new_new_n4436__ = ~new_new_n4433__ & ~new_new_n4435__;
  assign new_new_n4437__ = pi11 & pi30;
  assign new_new_n4438__ = pi05 & pi36;
  assign new_new_n4439__ = pi06 & pi35;
  assign new_new_n4440__ = ~new_new_n4438__ & ~new_new_n4439__;
  assign new_new_n4441__ = new_new_n4438__ & new_new_n4439__;
  assign new_new_n4442__ = ~new_new_n4440__ & ~new_new_n4441__;
  assign new_new_n4443__ = new_new_n4437__ & ~new_new_n4442__;
  assign new_new_n4444__ = ~new_new_n4437__ & new_new_n4442__;
  assign new_new_n4445__ = ~new_new_n4443__ & ~new_new_n4444__;
  assign new_new_n4446__ = new_new_n4436__ & new_new_n4445__;
  assign new_new_n4447__ = ~new_new_n4436__ & ~new_new_n4445__;
  assign new_new_n4448__ = ~new_new_n4446__ & ~new_new_n4447__;
  assign new_new_n4449__ = pi20 & pi21;
  assign new_new_n4450__ = pi08 & pi33;
  assign new_new_n4451__ = pi19 & pi22;
  assign new_new_n4452__ = new_new_n4450__ & ~new_new_n4451__;
  assign new_new_n4453__ = ~new_new_n4450__ & new_new_n4451__;
  assign new_new_n4454__ = ~new_new_n4452__ & ~new_new_n4453__;
  assign new_new_n4455__ = new_new_n4449__ & new_new_n4454__;
  assign new_new_n4456__ = ~new_new_n4449__ & ~new_new_n4454__;
  assign new_new_n4457__ = ~new_new_n4455__ & ~new_new_n4456__;
  assign new_new_n4458__ = new_new_n4448__ & ~new_new_n4457__;
  assign new_new_n4459__ = ~new_new_n4448__ & new_new_n4457__;
  assign new_new_n4460__ = ~new_new_n4458__ & ~new_new_n4459__;
  assign new_new_n4461__ = ~new_new_n4425__ & ~new_new_n4460__;
  assign new_new_n4462__ = new_new_n4425__ & new_new_n4460__;
  assign new_new_n4463__ = ~new_new_n4461__ & ~new_new_n4462__;
  assign new_new_n4464__ = pi18 & pi23;
  assign new_new_n4465__ = pi16 & pi25;
  assign new_new_n4466__ = pi17 & pi24;
  assign new_new_n4467__ = ~new_new_n4465__ & ~new_new_n4466__;
  assign new_new_n4468__ = new_new_n4465__ & new_new_n4466__;
  assign new_new_n4469__ = ~new_new_n4467__ & ~new_new_n4468__;
  assign new_new_n4470__ = new_new_n4464__ & ~new_new_n4469__;
  assign new_new_n4471__ = ~new_new_n4464__ & new_new_n4469__;
  assign new_new_n4472__ = ~new_new_n4470__ & ~new_new_n4471__;
  assign new_new_n4473__ = pi14 & pi27;
  assign new_new_n4474__ = pi12 & pi29;
  assign new_new_n4475__ = pi04 & pi37;
  assign new_new_n4476__ = ~new_new_n4474__ & ~new_new_n4475__;
  assign new_new_n4477__ = new_new_n4474__ & new_new_n4475__;
  assign new_new_n4478__ = ~new_new_n4476__ & ~new_new_n4477__;
  assign new_new_n4479__ = new_new_n4473__ & ~new_new_n4478__;
  assign new_new_n4480__ = ~new_new_n4473__ & new_new_n4478__;
  assign new_new_n4481__ = ~new_new_n4479__ & ~new_new_n4480__;
  assign new_new_n4482__ = new_new_n4472__ & new_new_n4481__;
  assign new_new_n4483__ = ~new_new_n4472__ & ~new_new_n4481__;
  assign new_new_n4484__ = ~new_new_n4482__ & ~new_new_n4483__;
  assign new_new_n4485__ = pi10 & pi31;
  assign new_new_n4486__ = pi09 & pi32;
  assign new_new_n4487__ = pi07 & pi34;
  assign new_new_n4488__ = ~new_new_n4486__ & ~new_new_n4487__;
  assign new_new_n4489__ = new_new_n4486__ & new_new_n4487__;
  assign new_new_n4490__ = ~new_new_n4488__ & ~new_new_n4489__;
  assign new_new_n4491__ = new_new_n4485__ & ~new_new_n4490__;
  assign new_new_n4492__ = ~new_new_n4485__ & new_new_n4490__;
  assign new_new_n4493__ = ~new_new_n4491__ & ~new_new_n4492__;
  assign new_new_n4494__ = new_new_n4484__ & ~new_new_n4493__;
  assign new_new_n4495__ = ~new_new_n4484__ & new_new_n4493__;
  assign new_new_n4496__ = ~new_new_n4494__ & ~new_new_n4495__;
  assign new_new_n4497__ = new_new_n4463__ & new_new_n4496__;
  assign new_new_n4498__ = ~new_new_n4463__ & ~new_new_n4496__;
  assign new_new_n4499__ = ~new_new_n4497__ & ~new_new_n4498__;
  assign new_new_n4500__ = new_new_n4423__ & ~new_new_n4499__;
  assign new_new_n4501__ = ~new_new_n4423__ & new_new_n4499__;
  assign new_new_n4502__ = ~new_new_n4500__ & ~new_new_n4501__;
  assign new_new_n4503__ = new_new_n4374__ & new_new_n4502__;
  assign new_new_n4504__ = ~new_new_n4374__ & ~new_new_n4502__;
  assign new_new_n4505__ = ~new_new_n4503__ & ~new_new_n4504__;
  assign new_new_n4506__ = ~new_new_n4315__ & ~new_new_n4349__;
  assign new_new_n4507__ = ~new_new_n4316__ & ~new_new_n4506__;
  assign new_new_n4508__ = ~new_new_n2379__ & ~new_new_n4342__;
  assign new_new_n4509__ = ~new_new_n4341__ & ~new_new_n4508__;
  assign new_new_n4510__ = ~new_new_n4252__ & ~new_new_n4256__;
  assign new_new_n4511__ = ~new_new_n4255__ & ~new_new_n4510__;
  assign new_new_n4512__ = ~new_new_n4509__ & ~new_new_n4511__;
  assign new_new_n4513__ = new_new_n4509__ & new_new_n4511__;
  assign new_new_n4514__ = ~new_new_n4512__ & ~new_new_n4513__;
  assign new_new_n4515__ = ~new_new_n4318__ & ~new_new_n4322__;
  assign new_new_n4516__ = ~new_new_n4321__ & ~new_new_n4515__;
  assign new_new_n4517__ = ~new_new_n4514__ & new_new_n4516__;
  assign new_new_n4518__ = ~new_new_n4513__ & ~new_new_n4516__;
  assign new_new_n4519__ = ~new_new_n4512__ & new_new_n4518__;
  assign new_new_n4520__ = ~new_new_n4517__ & ~new_new_n4519__;
  assign new_new_n4521__ = ~new_new_n4249__ & ~new_new_n4260__;
  assign new_new_n4522__ = ~new_new_n4250__ & ~new_new_n4521__;
  assign new_new_n4523__ = pi01 & pi40;
  assign new_new_n4524__ = pi21 & new_new_n4523__;
  assign new_new_n4525__ = ~pi21 & ~new_new_n4523__;
  assign new_new_n4526__ = ~new_new_n4524__ & ~new_new_n4525__;
  assign new_new_n4527__ = ~new_new_n4327__ & ~new_new_n4331__;
  assign new_new_n4528__ = ~new_new_n4330__ & ~new_new_n4527__;
  assign new_new_n4529__ = ~new_new_n4240__ & ~new_new_n4244__;
  assign new_new_n4530__ = ~new_new_n4243__ & ~new_new_n4529__;
  assign new_new_n4531__ = ~new_new_n4528__ & ~new_new_n4530__;
  assign new_new_n4532__ = new_new_n4528__ & new_new_n4530__;
  assign new_new_n4533__ = ~new_new_n4531__ & ~new_new_n4532__;
  assign new_new_n4534__ = new_new_n4526__ & ~new_new_n4533__;
  assign new_new_n4535__ = ~new_new_n4526__ & new_new_n4533__;
  assign new_new_n4536__ = ~new_new_n4534__ & ~new_new_n4535__;
  assign new_new_n4537__ = new_new_n4522__ & new_new_n4536__;
  assign new_new_n4538__ = ~new_new_n4522__ & ~new_new_n4536__;
  assign new_new_n4539__ = ~new_new_n4537__ & ~new_new_n4538__;
  assign new_new_n4540__ = new_new_n4520__ & new_new_n4539__;
  assign new_new_n4541__ = ~new_new_n4520__ & ~new_new_n4539__;
  assign new_new_n4542__ = ~new_new_n4540__ & ~new_new_n4541__;
  assign new_new_n4543__ = new_new_n4507__ & ~new_new_n4542__;
  assign new_new_n4544__ = ~new_new_n4507__ & new_new_n4542__;
  assign new_new_n4545__ = ~new_new_n4543__ & ~new_new_n4544__;
  assign new_new_n4546__ = ~new_new_n4266__ & ~new_new_n4285__;
  assign new_new_n4547__ = ~new_new_n4267__ & ~new_new_n4546__;
  assign new_new_n4548__ = new_new_n4545__ & ~new_new_n4547__;
  assign new_new_n4549__ = ~new_new_n4545__ & new_new_n4547__;
  assign new_new_n4550__ = ~new_new_n4548__ & ~new_new_n4549__;
  assign new_new_n4551__ = new_new_n4505__ & ~new_new_n4550__;
  assign new_new_n4552__ = ~new_new_n4505__ & new_new_n4550__;
  assign new_new_n4553__ = ~new_new_n4551__ & ~new_new_n4552__;
  assign new_new_n4554__ = new_new_n4194__ & ~new_new_n4553__;
  assign new_new_n4555__ = ~new_new_n4372__ & new_new_n4554__;
  assign new_new_n4556__ = ~new_new_n4194__ & new_new_n4553__;
  assign new_new_n4557__ = ~new_new_n4195__ & new_new_n4365__;
  assign new_new_n4558__ = new_new_n4191__ & ~new_new_n4361__;
  assign new_new_n4559__ = new_new_n4556__ & ~new_new_n4558__;
  assign new_new_n4560__ = ~new_new_n4557__ & new_new_n4559__;
  assign new_new_n4561__ = ~new_new_n4555__ & ~new_new_n4560__;
  assign new_new_n4562__ = ~new_new_n4362__ & ~new_new_n4561__;
  assign new_new_n4563__ = ~new_new_n4193__ & new_new_n4365__;
  assign new_new_n4564__ = ~new_new_n4191__ & ~new_new_n4362__;
  assign new_new_n4565__ = new_new_n4563__ & new_new_n4564__;
  assign new_new_n4566__ = new_new_n4553__ & ~new_new_n4565__;
  assign new_new_n4567__ = new_new_n4362__ & ~new_new_n4563__;
  assign new_new_n4568__ = new_new_n4191__ & new_new_n4567__;
  assign new_new_n4569__ = new_new_n4193__ & ~new_new_n4365__;
  assign new_new_n4570__ = ~new_new_n4564__ & new_new_n4569__;
  assign new_new_n4571__ = ~new_new_n4568__ & ~new_new_n4570__;
  assign new_new_n4572__ = ~new_new_n4566__ & new_new_n4571__;
  assign new_new_n4573__ = new_new_n4553__ & ~new_new_n4571__;
  assign new_new_n4574__ = ~new_new_n4361__ & ~new_new_n4572__;
  assign new_new_n4575__ = ~new_new_n4573__ & new_new_n4574__;
  assign new_new_n4576__ = new_new_n4361__ & new_new_n4365__;
  assign new_new_n4577__ = ~new_new_n4553__ & new_new_n4576__;
  assign new_new_n4578__ = new_new_n4196__ & new_new_n4577__;
  assign new_new_n4579__ = ~new_new_n4562__ & ~new_new_n4578__;
  assign po042 = ~new_new_n4575__ & new_new_n4579__;
  assign new_new_n4581__ = ~new_new_n4421__ & ~new_new_n4499__;
  assign new_new_n4582__ = ~new_new_n4422__ & ~new_new_n4581__;
  assign new_new_n4583__ = ~new_new_n4544__ & new_new_n4547__;
  assign new_new_n4584__ = ~new_new_n4543__ & ~new_new_n4583__;
  assign new_new_n4585__ = ~new_new_n4378__ & ~new_new_n4381__;
  assign new_new_n4586__ = ~new_new_n4382__ & ~new_new_n4585__;
  assign new_new_n4587__ = ~new_new_n4485__ & ~new_new_n4489__;
  assign new_new_n4588__ = ~new_new_n4488__ & ~new_new_n4587__;
  assign new_new_n4589__ = pi10 & pi32;
  assign new_new_n4590__ = pi09 & pi33;
  assign new_new_n4591__ = pi08 & pi34;
  assign new_new_n4592__ = ~new_new_n4590__ & ~new_new_n4591__;
  assign new_new_n4593__ = new_new_n4590__ & new_new_n4591__;
  assign new_new_n4594__ = ~new_new_n4592__ & ~new_new_n4593__;
  assign new_new_n4595__ = new_new_n4589__ & ~new_new_n4594__;
  assign new_new_n4596__ = ~new_new_n4589__ & new_new_n4594__;
  assign new_new_n4597__ = ~new_new_n4595__ & ~new_new_n4596__;
  assign new_new_n4598__ = ~new_new_n4588__ & new_new_n4597__;
  assign new_new_n4599__ = new_new_n4588__ & ~new_new_n4597__;
  assign new_new_n4600__ = ~new_new_n4598__ & ~new_new_n4599__;
  assign new_new_n4601__ = pi11 & pi31;
  assign new_new_n4602__ = pi06 & pi36;
  assign new_new_n4603__ = pi07 & pi35;
  assign new_new_n4604__ = ~new_new_n4602__ & ~new_new_n4603__;
  assign new_new_n4605__ = new_new_n4602__ & new_new_n4603__;
  assign new_new_n4606__ = ~new_new_n4604__ & ~new_new_n4605__;
  assign new_new_n4607__ = new_new_n4601__ & ~new_new_n4606__;
  assign new_new_n4608__ = ~new_new_n4601__ & new_new_n4606__;
  assign new_new_n4609__ = ~new_new_n4607__ & ~new_new_n4608__;
  assign new_new_n4610__ = new_new_n4600__ & new_new_n4609__;
  assign new_new_n4611__ = ~new_new_n4600__ & ~new_new_n4609__;
  assign new_new_n4612__ = ~new_new_n4610__ & ~new_new_n4611__;
  assign new_new_n4613__ = pi19 & pi23;
  assign new_new_n4614__ = pi17 & pi25;
  assign new_new_n4615__ = pi18 & pi24;
  assign new_new_n4616__ = ~new_new_n4614__ & ~new_new_n4615__;
  assign new_new_n4617__ = new_new_n4614__ & new_new_n4615__;
  assign new_new_n4618__ = ~new_new_n4616__ & ~new_new_n4617__;
  assign new_new_n4619__ = new_new_n4613__ & ~new_new_n4618__;
  assign new_new_n4620__ = ~new_new_n4613__ & new_new_n4618__;
  assign new_new_n4621__ = ~new_new_n4619__ & ~new_new_n4620__;
  assign new_new_n4622__ = pi15 & pi27;
  assign new_new_n4623__ = pi14 & pi28;
  assign new_new_n4624__ = pi04 & pi38;
  assign new_new_n4625__ = ~new_new_n4623__ & ~new_new_n4624__;
  assign new_new_n4626__ = new_new_n4623__ & new_new_n4624__;
  assign new_new_n4627__ = ~new_new_n4625__ & ~new_new_n4626__;
  assign new_new_n4628__ = new_new_n4622__ & ~new_new_n4627__;
  assign new_new_n4629__ = ~new_new_n4622__ & new_new_n4627__;
  assign new_new_n4630__ = ~new_new_n4628__ & ~new_new_n4629__;
  assign new_new_n4631__ = new_new_n4621__ & new_new_n4630__;
  assign new_new_n4632__ = ~new_new_n4621__ & ~new_new_n4630__;
  assign new_new_n4633__ = ~new_new_n4631__ & ~new_new_n4632__;
  assign new_new_n4634__ = pi16 & pi26;
  assign new_new_n4635__ = pi02 & pi40;
  assign new_new_n4636__ = pi03 & pi39;
  assign new_new_n4637__ = ~new_new_n4635__ & ~new_new_n4636__;
  assign new_new_n4638__ = new_new_n4635__ & new_new_n4636__;
  assign new_new_n4639__ = ~new_new_n4637__ & ~new_new_n4638__;
  assign new_new_n4640__ = new_new_n4634__ & ~new_new_n4639__;
  assign new_new_n4641__ = ~new_new_n4634__ & new_new_n4639__;
  assign new_new_n4642__ = ~new_new_n4640__ & ~new_new_n4641__;
  assign new_new_n4643__ = new_new_n4633__ & ~new_new_n4642__;
  assign new_new_n4644__ = ~new_new_n4633__ & new_new_n4642__;
  assign new_new_n4645__ = ~new_new_n4643__ & ~new_new_n4644__;
  assign new_new_n4646__ = ~new_new_n4612__ & ~new_new_n4645__;
  assign new_new_n4647__ = new_new_n4612__ & new_new_n4645__;
  assign new_new_n4648__ = ~new_new_n4646__ & ~new_new_n4647__;
  assign new_new_n4649__ = new_new_n4586__ & new_new_n4648__;
  assign new_new_n4650__ = ~new_new_n4586__ & ~new_new_n4648__;
  assign new_new_n4651__ = ~new_new_n4649__ & ~new_new_n4650__;
  assign new_new_n4652__ = ~new_new_n4584__ & new_new_n4651__;
  assign new_new_n4653__ = new_new_n4584__ & ~new_new_n4651__;
  assign new_new_n4654__ = ~new_new_n4652__ & ~new_new_n4653__;
  assign new_new_n4655__ = ~new_new_n4401__ & ~new_new_n4405__;
  assign new_new_n4656__ = new_new_n4404__ & ~new_new_n4655__;
  assign new_new_n4657__ = ~new_new_n4464__ & ~new_new_n4468__;
  assign new_new_n4658__ = ~new_new_n4467__ & ~new_new_n4657__;
  assign new_new_n4659__ = new_new_n4656__ & new_new_n4658__;
  assign new_new_n4660__ = ~new_new_n4656__ & ~new_new_n4658__;
  assign new_new_n4661__ = ~new_new_n4659__ & ~new_new_n4660__;
  assign new_new_n4662__ = ~new_new_n4392__ & ~new_new_n4396__;
  assign new_new_n4663__ = ~new_new_n4395__ & ~new_new_n4662__;
  assign new_new_n4664__ = ~new_new_n4661__ & new_new_n4663__;
  assign new_new_n4665__ = ~new_new_n4659__ & ~new_new_n4663__;
  assign new_new_n4666__ = ~new_new_n4660__ & new_new_n4665__;
  assign new_new_n4667__ = ~new_new_n4664__ & ~new_new_n4666__;
  assign new_new_n4668__ = ~new_new_n4473__ & ~new_new_n4477__;
  assign new_new_n4669__ = ~new_new_n4476__ & ~new_new_n4668__;
  assign new_new_n4670__ = ~new_new_n4437__ & ~new_new_n4441__;
  assign new_new_n4671__ = ~new_new_n4440__ & ~new_new_n4670__;
  assign new_new_n4672__ = ~new_new_n4669__ & ~new_new_n4671__;
  assign new_new_n4673__ = new_new_n4669__ & new_new_n4671__;
  assign new_new_n4674__ = ~new_new_n4672__ & ~new_new_n4673__;
  assign new_new_n4675__ = new_new_n4449__ & new_new_n4450__;
  assign new_new_n4676__ = ~new_new_n4451__ & ~new_new_n4675__;
  assign new_new_n4677__ = ~new_new_n4449__ & ~new_new_n4450__;
  assign new_new_n4678__ = ~new_new_n4676__ & ~new_new_n4677__;
  assign new_new_n4679__ = ~new_new_n4674__ & new_new_n4678__;
  assign new_new_n4680__ = new_new_n4674__ & ~new_new_n4678__;
  assign new_new_n4681__ = ~new_new_n4679__ & ~new_new_n4680__;
  assign new_new_n4682__ = ~new_new_n4447__ & new_new_n4457__;
  assign new_new_n4683__ = ~new_new_n4446__ & ~new_new_n4682__;
  assign new_new_n4684__ = new_new_n4681__ & ~new_new_n4683__;
  assign new_new_n4685__ = ~new_new_n4681__ & new_new_n4683__;
  assign new_new_n4686__ = ~new_new_n4684__ & ~new_new_n4685__;
  assign new_new_n4687__ = ~new_new_n4667__ & new_new_n4686__;
  assign new_new_n4688__ = new_new_n4667__ & ~new_new_n4686__;
  assign new_new_n4689__ = ~new_new_n4687__ & ~new_new_n4688__;
  assign new_new_n4690__ = pi13 & pi29;
  assign new_new_n4691__ = pi12 & pi30;
  assign new_new_n4692__ = pi05 & pi37;
  assign new_new_n4693__ = ~new_new_n4691__ & ~new_new_n4692__;
  assign new_new_n4694__ = new_new_n4691__ & new_new_n4692__;
  assign new_new_n4695__ = ~new_new_n4693__ & ~new_new_n4694__;
  assign new_new_n4696__ = new_new_n4690__ & ~new_new_n4695__;
  assign new_new_n4697__ = ~new_new_n4690__ & new_new_n4695__;
  assign new_new_n4698__ = ~new_new_n4696__ & ~new_new_n4697__;
  assign new_new_n4699__ = pi00 & pi42;
  assign new_new_n4700__ = pi20 & pi22;
  assign new_new_n4701__ = pi21 & pi40;
  assign new_new_n4702__ = ~pi41 & ~new_new_n4701__;
  assign new_new_n4703__ = pi41 & new_new_n4701__;
  assign new_new_n4704__ = pi01 & ~new_new_n4702__;
  assign new_new_n4705__ = ~new_new_n4703__ & new_new_n4704__;
  assign new_new_n4706__ = new_new_n4700__ & ~new_new_n4705__;
  assign new_new_n4707__ = ~new_new_n4700__ & new_new_n4705__;
  assign new_new_n4708__ = ~new_new_n4706__ & ~new_new_n4707__;
  assign new_new_n4709__ = new_new_n4699__ & new_new_n4708__;
  assign new_new_n4710__ = ~new_new_n4699__ & ~new_new_n4708__;
  assign new_new_n4711__ = ~new_new_n4709__ & ~new_new_n4710__;
  assign new_new_n4712__ = new_new_n4698__ & new_new_n4711__;
  assign new_new_n4713__ = ~new_new_n4698__ & ~new_new_n4711__;
  assign new_new_n4714__ = ~new_new_n4712__ & ~new_new_n4713__;
  assign new_new_n4715__ = new_new_n4526__ & ~new_new_n4531__;
  assign new_new_n4716__ = ~new_new_n4532__ & ~new_new_n4715__;
  assign new_new_n4717__ = new_new_n4714__ & ~new_new_n4716__;
  assign new_new_n4718__ = ~new_new_n4714__ & new_new_n4716__;
  assign new_new_n4719__ = ~new_new_n4717__ & ~new_new_n4718__;
  assign new_new_n4720__ = new_new_n4689__ & new_new_n4719__;
  assign new_new_n4721__ = ~new_new_n4689__ & ~new_new_n4719__;
  assign new_new_n4722__ = ~new_new_n4720__ & ~new_new_n4721__;
  assign new_new_n4723__ = ~new_new_n4520__ & ~new_new_n4537__;
  assign new_new_n4724__ = ~new_new_n4538__ & ~new_new_n4723__;
  assign new_new_n4725__ = new_new_n4722__ & new_new_n4724__;
  assign new_new_n4726__ = ~new_new_n4722__ & ~new_new_n4724__;
  assign new_new_n4727__ = ~new_new_n4725__ & ~new_new_n4726__;
  assign new_new_n4728__ = new_new_n4654__ & new_new_n4727__;
  assign new_new_n4729__ = ~new_new_n4654__ & ~new_new_n4727__;
  assign new_new_n4730__ = ~new_new_n4728__ & ~new_new_n4729__;
  assign new_new_n4731__ = new_new_n4582__ & new_new_n4730__;
  assign new_new_n4732__ = ~new_new_n4582__ & ~new_new_n4730__;
  assign new_new_n4733__ = ~new_new_n4731__ & ~new_new_n4732__;
  assign new_new_n4734__ = ~new_new_n4362__ & ~new_new_n4372__;
  assign new_new_n4735__ = ~new_new_n4556__ & new_new_n4734__;
  assign new_new_n4736__ = new_new_n4362__ & ~new_new_n4365__;
  assign new_new_n4737__ = ~new_new_n4553__ & ~new_new_n4736__;
  assign new_new_n4738__ = ~new_new_n4576__ & ~new_new_n4737__;
  assign new_new_n4739__ = ~new_new_n4195__ & ~new_new_n4738__;
  assign new_new_n4740__ = ~new_new_n4554__ & ~new_new_n4739__;
  assign new_new_n4741__ = ~new_new_n4735__ & new_new_n4740__;
  assign new_new_n4742__ = ~new_new_n4503__ & ~new_new_n4550__;
  assign new_new_n4743__ = ~new_new_n4504__ & ~new_new_n4742__;
  assign new_new_n4744__ = new_new_n4741__ & ~new_new_n4743__;
  assign new_new_n4745__ = ~new_new_n4741__ & new_new_n4743__;
  assign new_new_n4746__ = ~new_new_n4744__ & ~new_new_n4745__;
  assign new_new_n4747__ = ~new_new_n4389__ & ~new_new_n4417__;
  assign new_new_n4748__ = ~new_new_n4390__ & ~new_new_n4747__;
  assign new_new_n4749__ = ~new_new_n4410__ & new_new_n4414__;
  assign new_new_n4750__ = ~new_new_n4411__ & ~new_new_n4749__;
  assign new_new_n4751__ = ~new_new_n4482__ & ~new_new_n4493__;
  assign new_new_n4752__ = ~new_new_n4483__ & ~new_new_n4751__;
  assign new_new_n4753__ = ~new_new_n4512__ & ~new_new_n4518__;
  assign new_new_n4754__ = ~new_new_n4752__ & new_new_n4753__;
  assign new_new_n4755__ = new_new_n4752__ & ~new_new_n4753__;
  assign new_new_n4756__ = ~new_new_n4754__ & ~new_new_n4755__;
  assign new_new_n4757__ = new_new_n4750__ & new_new_n4756__;
  assign new_new_n4758__ = ~new_new_n4750__ & ~new_new_n4756__;
  assign new_new_n4759__ = ~new_new_n4757__ & ~new_new_n4758__;
  assign new_new_n4760__ = ~new_new_n4748__ & ~new_new_n4759__;
  assign new_new_n4761__ = new_new_n4748__ & new_new_n4759__;
  assign new_new_n4762__ = ~new_new_n4760__ & ~new_new_n4761__;
  assign new_new_n4763__ = ~new_new_n4462__ & ~new_new_n4496__;
  assign new_new_n4764__ = ~new_new_n4461__ & ~new_new_n4763__;
  assign new_new_n4765__ = new_new_n4762__ & ~new_new_n4764__;
  assign new_new_n4766__ = ~new_new_n4762__ & new_new_n4764__;
  assign new_new_n4767__ = ~new_new_n4765__ & ~new_new_n4766__;
  assign new_new_n4768__ = new_new_n4746__ & ~new_new_n4767__;
  assign new_new_n4769__ = ~new_new_n4746__ & new_new_n4767__;
  assign new_new_n4770__ = ~new_new_n4768__ & ~new_new_n4769__;
  assign new_new_n4771__ = new_new_n4733__ & new_new_n4770__;
  assign new_new_n4772__ = ~new_new_n4733__ & ~new_new_n4770__;
  assign po043 = new_new_n4771__ | new_new_n4772__;
  assign new_new_n4774__ = ~new_new_n4653__ & ~new_new_n4727__;
  assign new_new_n4775__ = ~new_new_n4652__ & ~new_new_n4774__;
  assign new_new_n4776__ = ~new_new_n4761__ & new_new_n4764__;
  assign new_new_n4777__ = ~new_new_n4760__ & ~new_new_n4776__;
  assign new_new_n4778__ = ~new_new_n4750__ & ~new_new_n4755__;
  assign new_new_n4779__ = ~new_new_n4754__ & ~new_new_n4778__;
  assign new_new_n4780__ = pi13 & pi30;
  assign new_new_n4781__ = pi05 & pi38;
  assign new_new_n4782__ = pi02 & pi41;
  assign new_new_n4783__ = ~new_new_n4781__ & ~new_new_n4782__;
  assign new_new_n4784__ = new_new_n4781__ & new_new_n4782__;
  assign new_new_n4785__ = ~new_new_n4783__ & ~new_new_n4784__;
  assign new_new_n4786__ = new_new_n4780__ & ~new_new_n4785__;
  assign new_new_n4787__ = ~new_new_n4780__ & new_new_n4785__;
  assign new_new_n4788__ = ~new_new_n4786__ & ~new_new_n4787__;
  assign new_new_n4789__ = pi21 & pi22;
  assign new_new_n4790__ = pi09 & pi34;
  assign new_new_n4791__ = pi20 & pi23;
  assign new_new_n4792__ = ~new_new_n4790__ & ~new_new_n4791__;
  assign new_new_n4793__ = new_new_n4790__ & new_new_n4791__;
  assign new_new_n4794__ = ~new_new_n4792__ & ~new_new_n4793__;
  assign new_new_n4795__ = new_new_n4789__ & ~new_new_n4794__;
  assign new_new_n4796__ = ~new_new_n4789__ & new_new_n4794__;
  assign new_new_n4797__ = ~new_new_n4795__ & ~new_new_n4796__;
  assign new_new_n4798__ = new_new_n4788__ & new_new_n4797__;
  assign new_new_n4799__ = ~new_new_n4788__ & ~new_new_n4797__;
  assign new_new_n4800__ = ~new_new_n4798__ & ~new_new_n4799__;
  assign new_new_n4801__ = pi10 & pi33;
  assign new_new_n4802__ = pi07 & pi36;
  assign new_new_n4803__ = pi08 & pi35;
  assign new_new_n4804__ = ~new_new_n4802__ & ~new_new_n4803__;
  assign new_new_n4805__ = new_new_n4802__ & new_new_n4803__;
  assign new_new_n4806__ = ~new_new_n4804__ & ~new_new_n4805__;
  assign new_new_n4807__ = new_new_n4801__ & ~new_new_n4806__;
  assign new_new_n4808__ = ~new_new_n4801__ & new_new_n4806__;
  assign new_new_n4809__ = ~new_new_n4807__ & ~new_new_n4808__;
  assign new_new_n4810__ = new_new_n4800__ & ~new_new_n4809__;
  assign new_new_n4811__ = ~new_new_n4800__ & new_new_n4809__;
  assign new_new_n4812__ = ~new_new_n4810__ & ~new_new_n4811__;
  assign new_new_n4813__ = ~new_new_n4779__ & new_new_n4812__;
  assign new_new_n4814__ = new_new_n4779__ & ~new_new_n4812__;
  assign new_new_n4815__ = ~new_new_n4813__ & ~new_new_n4814__;
  assign new_new_n4816__ = pi19 & pi24;
  assign new_new_n4817__ = pi18 & pi25;
  assign new_new_n4818__ = pi17 & pi26;
  assign new_new_n4819__ = ~new_new_n4817__ & ~new_new_n4818__;
  assign new_new_n4820__ = new_new_n4817__ & new_new_n4818__;
  assign new_new_n4821__ = ~new_new_n4819__ & ~new_new_n4820__;
  assign new_new_n4822__ = new_new_n4816__ & ~new_new_n4821__;
  assign new_new_n4823__ = ~new_new_n4816__ & new_new_n4821__;
  assign new_new_n4824__ = ~new_new_n4822__ & ~new_new_n4823__;
  assign new_new_n4825__ = pi04 & pi39;
  assign new_new_n4826__ = pi03 & pi40;
  assign new_new_n4827__ = pi00 & pi43;
  assign new_new_n4828__ = ~new_new_n4826__ & ~new_new_n4827__;
  assign new_new_n4829__ = new_new_n4826__ & new_new_n4827__;
  assign new_new_n4830__ = ~new_new_n4828__ & ~new_new_n4829__;
  assign new_new_n4831__ = new_new_n4825__ & ~new_new_n4830__;
  assign new_new_n4832__ = ~new_new_n4825__ & new_new_n4830__;
  assign new_new_n4833__ = ~new_new_n4831__ & ~new_new_n4832__;
  assign new_new_n4834__ = new_new_n4824__ & new_new_n4833__;
  assign new_new_n4835__ = ~new_new_n4824__ & ~new_new_n4833__;
  assign new_new_n4836__ = ~new_new_n4834__ & ~new_new_n4835__;
  assign new_new_n4837__ = pi16 & pi27;
  assign new_new_n4838__ = pi15 & pi28;
  assign new_new_n4839__ = ~new_new_n2730__ & ~new_new_n4838__;
  assign new_new_n4840__ = new_new_n2730__ & new_new_n4838__;
  assign new_new_n4841__ = ~new_new_n4839__ & ~new_new_n4840__;
  assign new_new_n4842__ = new_new_n4837__ & ~new_new_n4841__;
  assign new_new_n4843__ = ~new_new_n4837__ & new_new_n4841__;
  assign new_new_n4844__ = ~new_new_n4842__ & ~new_new_n4843__;
  assign new_new_n4845__ = new_new_n4836__ & ~new_new_n4844__;
  assign new_new_n4846__ = ~new_new_n4836__ & new_new_n4844__;
  assign new_new_n4847__ = ~new_new_n4845__ & ~new_new_n4846__;
  assign new_new_n4848__ = new_new_n4815__ & ~new_new_n4847__;
  assign new_new_n4849__ = ~new_new_n4815__ & new_new_n4847__;
  assign new_new_n4850__ = ~new_new_n4848__ & ~new_new_n4849__;
  assign new_new_n4851__ = ~new_new_n4777__ & ~new_new_n4850__;
  assign new_new_n4852__ = new_new_n4777__ & new_new_n4850__;
  assign new_new_n4853__ = ~new_new_n4851__ & ~new_new_n4852__;
  assign new_new_n4854__ = ~new_new_n4660__ & ~new_new_n4665__;
  assign new_new_n4855__ = ~new_new_n4673__ & ~new_new_n4678__;
  assign new_new_n4856__ = ~new_new_n4672__ & ~new_new_n4855__;
  assign new_new_n4857__ = pi12 & pi31;
  assign new_new_n4858__ = pi11 & pi32;
  assign new_new_n4859__ = pi06 & pi37;
  assign new_new_n4860__ = ~new_new_n4858__ & ~new_new_n4859__;
  assign new_new_n4861__ = new_new_n4858__ & new_new_n4859__;
  assign new_new_n4862__ = ~new_new_n4860__ & ~new_new_n4861__;
  assign new_new_n4863__ = new_new_n4857__ & ~new_new_n4862__;
  assign new_new_n4864__ = ~new_new_n4857__ & new_new_n4862__;
  assign new_new_n4865__ = ~new_new_n4863__ & ~new_new_n4864__;
  assign new_new_n4866__ = ~new_new_n4856__ & new_new_n4865__;
  assign new_new_n4867__ = new_new_n4856__ & ~new_new_n4865__;
  assign new_new_n4868__ = ~new_new_n4866__ & ~new_new_n4867__;
  assign new_new_n4869__ = new_new_n4854__ & ~new_new_n4868__;
  assign new_new_n4870__ = ~new_new_n4854__ & new_new_n4868__;
  assign new_new_n4871__ = ~new_new_n4869__ & ~new_new_n4870__;
  assign new_new_n4872__ = ~new_new_n4690__ & ~new_new_n4694__;
  assign new_new_n4873__ = ~new_new_n4693__ & ~new_new_n4872__;
  assign new_new_n4874__ = ~pi41 & new_new_n4700__;
  assign new_new_n4875__ = ~new_new_n4699__ & ~new_new_n4874__;
  assign new_new_n4876__ = new_new_n4701__ & ~new_new_n4875__;
  assign new_new_n4877__ = ~new_new_n4699__ & ~new_new_n4701__;
  assign new_new_n4878__ = pi41 & ~new_new_n4700__;
  assign new_new_n4879__ = ~new_new_n4877__ & new_new_n4878__;
  assign new_new_n4880__ = ~new_new_n4876__ & ~new_new_n4879__;
  assign new_new_n4881__ = pi01 & ~new_new_n4880__;
  assign new_new_n4882__ = pi20 & pi42;
  assign new_new_n4883__ = pi01 & pi41;
  assign new_new_n4884__ = new_new_n1474__ & new_new_n4882__;
  assign new_new_n4885__ = ~new_new_n4883__ & new_new_n4884__;
  assign new_new_n4886__ = ~new_new_n4881__ & ~new_new_n4885__;
  assign new_new_n4887__ = ~new_new_n4873__ & new_new_n4886__;
  assign new_new_n4888__ = new_new_n4873__ & ~new_new_n4886__;
  assign new_new_n4889__ = ~new_new_n4887__ & ~new_new_n4888__;
  assign new_new_n4890__ = ~new_new_n4634__ & ~new_new_n4638__;
  assign new_new_n4891__ = ~new_new_n4637__ & ~new_new_n4890__;
  assign new_new_n4892__ = new_new_n4889__ & ~new_new_n4891__;
  assign new_new_n4893__ = ~new_new_n4889__ & new_new_n4891__;
  assign new_new_n4894__ = ~new_new_n4892__ & ~new_new_n4893__;
  assign new_new_n4895__ = ~new_new_n4712__ & ~new_new_n4716__;
  assign new_new_n4896__ = ~new_new_n4713__ & ~new_new_n4895__;
  assign new_new_n4897__ = ~new_new_n4894__ & ~new_new_n4896__;
  assign new_new_n4898__ = new_new_n4894__ & new_new_n4896__;
  assign new_new_n4899__ = ~new_new_n4897__ & ~new_new_n4898__;
  assign new_new_n4900__ = ~new_new_n4622__ & ~new_new_n4626__;
  assign new_new_n4901__ = ~new_new_n4625__ & ~new_new_n4900__;
  assign new_new_n4902__ = ~new_new_n4613__ & ~new_new_n4617__;
  assign new_new_n4903__ = ~new_new_n4616__ & ~new_new_n4902__;
  assign new_new_n4904__ = ~new_new_n4601__ & ~new_new_n4605__;
  assign new_new_n4905__ = ~new_new_n4604__ & ~new_new_n4904__;
  assign new_new_n4906__ = new_new_n4903__ & new_new_n4905__;
  assign new_new_n4907__ = ~new_new_n4903__ & ~new_new_n4905__;
  assign new_new_n4908__ = ~new_new_n4901__ & ~new_new_n4906__;
  assign new_new_n4909__ = ~new_new_n4907__ & ~new_new_n4908__;
  assign new_new_n4910__ = ~new_new_n4906__ & new_new_n4909__;
  assign new_new_n4911__ = new_new_n4901__ & ~new_new_n4910__;
  assign new_new_n4912__ = ~new_new_n4907__ & new_new_n4908__;
  assign new_new_n4913__ = ~new_new_n4911__ & ~new_new_n4912__;
  assign new_new_n4914__ = new_new_n4899__ & ~new_new_n4913__;
  assign new_new_n4915__ = ~new_new_n4899__ & new_new_n4913__;
  assign new_new_n4916__ = ~new_new_n4914__ & ~new_new_n4915__;
  assign new_new_n4917__ = new_new_n4871__ & ~new_new_n4916__;
  assign new_new_n4918__ = ~new_new_n4871__ & new_new_n4916__;
  assign new_new_n4919__ = ~new_new_n4917__ & ~new_new_n4918__;
  assign new_new_n4920__ = new_new_n4667__ & ~new_new_n4685__;
  assign new_new_n4921__ = ~new_new_n4684__ & ~new_new_n4920__;
  assign new_new_n4922__ = new_new_n4919__ & new_new_n4921__;
  assign new_new_n4923__ = ~new_new_n4919__ & ~new_new_n4921__;
  assign new_new_n4924__ = ~new_new_n4922__ & ~new_new_n4923__;
  assign new_new_n4925__ = new_new_n4853__ & ~new_new_n4924__;
  assign new_new_n4926__ = ~new_new_n4853__ & new_new_n4924__;
  assign new_new_n4927__ = ~new_new_n4925__ & ~new_new_n4926__;
  assign new_new_n4928__ = ~new_new_n4775__ & ~new_new_n4927__;
  assign new_new_n4929__ = new_new_n4775__ & new_new_n4927__;
  assign new_new_n4930__ = ~new_new_n4928__ & ~new_new_n4929__;
  assign new_new_n4931__ = ~new_new_n4720__ & new_new_n4724__;
  assign new_new_n4932__ = ~new_new_n4721__ & ~new_new_n4931__;
  assign new_new_n4933__ = new_new_n4586__ & new_new_n4612__;
  assign new_new_n4934__ = ~new_new_n4586__ & ~new_new_n4612__;
  assign new_new_n4935__ = ~new_new_n4645__ & ~new_new_n4934__;
  assign new_new_n4936__ = ~new_new_n4933__ & ~new_new_n4935__;
  assign new_new_n4937__ = ~new_new_n4932__ & ~new_new_n4936__;
  assign new_new_n4938__ = new_new_n4932__ & new_new_n4936__;
  assign new_new_n4939__ = ~new_new_n4937__ & ~new_new_n4938__;
  assign new_new_n4940__ = ~new_new_n4631__ & ~new_new_n4642__;
  assign new_new_n4941__ = ~new_new_n4632__ & ~new_new_n4940__;
  assign new_new_n4942__ = ~new_new_n4589__ & ~new_new_n4593__;
  assign new_new_n4943__ = ~new_new_n4592__ & ~new_new_n4942__;
  assign new_new_n4944__ = pi22 & pi42;
  assign new_new_n4945__ = ~new_new_n4943__ & ~new_new_n4944__;
  assign new_new_n4946__ = pi20 & pi41;
  assign new_new_n4947__ = pi01 & ~pi42;
  assign new_new_n4948__ = new_new_n4943__ & ~new_new_n4947__;
  assign new_new_n4949__ = ~new_new_n4945__ & new_new_n4946__;
  assign new_new_n4950__ = ~new_new_n4948__ & new_new_n4949__;
  assign new_new_n4951__ = new_new_n4700__ & new_new_n4883__;
  assign new_new_n4952__ = pi01 & pi42;
  assign new_new_n4953__ = ~new_new_n4943__ & new_new_n4952__;
  assign new_new_n4954__ = new_new_n4943__ & ~new_new_n4952__;
  assign new_new_n4955__ = ~new_new_n4953__ & ~new_new_n4954__;
  assign new_new_n4956__ = pi22 & ~new_new_n4955__;
  assign new_new_n4957__ = ~pi22 & new_new_n4955__;
  assign new_new_n4958__ = ~new_new_n4951__ & ~new_new_n4956__;
  assign new_new_n4959__ = ~new_new_n4957__ & new_new_n4958__;
  assign new_new_n4960__ = ~new_new_n4950__ & ~new_new_n4959__;
  assign new_new_n4961__ = ~new_new_n4598__ & ~new_new_n4609__;
  assign new_new_n4962__ = ~new_new_n4599__ & ~new_new_n4961__;
  assign new_new_n4963__ = ~new_new_n4960__ & ~new_new_n4962__;
  assign new_new_n4964__ = new_new_n4960__ & new_new_n4962__;
  assign new_new_n4965__ = ~new_new_n4963__ & ~new_new_n4964__;
  assign new_new_n4966__ = ~new_new_n4941__ & new_new_n4965__;
  assign new_new_n4967__ = new_new_n4941__ & ~new_new_n4965__;
  assign new_new_n4968__ = ~new_new_n4966__ & ~new_new_n4967__;
  assign new_new_n4969__ = new_new_n4939__ & new_new_n4968__;
  assign new_new_n4970__ = ~new_new_n4939__ & ~new_new_n4968__;
  assign new_new_n4971__ = ~new_new_n4969__ & ~new_new_n4970__;
  assign new_new_n4972__ = new_new_n4930__ & ~new_new_n4971__;
  assign new_new_n4973__ = ~new_new_n4930__ & new_new_n4971__;
  assign new_new_n4974__ = ~new_new_n4972__ & ~new_new_n4973__;
  assign new_new_n4975__ = new_new_n4582__ & ~new_new_n4767__;
  assign new_new_n4976__ = ~new_new_n4582__ & new_new_n4767__;
  assign new_new_n4977__ = ~new_new_n4730__ & ~new_new_n4976__;
  assign new_new_n4978__ = ~new_new_n4975__ & ~new_new_n4977__;
  assign new_new_n4979__ = new_new_n4744__ & new_new_n4978__;
  assign new_new_n4980__ = ~new_new_n4975__ & ~new_new_n4976__;
  assign new_new_n4981__ = new_new_n4733__ & ~new_new_n4980__;
  assign new_new_n4982__ = new_new_n4746__ & ~new_new_n4981__;
  assign new_new_n4983__ = new_new_n4745__ & ~new_new_n4978__;
  assign new_new_n4984__ = new_new_n4974__ & ~new_new_n4979__;
  assign new_new_n4985__ = ~new_new_n4983__ & new_new_n4984__;
  assign new_new_n4986__ = ~new_new_n4982__ & new_new_n4985__;
  assign new_new_n4987__ = new_new_n4745__ & ~new_new_n4975__;
  assign new_new_n4988__ = ~new_new_n4744__ & new_new_n4976__;
  assign new_new_n4989__ = ~new_new_n4987__ & ~new_new_n4988__;
  assign new_new_n4990__ = new_new_n4730__ & ~new_new_n4989__;
  assign new_new_n4991__ = ~new_new_n4745__ & ~new_new_n4975__;
  assign new_new_n4992__ = ~new_new_n4744__ & ~new_new_n4976__;
  assign new_new_n4993__ = ~new_new_n4991__ & ~new_new_n4992__;
  assign new_new_n4994__ = new_new_n4582__ & ~new_new_n4745__;
  assign new_new_n4995__ = new_new_n4744__ & new_new_n4994__;
  assign new_new_n4996__ = new_new_n4767__ & ~new_new_n4995__;
  assign new_new_n4997__ = ~new_new_n4744__ & ~new_new_n4994__;
  assign new_new_n4998__ = ~new_new_n4730__ & ~new_new_n4997__;
  assign new_new_n4999__ = ~new_new_n4996__ & new_new_n4998__;
  assign new_new_n5000__ = ~new_new_n4974__ & ~new_new_n4993__;
  assign new_new_n5001__ = ~new_new_n4990__ & new_new_n5000__;
  assign new_new_n5002__ = ~new_new_n4999__ & new_new_n5001__;
  assign po044 = ~new_new_n4986__ & ~new_new_n5002__;
  assign new_new_n5004__ = ~new_new_n4813__ & ~new_new_n4847__;
  assign new_new_n5005__ = ~new_new_n4814__ & ~new_new_n5004__;
  assign new_new_n5006__ = ~new_new_n4834__ & ~new_new_n4844__;
  assign new_new_n5007__ = ~new_new_n4835__ & ~new_new_n5006__;
  assign new_new_n5008__ = ~new_new_n4798__ & ~new_new_n4809__;
  assign new_new_n5009__ = ~new_new_n4799__ & ~new_new_n5008__;
  assign new_new_n5010__ = new_new_n5007__ & new_new_n5009__;
  assign new_new_n5011__ = ~new_new_n5007__ & ~new_new_n5009__;
  assign new_new_n5012__ = ~new_new_n5010__ & ~new_new_n5011__;
  assign new_new_n5013__ = ~new_new_n4825__ & ~new_new_n4829__;
  assign new_new_n5014__ = ~new_new_n4828__ & ~new_new_n5013__;
  assign new_new_n5015__ = ~new_new_n4780__ & ~new_new_n4784__;
  assign new_new_n5016__ = ~new_new_n4783__ & ~new_new_n5015__;
  assign new_new_n5017__ = ~new_new_n4816__ & ~new_new_n4820__;
  assign new_new_n5018__ = ~new_new_n4819__ & ~new_new_n5017__;
  assign new_new_n5019__ = new_new_n5016__ & new_new_n5018__;
  assign new_new_n5020__ = ~new_new_n5016__ & ~new_new_n5018__;
  assign new_new_n5021__ = ~new_new_n5019__ & ~new_new_n5020__;
  assign new_new_n5022__ = new_new_n5014__ & ~new_new_n5021__;
  assign new_new_n5023__ = ~new_new_n5014__ & new_new_n5021__;
  assign new_new_n5024__ = ~new_new_n5022__ & ~new_new_n5023__;
  assign new_new_n5025__ = new_new_n5012__ & ~new_new_n5024__;
  assign new_new_n5026__ = ~new_new_n5012__ & new_new_n5024__;
  assign new_new_n5027__ = ~new_new_n5025__ & ~new_new_n5026__;
  assign new_new_n5028__ = new_new_n5005__ & new_new_n5027__;
  assign new_new_n5029__ = ~new_new_n5005__ & ~new_new_n5027__;
  assign new_new_n5030__ = ~new_new_n5028__ & ~new_new_n5029__;
  assign new_new_n5031__ = ~new_new_n4918__ & ~new_new_n4921__;
  assign new_new_n5032__ = ~new_new_n4917__ & ~new_new_n5031__;
  assign new_new_n5033__ = new_new_n5030__ & ~new_new_n5032__;
  assign new_new_n5034__ = ~new_new_n5030__ & new_new_n5032__;
  assign new_new_n5035__ = ~new_new_n5033__ & ~new_new_n5034__;
  assign new_new_n5036__ = ~new_new_n4852__ & new_new_n4924__;
  assign new_new_n5037__ = ~new_new_n4851__ & ~new_new_n5036__;
  assign new_new_n5038__ = ~new_new_n4898__ & ~new_new_n4913__;
  assign new_new_n5039__ = ~new_new_n4897__ & ~new_new_n5038__;
  assign new_new_n5040__ = ~new_new_n4943__ & ~new_new_n4947__;
  assign new_new_n5041__ = new_new_n4946__ & ~new_new_n5040__;
  assign new_new_n5042__ = ~new_new_n4954__ & ~new_new_n5041__;
  assign new_new_n5043__ = pi22 & ~new_new_n5042__;
  assign new_new_n5044__ = ~pi22 & new_new_n4952__;
  assign new_new_n5045__ = new_new_n4943__ & new_new_n5044__;
  assign new_new_n5046__ = ~new_new_n5043__ & ~new_new_n5045__;
  assign new_new_n5047__ = new_new_n4909__ & ~new_new_n5046__;
  assign new_new_n5048__ = ~new_new_n4909__ & new_new_n5046__;
  assign new_new_n5049__ = ~new_new_n5047__ & ~new_new_n5048__;
  assign new_new_n5050__ = ~new_new_n4887__ & new_new_n4891__;
  assign new_new_n5051__ = ~new_new_n4888__ & ~new_new_n5050__;
  assign new_new_n5052__ = new_new_n5049__ & new_new_n5051__;
  assign new_new_n5053__ = ~new_new_n5049__ & ~new_new_n5051__;
  assign new_new_n5054__ = ~new_new_n5052__ & ~new_new_n5053__;
  assign new_new_n5055__ = ~new_new_n5039__ & ~new_new_n5054__;
  assign new_new_n5056__ = new_new_n5039__ & new_new_n5054__;
  assign new_new_n5057__ = ~new_new_n5055__ & ~new_new_n5056__;
  assign new_new_n5058__ = new_new_n4854__ & ~new_new_n4866__;
  assign new_new_n5059__ = ~new_new_n4867__ & ~new_new_n5058__;
  assign new_new_n5060__ = ~new_new_n4789__ & ~new_new_n4793__;
  assign new_new_n5061__ = ~new_new_n4792__ & ~new_new_n5060__;
  assign new_new_n5062__ = ~new_new_n4801__ & ~new_new_n4805__;
  assign new_new_n5063__ = ~new_new_n4804__ & ~new_new_n5062__;
  assign new_new_n5064__ = ~new_new_n5061__ & ~new_new_n5063__;
  assign new_new_n5065__ = new_new_n5061__ & new_new_n5063__;
  assign new_new_n5066__ = ~new_new_n5064__ & ~new_new_n5065__;
  assign new_new_n5067__ = pi01 & pi43;
  assign new_new_n5068__ = pi21 & pi23;
  assign new_new_n5069__ = new_new_n5067__ & ~new_new_n5068__;
  assign new_new_n5070__ = ~new_new_n5067__ & new_new_n5068__;
  assign new_new_n5071__ = ~new_new_n5069__ & ~new_new_n5070__;
  assign new_new_n5072__ = new_new_n5066__ & new_new_n5071__;
  assign new_new_n5073__ = ~new_new_n5066__ & ~new_new_n5071__;
  assign new_new_n5074__ = ~new_new_n5072__ & ~new_new_n5073__;
  assign new_new_n5075__ = ~new_new_n5059__ & ~new_new_n5074__;
  assign new_new_n5076__ = new_new_n5059__ & new_new_n5074__;
  assign new_new_n5077__ = ~new_new_n5075__ & ~new_new_n5076__;
  assign new_new_n5078__ = ~new_new_n4837__ & ~new_new_n4840__;
  assign new_new_n5079__ = ~new_new_n4839__ & ~new_new_n5078__;
  assign new_new_n5080__ = ~new_new_n4857__ & ~new_new_n4861__;
  assign new_new_n5081__ = ~new_new_n4860__ & ~new_new_n5080__;
  assign new_new_n5082__ = ~new_new_n5079__ & ~new_new_n5081__;
  assign new_new_n5083__ = new_new_n5079__ & new_new_n5081__;
  assign new_new_n5084__ = ~new_new_n5082__ & ~new_new_n5083__;
  assign new_new_n5085__ = pi00 & pi44;
  assign new_new_n5086__ = pi02 & new_new_n1535__;
  assign new_new_n5087__ = ~pi02 & ~new_new_n1535__;
  assign new_new_n5088__ = pi42 & ~new_new_n5087__;
  assign new_new_n5089__ = ~new_new_n5086__ & new_new_n5088__;
  assign new_new_n5090__ = new_new_n5085__ & ~new_new_n5089__;
  assign new_new_n5091__ = ~new_new_n5085__ & new_new_n5089__;
  assign new_new_n5092__ = ~new_new_n5090__ & ~new_new_n5091__;
  assign new_new_n5093__ = new_new_n5084__ & ~new_new_n5092__;
  assign new_new_n5094__ = ~new_new_n5084__ & new_new_n5092__;
  assign new_new_n5095__ = ~new_new_n5093__ & ~new_new_n5094__;
  assign new_new_n5096__ = new_new_n5077__ & ~new_new_n5095__;
  assign new_new_n5097__ = ~new_new_n5077__ & new_new_n5095__;
  assign new_new_n5098__ = ~new_new_n5096__ & ~new_new_n5097__;
  assign new_new_n5099__ = new_new_n5057__ & ~new_new_n5098__;
  assign new_new_n5100__ = ~new_new_n5057__ & new_new_n5098__;
  assign new_new_n5101__ = ~new_new_n5099__ & ~new_new_n5100__;
  assign new_new_n5102__ = ~new_new_n4963__ & ~new_new_n4966__;
  assign new_new_n5103__ = pi16 & pi28;
  assign new_new_n5104__ = pi14 & pi30;
  assign new_new_n5105__ = pi04 & pi40;
  assign new_new_n5106__ = ~new_new_n5104__ & ~new_new_n5105__;
  assign new_new_n5107__ = new_new_n5104__ & new_new_n5105__;
  assign new_new_n5108__ = ~new_new_n5106__ & ~new_new_n5107__;
  assign new_new_n5109__ = new_new_n5103__ & ~new_new_n5108__;
  assign new_new_n5110__ = ~new_new_n5103__ & new_new_n5108__;
  assign new_new_n5111__ = ~new_new_n5109__ & ~new_new_n5110__;
  assign new_new_n5112__ = pi10 & pi34;
  assign new_new_n5113__ = pi08 & pi36;
  assign new_new_n5114__ = pi09 & pi35;
  assign new_new_n5115__ = ~new_new_n5113__ & ~new_new_n5114__;
  assign new_new_n5116__ = new_new_n5113__ & new_new_n5114__;
  assign new_new_n5117__ = ~new_new_n5115__ & ~new_new_n5116__;
  assign new_new_n5118__ = new_new_n5112__ & ~new_new_n5117__;
  assign new_new_n5119__ = ~new_new_n5112__ & new_new_n5117__;
  assign new_new_n5120__ = ~new_new_n5118__ & ~new_new_n5119__;
  assign new_new_n5121__ = new_new_n5111__ & new_new_n5120__;
  assign new_new_n5122__ = ~new_new_n5111__ & ~new_new_n5120__;
  assign new_new_n5123__ = ~new_new_n5121__ & ~new_new_n5122__;
  assign new_new_n5124__ = pi13 & pi31;
  assign new_new_n5125__ = pi12 & pi32;
  assign new_new_n5126__ = pi05 & pi39;
  assign new_new_n5127__ = ~new_new_n5125__ & ~new_new_n5126__;
  assign new_new_n5128__ = new_new_n5125__ & new_new_n5126__;
  assign new_new_n5129__ = ~new_new_n5127__ & ~new_new_n5128__;
  assign new_new_n5130__ = new_new_n5124__ & ~new_new_n5129__;
  assign new_new_n5131__ = ~new_new_n5124__ & new_new_n5129__;
  assign new_new_n5132__ = ~new_new_n5130__ & ~new_new_n5131__;
  assign new_new_n5133__ = new_new_n5123__ & ~new_new_n5132__;
  assign new_new_n5134__ = ~new_new_n5123__ & new_new_n5132__;
  assign new_new_n5135__ = ~new_new_n5133__ & ~new_new_n5134__;
  assign new_new_n5136__ = new_new_n5102__ & ~new_new_n5135__;
  assign new_new_n5137__ = ~new_new_n5102__ & new_new_n5135__;
  assign new_new_n5138__ = ~new_new_n5136__ & ~new_new_n5137__;
  assign new_new_n5139__ = pi11 & pi33;
  assign new_new_n5140__ = pi07 & pi37;
  assign new_new_n5141__ = pi06 & pi38;
  assign new_new_n5142__ = ~new_new_n5140__ & ~new_new_n5141__;
  assign new_new_n5143__ = new_new_n5140__ & new_new_n5141__;
  assign new_new_n5144__ = ~new_new_n5142__ & ~new_new_n5143__;
  assign new_new_n5145__ = new_new_n5139__ & ~new_new_n5144__;
  assign new_new_n5146__ = ~new_new_n5139__ & new_new_n5144__;
  assign new_new_n5147__ = ~new_new_n5145__ & ~new_new_n5146__;
  assign new_new_n5148__ = pi20 & pi24;
  assign new_new_n5149__ = pi18 & pi26;
  assign new_new_n5150__ = pi19 & pi25;
  assign new_new_n5151__ = ~new_new_n5149__ & ~new_new_n5150__;
  assign new_new_n5152__ = new_new_n5149__ & new_new_n5150__;
  assign new_new_n5153__ = ~new_new_n5151__ & ~new_new_n5152__;
  assign new_new_n5154__ = new_new_n5148__ & ~new_new_n5153__;
  assign new_new_n5155__ = ~new_new_n5148__ & new_new_n5153__;
  assign new_new_n5156__ = ~new_new_n5154__ & ~new_new_n5155__;
  assign new_new_n5157__ = new_new_n5147__ & new_new_n5156__;
  assign new_new_n5158__ = ~new_new_n5147__ & ~new_new_n5156__;
  assign new_new_n5159__ = ~new_new_n5157__ & ~new_new_n5158__;
  assign new_new_n5160__ = pi17 & pi27;
  assign new_new_n5161__ = pi15 & pi29;
  assign new_new_n5162__ = pi03 & pi41;
  assign new_new_n5163__ = ~new_new_n5161__ & ~new_new_n5162__;
  assign new_new_n5164__ = new_new_n5161__ & new_new_n5162__;
  assign new_new_n5165__ = ~new_new_n5163__ & ~new_new_n5164__;
  assign new_new_n5166__ = new_new_n5160__ & ~new_new_n5165__;
  assign new_new_n5167__ = ~new_new_n5160__ & new_new_n5165__;
  assign new_new_n5168__ = ~new_new_n5166__ & ~new_new_n5167__;
  assign new_new_n5169__ = ~new_new_n5159__ & new_new_n5168__;
  assign new_new_n5170__ = new_new_n5159__ & ~new_new_n5168__;
  assign new_new_n5171__ = ~new_new_n5169__ & ~new_new_n5170__;
  assign new_new_n5172__ = new_new_n5138__ & new_new_n5171__;
  assign new_new_n5173__ = ~new_new_n5138__ & ~new_new_n5171__;
  assign new_new_n5174__ = ~new_new_n5172__ & ~new_new_n5173__;
  assign new_new_n5175__ = ~new_new_n5101__ & ~new_new_n5174__;
  assign new_new_n5176__ = new_new_n5101__ & new_new_n5174__;
  assign new_new_n5177__ = ~new_new_n5175__ & ~new_new_n5176__;
  assign new_new_n5178__ = ~new_new_n4938__ & ~new_new_n4968__;
  assign new_new_n5179__ = ~new_new_n4937__ & ~new_new_n5178__;
  assign new_new_n5180__ = new_new_n5177__ & new_new_n5179__;
  assign new_new_n5181__ = ~new_new_n5177__ & ~new_new_n5179__;
  assign new_new_n5182__ = ~new_new_n5180__ & ~new_new_n5181__;
  assign new_new_n5183__ = ~new_new_n5037__ & new_new_n5182__;
  assign new_new_n5184__ = new_new_n5037__ & ~new_new_n5182__;
  assign new_new_n5185__ = ~new_new_n5183__ & ~new_new_n5184__;
  assign new_new_n5186__ = ~new_new_n4929__ & new_new_n4971__;
  assign new_new_n5187__ = ~new_new_n4928__ & ~new_new_n5186__;
  assign new_new_n5188__ = ~new_new_n4745__ & ~new_new_n4978__;
  assign new_new_n5189__ = new_new_n4974__ & ~new_new_n5188__;
  assign new_new_n5190__ = ~new_new_n4730__ & new_new_n4975__;
  assign new_new_n5191__ = new_new_n4974__ & ~new_new_n5190__;
  assign new_new_n5192__ = new_new_n4730__ & new_new_n4976__;
  assign new_new_n5193__ = ~new_new_n5191__ & ~new_new_n5192__;
  assign new_new_n5194__ = ~new_new_n4744__ & ~new_new_n5193__;
  assign new_new_n5195__ = new_new_n4745__ & new_new_n4978__;
  assign new_new_n5196__ = ~new_new_n5194__ & ~new_new_n5195__;
  assign new_new_n5197__ = ~new_new_n5189__ & new_new_n5196__;
  assign new_new_n5198__ = ~new_new_n5187__ & new_new_n5197__;
  assign new_new_n5199__ = new_new_n5187__ & ~new_new_n5197__;
  assign new_new_n5200__ = ~new_new_n5198__ & ~new_new_n5199__;
  assign new_new_n5201__ = new_new_n5185__ & ~new_new_n5200__;
  assign new_new_n5202__ = ~new_new_n5185__ & new_new_n5200__;
  assign new_new_n5203__ = ~new_new_n5201__ & ~new_new_n5202__;
  assign new_new_n5204__ = new_new_n5035__ & new_new_n5203__;
  assign new_new_n5205__ = ~new_new_n5035__ & ~new_new_n5203__;
  assign po045 = ~new_new_n5204__ & ~new_new_n5205__;
  assign new_new_n5207__ = ~new_new_n5037__ & new_new_n5197__;
  assign new_new_n5208__ = new_new_n5182__ & ~new_new_n5187__;
  assign new_new_n5209__ = new_new_n5207__ & new_new_n5208__;
  assign new_new_n5210__ = ~new_new_n5048__ & ~new_new_n5051__;
  assign new_new_n5211__ = ~new_new_n5047__ & ~new_new_n5210__;
  assign new_new_n5212__ = ~new_new_n5148__ & ~new_new_n5152__;
  assign new_new_n5213__ = ~new_new_n5151__ & ~new_new_n5212__;
  assign new_new_n5214__ = ~new_new_n5085__ & ~new_new_n5086__;
  assign new_new_n5215__ = new_new_n5088__ & ~new_new_n5214__;
  assign new_new_n5216__ = ~new_new_n5160__ & ~new_new_n5164__;
  assign new_new_n5217__ = ~new_new_n5163__ & ~new_new_n5216__;
  assign new_new_n5218__ = ~new_new_n5215__ & ~new_new_n5217__;
  assign new_new_n5219__ = new_new_n5215__ & new_new_n5217__;
  assign new_new_n5220__ = ~new_new_n5218__ & ~new_new_n5219__;
  assign new_new_n5221__ = new_new_n5213__ & ~new_new_n5220__;
  assign new_new_n5222__ = ~new_new_n5213__ & new_new_n5220__;
  assign new_new_n5223__ = ~new_new_n5221__ & ~new_new_n5222__;
  assign new_new_n5224__ = ~new_new_n5211__ & ~new_new_n5223__;
  assign new_new_n5225__ = new_new_n5211__ & new_new_n5223__;
  assign new_new_n5226__ = ~new_new_n5224__ & ~new_new_n5225__;
  assign new_new_n5227__ = pi12 & pi33;
  assign new_new_n5228__ = pi11 & pi34;
  assign new_new_n5229__ = pi06 & pi39;
  assign new_new_n5230__ = ~new_new_n5228__ & ~new_new_n5229__;
  assign new_new_n5231__ = new_new_n5228__ & new_new_n5229__;
  assign new_new_n5232__ = ~new_new_n5230__ & ~new_new_n5231__;
  assign new_new_n5233__ = new_new_n5227__ & ~new_new_n5232__;
  assign new_new_n5234__ = ~new_new_n5227__ & new_new_n5232__;
  assign new_new_n5235__ = ~new_new_n5233__ & ~new_new_n5234__;
  assign new_new_n5236__ = pi21 & pi43;
  assign new_new_n5237__ = pi01 & new_new_n5236__;
  assign new_new_n5238__ = pi23 & ~new_new_n5237__;
  assign new_new_n5239__ = pi03 & pi42;
  assign new_new_n5240__ = pi01 & pi44;
  assign new_new_n5241__ = new_new_n5239__ & ~new_new_n5240__;
  assign new_new_n5242__ = ~new_new_n5239__ & new_new_n5240__;
  assign new_new_n5243__ = ~new_new_n5241__ & ~new_new_n5242__;
  assign new_new_n5244__ = new_new_n5238__ & new_new_n5243__;
  assign new_new_n5245__ = ~new_new_n5238__ & ~new_new_n5243__;
  assign new_new_n5246__ = ~new_new_n5244__ & ~new_new_n5245__;
  assign new_new_n5247__ = ~new_new_n5235__ & ~new_new_n5246__;
  assign new_new_n5248__ = new_new_n5235__ & new_new_n5246__;
  assign new_new_n5249__ = ~new_new_n5247__ & ~new_new_n5248__;
  assign new_new_n5250__ = pi17 & pi28;
  assign new_new_n5251__ = pi16 & pi29;
  assign new_new_n5252__ = pi15 & pi30;
  assign new_new_n5253__ = ~new_new_n5251__ & ~new_new_n5252__;
  assign new_new_n5254__ = new_new_n5251__ & new_new_n5252__;
  assign new_new_n5255__ = ~new_new_n5253__ & ~new_new_n5254__;
  assign new_new_n5256__ = new_new_n5250__ & ~new_new_n5255__;
  assign new_new_n5257__ = ~new_new_n5250__ & new_new_n5255__;
  assign new_new_n5258__ = ~new_new_n5256__ & ~new_new_n5257__;
  assign new_new_n5259__ = new_new_n5249__ & ~new_new_n5258__;
  assign new_new_n5260__ = ~new_new_n5249__ & new_new_n5258__;
  assign new_new_n5261__ = ~new_new_n5259__ & ~new_new_n5260__;
  assign new_new_n5262__ = new_new_n5226__ & ~new_new_n5261__;
  assign new_new_n5263__ = ~new_new_n5226__ & new_new_n5261__;
  assign new_new_n5264__ = ~new_new_n5262__ & ~new_new_n5263__;
  assign new_new_n5265__ = ~new_new_n5137__ & ~new_new_n5171__;
  assign new_new_n5266__ = ~new_new_n5136__ & ~new_new_n5265__;
  assign new_new_n5267__ = new_new_n5264__ & ~new_new_n5266__;
  assign new_new_n5268__ = ~new_new_n5264__ & new_new_n5266__;
  assign new_new_n5269__ = ~new_new_n5267__ & ~new_new_n5268__;
  assign new_new_n5270__ = ~new_new_n5056__ & ~new_new_n5098__;
  assign new_new_n5271__ = ~new_new_n5055__ & ~new_new_n5270__;
  assign new_new_n5272__ = new_new_n5269__ & ~new_new_n5271__;
  assign new_new_n5273__ = ~new_new_n5269__ & new_new_n5271__;
  assign new_new_n5274__ = ~new_new_n5272__ & ~new_new_n5273__;
  assign new_new_n5275__ = ~new_new_n5176__ & ~new_new_n5179__;
  assign new_new_n5276__ = ~new_new_n5175__ & ~new_new_n5275__;
  assign new_new_n5277__ = ~new_new_n5274__ & ~new_new_n5276__;
  assign new_new_n5278__ = new_new_n5274__ & new_new_n5276__;
  assign new_new_n5279__ = ~new_new_n5277__ & ~new_new_n5278__;
  assign new_new_n5280__ = ~new_new_n5028__ & ~new_new_n5032__;
  assign new_new_n5281__ = ~new_new_n5029__ & ~new_new_n5280__;
  assign new_new_n5282__ = ~new_new_n5157__ & ~new_new_n5168__;
  assign new_new_n5283__ = ~new_new_n5158__ & ~new_new_n5282__;
  assign new_new_n5284__ = ~new_new_n5121__ & ~new_new_n5132__;
  assign new_new_n5285__ = ~new_new_n5122__ & ~new_new_n5284__;
  assign new_new_n5286__ = new_new_n5283__ & new_new_n5285__;
  assign new_new_n5287__ = ~new_new_n5283__ & ~new_new_n5285__;
  assign new_new_n5288__ = ~new_new_n5286__ & ~new_new_n5287__;
  assign new_new_n5289__ = ~new_new_n5139__ & ~new_new_n5143__;
  assign new_new_n5290__ = ~new_new_n5142__ & ~new_new_n5289__;
  assign new_new_n5291__ = ~new_new_n5103__ & ~new_new_n5107__;
  assign new_new_n5292__ = ~new_new_n5106__ & ~new_new_n5291__;
  assign new_new_n5293__ = ~new_new_n5124__ & ~new_new_n5128__;
  assign new_new_n5294__ = ~new_new_n5127__ & ~new_new_n5293__;
  assign new_new_n5295__ = ~new_new_n5292__ & ~new_new_n5294__;
  assign new_new_n5296__ = new_new_n5292__ & new_new_n5294__;
  assign new_new_n5297__ = ~new_new_n5295__ & ~new_new_n5296__;
  assign new_new_n5298__ = new_new_n5290__ & ~new_new_n5297__;
  assign new_new_n5299__ = ~new_new_n5290__ & new_new_n5297__;
  assign new_new_n5300__ = ~new_new_n5298__ & ~new_new_n5299__;
  assign new_new_n5301__ = new_new_n5288__ & ~new_new_n5300__;
  assign new_new_n5302__ = ~new_new_n5288__ & new_new_n5300__;
  assign new_new_n5303__ = ~new_new_n5301__ & ~new_new_n5302__;
  assign new_new_n5304__ = ~new_new_n5014__ & ~new_new_n5019__;
  assign new_new_n5305__ = ~new_new_n5020__ & ~new_new_n5304__;
  assign new_new_n5306__ = ~new_new_n5083__ & new_new_n5092__;
  assign new_new_n5307__ = ~new_new_n5082__ & ~new_new_n5306__;
  assign new_new_n5308__ = ~new_new_n5064__ & ~new_new_n5071__;
  assign new_new_n5309__ = ~new_new_n5065__ & ~new_new_n5308__;
  assign new_new_n5310__ = ~new_new_n5307__ & new_new_n5309__;
  assign new_new_n5311__ = new_new_n5307__ & ~new_new_n5309__;
  assign new_new_n5312__ = ~new_new_n5310__ & ~new_new_n5311__;
  assign new_new_n5313__ = new_new_n5305__ & ~new_new_n5312__;
  assign new_new_n5314__ = ~new_new_n5305__ & new_new_n5312__;
  assign new_new_n5315__ = ~new_new_n5313__ & ~new_new_n5314__;
  assign new_new_n5316__ = new_new_n5303__ & ~new_new_n5315__;
  assign new_new_n5317__ = ~new_new_n5303__ & new_new_n5315__;
  assign new_new_n5318__ = ~new_new_n5316__ & ~new_new_n5317__;
  assign new_new_n5319__ = ~new_new_n5076__ & new_new_n5095__;
  assign new_new_n5320__ = ~new_new_n5075__ & ~new_new_n5319__;
  assign new_new_n5321__ = new_new_n5318__ & new_new_n5320__;
  assign new_new_n5322__ = ~new_new_n5318__ & ~new_new_n5320__;
  assign new_new_n5323__ = ~new_new_n5321__ & ~new_new_n5322__;
  assign new_new_n5324__ = ~new_new_n5010__ & ~new_new_n5024__;
  assign new_new_n5325__ = ~new_new_n5011__ & ~new_new_n5324__;
  assign new_new_n5326__ = pi22 & pi23;
  assign new_new_n5327__ = pi21 & pi24;
  assign new_new_n5328__ = pi10 & pi35;
  assign new_new_n5329__ = ~new_new_n5327__ & ~new_new_n5328__;
  assign new_new_n5330__ = new_new_n5327__ & new_new_n5328__;
  assign new_new_n5331__ = ~new_new_n5329__ & ~new_new_n5330__;
  assign new_new_n5332__ = new_new_n5326__ & ~new_new_n5331__;
  assign new_new_n5333__ = ~new_new_n5326__ & new_new_n5331__;
  assign new_new_n5334__ = ~new_new_n5332__ & ~new_new_n5333__;
  assign new_new_n5335__ = pi04 & pi41;
  assign new_new_n5336__ = pi02 & pi43;
  assign new_new_n5337__ = pi00 & pi45;
  assign new_new_n5338__ = ~new_new_n5336__ & ~new_new_n5337__;
  assign new_new_n5339__ = new_new_n5336__ & new_new_n5337__;
  assign new_new_n5340__ = ~new_new_n5338__ & ~new_new_n5339__;
  assign new_new_n5341__ = new_new_n5335__ & ~new_new_n5340__;
  assign new_new_n5342__ = ~new_new_n5335__ & new_new_n5340__;
  assign new_new_n5343__ = ~new_new_n5341__ & ~new_new_n5342__;
  assign new_new_n5344__ = new_new_n5334__ & new_new_n5343__;
  assign new_new_n5345__ = ~new_new_n5334__ & ~new_new_n5343__;
  assign new_new_n5346__ = ~new_new_n5344__ & ~new_new_n5345__;
  assign new_new_n5347__ = pi09 & pi36;
  assign new_new_n5348__ = pi07 & pi38;
  assign new_new_n5349__ = pi08 & pi37;
  assign new_new_n5350__ = ~new_new_n5348__ & ~new_new_n5349__;
  assign new_new_n5351__ = new_new_n5348__ & new_new_n5349__;
  assign new_new_n5352__ = ~new_new_n5350__ & ~new_new_n5351__;
  assign new_new_n5353__ = new_new_n5347__ & ~new_new_n5352__;
  assign new_new_n5354__ = ~new_new_n5347__ & new_new_n5352__;
  assign new_new_n5355__ = ~new_new_n5353__ & ~new_new_n5354__;
  assign new_new_n5356__ = new_new_n5346__ & ~new_new_n5355__;
  assign new_new_n5357__ = ~new_new_n5346__ & new_new_n5355__;
  assign new_new_n5358__ = ~new_new_n5356__ & ~new_new_n5357__;
  assign new_new_n5359__ = ~new_new_n5325__ & new_new_n5358__;
  assign new_new_n5360__ = new_new_n5325__ & ~new_new_n5358__;
  assign new_new_n5361__ = ~new_new_n5359__ & ~new_new_n5360__;
  assign new_new_n5362__ = ~new_new_n5112__ & ~new_new_n5116__;
  assign new_new_n5363__ = ~new_new_n5115__ & ~new_new_n5362__;
  assign new_new_n5364__ = pi20 & pi25;
  assign new_new_n5365__ = pi19 & pi26;
  assign new_new_n5366__ = pi18 & pi27;
  assign new_new_n5367__ = ~new_new_n5365__ & ~new_new_n5366__;
  assign new_new_n5368__ = new_new_n5365__ & new_new_n5366__;
  assign new_new_n5369__ = ~new_new_n5367__ & ~new_new_n5368__;
  assign new_new_n5370__ = new_new_n5364__ & ~new_new_n5369__;
  assign new_new_n5371__ = ~new_new_n5364__ & new_new_n5369__;
  assign new_new_n5372__ = ~new_new_n5370__ & ~new_new_n5371__;
  assign new_new_n5373__ = pi14 & pi31;
  assign new_new_n5374__ = pi13 & pi32;
  assign new_new_n5375__ = pi05 & pi40;
  assign new_new_n5376__ = ~new_new_n5374__ & ~new_new_n5375__;
  assign new_new_n5377__ = new_new_n5374__ & new_new_n5375__;
  assign new_new_n5378__ = ~new_new_n5376__ & ~new_new_n5377__;
  assign new_new_n5379__ = new_new_n5373__ & ~new_new_n5378__;
  assign new_new_n5380__ = ~new_new_n5373__ & new_new_n5378__;
  assign new_new_n5381__ = ~new_new_n5379__ & ~new_new_n5380__;
  assign new_new_n5382__ = new_new_n5372__ & new_new_n5381__;
  assign new_new_n5383__ = ~new_new_n5372__ & ~new_new_n5381__;
  assign new_new_n5384__ = ~new_new_n5382__ & ~new_new_n5383__;
  assign new_new_n5385__ = new_new_n5363__ & new_new_n5384__;
  assign new_new_n5386__ = ~new_new_n5363__ & ~new_new_n5384__;
  assign new_new_n5387__ = ~new_new_n5385__ & ~new_new_n5386__;
  assign new_new_n5388__ = new_new_n5361__ & ~new_new_n5387__;
  assign new_new_n5389__ = ~new_new_n5361__ & new_new_n5387__;
  assign new_new_n5390__ = ~new_new_n5388__ & ~new_new_n5389__;
  assign new_new_n5391__ = ~new_new_n5323__ & ~new_new_n5390__;
  assign new_new_n5392__ = new_new_n5323__ & new_new_n5390__;
  assign new_new_n5393__ = ~new_new_n5391__ & ~new_new_n5392__;
  assign new_new_n5394__ = ~new_new_n5281__ & new_new_n5393__;
  assign new_new_n5395__ = new_new_n5281__ & ~new_new_n5393__;
  assign new_new_n5396__ = ~new_new_n5394__ & ~new_new_n5395__;
  assign new_new_n5397__ = new_new_n5279__ & ~new_new_n5396__;
  assign new_new_n5398__ = ~new_new_n5279__ & new_new_n5396__;
  assign new_new_n5399__ = ~new_new_n5397__ & ~new_new_n5398__;
  assign new_new_n5400__ = ~new_new_n5037__ & new_new_n5198__;
  assign new_new_n5401__ = ~new_new_n5037__ & ~new_new_n5199__;
  assign new_new_n5402__ = ~new_new_n5198__ & ~new_new_n5401__;
  assign new_new_n5403__ = new_new_n5182__ & ~new_new_n5402__;
  assign new_new_n5404__ = ~new_new_n5035__ & ~new_new_n5400__;
  assign new_new_n5405__ = ~new_new_n5403__ & new_new_n5404__;
  assign new_new_n5406__ = new_new_n5037__ & new_new_n5199__;
  assign new_new_n5407__ = ~new_new_n5182__ & new_new_n5402__;
  assign new_new_n5408__ = new_new_n5035__ & ~new_new_n5406__;
  assign new_new_n5409__ = ~new_new_n5407__ & new_new_n5408__;
  assign new_new_n5410__ = ~new_new_n5405__ & ~new_new_n5409__;
  assign new_new_n5411__ = ~new_new_n5182__ & new_new_n5187__;
  assign new_new_n5412__ = new_new_n5037__ & ~new_new_n5197__;
  assign new_new_n5413__ = new_new_n5411__ & new_new_n5412__;
  assign new_new_n5414__ = ~new_new_n5209__ & new_new_n5399__;
  assign new_new_n5415__ = ~new_new_n5413__ & new_new_n5414__;
  assign new_new_n5416__ = ~new_new_n5410__ & new_new_n5415__;
  assign new_new_n5417__ = ~new_new_n5035__ & ~new_new_n5184__;
  assign new_new_n5418__ = ~new_new_n5183__ & ~new_new_n5417__;
  assign new_new_n5419__ = new_new_n5198__ & new_new_n5418__;
  assign new_new_n5420__ = new_new_n5035__ & new_new_n5184__;
  assign new_new_n5421__ = ~new_new_n5035__ & new_new_n5183__;
  assign new_new_n5422__ = ~new_new_n5420__ & ~new_new_n5421__;
  assign new_new_n5423__ = new_new_n5200__ & new_new_n5422__;
  assign new_new_n5424__ = new_new_n5199__ & ~new_new_n5418__;
  assign new_new_n5425__ = ~new_new_n5399__ & ~new_new_n5419__;
  assign new_new_n5426__ = ~new_new_n5424__ & new_new_n5425__;
  assign new_new_n5427__ = ~new_new_n5423__ & new_new_n5426__;
  assign po046 = ~new_new_n5416__ & ~new_new_n5427__;
  assign new_new_n5429__ = new_new_n5035__ & ~new_new_n5208__;
  assign new_new_n5430__ = ~new_new_n5411__ & ~new_new_n5429__;
  assign new_new_n5431__ = ~new_new_n5399__ & ~new_new_n5430__;
  assign new_new_n5432__ = new_new_n5207__ & ~new_new_n5431__;
  assign new_new_n5433__ = new_new_n5399__ & new_new_n5430__;
  assign new_new_n5434__ = ~new_new_n5208__ & ~new_new_n5399__;
  assign new_new_n5435__ = new_new_n5399__ & ~new_new_n5411__;
  assign new_new_n5436__ = new_new_n5035__ & ~new_new_n5435__;
  assign new_new_n5437__ = ~new_new_n5434__ & ~new_new_n5436__;
  assign new_new_n5438__ = ~new_new_n5412__ & new_new_n5437__;
  assign new_new_n5439__ = ~new_new_n5432__ & ~new_new_n5433__;
  assign new_new_n5440__ = ~new_new_n5438__ & new_new_n5439__;
  assign new_new_n5441__ = ~new_new_n5278__ & new_new_n5396__;
  assign new_new_n5442__ = ~new_new_n5277__ & ~new_new_n5441__;
  assign new_new_n5443__ = ~new_new_n5440__ & new_new_n5442__;
  assign new_new_n5444__ = new_new_n5440__ & ~new_new_n5442__;
  assign new_new_n5445__ = ~new_new_n5443__ & ~new_new_n5444__;
  assign new_new_n5446__ = ~new_new_n5281__ & ~new_new_n5391__;
  assign new_new_n5447__ = ~new_new_n5392__ & ~new_new_n5446__;
  assign new_new_n5448__ = ~new_new_n5359__ & ~new_new_n5387__;
  assign new_new_n5449__ = ~new_new_n5360__ & ~new_new_n5448__;
  assign new_new_n5450__ = ~new_new_n5317__ & ~new_new_n5320__;
  assign new_new_n5451__ = ~new_new_n5316__ & ~new_new_n5450__;
  assign new_new_n5452__ = ~new_new_n5449__ & new_new_n5451__;
  assign new_new_n5453__ = new_new_n5449__ & ~new_new_n5451__;
  assign new_new_n5454__ = ~new_new_n5452__ & ~new_new_n5453__;
  assign new_new_n5455__ = new_new_n5305__ & ~new_new_n5310__;
  assign new_new_n5456__ = ~new_new_n5311__ & ~new_new_n5455__;
  assign new_new_n5457__ = ~new_new_n5290__ & ~new_new_n5296__;
  assign new_new_n5458__ = ~new_new_n5295__ & ~new_new_n5457__;
  assign new_new_n5459__ = pi14 & pi32;
  assign new_new_n5460__ = pi13 & pi33;
  assign new_new_n5461__ = pi06 & pi40;
  assign new_new_n5462__ = ~new_new_n5460__ & ~new_new_n5461__;
  assign new_new_n5463__ = new_new_n5460__ & new_new_n5461__;
  assign new_new_n5464__ = ~new_new_n5462__ & ~new_new_n5463__;
  assign new_new_n5465__ = new_new_n5459__ & ~new_new_n5464__;
  assign new_new_n5466__ = ~new_new_n5459__ & new_new_n5464__;
  assign new_new_n5467__ = ~new_new_n5465__ & ~new_new_n5466__;
  assign new_new_n5468__ = pi05 & pi41;
  assign new_new_n5469__ = pi02 & pi44;
  assign new_new_n5470__ = ~new_new_n5468__ & ~new_new_n5469__;
  assign new_new_n5471__ = new_new_n5468__ & new_new_n5469__;
  assign new_new_n5472__ = ~new_new_n5470__ & ~new_new_n5471__;
  assign new_new_n5473__ = new_new_n3016__ & ~new_new_n5472__;
  assign new_new_n5474__ = ~new_new_n3016__ & new_new_n5472__;
  assign new_new_n5475__ = ~new_new_n5473__ & ~new_new_n5474__;
  assign new_new_n5476__ = ~new_new_n5467__ & ~new_new_n5475__;
  assign new_new_n5477__ = new_new_n5467__ & new_new_n5475__;
  assign new_new_n5478__ = ~new_new_n5476__ & ~new_new_n5477__;
  assign new_new_n5479__ = new_new_n5458__ & ~new_new_n5478__;
  assign new_new_n5480__ = ~new_new_n5458__ & new_new_n5478__;
  assign new_new_n5481__ = ~new_new_n5479__ & ~new_new_n5480__;
  assign new_new_n5482__ = ~new_new_n5456__ & ~new_new_n5481__;
  assign new_new_n5483__ = new_new_n5456__ & new_new_n5481__;
  assign new_new_n5484__ = ~new_new_n5482__ & ~new_new_n5483__;
  assign new_new_n5485__ = ~new_new_n5364__ & ~new_new_n5368__;
  assign new_new_n5486__ = ~new_new_n5367__ & ~new_new_n5485__;
  assign new_new_n5487__ = ~new_new_n5227__ & ~new_new_n5231__;
  assign new_new_n5488__ = ~new_new_n5230__ & ~new_new_n5487__;
  assign new_new_n5489__ = ~new_new_n5250__ & ~new_new_n5254__;
  assign new_new_n5490__ = ~new_new_n5253__ & ~new_new_n5489__;
  assign new_new_n5491__ = new_new_n5488__ & new_new_n5490__;
  assign new_new_n5492__ = ~new_new_n5488__ & ~new_new_n5490__;
  assign new_new_n5493__ = ~new_new_n5491__ & ~new_new_n5492__;
  assign new_new_n5494__ = new_new_n5486__ & ~new_new_n5493__;
  assign new_new_n5495__ = ~new_new_n5486__ & new_new_n5493__;
  assign new_new_n5496__ = ~new_new_n5494__ & ~new_new_n5495__;
  assign new_new_n5497__ = new_new_n5484__ & new_new_n5496__;
  assign new_new_n5498__ = ~new_new_n5484__ & ~new_new_n5496__;
  assign new_new_n5499__ = ~new_new_n5497__ & ~new_new_n5498__;
  assign new_new_n5500__ = new_new_n5454__ & ~new_new_n5499__;
  assign new_new_n5501__ = ~new_new_n5454__ & new_new_n5499__;
  assign new_new_n5502__ = ~new_new_n5500__ & ~new_new_n5501__;
  assign new_new_n5503__ = ~new_new_n5286__ & ~new_new_n5300__;
  assign new_new_n5504__ = ~new_new_n5287__ & ~new_new_n5503__;
  assign new_new_n5505__ = pi11 & pi35;
  assign new_new_n5506__ = pi10 & pi36;
  assign new_new_n5507__ = pi09 & pi37;
  assign new_new_n5508__ = ~new_new_n5506__ & ~new_new_n5507__;
  assign new_new_n5509__ = new_new_n5506__ & new_new_n5507__;
  assign new_new_n5510__ = ~new_new_n5508__ & ~new_new_n5509__;
  assign new_new_n5511__ = new_new_n5505__ & ~new_new_n5510__;
  assign new_new_n5512__ = ~new_new_n5505__ & new_new_n5510__;
  assign new_new_n5513__ = ~new_new_n5511__ & ~new_new_n5512__;
  assign new_new_n5514__ = pi21 & pi25;
  assign new_new_n5515__ = pi19 & pi27;
  assign new_new_n5516__ = pi20 & pi26;
  assign new_new_n5517__ = ~new_new_n5515__ & ~new_new_n5516__;
  assign new_new_n5518__ = new_new_n5515__ & new_new_n5516__;
  assign new_new_n5519__ = ~new_new_n5517__ & ~new_new_n5518__;
  assign new_new_n5520__ = new_new_n5514__ & ~new_new_n5519__;
  assign new_new_n5521__ = ~new_new_n5514__ & new_new_n5519__;
  assign new_new_n5522__ = ~new_new_n5520__ & ~new_new_n5521__;
  assign new_new_n5523__ = new_new_n5513__ & new_new_n5522__;
  assign new_new_n5524__ = ~new_new_n5513__ & ~new_new_n5522__;
  assign new_new_n5525__ = ~new_new_n5523__ & ~new_new_n5524__;
  assign new_new_n5526__ = pi04 & pi42;
  assign new_new_n5527__ = pi03 & pi43;
  assign new_new_n5528__ = pi00 & pi46;
  assign new_new_n5529__ = ~new_new_n5527__ & ~new_new_n5528__;
  assign new_new_n5530__ = new_new_n5527__ & new_new_n5528__;
  assign new_new_n5531__ = ~new_new_n5529__ & ~new_new_n5530__;
  assign new_new_n5532__ = new_new_n5526__ & ~new_new_n5531__;
  assign new_new_n5533__ = ~new_new_n5526__ & new_new_n5531__;
  assign new_new_n5534__ = ~new_new_n5532__ & ~new_new_n5533__;
  assign new_new_n5535__ = new_new_n5525__ & ~new_new_n5534__;
  assign new_new_n5536__ = ~new_new_n5525__ & new_new_n5534__;
  assign new_new_n5537__ = ~new_new_n5535__ & ~new_new_n5536__;
  assign new_new_n5538__ = new_new_n5504__ & ~new_new_n5537__;
  assign new_new_n5539__ = ~new_new_n5504__ & new_new_n5537__;
  assign new_new_n5540__ = ~new_new_n5538__ & ~new_new_n5539__;
  assign new_new_n5541__ = pi18 & pi28;
  assign new_new_n5542__ = pi17 & pi29;
  assign new_new_n5543__ = ~new_new_n2728__ & ~new_new_n5542__;
  assign new_new_n5544__ = new_new_n2728__ & new_new_n5542__;
  assign new_new_n5545__ = ~new_new_n5543__ & ~new_new_n5544__;
  assign new_new_n5546__ = new_new_n5541__ & ~new_new_n5545__;
  assign new_new_n5547__ = ~new_new_n5541__ & new_new_n5545__;
  assign new_new_n5548__ = ~new_new_n5546__ & ~new_new_n5547__;
  assign new_new_n5549__ = pi12 & pi34;
  assign new_new_n5550__ = pi08 & pi38;
  assign new_new_n5551__ = pi07 & pi39;
  assign new_new_n5552__ = ~new_new_n5550__ & ~new_new_n5551__;
  assign new_new_n5553__ = new_new_n5550__ & new_new_n5551__;
  assign new_new_n5554__ = ~new_new_n5552__ & ~new_new_n5553__;
  assign new_new_n5555__ = new_new_n5549__ & ~new_new_n5554__;
  assign new_new_n5556__ = ~new_new_n5549__ & new_new_n5554__;
  assign new_new_n5557__ = ~new_new_n5555__ & ~new_new_n5556__;
  assign new_new_n5558__ = pi44 & ~new_new_n5239__;
  assign new_new_n5559__ = new_new_n5237__ & ~new_new_n5558__;
  assign new_new_n5560__ = ~new_new_n5241__ & ~new_new_n5559__;
  assign new_new_n5561__ = pi23 & ~new_new_n5560__;
  assign new_new_n5562__ = ~pi23 & new_new_n5239__;
  assign new_new_n5563__ = new_new_n5240__ & new_new_n5562__;
  assign new_new_n5564__ = ~new_new_n5561__ & ~new_new_n5563__;
  assign new_new_n5565__ = new_new_n5557__ & new_new_n5564__;
  assign new_new_n5566__ = ~new_new_n5557__ & ~new_new_n5564__;
  assign new_new_n5567__ = ~new_new_n5548__ & ~new_new_n5565__;
  assign new_new_n5568__ = ~new_new_n5566__ & ~new_new_n5567__;
  assign new_new_n5569__ = ~new_new_n5565__ & new_new_n5568__;
  assign new_new_n5570__ = new_new_n5548__ & ~new_new_n5569__;
  assign new_new_n5571__ = ~new_new_n5566__ & new_new_n5567__;
  assign new_new_n5572__ = ~new_new_n5570__ & ~new_new_n5571__;
  assign new_new_n5573__ = new_new_n5540__ & ~new_new_n5572__;
  assign new_new_n5574__ = ~new_new_n5540__ & new_new_n5572__;
  assign new_new_n5575__ = ~new_new_n5573__ & ~new_new_n5574__;
  assign new_new_n5576__ = ~new_new_n5225__ & new_new_n5261__;
  assign new_new_n5577__ = ~new_new_n5224__ & ~new_new_n5576__;
  assign new_new_n5578__ = ~new_new_n5248__ & ~new_new_n5258__;
  assign new_new_n5579__ = ~new_new_n5247__ & ~new_new_n5578__;
  assign new_new_n5580__ = new_new_n5363__ & ~new_new_n5382__;
  assign new_new_n5581__ = ~new_new_n5383__ & ~new_new_n5580__;
  assign new_new_n5582__ = ~new_new_n5344__ & ~new_new_n5355__;
  assign new_new_n5583__ = ~new_new_n5345__ & ~new_new_n5582__;
  assign new_new_n5584__ = ~new_new_n5581__ & ~new_new_n5583__;
  assign new_new_n5585__ = new_new_n5581__ & new_new_n5583__;
  assign new_new_n5586__ = ~new_new_n5584__ & ~new_new_n5585__;
  assign new_new_n5587__ = new_new_n5579__ & ~new_new_n5586__;
  assign new_new_n5588__ = ~new_new_n5579__ & new_new_n5586__;
  assign new_new_n5589__ = ~new_new_n5587__ & ~new_new_n5588__;
  assign new_new_n5590__ = new_new_n5577__ & ~new_new_n5589__;
  assign new_new_n5591__ = ~new_new_n5577__ & new_new_n5589__;
  assign new_new_n5592__ = ~new_new_n5590__ & ~new_new_n5591__;
  assign new_new_n5593__ = ~new_new_n5213__ & ~new_new_n5219__;
  assign new_new_n5594__ = ~new_new_n5218__ & ~new_new_n5593__;
  assign new_new_n5595__ = pi22 & pi24;
  assign new_new_n5596__ = ~new_new_n5326__ & ~new_new_n5330__;
  assign new_new_n5597__ = ~new_new_n5329__ & ~new_new_n5596__;
  assign new_new_n5598__ = new_new_n5595__ & new_new_n5597__;
  assign new_new_n5599__ = ~new_new_n5595__ & ~new_new_n5597__;
  assign new_new_n5600__ = ~new_new_n5598__ & ~new_new_n5599__;
  assign new_new_n5601__ = pi23 & pi44;
  assign new_new_n5602__ = ~pi45 & ~new_new_n5601__;
  assign new_new_n5603__ = pi23 & pi45;
  assign new_new_n5604__ = pi44 & new_new_n5603__;
  assign new_new_n5605__ = pi01 & ~new_new_n5602__;
  assign new_new_n5606__ = ~new_new_n5604__ & new_new_n5605__;
  assign new_new_n5607__ = ~new_new_n5600__ & new_new_n5606__;
  assign new_new_n5608__ = new_new_n5600__ & ~new_new_n5606__;
  assign new_new_n5609__ = ~new_new_n5607__ & ~new_new_n5608__;
  assign new_new_n5610__ = ~new_new_n5373__ & ~new_new_n5377__;
  assign new_new_n5611__ = ~new_new_n5376__ & ~new_new_n5610__;
  assign new_new_n5612__ = ~new_new_n5347__ & ~new_new_n5351__;
  assign new_new_n5613__ = ~new_new_n5350__ & ~new_new_n5612__;
  assign new_new_n5614__ = ~new_new_n5611__ & ~new_new_n5613__;
  assign new_new_n5615__ = new_new_n5611__ & new_new_n5613__;
  assign new_new_n5616__ = ~new_new_n5614__ & ~new_new_n5615__;
  assign new_new_n5617__ = ~new_new_n5335__ & ~new_new_n5339__;
  assign new_new_n5618__ = ~new_new_n5338__ & ~new_new_n5617__;
  assign new_new_n5619__ = ~new_new_n5616__ & new_new_n5618__;
  assign new_new_n5620__ = new_new_n5616__ & ~new_new_n5618__;
  assign new_new_n5621__ = ~new_new_n5619__ & ~new_new_n5620__;
  assign new_new_n5622__ = ~new_new_n5609__ & ~new_new_n5621__;
  assign new_new_n5623__ = new_new_n5609__ & new_new_n5621__;
  assign new_new_n5624__ = ~new_new_n5622__ & ~new_new_n5623__;
  assign new_new_n5625__ = new_new_n5594__ & new_new_n5624__;
  assign new_new_n5626__ = ~new_new_n5594__ & ~new_new_n5624__;
  assign new_new_n5627__ = ~new_new_n5625__ & ~new_new_n5626__;
  assign new_new_n5628__ = new_new_n5592__ & ~new_new_n5627__;
  assign new_new_n5629__ = ~new_new_n5592__ & new_new_n5627__;
  assign new_new_n5630__ = ~new_new_n5628__ & ~new_new_n5629__;
  assign new_new_n5631__ = new_new_n5575__ & new_new_n5630__;
  assign new_new_n5632__ = ~new_new_n5575__ & ~new_new_n5630__;
  assign new_new_n5633__ = ~new_new_n5631__ & ~new_new_n5632__;
  assign new_new_n5634__ = ~new_new_n5267__ & ~new_new_n5271__;
  assign new_new_n5635__ = ~new_new_n5268__ & ~new_new_n5634__;
  assign new_new_n5636__ = new_new_n5633__ & new_new_n5635__;
  assign new_new_n5637__ = ~new_new_n5633__ & ~new_new_n5635__;
  assign new_new_n5638__ = ~new_new_n5636__ & ~new_new_n5637__;
  assign new_new_n5639__ = new_new_n5502__ & ~new_new_n5638__;
  assign new_new_n5640__ = ~new_new_n5502__ & new_new_n5638__;
  assign new_new_n5641__ = ~new_new_n5639__ & ~new_new_n5640__;
  assign new_new_n5642__ = new_new_n5447__ & ~new_new_n5641__;
  assign new_new_n5643__ = ~new_new_n5447__ & new_new_n5641__;
  assign new_new_n5644__ = ~new_new_n5642__ & ~new_new_n5643__;
  assign new_new_n5645__ = new_new_n5445__ & new_new_n5644__;
  assign new_new_n5646__ = ~new_new_n5445__ & ~new_new_n5644__;
  assign po047 = new_new_n5645__ | new_new_n5646__;
  assign new_new_n5648__ = ~new_new_n5452__ & ~new_new_n5499__;
  assign new_new_n5649__ = ~new_new_n5453__ & ~new_new_n5648__;
  assign new_new_n5650__ = ~new_new_n5539__ & ~new_new_n5572__;
  assign new_new_n5651__ = ~new_new_n5538__ & ~new_new_n5650__;
  assign new_new_n5652__ = ~new_new_n5523__ & ~new_new_n5534__;
  assign new_new_n5653__ = ~new_new_n5524__ & ~new_new_n5652__;
  assign new_new_n5654__ = ~new_new_n5514__ & ~new_new_n5518__;
  assign new_new_n5655__ = ~new_new_n5517__ & ~new_new_n5654__;
  assign new_new_n5656__ = ~new_new_n5526__ & ~new_new_n5530__;
  assign new_new_n5657__ = ~new_new_n5529__ & ~new_new_n5656__;
  assign new_new_n5658__ = ~new_new_n5655__ & ~new_new_n5657__;
  assign new_new_n5659__ = new_new_n5655__ & new_new_n5657__;
  assign new_new_n5660__ = ~new_new_n5658__ & ~new_new_n5659__;
  assign new_new_n5661__ = new_new_n5653__ & ~new_new_n5660__;
  assign new_new_n5662__ = ~new_new_n5653__ & new_new_n5660__;
  assign new_new_n5663__ = ~new_new_n5661__ & ~new_new_n5662__;
  assign new_new_n5664__ = ~new_new_n3016__ & ~new_new_n5471__;
  assign new_new_n5665__ = ~new_new_n5470__ & ~new_new_n5664__;
  assign new_new_n5666__ = new_new_n5458__ & ~new_new_n5477__;
  assign new_new_n5667__ = ~new_new_n5476__ & ~new_new_n5666__;
  assign new_new_n5668__ = new_new_n5665__ & ~new_new_n5667__;
  assign new_new_n5669__ = ~new_new_n5665__ & new_new_n5667__;
  assign new_new_n5670__ = ~new_new_n5668__ & ~new_new_n5669__;
  assign new_new_n5671__ = new_new_n5663__ & new_new_n5670__;
  assign new_new_n5672__ = ~new_new_n5663__ & ~new_new_n5670__;
  assign new_new_n5673__ = ~new_new_n5671__ & ~new_new_n5672__;
  assign new_new_n5674__ = ~new_new_n5651__ & ~new_new_n5673__;
  assign new_new_n5675__ = new_new_n5651__ & new_new_n5673__;
  assign new_new_n5676__ = ~new_new_n5674__ & ~new_new_n5675__;
  assign new_new_n5677__ = ~new_new_n5483__ & ~new_new_n5496__;
  assign new_new_n5678__ = ~new_new_n5482__ & ~new_new_n5677__;
  assign new_new_n5679__ = new_new_n5676__ & ~new_new_n5678__;
  assign new_new_n5680__ = ~new_new_n5676__ & new_new_n5678__;
  assign new_new_n5681__ = ~new_new_n5679__ & ~new_new_n5680__;
  assign new_new_n5682__ = ~new_new_n5649__ & new_new_n5681__;
  assign new_new_n5683__ = new_new_n5649__ & ~new_new_n5681__;
  assign new_new_n5684__ = ~new_new_n5682__ & ~new_new_n5683__;
  assign new_new_n5685__ = ~new_new_n5591__ & ~new_new_n5627__;
  assign new_new_n5686__ = ~new_new_n5590__ & ~new_new_n5685__;
  assign new_new_n5687__ = new_new_n5684__ & ~new_new_n5686__;
  assign new_new_n5688__ = ~new_new_n5684__ & new_new_n5686__;
  assign new_new_n5689__ = ~new_new_n5687__ & ~new_new_n5688__;
  assign new_new_n5690__ = pi11 & pi36;
  assign new_new_n5691__ = pi08 & pi39;
  assign new_new_n5692__ = pi09 & pi38;
  assign new_new_n5693__ = ~new_new_n5691__ & ~new_new_n5692__;
  assign new_new_n5694__ = new_new_n5691__ & new_new_n5692__;
  assign new_new_n5695__ = ~new_new_n5693__ & ~new_new_n5694__;
  assign new_new_n5696__ = new_new_n5690__ & ~new_new_n5695__;
  assign new_new_n5697__ = ~new_new_n5690__ & new_new_n5695__;
  assign new_new_n5698__ = ~new_new_n5696__ & ~new_new_n5697__;
  assign new_new_n5699__ = pi14 & pi33;
  assign new_new_n5700__ = pi06 & pi41;
  assign new_new_n5701__ = pi05 & pi42;
  assign new_new_n5702__ = ~new_new_n5700__ & ~new_new_n5701__;
  assign new_new_n5703__ = new_new_n5700__ & new_new_n5701__;
  assign new_new_n5704__ = ~new_new_n5702__ & ~new_new_n5703__;
  assign new_new_n5705__ = new_new_n5699__ & ~new_new_n5704__;
  assign new_new_n5706__ = ~new_new_n5699__ & new_new_n5704__;
  assign new_new_n5707__ = ~new_new_n5705__ & ~new_new_n5706__;
  assign new_new_n5708__ = new_new_n5698__ & new_new_n5707__;
  assign new_new_n5709__ = ~new_new_n5698__ & ~new_new_n5707__;
  assign new_new_n5710__ = ~new_new_n5708__ & ~new_new_n5709__;
  assign new_new_n5711__ = pi23 & pi24;
  assign new_new_n5712__ = pi10 & pi37;
  assign new_new_n5713__ = pi22 & pi25;
  assign new_new_n5714__ = ~new_new_n5712__ & ~new_new_n5713__;
  assign new_new_n5715__ = new_new_n5712__ & new_new_n5713__;
  assign new_new_n5716__ = ~new_new_n5714__ & ~new_new_n5715__;
  assign new_new_n5717__ = new_new_n5711__ & ~new_new_n5716__;
  assign new_new_n5718__ = ~new_new_n5711__ & new_new_n5716__;
  assign new_new_n5719__ = ~new_new_n5717__ & ~new_new_n5718__;
  assign new_new_n5720__ = new_new_n5710__ & ~new_new_n5719__;
  assign new_new_n5721__ = ~new_new_n5710__ & new_new_n5719__;
  assign new_new_n5722__ = ~new_new_n5720__ & ~new_new_n5721__;
  assign new_new_n5723__ = ~new_new_n5459__ & ~new_new_n5463__;
  assign new_new_n5724__ = ~new_new_n5462__ & ~new_new_n5723__;
  assign new_new_n5725__ = pi15 & pi32;
  assign new_new_n5726__ = pi04 & pi43;
  assign new_new_n5727__ = pi03 & pi44;
  assign new_new_n5728__ = ~new_new_n5726__ & ~new_new_n5727__;
  assign new_new_n5729__ = new_new_n5726__ & new_new_n5727__;
  assign new_new_n5730__ = ~new_new_n5728__ & ~new_new_n5729__;
  assign new_new_n5731__ = new_new_n5725__ & ~new_new_n5730__;
  assign new_new_n5732__ = ~new_new_n5725__ & new_new_n5730__;
  assign new_new_n5733__ = ~new_new_n5731__ & ~new_new_n5732__;
  assign new_new_n5734__ = ~new_new_n5724__ & new_new_n5733__;
  assign new_new_n5735__ = new_new_n5724__ & ~new_new_n5733__;
  assign new_new_n5736__ = ~new_new_n5734__ & ~new_new_n5735__;
  assign new_new_n5737__ = ~new_new_n5541__ & ~new_new_n5544__;
  assign new_new_n5738__ = ~new_new_n5543__ & ~new_new_n5737__;
  assign new_new_n5739__ = new_new_n5736__ & ~new_new_n5738__;
  assign new_new_n5740__ = ~new_new_n5736__ & new_new_n5738__;
  assign new_new_n5741__ = ~new_new_n5739__ & ~new_new_n5740__;
  assign new_new_n5742__ = ~new_new_n5722__ & new_new_n5741__;
  assign new_new_n5743__ = new_new_n5722__ & ~new_new_n5741__;
  assign new_new_n5744__ = ~new_new_n5742__ & ~new_new_n5743__;
  assign new_new_n5745__ = pi00 & pi47;
  assign new_new_n5746__ = pi22 & new_new_n1844__;
  assign new_new_n5747__ = ~pi02 & ~new_new_n5746__;
  assign new_new_n5748__ = pi45 & ~new_new_n5747__;
  assign new_new_n5749__ = new_new_n1717__ & new_new_n1844__;
  assign new_new_n5750__ = new_new_n5748__ & ~new_new_n5749__;
  assign new_new_n5751__ = new_new_n5745__ & ~new_new_n5750__;
  assign new_new_n5752__ = ~new_new_n5745__ & new_new_n5750__;
  assign new_new_n5753__ = ~new_new_n5751__ & ~new_new_n5752__;
  assign new_new_n5754__ = pi21 & pi26;
  assign new_new_n5755__ = pi20 & pi27;
  assign new_new_n5756__ = pi19 & pi28;
  assign new_new_n5757__ = ~new_new_n5755__ & ~new_new_n5756__;
  assign new_new_n5758__ = new_new_n5755__ & new_new_n5756__;
  assign new_new_n5759__ = ~new_new_n5757__ & ~new_new_n5758__;
  assign new_new_n5760__ = new_new_n5754__ & ~new_new_n5759__;
  assign new_new_n5761__ = ~new_new_n5754__ & new_new_n5759__;
  assign new_new_n5762__ = ~new_new_n5760__ & ~new_new_n5761__;
  assign new_new_n5763__ = new_new_n5753__ & new_new_n5762__;
  assign new_new_n5764__ = ~new_new_n5753__ & ~new_new_n5762__;
  assign new_new_n5765__ = ~new_new_n5763__ & ~new_new_n5764__;
  assign new_new_n5766__ = pi18 & pi29;
  assign new_new_n5767__ = pi17 & pi30;
  assign new_new_n5768__ = pi16 & pi31;
  assign new_new_n5769__ = ~new_new_n5767__ & ~new_new_n5768__;
  assign new_new_n5770__ = new_new_n5767__ & new_new_n5768__;
  assign new_new_n5771__ = ~new_new_n5769__ & ~new_new_n5770__;
  assign new_new_n5772__ = new_new_n5766__ & ~new_new_n5771__;
  assign new_new_n5773__ = ~new_new_n5766__ & new_new_n5771__;
  assign new_new_n5774__ = ~new_new_n5772__ & ~new_new_n5773__;
  assign new_new_n5775__ = ~new_new_n5765__ & new_new_n5774__;
  assign new_new_n5776__ = new_new_n5765__ & ~new_new_n5774__;
  assign new_new_n5777__ = ~new_new_n5775__ & ~new_new_n5776__;
  assign new_new_n5778__ = new_new_n5744__ & new_new_n5777__;
  assign new_new_n5779__ = ~new_new_n5744__ & ~new_new_n5777__;
  assign new_new_n5780__ = ~new_new_n5778__ & ~new_new_n5779__;
  assign new_new_n5781__ = ~new_new_n5615__ & ~new_new_n5618__;
  assign new_new_n5782__ = ~new_new_n5614__ & ~new_new_n5781__;
  assign new_new_n5783__ = pi24 & pi46;
  assign new_new_n5784__ = pi01 & new_new_n5783__;
  assign new_new_n5785__ = pi01 & pi46;
  assign new_new_n5786__ = ~pi24 & ~new_new_n5785__;
  assign new_new_n5787__ = ~new_new_n5784__ & ~new_new_n5786__;
  assign new_new_n5788__ = ~new_new_n5549__ & ~new_new_n5553__;
  assign new_new_n5789__ = ~new_new_n5552__ & ~new_new_n5788__;
  assign new_new_n5790__ = ~new_new_n5505__ & ~new_new_n5509__;
  assign new_new_n5791__ = ~new_new_n5508__ & ~new_new_n5790__;
  assign new_new_n5792__ = new_new_n5789__ & new_new_n5791__;
  assign new_new_n5793__ = ~new_new_n5789__ & ~new_new_n5791__;
  assign new_new_n5794__ = ~new_new_n5792__ & ~new_new_n5793__;
  assign new_new_n5795__ = new_new_n5787__ & ~new_new_n5794__;
  assign new_new_n5796__ = ~new_new_n5787__ & new_new_n5794__;
  assign new_new_n5797__ = ~new_new_n5795__ & ~new_new_n5796__;
  assign new_new_n5798__ = ~new_new_n5568__ & ~new_new_n5797__;
  assign new_new_n5799__ = new_new_n5568__ & new_new_n5797__;
  assign new_new_n5800__ = ~new_new_n5798__ & ~new_new_n5799__;
  assign new_new_n5801__ = new_new_n5782__ & new_new_n5800__;
  assign new_new_n5802__ = ~new_new_n5782__ & ~new_new_n5800__;
  assign new_new_n5803__ = ~new_new_n5801__ & ~new_new_n5802__;
  assign new_new_n5804__ = new_new_n5780__ & new_new_n5803__;
  assign new_new_n5805__ = ~new_new_n5780__ & ~new_new_n5803__;
  assign new_new_n5806__ = ~new_new_n5804__ & ~new_new_n5805__;
  assign new_new_n5807__ = ~new_new_n5579__ & ~new_new_n5585__;
  assign new_new_n5808__ = ~new_new_n5584__ & ~new_new_n5807__;
  assign new_new_n5809__ = new_new_n5594__ & ~new_new_n5623__;
  assign new_new_n5810__ = ~new_new_n5622__ & ~new_new_n5809__;
  assign new_new_n5811__ = ~new_new_n5597__ & ~new_new_n5601__;
  assign new_new_n5812__ = pi45 & ~new_new_n5595__;
  assign new_new_n5813__ = ~new_new_n5811__ & new_new_n5812__;
  assign new_new_n5814__ = ~pi45 & new_new_n5595__;
  assign new_new_n5815__ = ~new_new_n5597__ & ~new_new_n5814__;
  assign new_new_n5816__ = new_new_n5601__ & ~new_new_n5815__;
  assign new_new_n5817__ = ~new_new_n5813__ & ~new_new_n5816__;
  assign new_new_n5818__ = pi01 & ~new_new_n5817__;
  assign new_new_n5819__ = pi01 & pi45;
  assign new_new_n5820__ = new_new_n5598__ & ~new_new_n5819__;
  assign new_new_n5821__ = ~new_new_n5818__ & ~new_new_n5820__;
  assign new_new_n5822__ = pi13 & pi34;
  assign new_new_n5823__ = pi12 & pi35;
  assign new_new_n5824__ = pi07 & pi40;
  assign new_new_n5825__ = ~new_new_n5823__ & ~new_new_n5824__;
  assign new_new_n5826__ = new_new_n5823__ & new_new_n5824__;
  assign new_new_n5827__ = ~new_new_n5825__ & ~new_new_n5826__;
  assign new_new_n5828__ = new_new_n5822__ & ~new_new_n5827__;
  assign new_new_n5829__ = ~new_new_n5822__ & new_new_n5827__;
  assign new_new_n5830__ = ~new_new_n5828__ & ~new_new_n5829__;
  assign new_new_n5831__ = new_new_n5821__ & new_new_n5830__;
  assign new_new_n5832__ = ~new_new_n5821__ & ~new_new_n5830__;
  assign new_new_n5833__ = ~new_new_n5831__ & ~new_new_n5832__;
  assign new_new_n5834__ = ~new_new_n5486__ & ~new_new_n5491__;
  assign new_new_n5835__ = ~new_new_n5492__ & ~new_new_n5834__;
  assign new_new_n5836__ = new_new_n5833__ & new_new_n5835__;
  assign new_new_n5837__ = ~new_new_n5833__ & ~new_new_n5835__;
  assign new_new_n5838__ = ~new_new_n5836__ & ~new_new_n5837__;
  assign new_new_n5839__ = new_new_n5810__ & ~new_new_n5838__;
  assign new_new_n5840__ = ~new_new_n5810__ & new_new_n5838__;
  assign new_new_n5841__ = ~new_new_n5808__ & ~new_new_n5839__;
  assign new_new_n5842__ = ~new_new_n5840__ & ~new_new_n5841__;
  assign new_new_n5843__ = ~new_new_n5839__ & new_new_n5842__;
  assign new_new_n5844__ = new_new_n5808__ & ~new_new_n5843__;
  assign new_new_n5845__ = ~new_new_n5840__ & new_new_n5841__;
  assign new_new_n5846__ = ~new_new_n5844__ & ~new_new_n5845__;
  assign new_new_n5847__ = new_new_n5806__ & ~new_new_n5846__;
  assign new_new_n5848__ = ~new_new_n5806__ & new_new_n5846__;
  assign new_new_n5849__ = ~new_new_n5847__ & ~new_new_n5848__;
  assign new_new_n5850__ = new_new_n5689__ & new_new_n5849__;
  assign new_new_n5851__ = ~new_new_n5689__ & ~new_new_n5849__;
  assign new_new_n5852__ = ~new_new_n5850__ & ~new_new_n5851__;
  assign new_new_n5853__ = ~new_new_n5631__ & ~new_new_n5635__;
  assign new_new_n5854__ = ~new_new_n5632__ & ~new_new_n5853__;
  assign new_new_n5855__ = new_new_n5852__ & new_new_n5854__;
  assign new_new_n5856__ = ~new_new_n5852__ & ~new_new_n5854__;
  assign new_new_n5857__ = ~new_new_n5855__ & ~new_new_n5856__;
  assign new_new_n5858__ = ~new_new_n5447__ & new_new_n5640__;
  assign new_new_n5859__ = new_new_n5447__ & new_new_n5639__;
  assign new_new_n5860__ = ~new_new_n5858__ & ~new_new_n5859__;
  assign new_new_n5861__ = new_new_n5445__ & new_new_n5860__;
  assign new_new_n5862__ = new_new_n5447__ & ~new_new_n5640__;
  assign new_new_n5863__ = ~new_new_n5639__ & ~new_new_n5862__;
  assign new_new_n5864__ = new_new_n5444__ & ~new_new_n5863__;
  assign new_new_n5865__ = new_new_n5443__ & new_new_n5863__;
  assign new_new_n5866__ = ~new_new_n5864__ & ~new_new_n5865__;
  assign new_new_n5867__ = ~new_new_n5861__ & new_new_n5866__;
  assign new_new_n5868__ = new_new_n5857__ & ~new_new_n5867__;
  assign new_new_n5869__ = ~new_new_n5443__ & new_new_n5638__;
  assign new_new_n5870__ = ~new_new_n5444__ & ~new_new_n5869__;
  assign new_new_n5871__ = new_new_n5502__ & new_new_n5870__;
  assign new_new_n5872__ = new_new_n5443__ & ~new_new_n5638__;
  assign new_new_n5873__ = ~new_new_n5871__ & ~new_new_n5872__;
  assign new_new_n5874__ = new_new_n5447__ & ~new_new_n5873__;
  assign new_new_n5875__ = ~new_new_n5502__ & ~new_new_n5870__;
  assign new_new_n5876__ = new_new_n5444__ & new_new_n5638__;
  assign new_new_n5877__ = ~new_new_n5875__ & ~new_new_n5876__;
  assign new_new_n5878__ = ~new_new_n5447__ & ~new_new_n5877__;
  assign new_new_n5879__ = new_new_n5440__ & new_new_n5638__;
  assign new_new_n5880__ = new_new_n5442__ & new_new_n5502__;
  assign new_new_n5881__ = ~new_new_n5879__ & ~new_new_n5880__;
  assign new_new_n5882__ = ~new_new_n5440__ & ~new_new_n5638__;
  assign new_new_n5883__ = ~new_new_n5442__ & ~new_new_n5502__;
  assign new_new_n5884__ = ~new_new_n5882__ & ~new_new_n5883__;
  assign new_new_n5885__ = ~new_new_n5881__ & ~new_new_n5884__;
  assign new_new_n5886__ = ~new_new_n5874__ & ~new_new_n5885__;
  assign new_new_n5887__ = ~new_new_n5878__ & new_new_n5886__;
  assign new_new_n5888__ = ~new_new_n5857__ & ~new_new_n5887__;
  assign po048 = new_new_n5868__ | new_new_n5888__;
  assign new_new_n5890__ = ~new_new_n5682__ & ~new_new_n5686__;
  assign new_new_n5891__ = ~new_new_n5683__ & ~new_new_n5890__;
  assign new_new_n5892__ = ~new_new_n5804__ & ~new_new_n5846__;
  assign new_new_n5893__ = ~new_new_n5805__ & ~new_new_n5892__;
  assign new_new_n5894__ = ~new_new_n5743__ & ~new_new_n5777__;
  assign new_new_n5895__ = ~new_new_n5742__ & ~new_new_n5894__;
  assign new_new_n5896__ = ~new_new_n5763__ & ~new_new_n5774__;
  assign new_new_n5897__ = ~new_new_n5764__ & ~new_new_n5896__;
  assign new_new_n5898__ = ~new_new_n5787__ & ~new_new_n5792__;
  assign new_new_n5899__ = ~new_new_n5793__ & ~new_new_n5898__;
  assign new_new_n5900__ = ~new_new_n5766__ & ~new_new_n5770__;
  assign new_new_n5901__ = ~new_new_n5769__ & ~new_new_n5900__;
  assign new_new_n5902__ = ~new_new_n5725__ & ~new_new_n5729__;
  assign new_new_n5903__ = ~new_new_n5728__ & ~new_new_n5902__;
  assign new_new_n5904__ = ~new_new_n5745__ & ~new_new_n5749__;
  assign new_new_n5905__ = new_new_n5748__ & ~new_new_n5904__;
  assign new_new_n5906__ = new_new_n5903__ & new_new_n5905__;
  assign new_new_n5907__ = ~new_new_n5903__ & ~new_new_n5905__;
  assign new_new_n5908__ = ~new_new_n5906__ & ~new_new_n5907__;
  assign new_new_n5909__ = ~new_new_n5901__ & ~new_new_n5908__;
  assign new_new_n5910__ = new_new_n5901__ & new_new_n5908__;
  assign new_new_n5911__ = ~new_new_n5909__ & ~new_new_n5910__;
  assign new_new_n5912__ = ~new_new_n5899__ & ~new_new_n5911__;
  assign new_new_n5913__ = new_new_n5899__ & new_new_n5911__;
  assign new_new_n5914__ = ~new_new_n5912__ & ~new_new_n5913__;
  assign new_new_n5915__ = new_new_n5897__ & ~new_new_n5914__;
  assign new_new_n5916__ = ~new_new_n5897__ & new_new_n5914__;
  assign new_new_n5917__ = ~new_new_n5915__ & ~new_new_n5916__;
  assign new_new_n5918__ = ~new_new_n5895__ & ~new_new_n5917__;
  assign new_new_n5919__ = new_new_n5895__ & new_new_n5917__;
  assign new_new_n5920__ = ~new_new_n5918__ & ~new_new_n5919__;
  assign new_new_n5921__ = ~new_new_n5690__ & ~new_new_n5694__;
  assign new_new_n5922__ = ~new_new_n5693__ & ~new_new_n5921__;
  assign new_new_n5923__ = ~new_new_n5754__ & ~new_new_n5758__;
  assign new_new_n5924__ = ~new_new_n5757__ & ~new_new_n5923__;
  assign new_new_n5925__ = new_new_n5922__ & new_new_n5924__;
  assign new_new_n5926__ = ~new_new_n5922__ & ~new_new_n5924__;
  assign new_new_n5927__ = ~new_new_n5925__ & ~new_new_n5926__;
  assign new_new_n5928__ = ~new_new_n5699__ & ~new_new_n5703__;
  assign new_new_n5929__ = ~new_new_n5702__ & ~new_new_n5928__;
  assign new_new_n5930__ = ~new_new_n5927__ & new_new_n5929__;
  assign new_new_n5931__ = ~new_new_n5925__ & ~new_new_n5929__;
  assign new_new_n5932__ = ~new_new_n5926__ & new_new_n5931__;
  assign new_new_n5933__ = ~new_new_n5930__ & ~new_new_n5932__;
  assign new_new_n5934__ = ~new_new_n5708__ & ~new_new_n5719__;
  assign new_new_n5935__ = ~new_new_n5709__ & ~new_new_n5934__;
  assign new_new_n5936__ = ~new_new_n5711__ & ~new_new_n5715__;
  assign new_new_n5937__ = ~new_new_n5714__ & ~new_new_n5936__;
  assign new_new_n5938__ = pi16 & pi32;
  assign new_new_n5939__ = pi03 & pi45;
  assign new_new_n5940__ = pi02 & pi46;
  assign new_new_n5941__ = ~new_new_n5939__ & ~new_new_n5940__;
  assign new_new_n5942__ = new_new_n5939__ & new_new_n5940__;
  assign new_new_n5943__ = ~new_new_n5941__ & ~new_new_n5942__;
  assign new_new_n5944__ = new_new_n5938__ & ~new_new_n5943__;
  assign new_new_n5945__ = ~new_new_n5938__ & new_new_n5943__;
  assign new_new_n5946__ = ~new_new_n5944__ & ~new_new_n5945__;
  assign new_new_n5947__ = ~new_new_n5937__ & new_new_n5946__;
  assign new_new_n5948__ = new_new_n5937__ & ~new_new_n5946__;
  assign new_new_n5949__ = ~new_new_n5947__ & ~new_new_n5948__;
  assign new_new_n5950__ = ~new_new_n5822__ & ~new_new_n5826__;
  assign new_new_n5951__ = ~new_new_n5825__ & ~new_new_n5950__;
  assign new_new_n5952__ = new_new_n5949__ & ~new_new_n5951__;
  assign new_new_n5953__ = ~new_new_n5949__ & new_new_n5951__;
  assign new_new_n5954__ = ~new_new_n5952__ & ~new_new_n5953__;
  assign new_new_n5955__ = new_new_n5935__ & ~new_new_n5954__;
  assign new_new_n5956__ = ~new_new_n5935__ & new_new_n5954__;
  assign new_new_n5957__ = ~new_new_n5955__ & ~new_new_n5956__;
  assign new_new_n5958__ = new_new_n5933__ & new_new_n5957__;
  assign new_new_n5959__ = ~new_new_n5933__ & ~new_new_n5957__;
  assign new_new_n5960__ = ~new_new_n5958__ & ~new_new_n5959__;
  assign new_new_n5961__ = new_new_n5920__ & new_new_n5960__;
  assign new_new_n5962__ = ~new_new_n5920__ & ~new_new_n5960__;
  assign new_new_n5963__ = ~new_new_n5961__ & ~new_new_n5962__;
  assign new_new_n5964__ = ~new_new_n5893__ & ~new_new_n5963__;
  assign new_new_n5965__ = new_new_n5893__ & new_new_n5963__;
  assign new_new_n5966__ = ~new_new_n5964__ & ~new_new_n5965__;
  assign new_new_n5967__ = ~new_new_n5659__ & ~new_new_n5665__;
  assign new_new_n5968__ = ~new_new_n5658__ & ~new_new_n5967__;
  assign new_new_n5969__ = pi00 & pi48;
  assign new_new_n5970__ = pi23 & pi25;
  assign new_new_n5971__ = pi01 & pi47;
  assign new_new_n5972__ = ~new_new_n5970__ & new_new_n5971__;
  assign new_new_n5973__ = new_new_n5970__ & ~new_new_n5971__;
  assign new_new_n5974__ = ~new_new_n5972__ & ~new_new_n5973__;
  assign new_new_n5975__ = ~new_new_n5969__ & new_new_n5974__;
  assign new_new_n5976__ = new_new_n5969__ & ~new_new_n5974__;
  assign new_new_n5977__ = ~new_new_n5975__ & ~new_new_n5976__;
  assign new_new_n5978__ = new_new_n5784__ & new_new_n5977__;
  assign new_new_n5979__ = ~new_new_n5784__ & ~new_new_n5977__;
  assign new_new_n5980__ = ~new_new_n5978__ & ~new_new_n5979__;
  assign new_new_n5981__ = ~new_new_n5968__ & ~new_new_n5980__;
  assign new_new_n5982__ = new_new_n5968__ & new_new_n5980__;
  assign new_new_n5983__ = ~new_new_n5981__ & ~new_new_n5982__;
  assign new_new_n5984__ = ~new_new_n5734__ & new_new_n5738__;
  assign new_new_n5985__ = ~new_new_n5735__ & ~new_new_n5984__;
  assign new_new_n5986__ = new_new_n5983__ & ~new_new_n5985__;
  assign new_new_n5987__ = ~new_new_n5983__ & new_new_n5985__;
  assign new_new_n5988__ = ~new_new_n5986__ & ~new_new_n5987__;
  assign new_new_n5989__ = ~new_new_n5782__ & ~new_new_n5798__;
  assign new_new_n5990__ = ~new_new_n5799__ & ~new_new_n5989__;
  assign new_new_n5991__ = new_new_n5988__ & new_new_n5990__;
  assign new_new_n5992__ = ~new_new_n5988__ & ~new_new_n5990__;
  assign new_new_n5993__ = ~new_new_n5991__ & ~new_new_n5992__;
  assign new_new_n5994__ = new_new_n5653__ & new_new_n5667__;
  assign new_new_n5995__ = ~new_new_n5653__ & ~new_new_n5667__;
  assign new_new_n5996__ = ~new_new_n5660__ & new_new_n5665__;
  assign new_new_n5997__ = new_new_n5660__ & ~new_new_n5665__;
  assign new_new_n5998__ = ~new_new_n5996__ & ~new_new_n5997__;
  assign new_new_n5999__ = ~new_new_n5995__ & new_new_n5998__;
  assign new_new_n6000__ = ~new_new_n5994__ & ~new_new_n5999__;
  assign new_new_n6001__ = new_new_n5993__ & ~new_new_n6000__;
  assign new_new_n6002__ = ~new_new_n5993__ & new_new_n6000__;
  assign new_new_n6003__ = ~new_new_n6001__ & ~new_new_n6002__;
  assign new_new_n6004__ = new_new_n5966__ & ~new_new_n6003__;
  assign new_new_n6005__ = ~new_new_n5966__ & new_new_n6003__;
  assign new_new_n6006__ = ~new_new_n6004__ & ~new_new_n6005__;
  assign new_new_n6007__ = ~new_new_n5891__ & ~new_new_n6006__;
  assign new_new_n6008__ = new_new_n5891__ & new_new_n6006__;
  assign new_new_n6009__ = ~new_new_n6007__ & ~new_new_n6008__;
  assign new_new_n6010__ = ~new_new_n5674__ & ~new_new_n5678__;
  assign new_new_n6011__ = ~new_new_n5675__ & ~new_new_n6010__;
  assign new_new_n6012__ = pi14 & pi34;
  assign new_new_n6013__ = pi13 & pi35;
  assign new_new_n6014__ = pi06 & pi42;
  assign new_new_n6015__ = ~new_new_n6013__ & ~new_new_n6014__;
  assign new_new_n6016__ = new_new_n6013__ & new_new_n6014__;
  assign new_new_n6017__ = ~new_new_n6015__ & ~new_new_n6016__;
  assign new_new_n6018__ = new_new_n6012__ & ~new_new_n6017__;
  assign new_new_n6019__ = ~new_new_n6012__ & new_new_n6017__;
  assign new_new_n6020__ = ~new_new_n6018__ & ~new_new_n6019__;
  assign new_new_n6021__ = pi11 & pi37;
  assign new_new_n6022__ = pi09 & pi39;
  assign new_new_n6023__ = pi10 & pi38;
  assign new_new_n6024__ = ~new_new_n6022__ & ~new_new_n6023__;
  assign new_new_n6025__ = new_new_n6022__ & new_new_n6023__;
  assign new_new_n6026__ = ~new_new_n6024__ & ~new_new_n6025__;
  assign new_new_n6027__ = new_new_n6021__ & ~new_new_n6026__;
  assign new_new_n6028__ = ~new_new_n6021__ & new_new_n6026__;
  assign new_new_n6029__ = ~new_new_n6027__ & ~new_new_n6028__;
  assign new_new_n6030__ = new_new_n6020__ & new_new_n6029__;
  assign new_new_n6031__ = ~new_new_n6020__ & ~new_new_n6029__;
  assign new_new_n6032__ = ~new_new_n6030__ & ~new_new_n6031__;
  assign new_new_n6033__ = pi12 & pi36;
  assign new_new_n6034__ = pi08 & pi40;
  assign new_new_n6035__ = pi07 & pi41;
  assign new_new_n6036__ = ~new_new_n6034__ & ~new_new_n6035__;
  assign new_new_n6037__ = new_new_n6034__ & new_new_n6035__;
  assign new_new_n6038__ = ~new_new_n6036__ & ~new_new_n6037__;
  assign new_new_n6039__ = new_new_n6033__ & ~new_new_n6038__;
  assign new_new_n6040__ = ~new_new_n6033__ & new_new_n6038__;
  assign new_new_n6041__ = ~new_new_n6039__ & ~new_new_n6040__;
  assign new_new_n6042__ = new_new_n6032__ & ~new_new_n6041__;
  assign new_new_n6043__ = ~new_new_n6032__ & new_new_n6041__;
  assign new_new_n6044__ = ~new_new_n6042__ & ~new_new_n6043__;
  assign new_new_n6045__ = ~new_new_n5831__ & new_new_n5835__;
  assign new_new_n6046__ = ~new_new_n5832__ & ~new_new_n6045__;
  assign new_new_n6047__ = ~new_new_n6044__ & new_new_n6046__;
  assign new_new_n6048__ = new_new_n6044__ & ~new_new_n6046__;
  assign new_new_n6049__ = ~new_new_n6047__ & ~new_new_n6048__;
  assign new_new_n6050__ = pi15 & pi33;
  assign new_new_n6051__ = pi04 & pi44;
  assign new_new_n6052__ = pi05 & pi43;
  assign new_new_n6053__ = ~new_new_n6051__ & ~new_new_n6052__;
  assign new_new_n6054__ = new_new_n6051__ & new_new_n6052__;
  assign new_new_n6055__ = ~new_new_n6053__ & ~new_new_n6054__;
  assign new_new_n6056__ = new_new_n6050__ & ~new_new_n6055__;
  assign new_new_n6057__ = ~new_new_n6050__ & new_new_n6055__;
  assign new_new_n6058__ = ~new_new_n6056__ & ~new_new_n6057__;
  assign new_new_n6059__ = pi19 & pi29;
  assign new_new_n6060__ = pi17 & pi31;
  assign new_new_n6061__ = pi18 & pi30;
  assign new_new_n6062__ = ~new_new_n6060__ & ~new_new_n6061__;
  assign new_new_n6063__ = new_new_n6060__ & new_new_n6061__;
  assign new_new_n6064__ = ~new_new_n6062__ & ~new_new_n6063__;
  assign new_new_n6065__ = new_new_n6059__ & ~new_new_n6064__;
  assign new_new_n6066__ = ~new_new_n6059__ & new_new_n6064__;
  assign new_new_n6067__ = ~new_new_n6065__ & ~new_new_n6066__;
  assign new_new_n6068__ = pi22 & pi26;
  assign new_new_n6069__ = pi20 & pi28;
  assign new_new_n6070__ = pi21 & pi27;
  assign new_new_n6071__ = ~new_new_n6069__ & ~new_new_n6070__;
  assign new_new_n6072__ = new_new_n6069__ & new_new_n6070__;
  assign new_new_n6073__ = ~new_new_n6071__ & ~new_new_n6072__;
  assign new_new_n6074__ = new_new_n6068__ & ~new_new_n6073__;
  assign new_new_n6075__ = ~new_new_n6068__ & new_new_n6073__;
  assign new_new_n6076__ = ~new_new_n6074__ & ~new_new_n6075__;
  assign new_new_n6077__ = new_new_n6067__ & new_new_n6076__;
  assign new_new_n6078__ = ~new_new_n6067__ & ~new_new_n6076__;
  assign new_new_n6079__ = ~new_new_n6077__ & ~new_new_n6078__;
  assign new_new_n6080__ = ~new_new_n6058__ & new_new_n6079__;
  assign new_new_n6081__ = new_new_n6058__ & ~new_new_n6079__;
  assign new_new_n6082__ = ~new_new_n6080__ & ~new_new_n6081__;
  assign new_new_n6083__ = new_new_n6049__ & ~new_new_n6082__;
  assign new_new_n6084__ = ~new_new_n6049__ & new_new_n6082__;
  assign new_new_n6085__ = ~new_new_n6083__ & ~new_new_n6084__;
  assign new_new_n6086__ = new_new_n6011__ & new_new_n6085__;
  assign new_new_n6087__ = ~new_new_n6011__ & ~new_new_n6085__;
  assign new_new_n6088__ = ~new_new_n6086__ & ~new_new_n6087__;
  assign new_new_n6089__ = new_new_n5842__ & new_new_n6088__;
  assign new_new_n6090__ = ~new_new_n5842__ & ~new_new_n6088__;
  assign new_new_n6091__ = ~new_new_n6089__ & ~new_new_n6090__;
  assign new_new_n6092__ = new_new_n6009__ & ~new_new_n6091__;
  assign new_new_n6093__ = ~new_new_n6009__ & new_new_n6091__;
  assign new_new_n6094__ = ~new_new_n6092__ & ~new_new_n6093__;
  assign new_new_n6095__ = ~new_new_n5447__ & ~new_new_n5880__;
  assign new_new_n6096__ = new_new_n5857__ & ~new_new_n5882__;
  assign new_new_n6097__ = ~new_new_n5883__ & ~new_new_n6095__;
  assign new_new_n6098__ = ~new_new_n6096__ & new_new_n6097__;
  assign new_new_n6099__ = ~new_new_n5857__ & ~new_new_n5883__;
  assign new_new_n6100__ = new_new_n5857__ & ~new_new_n5880__;
  assign new_new_n6101__ = new_new_n5447__ & ~new_new_n6100__;
  assign new_new_n6102__ = ~new_new_n6099__ & ~new_new_n6101__;
  assign new_new_n6103__ = ~new_new_n5879__ & ~new_new_n6102__;
  assign new_new_n6104__ = ~new_new_n5857__ & new_new_n5882__;
  assign new_new_n6105__ = ~new_new_n6103__ & ~new_new_n6104__;
  assign new_new_n6106__ = ~new_new_n6098__ & new_new_n6105__;
  assign new_new_n6107__ = ~new_new_n6094__ & new_new_n6106__;
  assign new_new_n6108__ = new_new_n6094__ & ~new_new_n6106__;
  assign new_new_n6109__ = ~new_new_n6107__ & ~new_new_n6108__;
  assign new_new_n6110__ = ~new_new_n5850__ & ~new_new_n5854__;
  assign new_new_n6111__ = ~new_new_n5851__ & ~new_new_n6110__;
  assign new_new_n6112__ = new_new_n6109__ & new_new_n6111__;
  assign new_new_n6113__ = ~new_new_n6109__ & ~new_new_n6111__;
  assign po049 = new_new_n6112__ | new_new_n6113__;
  assign new_new_n6115__ = ~new_new_n5965__ & new_new_n6003__;
  assign new_new_n6116__ = ~new_new_n5964__ & ~new_new_n6115__;
  assign new_new_n6117__ = ~new_new_n5935__ & ~new_new_n5954__;
  assign new_new_n6118__ = ~new_new_n5906__ & ~new_new_n5910__;
  assign new_new_n6119__ = ~new_new_n5926__ & ~new_new_n5931__;
  assign new_new_n6120__ = ~new_new_n6118__ & new_new_n6119__;
  assign new_new_n6121__ = new_new_n6118__ & ~new_new_n6119__;
  assign new_new_n6122__ = ~new_new_n6120__ & ~new_new_n6121__;
  assign new_new_n6123__ = ~new_new_n5947__ & new_new_n5951__;
  assign new_new_n6124__ = ~new_new_n5948__ & ~new_new_n6123__;
  assign new_new_n6125__ = new_new_n6122__ & ~new_new_n6124__;
  assign new_new_n6126__ = ~new_new_n6122__ & new_new_n6124__;
  assign new_new_n6127__ = ~new_new_n6125__ & ~new_new_n6126__;
  assign new_new_n6128__ = new_new_n6117__ & new_new_n6127__;
  assign new_new_n6129__ = new_new_n5935__ & new_new_n5954__;
  assign new_new_n6130__ = new_new_n6127__ & ~new_new_n6129__;
  assign new_new_n6131__ = ~new_new_n5929__ & ~new_new_n6130__;
  assign new_new_n6132__ = ~new_new_n6117__ & ~new_new_n6127__;
  assign new_new_n6133__ = new_new_n5929__ & ~new_new_n6132__;
  assign new_new_n6134__ = new_new_n5927__ & ~new_new_n6131__;
  assign new_new_n6135__ = ~new_new_n6133__ & new_new_n6134__;
  assign new_new_n6136__ = ~new_new_n5929__ & ~new_new_n6132__;
  assign new_new_n6137__ = new_new_n5929__ & ~new_new_n6130__;
  assign new_new_n6138__ = ~new_new_n5927__ & ~new_new_n6136__;
  assign new_new_n6139__ = ~new_new_n6137__ & new_new_n6138__;
  assign new_new_n6140__ = ~new_new_n6127__ & new_new_n6129__;
  assign new_new_n6141__ = ~new_new_n6128__ & ~new_new_n6140__;
  assign new_new_n6142__ = ~new_new_n6135__ & new_new_n6141__;
  assign new_new_n6143__ = ~new_new_n6139__ & new_new_n6142__;
  assign new_new_n6144__ = new_new_n5897__ & ~new_new_n5913__;
  assign new_new_n6145__ = ~new_new_n5912__ & ~new_new_n6144__;
  assign new_new_n6146__ = new_new_n6143__ & ~new_new_n6145__;
  assign new_new_n6147__ = ~new_new_n6143__ & new_new_n6145__;
  assign new_new_n6148__ = ~new_new_n6146__ & ~new_new_n6147__;
  assign new_new_n6149__ = ~new_new_n6047__ & new_new_n6082__;
  assign new_new_n6150__ = ~new_new_n6048__ & ~new_new_n6149__;
  assign new_new_n6151__ = ~new_new_n6050__ & ~new_new_n6054__;
  assign new_new_n6152__ = ~new_new_n6053__ & ~new_new_n6151__;
  assign new_new_n6153__ = ~new_new_n6068__ & ~new_new_n6072__;
  assign new_new_n6154__ = ~new_new_n6071__ & ~new_new_n6153__;
  assign new_new_n6155__ = ~new_new_n6152__ & ~new_new_n6154__;
  assign new_new_n6156__ = new_new_n6152__ & new_new_n6154__;
  assign new_new_n6157__ = ~new_new_n6155__ & ~new_new_n6156__;
  assign new_new_n6158__ = ~new_new_n5938__ & ~new_new_n5942__;
  assign new_new_n6159__ = ~new_new_n5941__ & ~new_new_n6158__;
  assign new_new_n6160__ = ~new_new_n6157__ & new_new_n6159__;
  assign new_new_n6161__ = ~new_new_n6156__ & ~new_new_n6159__;
  assign new_new_n6162__ = ~new_new_n6155__ & new_new_n6161__;
  assign new_new_n6163__ = ~new_new_n6160__ & ~new_new_n6162__;
  assign new_new_n6164__ = pi23 & pi47;
  assign new_new_n6165__ = ~new_new_n6021__ & ~new_new_n6025__;
  assign new_new_n6166__ = ~new_new_n6024__ & ~new_new_n6165__;
  assign new_new_n6167__ = pi01 & ~pi48;
  assign new_new_n6168__ = ~new_new_n6166__ & ~new_new_n6167__;
  assign new_new_n6169__ = new_new_n6164__ & ~new_new_n6168__;
  assign new_new_n6170__ = pi25 & pi48;
  assign new_new_n6171__ = new_new_n6166__ & ~new_new_n6170__;
  assign new_new_n6172__ = new_new_n6169__ & ~new_new_n6171__;
  assign new_new_n6173__ = new_new_n5970__ & new_new_n5971__;
  assign new_new_n6174__ = pi01 & pi48;
  assign new_new_n6175__ = new_new_n6166__ & ~new_new_n6174__;
  assign new_new_n6176__ = ~new_new_n6166__ & new_new_n6174__;
  assign new_new_n6177__ = ~new_new_n6175__ & ~new_new_n6176__;
  assign new_new_n6178__ = pi25 & new_new_n6177__;
  assign new_new_n6179__ = ~pi25 & ~new_new_n6177__;
  assign new_new_n6180__ = ~new_new_n6173__ & ~new_new_n6178__;
  assign new_new_n6181__ = ~new_new_n6179__ & new_new_n6180__;
  assign new_new_n6182__ = ~new_new_n6172__ & ~new_new_n6181__;
  assign new_new_n6183__ = ~new_new_n6030__ & ~new_new_n6041__;
  assign new_new_n6184__ = ~new_new_n6031__ & ~new_new_n6183__;
  assign new_new_n6185__ = ~new_new_n6182__ & new_new_n6184__;
  assign new_new_n6186__ = new_new_n6182__ & ~new_new_n6184__;
  assign new_new_n6187__ = ~new_new_n6185__ & ~new_new_n6186__;
  assign new_new_n6188__ = ~new_new_n6163__ & new_new_n6187__;
  assign new_new_n6189__ = new_new_n6163__ & ~new_new_n6187__;
  assign new_new_n6190__ = ~new_new_n6188__ & ~new_new_n6189__;
  assign new_new_n6191__ = ~new_new_n6150__ & new_new_n6190__;
  assign new_new_n6192__ = new_new_n6150__ & ~new_new_n6190__;
  assign new_new_n6193__ = ~new_new_n6191__ & ~new_new_n6192__;
  assign new_new_n6194__ = ~new_new_n6058__ & ~new_new_n6077__;
  assign new_new_n6195__ = ~new_new_n6078__ & ~new_new_n6194__;
  assign new_new_n6196__ = ~new_new_n6012__ & ~new_new_n6016__;
  assign new_new_n6197__ = ~new_new_n6015__ & ~new_new_n6196__;
  assign new_new_n6198__ = ~new_new_n6033__ & ~new_new_n6037__;
  assign new_new_n6199__ = ~new_new_n6036__ & ~new_new_n6198__;
  assign new_new_n6200__ = ~new_new_n6197__ & ~new_new_n6199__;
  assign new_new_n6201__ = new_new_n6197__ & new_new_n6199__;
  assign new_new_n6202__ = ~new_new_n6200__ & ~new_new_n6201__;
  assign new_new_n6203__ = new_new_n6195__ & ~new_new_n6202__;
  assign new_new_n6204__ = ~new_new_n6195__ & new_new_n6202__;
  assign new_new_n6205__ = ~new_new_n6203__ & ~new_new_n6204__;
  assign new_new_n6206__ = ~new_new_n6059__ & ~new_new_n6063__;
  assign new_new_n6207__ = ~new_new_n6062__ & ~new_new_n6206__;
  assign new_new_n6208__ = ~new_new_n5981__ & ~new_new_n5985__;
  assign new_new_n6209__ = ~new_new_n5982__ & ~new_new_n6208__;
  assign new_new_n6210__ = new_new_n6207__ & ~new_new_n6209__;
  assign new_new_n6211__ = ~new_new_n6207__ & new_new_n6209__;
  assign new_new_n6212__ = ~new_new_n6210__ & ~new_new_n6211__;
  assign new_new_n6213__ = new_new_n6205__ & new_new_n6212__;
  assign new_new_n6214__ = ~new_new_n6205__ & ~new_new_n6212__;
  assign new_new_n6215__ = ~new_new_n6213__ & ~new_new_n6214__;
  assign new_new_n6216__ = new_new_n6193__ & ~new_new_n6215__;
  assign new_new_n6217__ = ~new_new_n6193__ & new_new_n6215__;
  assign new_new_n6218__ = ~new_new_n6216__ & ~new_new_n6217__;
  assign new_new_n6219__ = ~new_new_n6148__ & ~new_new_n6218__;
  assign new_new_n6220__ = new_new_n6148__ & new_new_n6218__;
  assign new_new_n6221__ = ~new_new_n6219__ & ~new_new_n6220__;
  assign new_new_n6222__ = ~new_new_n5842__ & ~new_new_n6086__;
  assign new_new_n6223__ = ~new_new_n6087__ & ~new_new_n6222__;
  assign new_new_n6224__ = new_new_n6221__ & new_new_n6223__;
  assign new_new_n6225__ = ~new_new_n6221__ & ~new_new_n6223__;
  assign new_new_n6226__ = ~new_new_n6224__ & ~new_new_n6225__;
  assign new_new_n6227__ = new_new_n6116__ & ~new_new_n6226__;
  assign new_new_n6228__ = ~new_new_n6116__ & new_new_n6226__;
  assign new_new_n6229__ = ~new_new_n6227__ & ~new_new_n6228__;
  assign new_new_n6230__ = ~new_new_n6008__ & new_new_n6091__;
  assign new_new_n6231__ = ~new_new_n6007__ & ~new_new_n6230__;
  assign new_new_n6232__ = ~new_new_n6108__ & new_new_n6111__;
  assign new_new_n6233__ = ~new_new_n6107__ & ~new_new_n6232__;
  assign new_new_n6234__ = ~new_new_n6231__ & ~new_new_n6233__;
  assign new_new_n6235__ = new_new_n6231__ & new_new_n6233__;
  assign new_new_n6236__ = ~new_new_n6234__ & ~new_new_n6235__;
  assign new_new_n6237__ = ~new_new_n5991__ & ~new_new_n6000__;
  assign new_new_n6238__ = ~new_new_n5992__ & ~new_new_n6237__;
  assign new_new_n6239__ = pi24 & pi25;
  assign new_new_n6240__ = pi23 & pi26;
  assign new_new_n6241__ = pi11 & pi38;
  assign new_new_n6242__ = ~new_new_n6240__ & ~new_new_n6241__;
  assign new_new_n6243__ = new_new_n6240__ & new_new_n6241__;
  assign new_new_n6244__ = ~new_new_n6242__ & ~new_new_n6243__;
  assign new_new_n6245__ = new_new_n6239__ & ~new_new_n6244__;
  assign new_new_n6246__ = ~new_new_n6239__ & new_new_n6244__;
  assign new_new_n6247__ = ~new_new_n6245__ & ~new_new_n6246__;
  assign new_new_n6248__ = pi13 & pi36;
  assign new_new_n6249__ = pi08 & pi41;
  assign new_new_n6250__ = pi07 & pi42;
  assign new_new_n6251__ = ~new_new_n6249__ & ~new_new_n6250__;
  assign new_new_n6252__ = new_new_n6249__ & new_new_n6250__;
  assign new_new_n6253__ = ~new_new_n6251__ & ~new_new_n6252__;
  assign new_new_n6254__ = new_new_n6248__ & ~new_new_n6253__;
  assign new_new_n6255__ = ~new_new_n6248__ & new_new_n6253__;
  assign new_new_n6256__ = ~new_new_n6254__ & ~new_new_n6255__;
  assign new_new_n6257__ = new_new_n6247__ & new_new_n6256__;
  assign new_new_n6258__ = ~new_new_n6247__ & ~new_new_n6256__;
  assign new_new_n6259__ = ~new_new_n6257__ & ~new_new_n6258__;
  assign new_new_n6260__ = pi15 & pi34;
  assign new_new_n6261__ = pi14 & pi35;
  assign new_new_n6262__ = pi06 & pi43;
  assign new_new_n6263__ = ~new_new_n6261__ & ~new_new_n6262__;
  assign new_new_n6264__ = new_new_n6261__ & new_new_n6262__;
  assign new_new_n6265__ = ~new_new_n6263__ & ~new_new_n6264__;
  assign new_new_n6266__ = new_new_n6260__ & ~new_new_n6265__;
  assign new_new_n6267__ = ~new_new_n6260__ & new_new_n6265__;
  assign new_new_n6268__ = ~new_new_n6266__ & ~new_new_n6267__;
  assign new_new_n6269__ = ~new_new_n6259__ & new_new_n6268__;
  assign new_new_n6270__ = new_new_n6259__ & ~new_new_n6268__;
  assign new_new_n6271__ = ~new_new_n6269__ & ~new_new_n6270__;
  assign new_new_n6272__ = pi05 & pi44;
  assign new_new_n6273__ = pi04 & pi45;
  assign new_new_n6274__ = pi00 & pi49;
  assign new_new_n6275__ = ~new_new_n6273__ & ~new_new_n6274__;
  assign new_new_n6276__ = new_new_n6273__ & new_new_n6274__;
  assign new_new_n6277__ = ~new_new_n6275__ & ~new_new_n6276__;
  assign new_new_n6278__ = new_new_n6272__ & ~new_new_n6277__;
  assign new_new_n6279__ = ~new_new_n6272__ & new_new_n6277__;
  assign new_new_n6280__ = ~new_new_n6278__ & ~new_new_n6279__;
  assign new_new_n6281__ = new_new_n5784__ & ~new_new_n5975__;
  assign new_new_n6282__ = ~new_new_n5976__ & ~new_new_n6281__;
  assign new_new_n6283__ = new_new_n6280__ & new_new_n6282__;
  assign new_new_n6284__ = ~new_new_n6280__ & ~new_new_n6282__;
  assign new_new_n6285__ = ~new_new_n6283__ & ~new_new_n6284__;
  assign new_new_n6286__ = pi18 & pi31;
  assign new_new_n6287__ = ~pi16 & ~new_new_n3207__;
  assign new_new_n6288__ = ~new_new_n3208__ & ~new_new_n6287__;
  assign new_new_n6289__ = pi32 & pi33;
  assign new_new_n6290__ = new_new_n2941__ & new_new_n6289__;
  assign new_new_n6291__ = new_new_n6288__ & ~new_new_n6290__;
  assign new_new_n6292__ = new_new_n6286__ & ~new_new_n6291__;
  assign new_new_n6293__ = ~new_new_n6286__ & new_new_n6291__;
  assign new_new_n6294__ = ~new_new_n6292__ & ~new_new_n6293__;
  assign new_new_n6295__ = ~new_new_n6285__ & new_new_n6294__;
  assign new_new_n6296__ = new_new_n6285__ & ~new_new_n6294__;
  assign new_new_n6297__ = ~new_new_n6295__ & ~new_new_n6296__;
  assign new_new_n6298__ = new_new_n6271__ & new_new_n6297__;
  assign new_new_n6299__ = ~new_new_n6271__ & ~new_new_n6297__;
  assign new_new_n6300__ = ~new_new_n6298__ & ~new_new_n6299__;
  assign new_new_n6301__ = pi12 & pi37;
  assign new_new_n6302__ = pi10 & pi39;
  assign new_new_n6303__ = pi09 & pi40;
  assign new_new_n6304__ = ~new_new_n6302__ & ~new_new_n6303__;
  assign new_new_n6305__ = new_new_n6302__ & new_new_n6303__;
  assign new_new_n6306__ = ~new_new_n6304__ & ~new_new_n6305__;
  assign new_new_n6307__ = new_new_n6301__ & ~new_new_n6306__;
  assign new_new_n6308__ = ~new_new_n6301__ & new_new_n6306__;
  assign new_new_n6309__ = ~new_new_n6307__ & ~new_new_n6308__;
  assign new_new_n6310__ = pi21 & pi28;
  assign new_new_n6311__ = pi20 & pi29;
  assign new_new_n6312__ = pi19 & pi30;
  assign new_new_n6313__ = ~new_new_n6311__ & ~new_new_n6312__;
  assign new_new_n6314__ = new_new_n6311__ & new_new_n6312__;
  assign new_new_n6315__ = ~new_new_n6313__ & ~new_new_n6314__;
  assign new_new_n6316__ = new_new_n6310__ & ~new_new_n6315__;
  assign new_new_n6317__ = ~new_new_n6310__ & new_new_n6315__;
  assign new_new_n6318__ = ~new_new_n6316__ & ~new_new_n6317__;
  assign new_new_n6319__ = pi22 & pi27;
  assign new_new_n6320__ = pi03 & pi46;
  assign new_new_n6321__ = pi02 & pi47;
  assign new_new_n6322__ = ~new_new_n6320__ & ~new_new_n6321__;
  assign new_new_n6323__ = new_new_n6320__ & new_new_n6321__;
  assign new_new_n6324__ = ~new_new_n6322__ & ~new_new_n6323__;
  assign new_new_n6325__ = new_new_n6319__ & ~new_new_n6324__;
  assign new_new_n6326__ = ~new_new_n6319__ & new_new_n6324__;
  assign new_new_n6327__ = ~new_new_n6325__ & ~new_new_n6326__;
  assign new_new_n6328__ = new_new_n6318__ & new_new_n6327__;
  assign new_new_n6329__ = ~new_new_n6318__ & ~new_new_n6327__;
  assign new_new_n6330__ = ~new_new_n6309__ & ~new_new_n6328__;
  assign new_new_n6331__ = ~new_new_n6329__ & ~new_new_n6330__;
  assign new_new_n6332__ = ~new_new_n6328__ & new_new_n6331__;
  assign new_new_n6333__ = new_new_n6309__ & ~new_new_n6332__;
  assign new_new_n6334__ = ~new_new_n6329__ & new_new_n6330__;
  assign new_new_n6335__ = ~new_new_n6333__ & ~new_new_n6334__;
  assign new_new_n6336__ = new_new_n6300__ & ~new_new_n6335__;
  assign new_new_n6337__ = ~new_new_n6300__ & new_new_n6335__;
  assign new_new_n6338__ = ~new_new_n6336__ & ~new_new_n6337__;
  assign new_new_n6339__ = ~new_new_n5919__ & ~new_new_n5960__;
  assign new_new_n6340__ = ~new_new_n5918__ & ~new_new_n6339__;
  assign new_new_n6341__ = new_new_n6338__ & ~new_new_n6340__;
  assign new_new_n6342__ = ~new_new_n6338__ & new_new_n6340__;
  assign new_new_n6343__ = ~new_new_n6341__ & ~new_new_n6342__;
  assign new_new_n6344__ = new_new_n6238__ & new_new_n6343__;
  assign new_new_n6345__ = ~new_new_n6238__ & ~new_new_n6343__;
  assign new_new_n6346__ = ~new_new_n6344__ & ~new_new_n6345__;
  assign new_new_n6347__ = new_new_n6236__ & ~new_new_n6346__;
  assign new_new_n6348__ = ~new_new_n6236__ & new_new_n6346__;
  assign new_new_n6349__ = ~new_new_n6347__ & ~new_new_n6348__;
  assign new_new_n6350__ = new_new_n6229__ & new_new_n6349__;
  assign new_new_n6351__ = ~new_new_n6229__ & ~new_new_n6349__;
  assign po050 = new_new_n6350__ | new_new_n6351__;
  assign new_new_n6353__ = ~new_new_n6238__ & ~new_new_n6342__;
  assign new_new_n6354__ = ~new_new_n6341__ & ~new_new_n6353__;
  assign new_new_n6355__ = ~new_new_n6298__ & ~new_new_n6335__;
  assign new_new_n6356__ = ~new_new_n6299__ & ~new_new_n6355__;
  assign new_new_n6357__ = pi24 & pi26;
  assign new_new_n6358__ = pi01 & pi49;
  assign new_new_n6359__ = ~new_new_n6357__ & new_new_n6358__;
  assign new_new_n6360__ = new_new_n6357__ & ~new_new_n6358__;
  assign new_new_n6361__ = ~new_new_n6359__ & ~new_new_n6360__;
  assign new_new_n6362__ = ~new_new_n6301__ & ~new_new_n6305__;
  assign new_new_n6363__ = ~new_new_n6304__ & ~new_new_n6362__;
  assign new_new_n6364__ = ~new_new_n6239__ & ~new_new_n6243__;
  assign new_new_n6365__ = ~new_new_n6242__ & ~new_new_n6364__;
  assign new_new_n6366__ = new_new_n6363__ & new_new_n6365__;
  assign new_new_n6367__ = ~new_new_n6363__ & ~new_new_n6365__;
  assign new_new_n6368__ = ~new_new_n6366__ & ~new_new_n6367__;
  assign new_new_n6369__ = new_new_n6361__ & new_new_n6368__;
  assign new_new_n6370__ = ~new_new_n6361__ & ~new_new_n6368__;
  assign new_new_n6371__ = ~new_new_n6369__ & ~new_new_n6370__;
  assign new_new_n6372__ = ~new_new_n6331__ & ~new_new_n6371__;
  assign new_new_n6373__ = new_new_n6331__ & new_new_n6371__;
  assign new_new_n6374__ = ~new_new_n6372__ & ~new_new_n6373__;
  assign new_new_n6375__ = ~new_new_n6283__ & ~new_new_n6294__;
  assign new_new_n6376__ = ~new_new_n6284__ & ~new_new_n6375__;
  assign new_new_n6377__ = new_new_n6374__ & ~new_new_n6376__;
  assign new_new_n6378__ = ~new_new_n6374__ & new_new_n6376__;
  assign new_new_n6379__ = ~new_new_n6377__ & ~new_new_n6378__;
  assign new_new_n6380__ = ~new_new_n6356__ & ~new_new_n6379__;
  assign new_new_n6381__ = new_new_n6356__ & new_new_n6379__;
  assign new_new_n6382__ = ~new_new_n6380__ & ~new_new_n6381__;
  assign new_new_n6383__ = ~new_new_n6310__ & ~new_new_n6314__;
  assign new_new_n6384__ = ~new_new_n6313__ & ~new_new_n6383__;
  assign new_new_n6385__ = ~new_new_n6248__ & ~new_new_n6252__;
  assign new_new_n6386__ = ~new_new_n6251__ & ~new_new_n6385__;
  assign new_new_n6387__ = new_new_n6384__ & new_new_n6386__;
  assign new_new_n6388__ = ~new_new_n6384__ & ~new_new_n6386__;
  assign new_new_n6389__ = ~new_new_n6387__ & ~new_new_n6388__;
  assign new_new_n6390__ = ~new_new_n6286__ & ~new_new_n6290__;
  assign new_new_n6391__ = new_new_n6288__ & ~new_new_n6390__;
  assign new_new_n6392__ = ~new_new_n6389__ & new_new_n6391__;
  assign new_new_n6393__ = new_new_n6389__ & ~new_new_n6391__;
  assign new_new_n6394__ = ~new_new_n6392__ & ~new_new_n6393__;
  assign new_new_n6395__ = ~new_new_n6257__ & ~new_new_n6268__;
  assign new_new_n6396__ = ~new_new_n6258__ & ~new_new_n6395__;
  assign new_new_n6397__ = ~new_new_n6121__ & ~new_new_n6124__;
  assign new_new_n6398__ = ~new_new_n6120__ & ~new_new_n6397__;
  assign new_new_n6399__ = ~new_new_n6396__ & ~new_new_n6398__;
  assign new_new_n6400__ = new_new_n6396__ & new_new_n6398__;
  assign new_new_n6401__ = ~new_new_n6399__ & ~new_new_n6400__;
  assign new_new_n6402__ = ~new_new_n6394__ & new_new_n6401__;
  assign new_new_n6403__ = new_new_n6394__ & ~new_new_n6401__;
  assign new_new_n6404__ = ~new_new_n6402__ & ~new_new_n6403__;
  assign new_new_n6405__ = new_new_n6382__ & new_new_n6404__;
  assign new_new_n6406__ = ~new_new_n6382__ & ~new_new_n6404__;
  assign new_new_n6407__ = ~new_new_n6405__ & ~new_new_n6406__;
  assign new_new_n6408__ = new_new_n6354__ & new_new_n6407__;
  assign new_new_n6409__ = ~new_new_n6354__ & ~new_new_n6407__;
  assign new_new_n6410__ = ~new_new_n6408__ & ~new_new_n6409__;
  assign new_new_n6411__ = ~new_new_n6155__ & ~new_new_n6161__;
  assign new_new_n6412__ = ~new_new_n6201__ & ~new_new_n6207__;
  assign new_new_n6413__ = ~new_new_n6200__ & ~new_new_n6412__;
  assign new_new_n6414__ = new_new_n6411__ & new_new_n6413__;
  assign new_new_n6415__ = ~new_new_n6411__ & ~new_new_n6413__;
  assign new_new_n6416__ = ~new_new_n6414__ & ~new_new_n6415__;
  assign new_new_n6417__ = ~new_new_n6319__ & ~new_new_n6323__;
  assign new_new_n6418__ = ~new_new_n6322__ & ~new_new_n6417__;
  assign new_new_n6419__ = ~new_new_n6260__ & ~new_new_n6264__;
  assign new_new_n6420__ = ~new_new_n6263__ & ~new_new_n6419__;
  assign new_new_n6421__ = ~new_new_n6272__ & ~new_new_n6276__;
  assign new_new_n6422__ = ~new_new_n6275__ & ~new_new_n6421__;
  assign new_new_n6423__ = new_new_n6420__ & new_new_n6422__;
  assign new_new_n6424__ = ~new_new_n6420__ & ~new_new_n6422__;
  assign new_new_n6425__ = ~new_new_n6423__ & ~new_new_n6424__;
  assign new_new_n6426__ = ~new_new_n6418__ & new_new_n6425__;
  assign new_new_n6427__ = new_new_n6418__ & ~new_new_n6425__;
  assign new_new_n6428__ = ~new_new_n6426__ & ~new_new_n6427__;
  assign new_new_n6429__ = new_new_n6416__ & ~new_new_n6428__;
  assign new_new_n6430__ = ~new_new_n6416__ & new_new_n6428__;
  assign new_new_n6431__ = ~new_new_n6429__ & ~new_new_n6430__;
  assign new_new_n6432__ = new_new_n6195__ & new_new_n6209__;
  assign new_new_n6433__ = ~new_new_n6195__ & ~new_new_n6209__;
  assign new_new_n6434__ = new_new_n6202__ & ~new_new_n6207__;
  assign new_new_n6435__ = ~new_new_n6202__ & new_new_n6207__;
  assign new_new_n6436__ = ~new_new_n6434__ & ~new_new_n6435__;
  assign new_new_n6437__ = ~new_new_n6433__ & new_new_n6436__;
  assign new_new_n6438__ = ~new_new_n6432__ & ~new_new_n6437__;
  assign new_new_n6439__ = ~new_new_n6431__ & ~new_new_n6438__;
  assign new_new_n6440__ = new_new_n6431__ & new_new_n6438__;
  assign new_new_n6441__ = ~new_new_n6439__ & ~new_new_n6440__;
  assign new_new_n6442__ = new_new_n6163__ & ~new_new_n6186__;
  assign new_new_n6443__ = ~new_new_n6185__ & ~new_new_n6442__;
  assign new_new_n6444__ = new_new_n6441__ & ~new_new_n6443__;
  assign new_new_n6445__ = ~new_new_n6441__ & new_new_n6443__;
  assign new_new_n6446__ = ~new_new_n6444__ & ~new_new_n6445__;
  assign new_new_n6447__ = new_new_n6410__ & ~new_new_n6446__;
  assign new_new_n6448__ = ~new_new_n6410__ & new_new_n6446__;
  assign new_new_n6449__ = ~new_new_n6447__ & ~new_new_n6448__;
  assign new_new_n6450__ = ~new_new_n6220__ & ~new_new_n6223__;
  assign new_new_n6451__ = ~new_new_n6219__ & ~new_new_n6450__;
  assign new_new_n6452__ = new_new_n6449__ & ~new_new_n6451__;
  assign new_new_n6453__ = ~new_new_n6449__ & new_new_n6451__;
  assign new_new_n6454__ = ~new_new_n6452__ & ~new_new_n6453__;
  assign new_new_n6455__ = ~new_new_n6191__ & ~new_new_n6215__;
  assign new_new_n6456__ = ~new_new_n6192__ & ~new_new_n6455__;
  assign new_new_n6457__ = ~new_new_n6127__ & ~new_new_n6145__;
  assign new_new_n6458__ = new_new_n6127__ & new_new_n6145__;
  assign new_new_n6459__ = new_new_n5933__ & ~new_new_n6117__;
  assign new_new_n6460__ = ~new_new_n6129__ & ~new_new_n6459__;
  assign new_new_n6461__ = ~new_new_n6458__ & ~new_new_n6460__;
  assign new_new_n6462__ = ~new_new_n6457__ & ~new_new_n6461__;
  assign new_new_n6463__ = new_new_n6456__ & new_new_n6462__;
  assign new_new_n6464__ = ~new_new_n6456__ & ~new_new_n6462__;
  assign new_new_n6465__ = pi23 & pi27;
  assign new_new_n6466__ = pi22 & pi28;
  assign new_new_n6467__ = pi18 & pi32;
  assign new_new_n6468__ = ~new_new_n6466__ & ~new_new_n6467__;
  assign new_new_n6469__ = new_new_n6466__ & new_new_n6467__;
  assign new_new_n6470__ = ~new_new_n6468__ & ~new_new_n6469__;
  assign new_new_n6471__ = new_new_n6465__ & ~new_new_n6470__;
  assign new_new_n6472__ = ~new_new_n6465__ & new_new_n6470__;
  assign new_new_n6473__ = ~new_new_n6471__ & ~new_new_n6472__;
  assign new_new_n6474__ = pi16 & pi34;
  assign new_new_n6475__ = pi15 & pi35;
  assign new_new_n6476__ = pi05 & pi45;
  assign new_new_n6477__ = ~new_new_n6475__ & ~new_new_n6476__;
  assign new_new_n6478__ = new_new_n6475__ & new_new_n6476__;
  assign new_new_n6479__ = ~new_new_n6477__ & ~new_new_n6478__;
  assign new_new_n6480__ = new_new_n6474__ & ~new_new_n6479__;
  assign new_new_n6481__ = ~new_new_n6474__ & new_new_n6479__;
  assign new_new_n6482__ = ~new_new_n6480__ & ~new_new_n6481__;
  assign new_new_n6483__ = new_new_n6473__ & new_new_n6482__;
  assign new_new_n6484__ = ~new_new_n6473__ & ~new_new_n6482__;
  assign new_new_n6485__ = ~new_new_n6483__ & ~new_new_n6484__;
  assign new_new_n6486__ = ~new_new_n6169__ & ~new_new_n6175__;
  assign new_new_n6487__ = pi25 & ~new_new_n6486__;
  assign new_new_n6488__ = ~pi25 & new_new_n6174__;
  assign new_new_n6489__ = new_new_n6166__ & new_new_n6488__;
  assign new_new_n6490__ = ~new_new_n6487__ & ~new_new_n6489__;
  assign new_new_n6491__ = new_new_n6485__ & ~new_new_n6490__;
  assign new_new_n6492__ = ~new_new_n6485__ & new_new_n6490__;
  assign new_new_n6493__ = ~new_new_n6491__ & ~new_new_n6492__;
  assign new_new_n6494__ = pi21 & pi29;
  assign new_new_n6495__ = pi20 & pi30;
  assign new_new_n6496__ = pi19 & pi31;
  assign new_new_n6497__ = ~new_new_n6495__ & ~new_new_n6496__;
  assign new_new_n6498__ = new_new_n6495__ & new_new_n6496__;
  assign new_new_n6499__ = ~new_new_n6497__ & ~new_new_n6498__;
  assign new_new_n6500__ = new_new_n6494__ & ~new_new_n6499__;
  assign new_new_n6501__ = ~new_new_n6494__ & new_new_n6499__;
  assign new_new_n6502__ = ~new_new_n6500__ & ~new_new_n6501__;
  assign new_new_n6503__ = pi00 & pi50;
  assign new_new_n6504__ = pi02 & new_new_n1907__;
  assign new_new_n6505__ = ~pi02 & ~new_new_n1907__;
  assign new_new_n6506__ = pi48 & ~new_new_n6505__;
  assign new_new_n6507__ = ~new_new_n6504__ & new_new_n6506__;
  assign new_new_n6508__ = new_new_n6503__ & ~new_new_n6507__;
  assign new_new_n6509__ = ~new_new_n6503__ & new_new_n6507__;
  assign new_new_n6510__ = ~new_new_n6508__ & ~new_new_n6509__;
  assign new_new_n6511__ = new_new_n6502__ & new_new_n6510__;
  assign new_new_n6512__ = ~new_new_n6502__ & ~new_new_n6510__;
  assign new_new_n6513__ = ~new_new_n6511__ & ~new_new_n6512__;
  assign new_new_n6514__ = pi17 & pi33;
  assign new_new_n6515__ = pi03 & pi47;
  assign new_new_n6516__ = pi04 & pi46;
  assign new_new_n6517__ = ~new_new_n6515__ & ~new_new_n6516__;
  assign new_new_n6518__ = new_new_n6515__ & new_new_n6516__;
  assign new_new_n6519__ = ~new_new_n6517__ & ~new_new_n6518__;
  assign new_new_n6520__ = new_new_n6514__ & ~new_new_n6519__;
  assign new_new_n6521__ = ~new_new_n6514__ & new_new_n6519__;
  assign new_new_n6522__ = ~new_new_n6520__ & ~new_new_n6521__;
  assign new_new_n6523__ = new_new_n6513__ & ~new_new_n6522__;
  assign new_new_n6524__ = ~new_new_n6513__ & new_new_n6522__;
  assign new_new_n6525__ = ~new_new_n6523__ & ~new_new_n6524__;
  assign new_new_n6526__ = pi14 & pi36;
  assign new_new_n6527__ = pi07 & pi43;
  assign new_new_n6528__ = pi06 & pi44;
  assign new_new_n6529__ = ~new_new_n6527__ & ~new_new_n6528__;
  assign new_new_n6530__ = new_new_n6527__ & new_new_n6528__;
  assign new_new_n6531__ = ~new_new_n6529__ & ~new_new_n6530__;
  assign new_new_n6532__ = new_new_n6526__ & ~new_new_n6531__;
  assign new_new_n6533__ = ~new_new_n6526__ & new_new_n6531__;
  assign new_new_n6534__ = ~new_new_n6532__ & ~new_new_n6533__;
  assign new_new_n6535__ = pi13 & pi37;
  assign new_new_n6536__ = pi08 & pi42;
  assign new_new_n6537__ = pi09 & pi41;
  assign new_new_n6538__ = ~new_new_n6536__ & ~new_new_n6537__;
  assign new_new_n6539__ = new_new_n6536__ & new_new_n6537__;
  assign new_new_n6540__ = ~new_new_n6538__ & ~new_new_n6539__;
  assign new_new_n6541__ = new_new_n6535__ & ~new_new_n6540__;
  assign new_new_n6542__ = ~new_new_n6535__ & new_new_n6540__;
  assign new_new_n6543__ = ~new_new_n6541__ & ~new_new_n6542__;
  assign new_new_n6544__ = new_new_n6534__ & new_new_n6543__;
  assign new_new_n6545__ = ~new_new_n6534__ & ~new_new_n6543__;
  assign new_new_n6546__ = ~new_new_n6544__ & ~new_new_n6545__;
  assign new_new_n6547__ = pi12 & pi38;
  assign new_new_n6548__ = pi11 & pi39;
  assign new_new_n6549__ = pi10 & pi40;
  assign new_new_n6550__ = ~new_new_n6548__ & ~new_new_n6549__;
  assign new_new_n6551__ = new_new_n6548__ & new_new_n6549__;
  assign new_new_n6552__ = ~new_new_n6550__ & ~new_new_n6551__;
  assign new_new_n6553__ = new_new_n6547__ & ~new_new_n6552__;
  assign new_new_n6554__ = ~new_new_n6547__ & new_new_n6552__;
  assign new_new_n6555__ = ~new_new_n6553__ & ~new_new_n6554__;
  assign new_new_n6556__ = new_new_n6546__ & ~new_new_n6555__;
  assign new_new_n6557__ = ~new_new_n6546__ & new_new_n6555__;
  assign new_new_n6558__ = ~new_new_n6556__ & ~new_new_n6557__;
  assign new_new_n6559__ = new_new_n6525__ & ~new_new_n6558__;
  assign new_new_n6560__ = ~new_new_n6525__ & new_new_n6558__;
  assign new_new_n6561__ = ~new_new_n6559__ & ~new_new_n6560__;
  assign new_new_n6562__ = new_new_n6493__ & new_new_n6561__;
  assign new_new_n6563__ = ~new_new_n6493__ & ~new_new_n6561__;
  assign new_new_n6564__ = ~new_new_n6562__ & ~new_new_n6563__;
  assign new_new_n6565__ = ~new_new_n6463__ & new_new_n6564__;
  assign new_new_n6566__ = ~new_new_n6464__ & ~new_new_n6565__;
  assign new_new_n6567__ = ~new_new_n6463__ & new_new_n6566__;
  assign new_new_n6568__ = ~new_new_n6464__ & new_new_n6565__;
  assign new_new_n6569__ = new_new_n6564__ & ~new_new_n6568__;
  assign new_new_n6570__ = ~new_new_n6567__ & ~new_new_n6569__;
  assign new_new_n6571__ = new_new_n6454__ & ~new_new_n6570__;
  assign new_new_n6572__ = ~new_new_n6454__ & new_new_n6570__;
  assign new_new_n6573__ = ~new_new_n6571__ & ~new_new_n6572__;
  assign new_new_n6574__ = new_new_n6227__ & new_new_n6346__;
  assign new_new_n6575__ = new_new_n6228__ & ~new_new_n6346__;
  assign new_new_n6576__ = ~new_new_n6574__ & ~new_new_n6575__;
  assign new_new_n6577__ = new_new_n6236__ & new_new_n6576__;
  assign new_new_n6578__ = ~new_new_n6227__ & ~new_new_n6346__;
  assign new_new_n6579__ = ~new_new_n6228__ & ~new_new_n6578__;
  assign new_new_n6580__ = new_new_n6235__ & ~new_new_n6579__;
  assign new_new_n6581__ = new_new_n6234__ & new_new_n6579__;
  assign new_new_n6582__ = new_new_n6573__ & ~new_new_n6580__;
  assign new_new_n6583__ = ~new_new_n6581__ & new_new_n6582__;
  assign new_new_n6584__ = ~new_new_n6577__ & new_new_n6583__;
  assign new_new_n6585__ = new_new_n6226__ & ~new_new_n6231__;
  assign new_new_n6586__ = ~new_new_n6233__ & new_new_n6585__;
  assign new_new_n6587__ = ~new_new_n6116__ & new_new_n6586__;
  assign new_new_n6588__ = new_new_n6116__ & ~new_new_n6586__;
  assign new_new_n6589__ = ~new_new_n6226__ & new_new_n6231__;
  assign new_new_n6590__ = ~new_new_n6233__ & ~new_new_n6589__;
  assign new_new_n6591__ = ~new_new_n6585__ & ~new_new_n6590__;
  assign new_new_n6592__ = ~new_new_n6346__ & ~new_new_n6588__;
  assign new_new_n6593__ = ~new_new_n6591__ & new_new_n6592__;
  assign new_new_n6594__ = new_new_n6116__ & new_new_n6591__;
  assign new_new_n6595__ = new_new_n6233__ & new_new_n6589__;
  assign new_new_n6596__ = ~new_new_n6594__ & ~new_new_n6595__;
  assign new_new_n6597__ = new_new_n6346__ & ~new_new_n6596__;
  assign new_new_n6598__ = new_new_n6116__ & new_new_n6233__;
  assign new_new_n6599__ = new_new_n6589__ & new_new_n6598__;
  assign new_new_n6600__ = ~new_new_n6573__ & ~new_new_n6587__;
  assign new_new_n6601__ = ~new_new_n6599__ & new_new_n6600__;
  assign new_new_n6602__ = ~new_new_n6593__ & new_new_n6601__;
  assign new_new_n6603__ = ~new_new_n6597__ & new_new_n6602__;
  assign po051 = ~new_new_n6584__ & ~new_new_n6603__;
  assign new_new_n6605__ = ~new_new_n6116__ & ~new_new_n6233__;
  assign new_new_n6606__ = ~new_new_n6573__ & ~new_new_n6605__;
  assign new_new_n6607__ = ~new_new_n6346__ & ~new_new_n6606__;
  assign new_new_n6608__ = new_new_n6573__ & ~new_new_n6598__;
  assign new_new_n6609__ = ~new_new_n6585__ & ~new_new_n6608__;
  assign new_new_n6610__ = ~new_new_n6607__ & new_new_n6609__;
  assign new_new_n6611__ = ~new_new_n6346__ & ~new_new_n6598__;
  assign new_new_n6612__ = new_new_n6573__ & ~new_new_n6589__;
  assign new_new_n6613__ = ~new_new_n6605__ & ~new_new_n6612__;
  assign new_new_n6614__ = ~new_new_n6611__ & new_new_n6613__;
  assign new_new_n6615__ = ~new_new_n6573__ & new_new_n6589__;
  assign new_new_n6616__ = ~new_new_n6614__ & ~new_new_n6615__;
  assign new_new_n6617__ = ~new_new_n6610__ & new_new_n6616__;
  assign new_new_n6618__ = ~new_new_n6453__ & new_new_n6570__;
  assign new_new_n6619__ = ~new_new_n6452__ & ~new_new_n6618__;
  assign new_new_n6620__ = ~new_new_n6617__ & ~new_new_n6619__;
  assign new_new_n6621__ = new_new_n6617__ & new_new_n6619__;
  assign new_new_n6622__ = ~new_new_n6620__ & ~new_new_n6621__;
  assign new_new_n6623__ = ~new_new_n6408__ & new_new_n6446__;
  assign new_new_n6624__ = ~new_new_n6409__ & ~new_new_n6623__;
  assign new_new_n6625__ = ~new_new_n6373__ & ~new_new_n6376__;
  assign new_new_n6626__ = ~new_new_n6372__ & ~new_new_n6625__;
  assign new_new_n6627__ = ~new_new_n6511__ & ~new_new_n6522__;
  assign new_new_n6628__ = ~new_new_n6512__ & ~new_new_n6627__;
  assign new_new_n6629__ = ~new_new_n6418__ & ~new_new_n6423__;
  assign new_new_n6630__ = ~new_new_n6424__ & ~new_new_n6629__;
  assign new_new_n6631__ = new_new_n6361__ & ~new_new_n6366__;
  assign new_new_n6632__ = ~new_new_n6367__ & ~new_new_n6631__;
  assign new_new_n6633__ = ~new_new_n6630__ & ~new_new_n6632__;
  assign new_new_n6634__ = new_new_n6630__ & new_new_n6632__;
  assign new_new_n6635__ = ~new_new_n6633__ & ~new_new_n6634__;
  assign new_new_n6636__ = new_new_n6628__ & ~new_new_n6635__;
  assign new_new_n6637__ = ~new_new_n6628__ & new_new_n6635__;
  assign new_new_n6638__ = ~new_new_n6636__ & ~new_new_n6637__;
  assign new_new_n6639__ = new_new_n6626__ & ~new_new_n6638__;
  assign new_new_n6640__ = ~new_new_n6626__ & new_new_n6638__;
  assign new_new_n6641__ = ~new_new_n6639__ & ~new_new_n6640__;
  assign new_new_n6642__ = ~new_new_n6394__ & ~new_new_n6400__;
  assign new_new_n6643__ = ~new_new_n6399__ & ~new_new_n6642__;
  assign new_new_n6644__ = new_new_n6641__ & ~new_new_n6643__;
  assign new_new_n6645__ = ~new_new_n6641__ & new_new_n6643__;
  assign new_new_n6646__ = ~new_new_n6644__ & ~new_new_n6645__;
  assign new_new_n6647__ = ~new_new_n6566__ & ~new_new_n6646__;
  assign new_new_n6648__ = new_new_n6566__ & new_new_n6646__;
  assign new_new_n6649__ = ~new_new_n6647__ & ~new_new_n6648__;
  assign new_new_n6650__ = ~new_new_n6526__ & ~new_new_n6530__;
  assign new_new_n6651__ = ~new_new_n6529__ & ~new_new_n6650__;
  assign new_new_n6652__ = ~new_new_n6535__ & ~new_new_n6539__;
  assign new_new_n6653__ = ~new_new_n6538__ & ~new_new_n6652__;
  assign new_new_n6654__ = ~new_new_n6651__ & ~new_new_n6653__;
  assign new_new_n6655__ = new_new_n6651__ & new_new_n6653__;
  assign new_new_n6656__ = ~new_new_n6654__ & ~new_new_n6655__;
  assign new_new_n6657__ = ~new_new_n6465__ & ~new_new_n6469__;
  assign new_new_n6658__ = ~new_new_n6468__ & ~new_new_n6657__;
  assign new_new_n6659__ = ~new_new_n6656__ & new_new_n6658__;
  assign new_new_n6660__ = ~new_new_n6655__ & ~new_new_n6658__;
  assign new_new_n6661__ = ~new_new_n6654__ & new_new_n6660__;
  assign new_new_n6662__ = ~new_new_n6659__ & ~new_new_n6661__;
  assign new_new_n6663__ = ~new_new_n6544__ & ~new_new_n6555__;
  assign new_new_n6664__ = ~new_new_n6545__ & ~new_new_n6663__;
  assign new_new_n6665__ = new_new_n6662__ & new_new_n6664__;
  assign new_new_n6666__ = ~new_new_n6662__ & ~new_new_n6664__;
  assign new_new_n6667__ = ~new_new_n6665__ & ~new_new_n6666__;
  assign new_new_n6668__ = ~new_new_n6503__ & ~new_new_n6504__;
  assign new_new_n6669__ = new_new_n6506__ & ~new_new_n6668__;
  assign new_new_n6670__ = ~new_new_n6494__ & ~new_new_n6498__;
  assign new_new_n6671__ = ~new_new_n6497__ & ~new_new_n6670__;
  assign new_new_n6672__ = ~new_new_n6514__ & ~new_new_n6518__;
  assign new_new_n6673__ = ~new_new_n6517__ & ~new_new_n6672__;
  assign new_new_n6674__ = ~new_new_n6671__ & ~new_new_n6673__;
  assign new_new_n6675__ = new_new_n6671__ & new_new_n6673__;
  assign new_new_n6676__ = ~new_new_n6674__ & ~new_new_n6675__;
  assign new_new_n6677__ = new_new_n6669__ & ~new_new_n6676__;
  assign new_new_n6678__ = ~new_new_n6669__ & new_new_n6676__;
  assign new_new_n6679__ = ~new_new_n6677__ & ~new_new_n6678__;
  assign new_new_n6680__ = new_new_n6667__ & ~new_new_n6679__;
  assign new_new_n6681__ = ~new_new_n6667__ & new_new_n6679__;
  assign new_new_n6682__ = ~new_new_n6680__ & ~new_new_n6681__;
  assign new_new_n6683__ = ~new_new_n6483__ & ~new_new_n6490__;
  assign new_new_n6684__ = ~new_new_n6484__ & ~new_new_n6683__;
  assign new_new_n6685__ = ~new_new_n6415__ & ~new_new_n6428__;
  assign new_new_n6686__ = ~new_new_n6414__ & ~new_new_n6685__;
  assign new_new_n6687__ = new_new_n6684__ & new_new_n6686__;
  assign new_new_n6688__ = ~new_new_n6684__ & ~new_new_n6686__;
  assign new_new_n6689__ = ~new_new_n6687__ & ~new_new_n6688__;
  assign new_new_n6690__ = ~new_new_n6474__ & ~new_new_n6478__;
  assign new_new_n6691__ = ~new_new_n6477__ & ~new_new_n6690__;
  assign new_new_n6692__ = ~new_new_n6547__ & ~new_new_n6551__;
  assign new_new_n6693__ = ~new_new_n6550__ & ~new_new_n6692__;
  assign new_new_n6694__ = ~new_new_n6691__ & ~new_new_n6693__;
  assign new_new_n6695__ = new_new_n6691__ & new_new_n6693__;
  assign new_new_n6696__ = ~new_new_n6694__ & ~new_new_n6695__;
  assign new_new_n6697__ = pi04 & pi47;
  assign new_new_n6698__ = pi03 & pi48;
  assign new_new_n6699__ = pi02 & pi49;
  assign new_new_n6700__ = ~new_new_n6698__ & ~new_new_n6699__;
  assign new_new_n6701__ = new_new_n6698__ & new_new_n6699__;
  assign new_new_n6702__ = ~new_new_n6700__ & ~new_new_n6701__;
  assign new_new_n6703__ = new_new_n6697__ & ~new_new_n6702__;
  assign new_new_n6704__ = ~new_new_n6697__ & new_new_n6702__;
  assign new_new_n6705__ = ~new_new_n6703__ & ~new_new_n6704__;
  assign new_new_n6706__ = ~new_new_n6696__ & new_new_n6705__;
  assign new_new_n6707__ = new_new_n6696__ & ~new_new_n6705__;
  assign new_new_n6708__ = ~new_new_n6706__ & ~new_new_n6707__;
  assign new_new_n6709__ = new_new_n6689__ & new_new_n6708__;
  assign new_new_n6710__ = ~new_new_n6689__ & ~new_new_n6708__;
  assign new_new_n6711__ = ~new_new_n6709__ & ~new_new_n6710__;
  assign new_new_n6712__ = new_new_n6682__ & new_new_n6711__;
  assign new_new_n6713__ = ~new_new_n6682__ & ~new_new_n6711__;
  assign new_new_n6714__ = ~new_new_n6712__ & ~new_new_n6713__;
  assign new_new_n6715__ = ~new_new_n6525__ & ~new_new_n6558__;
  assign new_new_n6716__ = new_new_n6525__ & new_new_n6558__;
  assign new_new_n6717__ = ~new_new_n6493__ & ~new_new_n6716__;
  assign new_new_n6718__ = ~new_new_n6715__ & ~new_new_n6717__;
  assign new_new_n6719__ = new_new_n6714__ & new_new_n6718__;
  assign new_new_n6720__ = ~new_new_n6714__ & ~new_new_n6718__;
  assign new_new_n6721__ = ~new_new_n6719__ & ~new_new_n6720__;
  assign new_new_n6722__ = new_new_n6649__ & ~new_new_n6721__;
  assign new_new_n6723__ = ~new_new_n6649__ & new_new_n6721__;
  assign new_new_n6724__ = ~new_new_n6722__ & ~new_new_n6723__;
  assign new_new_n6725__ = pi12 & pi39;
  assign new_new_n6726__ = pi09 & pi42;
  assign new_new_n6727__ = pi10 & pi41;
  assign new_new_n6728__ = ~new_new_n6726__ & ~new_new_n6727__;
  assign new_new_n6729__ = new_new_n6726__ & new_new_n6727__;
  assign new_new_n6730__ = ~new_new_n6728__ & ~new_new_n6729__;
  assign new_new_n6731__ = new_new_n6725__ & ~new_new_n6730__;
  assign new_new_n6732__ = ~new_new_n6725__ & new_new_n6730__;
  assign new_new_n6733__ = ~new_new_n6731__ & ~new_new_n6732__;
  assign new_new_n6734__ = pi25 & pi26;
  assign new_new_n6735__ = pi11 & pi40;
  assign new_new_n6736__ = pi24 & pi27;
  assign new_new_n6737__ = ~new_new_n6735__ & ~new_new_n6736__;
  assign new_new_n6738__ = new_new_n6735__ & new_new_n6736__;
  assign new_new_n6739__ = ~new_new_n6737__ & ~new_new_n6738__;
  assign new_new_n6740__ = new_new_n6734__ & ~new_new_n6739__;
  assign new_new_n6741__ = ~new_new_n6734__ & new_new_n6739__;
  assign new_new_n6742__ = ~new_new_n6740__ & ~new_new_n6741__;
  assign new_new_n6743__ = new_new_n6733__ & new_new_n6742__;
  assign new_new_n6744__ = ~new_new_n6733__ & ~new_new_n6742__;
  assign new_new_n6745__ = ~new_new_n6743__ & ~new_new_n6744__;
  assign new_new_n6746__ = pi13 & pi38;
  assign new_new_n6747__ = pi07 & pi44;
  assign new_new_n6748__ = pi08 & pi43;
  assign new_new_n6749__ = ~new_new_n6747__ & ~new_new_n6748__;
  assign new_new_n6750__ = new_new_n6747__ & new_new_n6748__;
  assign new_new_n6751__ = ~new_new_n6749__ & ~new_new_n6750__;
  assign new_new_n6752__ = new_new_n6746__ & ~new_new_n6751__;
  assign new_new_n6753__ = ~new_new_n6746__ & new_new_n6751__;
  assign new_new_n6754__ = ~new_new_n6752__ & ~new_new_n6753__;
  assign new_new_n6755__ = ~new_new_n6745__ & new_new_n6754__;
  assign new_new_n6756__ = new_new_n6745__ & ~new_new_n6754__;
  assign new_new_n6757__ = ~new_new_n6755__ & ~new_new_n6756__;
  assign new_new_n6758__ = pi15 & pi36;
  assign new_new_n6759__ = pi14 & pi37;
  assign new_new_n6760__ = pi06 & pi45;
  assign new_new_n6761__ = ~new_new_n6759__ & ~new_new_n6760__;
  assign new_new_n6762__ = new_new_n6759__ & new_new_n6760__;
  assign new_new_n6763__ = ~new_new_n6761__ & ~new_new_n6762__;
  assign new_new_n6764__ = new_new_n6758__ & ~new_new_n6763__;
  assign new_new_n6765__ = ~new_new_n6758__ & new_new_n6763__;
  assign new_new_n6766__ = ~new_new_n6764__ & ~new_new_n6765__;
  assign new_new_n6767__ = pi18 & pi33;
  assign new_new_n6768__ = pi16 & pi35;
  assign new_new_n6769__ = pi05 & pi46;
  assign new_new_n6770__ = ~new_new_n6768__ & ~new_new_n6769__;
  assign new_new_n6771__ = new_new_n6768__ & new_new_n6769__;
  assign new_new_n6772__ = ~new_new_n6770__ & ~new_new_n6771__;
  assign new_new_n6773__ = new_new_n6767__ & ~new_new_n6772__;
  assign new_new_n6774__ = ~new_new_n6767__ & new_new_n6772__;
  assign new_new_n6775__ = ~new_new_n6773__ & ~new_new_n6774__;
  assign new_new_n6776__ = new_new_n6766__ & new_new_n6775__;
  assign new_new_n6777__ = ~new_new_n6766__ & ~new_new_n6775__;
  assign new_new_n6778__ = ~new_new_n6776__ & ~new_new_n6777__;
  assign new_new_n6779__ = pi23 & pi28;
  assign new_new_n6780__ = pi22 & pi29;
  assign new_new_n6781__ = pi21 & pi30;
  assign new_new_n6782__ = ~new_new_n6780__ & ~new_new_n6781__;
  assign new_new_n6783__ = new_new_n6780__ & new_new_n6781__;
  assign new_new_n6784__ = ~new_new_n6782__ & ~new_new_n6783__;
  assign new_new_n6785__ = new_new_n6779__ & ~new_new_n6784__;
  assign new_new_n6786__ = ~new_new_n6779__ & new_new_n6784__;
  assign new_new_n6787__ = ~new_new_n6785__ & ~new_new_n6786__;
  assign new_new_n6788__ = new_new_n6778__ & ~new_new_n6787__;
  assign new_new_n6789__ = ~new_new_n6778__ & new_new_n6787__;
  assign new_new_n6790__ = ~new_new_n6788__ & ~new_new_n6789__;
  assign new_new_n6791__ = ~new_new_n6757__ & ~new_new_n6790__;
  assign new_new_n6792__ = new_new_n6757__ & new_new_n6790__;
  assign new_new_n6793__ = ~new_new_n6791__ & ~new_new_n6792__;
  assign new_new_n6794__ = pi24 & pi49;
  assign new_new_n6795__ = pi00 & pi51;
  assign new_new_n6796__ = pi01 & ~pi50;
  assign new_new_n6797__ = ~new_new_n6795__ & ~new_new_n6796__;
  assign new_new_n6798__ = new_new_n6794__ & ~new_new_n6797__;
  assign new_new_n6799__ = pi26 & pi50;
  assign new_new_n6800__ = new_new_n6795__ & ~new_new_n6799__;
  assign new_new_n6801__ = new_new_n6798__ & ~new_new_n6800__;
  assign new_new_n6802__ = new_new_n6357__ & new_new_n6358__;
  assign new_new_n6803__ = pi01 & pi50;
  assign new_new_n6804__ = new_new_n6795__ & ~new_new_n6803__;
  assign new_new_n6805__ = ~new_new_n6795__ & new_new_n6803__;
  assign new_new_n6806__ = ~new_new_n6804__ & ~new_new_n6805__;
  assign new_new_n6807__ = pi26 & new_new_n6806__;
  assign new_new_n6808__ = ~pi26 & ~new_new_n6806__;
  assign new_new_n6809__ = ~new_new_n6802__ & ~new_new_n6807__;
  assign new_new_n6810__ = ~new_new_n6808__ & new_new_n6809__;
  assign new_new_n6811__ = ~new_new_n6801__ & ~new_new_n6810__;
  assign new_new_n6812__ = ~new_new_n6387__ & ~new_new_n6391__;
  assign new_new_n6813__ = ~new_new_n6388__ & ~new_new_n6812__;
  assign new_new_n6814__ = pi20 & pi31;
  assign new_new_n6815__ = pi19 & pi32;
  assign new_new_n6816__ = pi17 & pi34;
  assign new_new_n6817__ = ~new_new_n6815__ & ~new_new_n6816__;
  assign new_new_n6818__ = new_new_n6815__ & new_new_n6816__;
  assign new_new_n6819__ = ~new_new_n6817__ & ~new_new_n6818__;
  assign new_new_n6820__ = new_new_n6814__ & ~new_new_n6819__;
  assign new_new_n6821__ = ~new_new_n6814__ & new_new_n6819__;
  assign new_new_n6822__ = ~new_new_n6820__ & ~new_new_n6821__;
  assign new_new_n6823__ = new_new_n6813__ & ~new_new_n6822__;
  assign new_new_n6824__ = ~new_new_n6813__ & new_new_n6822__;
  assign new_new_n6825__ = ~new_new_n6823__ & ~new_new_n6824__;
  assign new_new_n6826__ = new_new_n6811__ & new_new_n6825__;
  assign new_new_n6827__ = ~new_new_n6811__ & ~new_new_n6825__;
  assign new_new_n6828__ = ~new_new_n6826__ & ~new_new_n6827__;
  assign new_new_n6829__ = new_new_n6793__ & ~new_new_n6828__;
  assign new_new_n6830__ = ~new_new_n6793__ & new_new_n6828__;
  assign new_new_n6831__ = ~new_new_n6829__ & ~new_new_n6830__;
  assign new_new_n6832__ = ~new_new_n6381__ & ~new_new_n6404__;
  assign new_new_n6833__ = ~new_new_n6380__ & ~new_new_n6832__;
  assign new_new_n6834__ = ~new_new_n6831__ & new_new_n6833__;
  assign new_new_n6835__ = new_new_n6831__ & ~new_new_n6833__;
  assign new_new_n6836__ = ~new_new_n6834__ & ~new_new_n6835__;
  assign new_new_n6837__ = ~new_new_n6440__ & ~new_new_n6443__;
  assign new_new_n6838__ = ~new_new_n6439__ & ~new_new_n6837__;
  assign new_new_n6839__ = new_new_n6836__ & ~new_new_n6838__;
  assign new_new_n6840__ = ~new_new_n6836__ & new_new_n6838__;
  assign new_new_n6841__ = ~new_new_n6839__ & ~new_new_n6840__;
  assign new_new_n6842__ = ~new_new_n6724__ & ~new_new_n6841__;
  assign new_new_n6843__ = new_new_n6724__ & new_new_n6841__;
  assign new_new_n6844__ = ~new_new_n6624__ & ~new_new_n6842__;
  assign new_new_n6845__ = ~new_new_n6843__ & ~new_new_n6844__;
  assign new_new_n6846__ = ~new_new_n6842__ & new_new_n6845__;
  assign new_new_n6847__ = new_new_n6624__ & ~new_new_n6846__;
  assign new_new_n6848__ = ~new_new_n6843__ & new_new_n6844__;
  assign new_new_n6849__ = ~new_new_n6847__ & ~new_new_n6848__;
  assign new_new_n6850__ = new_new_n6622__ & ~new_new_n6849__;
  assign new_new_n6851__ = ~new_new_n6622__ & new_new_n6849__;
  assign po052 = ~new_new_n6850__ & ~new_new_n6851__;
  assign new_new_n6853__ = ~new_new_n6621__ & ~new_new_n6849__;
  assign new_new_n6854__ = ~new_new_n6620__ & ~new_new_n6853__;
  assign new_new_n6855__ = new_new_n6845__ & ~new_new_n6854__;
  assign new_new_n6856__ = ~new_new_n6845__ & new_new_n6854__;
  assign new_new_n6857__ = ~new_new_n6855__ & ~new_new_n6856__;
  assign new_new_n6858__ = ~new_new_n6647__ & new_new_n6721__;
  assign new_new_n6859__ = ~new_new_n6648__ & ~new_new_n6858__;
  assign new_new_n6860__ = ~new_new_n6798__ & ~new_new_n6804__;
  assign new_new_n6861__ = pi26 & ~new_new_n6860__;
  assign new_new_n6862__ = ~pi26 & new_new_n6795__;
  assign new_new_n6863__ = new_new_n6803__ & new_new_n6862__;
  assign new_new_n6864__ = ~new_new_n6861__ & ~new_new_n6863__;
  assign new_new_n6865__ = pi04 & pi48;
  assign new_new_n6866__ = pi00 & pi52;
  assign new_new_n6867__ = ~new_new_n6865__ & ~new_new_n6866__;
  assign new_new_n6868__ = new_new_n6865__ & new_new_n6866__;
  assign new_new_n6869__ = ~new_new_n6867__ & ~new_new_n6868__;
  assign new_new_n6870__ = new_new_n3722__ & ~new_new_n6869__;
  assign new_new_n6871__ = ~new_new_n3722__ & new_new_n6869__;
  assign new_new_n6872__ = ~new_new_n6870__ & ~new_new_n6871__;
  assign new_new_n6873__ = new_new_n6864__ & new_new_n6872__;
  assign new_new_n6874__ = ~new_new_n6864__ & ~new_new_n6872__;
  assign new_new_n6875__ = ~new_new_n6873__ & ~new_new_n6874__;
  assign new_new_n6876__ = ~new_new_n6725__ & ~new_new_n6729__;
  assign new_new_n6877__ = ~new_new_n6728__ & ~new_new_n6876__;
  assign new_new_n6878__ = new_new_n6875__ & new_new_n6877__;
  assign new_new_n6879__ = ~new_new_n6875__ & ~new_new_n6877__;
  assign new_new_n6880__ = ~new_new_n6878__ & ~new_new_n6879__;
  assign new_new_n6881__ = ~new_new_n6811__ & ~new_new_n6823__;
  assign new_new_n6882__ = ~new_new_n6824__ & ~new_new_n6881__;
  assign new_new_n6883__ = new_new_n6880__ & ~new_new_n6882__;
  assign new_new_n6884__ = ~new_new_n6880__ & new_new_n6882__;
  assign new_new_n6885__ = ~new_new_n6883__ & ~new_new_n6884__;
  assign new_new_n6886__ = new_new_n6628__ & ~new_new_n6634__;
  assign new_new_n6887__ = ~new_new_n6633__ & ~new_new_n6886__;
  assign new_new_n6888__ = ~new_new_n6746__ & ~new_new_n6750__;
  assign new_new_n6889__ = ~new_new_n6749__ & ~new_new_n6888__;
  assign new_new_n6890__ = ~new_new_n6776__ & ~new_new_n6787__;
  assign new_new_n6891__ = ~new_new_n6777__ & ~new_new_n6890__;
  assign new_new_n6892__ = new_new_n6889__ & ~new_new_n6891__;
  assign new_new_n6893__ = ~new_new_n6889__ & new_new_n6891__;
  assign new_new_n6894__ = ~new_new_n6892__ & ~new_new_n6893__;
  assign new_new_n6895__ = ~new_new_n6814__ & ~new_new_n6818__;
  assign new_new_n6896__ = ~new_new_n6817__ & ~new_new_n6895__;
  assign new_new_n6897__ = ~new_new_n6697__ & ~new_new_n6701__;
  assign new_new_n6898__ = ~new_new_n6700__ & ~new_new_n6897__;
  assign new_new_n6899__ = ~new_new_n6896__ & ~new_new_n6898__;
  assign new_new_n6900__ = new_new_n6896__ & new_new_n6898__;
  assign new_new_n6901__ = ~new_new_n6899__ & ~new_new_n6900__;
  assign new_new_n6902__ = ~new_new_n6758__ & ~new_new_n6762__;
  assign new_new_n6903__ = ~new_new_n6761__ & ~new_new_n6902__;
  assign new_new_n6904__ = ~new_new_n6767__ & ~new_new_n6771__;
  assign new_new_n6905__ = ~new_new_n6770__ & ~new_new_n6904__;
  assign new_new_n6906__ = ~new_new_n6779__ & ~new_new_n6783__;
  assign new_new_n6907__ = ~new_new_n6782__ & ~new_new_n6906__;
  assign new_new_n6908__ = new_new_n6905__ & ~new_new_n6907__;
  assign new_new_n6909__ = ~new_new_n6905__ & new_new_n6907__;
  assign new_new_n6910__ = ~new_new_n6908__ & ~new_new_n6909__;
  assign new_new_n6911__ = new_new_n6903__ & new_new_n6910__;
  assign new_new_n6912__ = ~new_new_n6903__ & ~new_new_n6910__;
  assign new_new_n6913__ = ~new_new_n6911__ & ~new_new_n6912__;
  assign new_new_n6914__ = new_new_n6901__ & ~new_new_n6913__;
  assign new_new_n6915__ = ~new_new_n6901__ & new_new_n6913__;
  assign new_new_n6916__ = ~new_new_n6914__ & ~new_new_n6915__;
  assign new_new_n6917__ = new_new_n6894__ & new_new_n6916__;
  assign new_new_n6918__ = ~new_new_n6894__ & ~new_new_n6916__;
  assign new_new_n6919__ = ~new_new_n6917__ & ~new_new_n6918__;
  assign new_new_n6920__ = new_new_n6887__ & new_new_n6919__;
  assign new_new_n6921__ = ~new_new_n6887__ & ~new_new_n6919__;
  assign new_new_n6922__ = ~new_new_n6920__ & ~new_new_n6921__;
  assign new_new_n6923__ = ~new_new_n6792__ & ~new_new_n6828__;
  assign new_new_n6924__ = ~new_new_n6791__ & ~new_new_n6923__;
  assign new_new_n6925__ = new_new_n6922__ & ~new_new_n6924__;
  assign new_new_n6926__ = ~new_new_n6922__ & new_new_n6924__;
  assign new_new_n6927__ = ~new_new_n6925__ & ~new_new_n6926__;
  assign new_new_n6928__ = new_new_n6885__ & new_new_n6927__;
  assign new_new_n6929__ = ~new_new_n6885__ & ~new_new_n6927__;
  assign new_new_n6930__ = ~new_new_n6928__ & ~new_new_n6929__;
  assign new_new_n6931__ = ~new_new_n6834__ & ~new_new_n6838__;
  assign new_new_n6932__ = ~new_new_n6835__ & ~new_new_n6931__;
  assign new_new_n6933__ = new_new_n6930__ & new_new_n6932__;
  assign new_new_n6934__ = ~new_new_n6930__ & ~new_new_n6932__;
  assign new_new_n6935__ = ~new_new_n6933__ & ~new_new_n6934__;
  assign new_new_n6936__ = ~new_new_n6744__ & new_new_n6754__;
  assign new_new_n6937__ = ~new_new_n6743__ & ~new_new_n6936__;
  assign new_new_n6938__ = ~new_new_n6734__ & ~new_new_n6738__;
  assign new_new_n6939__ = ~new_new_n6737__ & ~new_new_n6938__;
  assign new_new_n6940__ = pi25 & pi27;
  assign new_new_n6941__ = ~pi51 & ~new_new_n6799__;
  assign new_new_n6942__ = pi26 & pi51;
  assign new_new_n6943__ = pi50 & new_new_n6942__;
  assign new_new_n6944__ = pi01 & ~new_new_n6941__;
  assign new_new_n6945__ = ~new_new_n6943__ & new_new_n6944__;
  assign new_new_n6946__ = new_new_n6940__ & ~new_new_n6945__;
  assign new_new_n6947__ = ~new_new_n6940__ & new_new_n6945__;
  assign new_new_n6948__ = ~new_new_n6946__ & ~new_new_n6947__;
  assign new_new_n6949__ = new_new_n6939__ & new_new_n6948__;
  assign new_new_n6950__ = ~new_new_n6939__ & ~new_new_n6948__;
  assign new_new_n6951__ = ~new_new_n6949__ & ~new_new_n6950__;
  assign new_new_n6952__ = ~new_new_n6937__ & new_new_n6951__;
  assign new_new_n6953__ = new_new_n6937__ & ~new_new_n6951__;
  assign new_new_n6954__ = ~new_new_n6952__ & ~new_new_n6953__;
  assign new_new_n6955__ = ~new_new_n6695__ & new_new_n6705__;
  assign new_new_n6956__ = ~new_new_n6694__ & ~new_new_n6955__;
  assign new_new_n6957__ = new_new_n6954__ & ~new_new_n6956__;
  assign new_new_n6958__ = ~new_new_n6954__ & new_new_n6956__;
  assign new_new_n6959__ = ~new_new_n6957__ & ~new_new_n6958__;
  assign new_new_n6960__ = ~new_new_n6669__ & ~new_new_n6675__;
  assign new_new_n6961__ = ~new_new_n6674__ & ~new_new_n6960__;
  assign new_new_n6962__ = ~new_new_n6654__ & ~new_new_n6660__;
  assign new_new_n6963__ = pi19 & pi33;
  assign new_new_n6964__ = pi03 & pi49;
  assign new_new_n6965__ = pi02 & pi50;
  assign new_new_n6966__ = ~new_new_n6964__ & ~new_new_n6965__;
  assign new_new_n6967__ = new_new_n6964__ & new_new_n6965__;
  assign new_new_n6968__ = ~new_new_n6966__ & ~new_new_n6967__;
  assign new_new_n6969__ = new_new_n6963__ & ~new_new_n6968__;
  assign new_new_n6970__ = ~new_new_n6963__ & new_new_n6968__;
  assign new_new_n6971__ = ~new_new_n6969__ & ~new_new_n6970__;
  assign new_new_n6972__ = new_new_n6962__ & ~new_new_n6971__;
  assign new_new_n6973__ = ~new_new_n6962__ & new_new_n6971__;
  assign new_new_n6974__ = ~new_new_n6972__ & ~new_new_n6973__;
  assign new_new_n6975__ = new_new_n6961__ & new_new_n6974__;
  assign new_new_n6976__ = ~new_new_n6961__ & ~new_new_n6974__;
  assign new_new_n6977__ = ~new_new_n6975__ & ~new_new_n6976__;
  assign new_new_n6978__ = new_new_n6959__ & ~new_new_n6977__;
  assign new_new_n6979__ = ~new_new_n6959__ & new_new_n6977__;
  assign new_new_n6980__ = ~new_new_n6978__ & ~new_new_n6979__;
  assign new_new_n6981__ = ~new_new_n6688__ & ~new_new_n6708__;
  assign new_new_n6982__ = ~new_new_n6687__ & ~new_new_n6981__;
  assign new_new_n6983__ = new_new_n6980__ & new_new_n6982__;
  assign new_new_n6984__ = ~new_new_n6980__ & ~new_new_n6982__;
  assign new_new_n6985__ = ~new_new_n6983__ & ~new_new_n6984__;
  assign new_new_n6986__ = new_new_n6935__ & ~new_new_n6985__;
  assign new_new_n6987__ = ~new_new_n6935__ & new_new_n6985__;
  assign new_new_n6988__ = ~new_new_n6986__ & ~new_new_n6987__;
  assign new_new_n6989__ = new_new_n6859__ & new_new_n6988__;
  assign new_new_n6990__ = ~new_new_n6859__ & ~new_new_n6988__;
  assign new_new_n6991__ = ~new_new_n6989__ & ~new_new_n6990__;
  assign new_new_n6992__ = ~new_new_n6712__ & ~new_new_n6718__;
  assign new_new_n6993__ = ~new_new_n6713__ & ~new_new_n6992__;
  assign new_new_n6994__ = ~new_new_n6639__ & ~new_new_n6643__;
  assign new_new_n6995__ = ~new_new_n6640__ & ~new_new_n6994__;
  assign new_new_n6996__ = ~new_new_n6665__ & ~new_new_n6679__;
  assign new_new_n6997__ = ~new_new_n6666__ & ~new_new_n6996__;
  assign new_new_n6998__ = pi24 & pi28;
  assign new_new_n6999__ = pi22 & pi30;
  assign new_new_n7000__ = pi23 & pi29;
  assign new_new_n7001__ = ~new_new_n6999__ & ~new_new_n7000__;
  assign new_new_n7002__ = new_new_n6999__ & new_new_n7000__;
  assign new_new_n7003__ = ~new_new_n7001__ & ~new_new_n7002__;
  assign new_new_n7004__ = new_new_n6998__ & ~new_new_n7003__;
  assign new_new_n7005__ = ~new_new_n6998__ & new_new_n7003__;
  assign new_new_n7006__ = ~new_new_n7004__ & ~new_new_n7005__;
  assign new_new_n7007__ = pi21 & pi31;
  assign new_new_n7008__ = pi20 & pi32;
  assign new_new_n7009__ = ~new_new_n3345__ & ~new_new_n7008__;
  assign new_new_n7010__ = new_new_n3345__ & new_new_n7008__;
  assign new_new_n7011__ = ~new_new_n7009__ & ~new_new_n7010__;
  assign new_new_n7012__ = new_new_n7007__ & ~new_new_n7011__;
  assign new_new_n7013__ = ~new_new_n7007__ & new_new_n7011__;
  assign new_new_n7014__ = ~new_new_n7012__ & ~new_new_n7013__;
  assign new_new_n7015__ = new_new_n7006__ & new_new_n7014__;
  assign new_new_n7016__ = ~new_new_n7006__ & ~new_new_n7014__;
  assign new_new_n7017__ = ~new_new_n7015__ & ~new_new_n7016__;
  assign new_new_n7018__ = pi14 & pi38;
  assign new_new_n7019__ = pi13 & pi39;
  assign new_new_n7020__ = pi09 & pi43;
  assign new_new_n7021__ = ~new_new_n7019__ & ~new_new_n7020__;
  assign new_new_n7022__ = new_new_n7019__ & new_new_n7020__;
  assign new_new_n7023__ = ~new_new_n7021__ & ~new_new_n7022__;
  assign new_new_n7024__ = new_new_n7018__ & ~new_new_n7023__;
  assign new_new_n7025__ = ~new_new_n7018__ & new_new_n7023__;
  assign new_new_n7026__ = ~new_new_n7024__ & ~new_new_n7025__;
  assign new_new_n7027__ = new_new_n7017__ & ~new_new_n7026__;
  assign new_new_n7028__ = ~new_new_n7017__ & new_new_n7026__;
  assign new_new_n7029__ = ~new_new_n7027__ & ~new_new_n7028__;
  assign new_new_n7030__ = ~new_new_n6997__ & new_new_n7029__;
  assign new_new_n7031__ = new_new_n6997__ & ~new_new_n7029__;
  assign new_new_n7032__ = ~new_new_n7030__ & ~new_new_n7031__;
  assign new_new_n7033__ = pi16 & pi36;
  assign new_new_n7034__ = pi06 & pi46;
  assign new_new_n7035__ = pi05 & pi47;
  assign new_new_n7036__ = ~new_new_n7034__ & ~new_new_n7035__;
  assign new_new_n7037__ = new_new_n7034__ & new_new_n7035__;
  assign new_new_n7038__ = ~new_new_n7036__ & ~new_new_n7037__;
  assign new_new_n7039__ = new_new_n7033__ & ~new_new_n7038__;
  assign new_new_n7040__ = ~new_new_n7033__ & new_new_n7038__;
  assign new_new_n7041__ = ~new_new_n7039__ & ~new_new_n7040__;
  assign new_new_n7042__ = pi12 & pi40;
  assign new_new_n7043__ = pi10 & pi42;
  assign new_new_n7044__ = pi11 & pi41;
  assign new_new_n7045__ = ~new_new_n7043__ & ~new_new_n7044__;
  assign new_new_n7046__ = new_new_n7043__ & new_new_n7044__;
  assign new_new_n7047__ = ~new_new_n7045__ & ~new_new_n7046__;
  assign new_new_n7048__ = new_new_n7042__ & ~new_new_n7047__;
  assign new_new_n7049__ = ~new_new_n7042__ & new_new_n7047__;
  assign new_new_n7050__ = ~new_new_n7048__ & ~new_new_n7049__;
  assign new_new_n7051__ = new_new_n7041__ & new_new_n7050__;
  assign new_new_n7052__ = ~new_new_n7041__ & ~new_new_n7050__;
  assign new_new_n7053__ = ~new_new_n7051__ & ~new_new_n7052__;
  assign new_new_n7054__ = pi15 & pi37;
  assign new_new_n7055__ = pi08 & pi44;
  assign new_new_n7056__ = pi07 & pi45;
  assign new_new_n7057__ = ~new_new_n7055__ & ~new_new_n7056__;
  assign new_new_n7058__ = new_new_n7055__ & new_new_n7056__;
  assign new_new_n7059__ = ~new_new_n7057__ & ~new_new_n7058__;
  assign new_new_n7060__ = new_new_n7054__ & ~new_new_n7059__;
  assign new_new_n7061__ = ~new_new_n7054__ & new_new_n7059__;
  assign new_new_n7062__ = ~new_new_n7060__ & ~new_new_n7061__;
  assign new_new_n7063__ = new_new_n7053__ & ~new_new_n7062__;
  assign new_new_n7064__ = ~new_new_n7053__ & new_new_n7062__;
  assign new_new_n7065__ = ~new_new_n7063__ & ~new_new_n7064__;
  assign new_new_n7066__ = new_new_n7032__ & ~new_new_n7065__;
  assign new_new_n7067__ = ~new_new_n7032__ & new_new_n7065__;
  assign new_new_n7068__ = ~new_new_n7066__ & ~new_new_n7067__;
  assign new_new_n7069__ = ~new_new_n6995__ & ~new_new_n7068__;
  assign new_new_n7070__ = new_new_n6995__ & new_new_n7068__;
  assign new_new_n7071__ = ~new_new_n7069__ & ~new_new_n7070__;
  assign new_new_n7072__ = new_new_n6993__ & ~new_new_n7071__;
  assign new_new_n7073__ = ~new_new_n6993__ & new_new_n7071__;
  assign new_new_n7074__ = ~new_new_n7072__ & ~new_new_n7073__;
  assign new_new_n7075__ = new_new_n6991__ & ~new_new_n7074__;
  assign new_new_n7076__ = ~new_new_n6991__ & new_new_n7074__;
  assign new_new_n7077__ = ~new_new_n7075__ & ~new_new_n7076__;
  assign new_new_n7078__ = new_new_n6857__ & new_new_n7077__;
  assign new_new_n7079__ = ~new_new_n6857__ & ~new_new_n7077__;
  assign po053 = ~new_new_n7078__ & ~new_new_n7079__;
  assign new_new_n7081__ = ~new_new_n6933__ & ~new_new_n6985__;
  assign new_new_n7082__ = ~new_new_n6934__ & ~new_new_n7081__;
  assign new_new_n7083__ = ~new_new_n6961__ & ~new_new_n6972__;
  assign new_new_n7084__ = ~new_new_n6973__ & ~new_new_n7083__;
  assign new_new_n7085__ = pi15 & pi38;
  assign new_new_n7086__ = pi06 & pi47;
  assign new_new_n7087__ = pi07 & pi46;
  assign new_new_n7088__ = ~new_new_n7086__ & ~new_new_n7087__;
  assign new_new_n7089__ = new_new_n7086__ & new_new_n7087__;
  assign new_new_n7090__ = ~new_new_n7088__ & ~new_new_n7089__;
  assign new_new_n7091__ = new_new_n7085__ & ~new_new_n7090__;
  assign new_new_n7092__ = ~new_new_n7085__ & new_new_n7090__;
  assign new_new_n7093__ = ~new_new_n7091__ & ~new_new_n7092__;
  assign new_new_n7094__ = pi14 & pi39;
  assign new_new_n7095__ = pi08 & pi45;
  assign new_new_n7096__ = pi09 & pi44;
  assign new_new_n7097__ = ~new_new_n7095__ & ~new_new_n7096__;
  assign new_new_n7098__ = new_new_n7095__ & new_new_n7096__;
  assign new_new_n7099__ = ~new_new_n7097__ & ~new_new_n7098__;
  assign new_new_n7100__ = new_new_n7094__ & ~new_new_n7099__;
  assign new_new_n7101__ = ~new_new_n7094__ & new_new_n7099__;
  assign new_new_n7102__ = ~new_new_n7100__ & ~new_new_n7101__;
  assign new_new_n7103__ = new_new_n7093__ & new_new_n7102__;
  assign new_new_n7104__ = ~new_new_n7093__ & ~new_new_n7102__;
  assign new_new_n7105__ = ~new_new_n7103__ & ~new_new_n7104__;
  assign new_new_n7106__ = pi16 & pi37;
  assign new_new_n7107__ = pi05 & pi48;
  assign new_new_n7108__ = pi00 & pi53;
  assign new_new_n7109__ = ~new_new_n7107__ & ~new_new_n7108__;
  assign new_new_n7110__ = new_new_n7107__ & new_new_n7108__;
  assign new_new_n7111__ = ~new_new_n7109__ & ~new_new_n7110__;
  assign new_new_n7112__ = new_new_n7106__ & ~new_new_n7111__;
  assign new_new_n7113__ = ~new_new_n7106__ & new_new_n7111__;
  assign new_new_n7114__ = ~new_new_n7112__ & ~new_new_n7113__;
  assign new_new_n7115__ = ~new_new_n7105__ & new_new_n7114__;
  assign new_new_n7116__ = new_new_n7105__ & ~new_new_n7114__;
  assign new_new_n7117__ = ~new_new_n7115__ & ~new_new_n7116__;
  assign new_new_n7118__ = ~new_new_n7084__ & ~new_new_n7117__;
  assign new_new_n7119__ = new_new_n7084__ & new_new_n7117__;
  assign new_new_n7120__ = ~new_new_n7118__ & ~new_new_n7119__;
  assign new_new_n7121__ = pi18 & pi35;
  assign new_new_n7122__ = pi04 & pi49;
  assign new_new_n7123__ = pi17 & pi36;
  assign new_new_n7124__ = ~new_new_n7122__ & ~new_new_n7123__;
  assign new_new_n7125__ = new_new_n7122__ & new_new_n7123__;
  assign new_new_n7126__ = ~new_new_n7124__ & ~new_new_n7125__;
  assign new_new_n7127__ = new_new_n7121__ & ~new_new_n7126__;
  assign new_new_n7128__ = ~new_new_n7121__ & new_new_n7126__;
  assign new_new_n7129__ = ~new_new_n7127__ & ~new_new_n7128__;
  assign new_new_n7130__ = pi03 & pi50;
  assign new_new_n7131__ = pi27 & new_new_n1907__;
  assign new_new_n7132__ = ~pi02 & ~new_new_n7131__;
  assign new_new_n7133__ = pi51 & ~new_new_n7132__;
  assign new_new_n7134__ = pi27 & new_new_n6504__;
  assign new_new_n7135__ = new_new_n7133__ & ~new_new_n7134__;
  assign new_new_n7136__ = new_new_n7130__ & ~new_new_n7135__;
  assign new_new_n7137__ = ~new_new_n7130__ & new_new_n7135__;
  assign new_new_n7138__ = ~new_new_n7136__ & ~new_new_n7137__;
  assign new_new_n7139__ = pi21 & pi32;
  assign new_new_n7140__ = pi19 & pi34;
  assign new_new_n7141__ = pi20 & pi33;
  assign new_new_n7142__ = ~new_new_n7140__ & ~new_new_n7141__;
  assign new_new_n7143__ = new_new_n7140__ & new_new_n7141__;
  assign new_new_n7144__ = ~new_new_n7142__ & ~new_new_n7143__;
  assign new_new_n7145__ = new_new_n7139__ & ~new_new_n7144__;
  assign new_new_n7146__ = ~new_new_n7139__ & new_new_n7144__;
  assign new_new_n7147__ = ~new_new_n7145__ & ~new_new_n7146__;
  assign new_new_n7148__ = new_new_n7138__ & new_new_n7147__;
  assign new_new_n7149__ = ~new_new_n7138__ & ~new_new_n7147__;
  assign new_new_n7150__ = ~new_new_n7148__ & ~new_new_n7149__;
  assign new_new_n7151__ = new_new_n7129__ & new_new_n7150__;
  assign new_new_n7152__ = ~new_new_n7129__ & ~new_new_n7150__;
  assign new_new_n7153__ = ~new_new_n7151__ & ~new_new_n7152__;
  assign new_new_n7154__ = new_new_n7120__ & ~new_new_n7153__;
  assign new_new_n7155__ = ~new_new_n7120__ & new_new_n7153__;
  assign new_new_n7156__ = ~new_new_n7154__ & ~new_new_n7155__;
  assign new_new_n7157__ = ~new_new_n6919__ & ~new_new_n6924__;
  assign new_new_n7158__ = new_new_n6919__ & new_new_n6924__;
  assign new_new_n7159__ = new_new_n6885__ & ~new_new_n6887__;
  assign new_new_n7160__ = ~new_new_n6885__ & new_new_n6887__;
  assign new_new_n7161__ = ~new_new_n7159__ & ~new_new_n7160__;
  assign new_new_n7162__ = ~new_new_n7158__ & ~new_new_n7161__;
  assign new_new_n7163__ = ~new_new_n7157__ & ~new_new_n7162__;
  assign new_new_n7164__ = new_new_n7156__ & new_new_n7163__;
  assign new_new_n7165__ = ~new_new_n7156__ & ~new_new_n7163__;
  assign new_new_n7166__ = ~new_new_n7164__ & ~new_new_n7165__;
  assign new_new_n7167__ = ~new_new_n6953__ & ~new_new_n6956__;
  assign new_new_n7168__ = ~new_new_n6952__ & ~new_new_n7167__;
  assign new_new_n7169__ = new_new_n6901__ & ~new_new_n6903__;
  assign new_new_n7170__ = ~new_new_n6901__ & new_new_n6903__;
  assign new_new_n7171__ = ~new_new_n7169__ & ~new_new_n7170__;
  assign new_new_n7172__ = new_new_n6891__ & new_new_n7171__;
  assign new_new_n7173__ = ~new_new_n6891__ & ~new_new_n7171__;
  assign new_new_n7174__ = new_new_n6889__ & new_new_n6910__;
  assign new_new_n7175__ = ~new_new_n6889__ & ~new_new_n6910__;
  assign new_new_n7176__ = ~new_new_n7174__ & ~new_new_n7175__;
  assign new_new_n7177__ = ~new_new_n7173__ & new_new_n7176__;
  assign new_new_n7178__ = ~new_new_n7172__ & ~new_new_n7177__;
  assign new_new_n7179__ = ~new_new_n7168__ & ~new_new_n7178__;
  assign new_new_n7180__ = new_new_n7168__ & new_new_n7178__;
  assign new_new_n7181__ = ~new_new_n7179__ & ~new_new_n7180__;
  assign new_new_n7182__ = pi24 & pi29;
  assign new_new_n7183__ = pi23 & pi30;
  assign new_new_n7184__ = pi22 & pi31;
  assign new_new_n7185__ = ~new_new_n7183__ & ~new_new_n7184__;
  assign new_new_n7186__ = new_new_n7183__ & new_new_n7184__;
  assign new_new_n7187__ = ~new_new_n7185__ & ~new_new_n7186__;
  assign new_new_n7188__ = new_new_n7182__ & ~new_new_n7187__;
  assign new_new_n7189__ = ~new_new_n7182__ & new_new_n7187__;
  assign new_new_n7190__ = ~new_new_n7188__ & ~new_new_n7189__;
  assign new_new_n7191__ = pi13 & pi40;
  assign new_new_n7192__ = pi12 & pi41;
  assign new_new_n7193__ = pi10 & pi43;
  assign new_new_n7194__ = ~new_new_n7192__ & ~new_new_n7193__;
  assign new_new_n7195__ = new_new_n7192__ & new_new_n7193__;
  assign new_new_n7196__ = ~new_new_n7194__ & ~new_new_n7195__;
  assign new_new_n7197__ = new_new_n7191__ & ~new_new_n7196__;
  assign new_new_n7198__ = ~new_new_n7191__ & new_new_n7196__;
  assign new_new_n7199__ = ~new_new_n7197__ & ~new_new_n7198__;
  assign new_new_n7200__ = new_new_n7190__ & new_new_n7199__;
  assign new_new_n7201__ = ~new_new_n7190__ & ~new_new_n7199__;
  assign new_new_n7202__ = ~new_new_n7200__ & ~new_new_n7201__;
  assign new_new_n7203__ = pi26 & pi27;
  assign new_new_n7204__ = pi11 & pi42;
  assign new_new_n7205__ = pi25 & pi28;
  assign new_new_n7206__ = ~new_new_n7204__ & ~new_new_n7205__;
  assign new_new_n7207__ = new_new_n7204__ & new_new_n7205__;
  assign new_new_n7208__ = ~new_new_n7206__ & ~new_new_n7207__;
  assign new_new_n7209__ = new_new_n7203__ & ~new_new_n7208__;
  assign new_new_n7210__ = ~new_new_n7203__ & new_new_n7208__;
  assign new_new_n7211__ = ~new_new_n7209__ & ~new_new_n7210__;
  assign new_new_n7212__ = new_new_n7202__ & ~new_new_n7211__;
  assign new_new_n7213__ = ~new_new_n7202__ & new_new_n7211__;
  assign new_new_n7214__ = ~new_new_n7212__ & ~new_new_n7213__;
  assign new_new_n7215__ = new_new_n7181__ & new_new_n7214__;
  assign new_new_n7216__ = ~new_new_n7181__ & ~new_new_n7214__;
  assign new_new_n7217__ = ~new_new_n7215__ & ~new_new_n7216__;
  assign new_new_n7218__ = new_new_n7166__ & ~new_new_n7217__;
  assign new_new_n7219__ = ~new_new_n7166__ & new_new_n7217__;
  assign new_new_n7220__ = ~new_new_n7218__ & ~new_new_n7219__;
  assign new_new_n7221__ = new_new_n7082__ & ~new_new_n7220__;
  assign new_new_n7222__ = ~new_new_n7082__ & new_new_n7220__;
  assign new_new_n7223__ = ~new_new_n7221__ & ~new_new_n7222__;
  assign new_new_n7224__ = new_new_n6993__ & ~new_new_n7070__;
  assign new_new_n7225__ = ~new_new_n7069__ & ~new_new_n7224__;
  assign new_new_n7226__ = ~new_new_n7015__ & ~new_new_n7026__;
  assign new_new_n7227__ = ~new_new_n7016__ & ~new_new_n7226__;
  assign new_new_n7228__ = ~new_new_n6874__ & ~new_new_n6877__;
  assign new_new_n7229__ = ~new_new_n6873__ & ~new_new_n7228__;
  assign new_new_n7230__ = ~new_new_n7227__ & new_new_n7229__;
  assign new_new_n7231__ = new_new_n7227__ & ~new_new_n7229__;
  assign new_new_n7232__ = ~new_new_n7230__ & ~new_new_n7231__;
  assign new_new_n7233__ = ~new_new_n3722__ & ~new_new_n6868__;
  assign new_new_n7234__ = ~new_new_n6867__ & ~new_new_n7233__;
  assign new_new_n7235__ = ~new_new_n6963__ & ~new_new_n6967__;
  assign new_new_n7236__ = ~new_new_n6966__ & ~new_new_n7235__;
  assign new_new_n7237__ = ~new_new_n6998__ & ~new_new_n7002__;
  assign new_new_n7238__ = ~new_new_n7001__ & ~new_new_n7237__;
  assign new_new_n7239__ = ~new_new_n7236__ & ~new_new_n7238__;
  assign new_new_n7240__ = new_new_n7236__ & new_new_n7238__;
  assign new_new_n7241__ = ~new_new_n7239__ & ~new_new_n7240__;
  assign new_new_n7242__ = new_new_n7234__ & ~new_new_n7241__;
  assign new_new_n7243__ = ~new_new_n7234__ & new_new_n7241__;
  assign new_new_n7244__ = ~new_new_n7242__ & ~new_new_n7243__;
  assign new_new_n7245__ = new_new_n7232__ & new_new_n7244__;
  assign new_new_n7246__ = ~new_new_n7232__ & ~new_new_n7244__;
  assign new_new_n7247__ = ~new_new_n7245__ & ~new_new_n7246__;
  assign new_new_n7248__ = ~new_new_n7007__ & ~new_new_n7010__;
  assign new_new_n7249__ = ~new_new_n7009__ & ~new_new_n7248__;
  assign new_new_n7250__ = ~new_new_n7054__ & ~new_new_n7058__;
  assign new_new_n7251__ = ~new_new_n7057__ & ~new_new_n7250__;
  assign new_new_n7252__ = new_new_n7249__ & new_new_n7251__;
  assign new_new_n7253__ = ~new_new_n7249__ & ~new_new_n7251__;
  assign new_new_n7254__ = ~new_new_n7252__ & ~new_new_n7253__;
  assign new_new_n7255__ = ~new_new_n7033__ & ~new_new_n7037__;
  assign new_new_n7256__ = ~new_new_n7036__ & ~new_new_n7255__;
  assign new_new_n7257__ = ~new_new_n7254__ & new_new_n7256__;
  assign new_new_n7258__ = ~new_new_n7252__ & ~new_new_n7256__;
  assign new_new_n7259__ = ~new_new_n7253__ & new_new_n7258__;
  assign new_new_n7260__ = ~new_new_n7257__ & ~new_new_n7259__;
  assign new_new_n7261__ = ~new_new_n7051__ & ~new_new_n7062__;
  assign new_new_n7262__ = ~new_new_n7052__ & ~new_new_n7261__;
  assign new_new_n7263__ = pi52 & new_new_n2384__;
  assign new_new_n7264__ = pi01 & pi52;
  assign new_new_n7265__ = ~pi27 & ~new_new_n7264__;
  assign new_new_n7266__ = ~new_new_n7263__ & ~new_new_n7265__;
  assign new_new_n7267__ = ~new_new_n7018__ & ~new_new_n7022__;
  assign new_new_n7268__ = ~new_new_n7021__ & ~new_new_n7267__;
  assign new_new_n7269__ = ~new_new_n7042__ & ~new_new_n7046__;
  assign new_new_n7270__ = ~new_new_n7045__ & ~new_new_n7269__;
  assign new_new_n7271__ = ~new_new_n7268__ & ~new_new_n7270__;
  assign new_new_n7272__ = new_new_n7268__ & new_new_n7270__;
  assign new_new_n7273__ = ~new_new_n7271__ & ~new_new_n7272__;
  assign new_new_n7274__ = new_new_n7266__ & ~new_new_n7273__;
  assign new_new_n7275__ = ~new_new_n7266__ & new_new_n7273__;
  assign new_new_n7276__ = ~new_new_n7274__ & ~new_new_n7275__;
  assign new_new_n7277__ = ~new_new_n7262__ & ~new_new_n7276__;
  assign new_new_n7278__ = new_new_n7262__ & new_new_n7276__;
  assign new_new_n7279__ = ~new_new_n7277__ & ~new_new_n7278__;
  assign new_new_n7280__ = ~new_new_n7260__ & new_new_n7279__;
  assign new_new_n7281__ = new_new_n7260__ & ~new_new_n7279__;
  assign new_new_n7282__ = ~new_new_n7280__ & ~new_new_n7281__;
  assign new_new_n7283__ = new_new_n7247__ & ~new_new_n7282__;
  assign new_new_n7284__ = ~new_new_n7247__ & new_new_n7282__;
  assign new_new_n7285__ = ~new_new_n7283__ & ~new_new_n7284__;
  assign new_new_n7286__ = ~new_new_n6979__ & ~new_new_n6982__;
  assign new_new_n7287__ = ~new_new_n6978__ & ~new_new_n7286__;
  assign new_new_n7288__ = new_new_n7285__ & new_new_n7287__;
  assign new_new_n7289__ = ~new_new_n7285__ & ~new_new_n7287__;
  assign new_new_n7290__ = ~new_new_n7288__ & ~new_new_n7289__;
  assign new_new_n7291__ = new_new_n7225__ & ~new_new_n7290__;
  assign new_new_n7292__ = ~new_new_n7225__ & new_new_n7290__;
  assign new_new_n7293__ = ~new_new_n7291__ & ~new_new_n7292__;
  assign new_new_n7294__ = ~new_new_n7030__ & ~new_new_n7065__;
  assign new_new_n7295__ = ~new_new_n7031__ & ~new_new_n7294__;
  assign new_new_n7296__ = ~new_new_n6900__ & ~new_new_n6903__;
  assign new_new_n7297__ = ~new_new_n6899__ & ~new_new_n7296__;
  assign new_new_n7298__ = ~new_new_n6799__ & ~new_new_n6939__;
  assign new_new_n7299__ = pi51 & ~new_new_n6940__;
  assign new_new_n7300__ = ~new_new_n7298__ & new_new_n7299__;
  assign new_new_n7301__ = ~pi51 & new_new_n6940__;
  assign new_new_n7302__ = ~new_new_n6939__ & ~new_new_n7301__;
  assign new_new_n7303__ = new_new_n6799__ & ~new_new_n7302__;
  assign new_new_n7304__ = ~new_new_n7300__ & ~new_new_n7303__;
  assign new_new_n7305__ = pi01 & ~new_new_n7304__;
  assign new_new_n7306__ = pi01 & pi51;
  assign new_new_n7307__ = new_new_n6940__ & ~new_new_n7306__;
  assign new_new_n7308__ = new_new_n6939__ & new_new_n7307__;
  assign new_new_n7309__ = ~new_new_n7305__ & ~new_new_n7308__;
  assign new_new_n7310__ = ~new_new_n7297__ & new_new_n7309__;
  assign new_new_n7311__ = new_new_n7297__ & ~new_new_n7309__;
  assign new_new_n7312__ = ~new_new_n7310__ & ~new_new_n7311__;
  assign new_new_n7313__ = ~new_new_n6889__ & ~new_new_n6907__;
  assign new_new_n7314__ = new_new_n6889__ & new_new_n6907__;
  assign new_new_n7315__ = ~new_new_n6905__ & ~new_new_n7314__;
  assign new_new_n7316__ = ~new_new_n7313__ & ~new_new_n7315__;
  assign new_new_n7317__ = ~new_new_n7312__ & new_new_n7316__;
  assign new_new_n7318__ = new_new_n7312__ & ~new_new_n7316__;
  assign new_new_n7319__ = ~new_new_n7317__ & ~new_new_n7318__;
  assign new_new_n7320__ = ~new_new_n7295__ & new_new_n7319__;
  assign new_new_n7321__ = new_new_n7295__ & ~new_new_n7319__;
  assign new_new_n7322__ = ~new_new_n7320__ & ~new_new_n7321__;
  assign new_new_n7323__ = new_new_n6882__ & new_new_n6887__;
  assign new_new_n7324__ = ~new_new_n6882__ & ~new_new_n6887__;
  assign new_new_n7325__ = new_new_n6880__ & ~new_new_n7324__;
  assign new_new_n7326__ = ~new_new_n7323__ & ~new_new_n7325__;
  assign new_new_n7327__ = new_new_n7322__ & ~new_new_n7326__;
  assign new_new_n7328__ = ~new_new_n7322__ & new_new_n7326__;
  assign new_new_n7329__ = ~new_new_n7327__ & ~new_new_n7328__;
  assign new_new_n7330__ = new_new_n7293__ & ~new_new_n7329__;
  assign new_new_n7331__ = ~new_new_n7293__ & new_new_n7329__;
  assign new_new_n7332__ = ~new_new_n7330__ & ~new_new_n7331__;
  assign new_new_n7333__ = new_new_n7223__ & new_new_n7332__;
  assign new_new_n7334__ = ~new_new_n7223__ & ~new_new_n7332__;
  assign new_new_n7335__ = ~new_new_n7333__ & ~new_new_n7334__;
  assign new_new_n7336__ = new_new_n6989__ & new_new_n7074__;
  assign new_new_n7337__ = new_new_n6990__ & ~new_new_n7074__;
  assign new_new_n7338__ = ~new_new_n7336__ & ~new_new_n7337__;
  assign new_new_n7339__ = new_new_n6857__ & new_new_n7338__;
  assign new_new_n7340__ = ~new_new_n6989__ & ~new_new_n7074__;
  assign new_new_n7341__ = ~new_new_n6990__ & ~new_new_n7340__;
  assign new_new_n7342__ = new_new_n6856__ & ~new_new_n7341__;
  assign new_new_n7343__ = new_new_n6855__ & new_new_n7341__;
  assign new_new_n7344__ = ~new_new_n7342__ & ~new_new_n7343__;
  assign new_new_n7345__ = ~new_new_n7339__ & new_new_n7344__;
  assign new_new_n7346__ = new_new_n7335__ & ~new_new_n7345__;
  assign new_new_n7347__ = ~new_new_n6856__ & ~new_new_n6988__;
  assign new_new_n7348__ = ~new_new_n6855__ & ~new_new_n7347__;
  assign new_new_n7349__ = ~new_new_n6859__ & ~new_new_n7348__;
  assign new_new_n7350__ = new_new_n6855__ & ~new_new_n6988__;
  assign new_new_n7351__ = ~new_new_n7349__ & ~new_new_n7350__;
  assign new_new_n7352__ = ~new_new_n7074__ & ~new_new_n7351__;
  assign new_new_n7353__ = new_new_n6859__ & new_new_n7348__;
  assign new_new_n7354__ = new_new_n6856__ & new_new_n6988__;
  assign new_new_n7355__ = ~new_new_n7353__ & ~new_new_n7354__;
  assign new_new_n7356__ = new_new_n7074__ & ~new_new_n7355__;
  assign new_new_n7357__ = new_new_n6845__ & ~new_new_n6859__;
  assign new_new_n7358__ = ~new_new_n6989__ & ~new_new_n7357__;
  assign new_new_n7359__ = ~new_new_n6854__ & ~new_new_n6988__;
  assign new_new_n7360__ = ~new_new_n6856__ & ~new_new_n7359__;
  assign new_new_n7361__ = ~new_new_n7358__ & ~new_new_n7360__;
  assign new_new_n7362__ = ~new_new_n7352__ & ~new_new_n7361__;
  assign new_new_n7363__ = ~new_new_n7356__ & new_new_n7362__;
  assign new_new_n7364__ = ~new_new_n7335__ & ~new_new_n7363__;
  assign po054 = new_new_n7346__ | new_new_n7364__;
  assign new_new_n7366__ = ~new_new_n7074__ & new_new_n7357__;
  assign new_new_n7367__ = new_new_n7335__ & ~new_new_n7366__;
  assign new_new_n7368__ = ~new_new_n6845__ & new_new_n6859__;
  assign new_new_n7369__ = new_new_n7074__ & new_new_n7368__;
  assign new_new_n7370__ = ~new_new_n7367__ & ~new_new_n7369__;
  assign new_new_n7371__ = ~new_new_n7359__ & ~new_new_n7370__;
  assign new_new_n7372__ = new_new_n7074__ & ~new_new_n7357__;
  assign new_new_n7373__ = ~new_new_n7368__ & ~new_new_n7372__;
  assign new_new_n7374__ = ~new_new_n7335__ & new_new_n7373__;
  assign new_new_n7375__ = new_new_n6988__ & ~new_new_n7374__;
  assign new_new_n7376__ = new_new_n6854__ & new_new_n7375__;
  assign new_new_n7377__ = new_new_n7335__ & ~new_new_n7373__;
  assign new_new_n7378__ = ~new_new_n7376__ & ~new_new_n7377__;
  assign new_new_n7379__ = ~new_new_n7371__ & new_new_n7378__;
  assign new_new_n7380__ = ~new_new_n7222__ & ~new_new_n7332__;
  assign new_new_n7381__ = ~new_new_n7221__ & ~new_new_n7380__;
  assign new_new_n7382__ = ~new_new_n7379__ & new_new_n7381__;
  assign new_new_n7383__ = new_new_n7379__ & ~new_new_n7381__;
  assign new_new_n7384__ = ~new_new_n7382__ & ~new_new_n7383__;
  assign new_new_n7385__ = ~new_new_n7260__ & ~new_new_n7278__;
  assign new_new_n7386__ = ~new_new_n7277__ & ~new_new_n7385__;
  assign new_new_n7387__ = ~new_new_n7230__ & new_new_n7244__;
  assign new_new_n7388__ = ~new_new_n7231__ & ~new_new_n7387__;
  assign new_new_n7389__ = new_new_n7386__ & ~new_new_n7388__;
  assign new_new_n7390__ = ~new_new_n7386__ & new_new_n7388__;
  assign new_new_n7391__ = ~new_new_n7389__ & ~new_new_n7390__;
  assign new_new_n7392__ = pi22 & pi32;
  assign new_new_n7393__ = pi19 & pi35;
  assign new_new_n7394__ = pi21 & pi33;
  assign new_new_n7395__ = ~new_new_n7393__ & ~new_new_n7394__;
  assign new_new_n7396__ = new_new_n7393__ & new_new_n7394__;
  assign new_new_n7397__ = ~new_new_n7395__ & ~new_new_n7396__;
  assign new_new_n7398__ = new_new_n7392__ & ~new_new_n7397__;
  assign new_new_n7399__ = ~new_new_n7392__ & new_new_n7397__;
  assign new_new_n7400__ = ~new_new_n7398__ & ~new_new_n7399__;
  assign new_new_n7401__ = pi00 & pi54;
  assign new_new_n7402__ = pi26 & pi28;
  assign new_new_n7403__ = pi01 & pi53;
  assign new_new_n7404__ = ~new_new_n7402__ & new_new_n7403__;
  assign new_new_n7405__ = new_new_n7402__ & ~new_new_n7403__;
  assign new_new_n7406__ = ~new_new_n7404__ & ~new_new_n7405__;
  assign new_new_n7407__ = new_new_n7263__ & ~new_new_n7406__;
  assign new_new_n7408__ = ~new_new_n7263__ & new_new_n7406__;
  assign new_new_n7409__ = ~new_new_n7407__ & ~new_new_n7408__;
  assign new_new_n7410__ = new_new_n7401__ & new_new_n7409__;
  assign new_new_n7411__ = ~new_new_n7401__ & ~new_new_n7409__;
  assign new_new_n7412__ = ~new_new_n7410__ & ~new_new_n7411__;
  assign new_new_n7413__ = new_new_n7400__ & ~new_new_n7412__;
  assign new_new_n7414__ = ~new_new_n7400__ & new_new_n7412__;
  assign new_new_n7415__ = ~new_new_n7413__ & ~new_new_n7414__;
  assign new_new_n7416__ = pi25 & pi29;
  assign new_new_n7417__ = pi23 & pi31;
  assign new_new_n7418__ = pi24 & pi30;
  assign new_new_n7419__ = ~new_new_n7417__ & ~new_new_n7418__;
  assign new_new_n7420__ = new_new_n7417__ & new_new_n7418__;
  assign new_new_n7421__ = ~new_new_n7419__ & ~new_new_n7420__;
  assign new_new_n7422__ = new_new_n7416__ & ~new_new_n7421__;
  assign new_new_n7423__ = ~new_new_n7416__ & new_new_n7421__;
  assign new_new_n7424__ = ~new_new_n7422__ & ~new_new_n7423__;
  assign new_new_n7425__ = ~new_new_n7415__ & new_new_n7424__;
  assign new_new_n7426__ = new_new_n7415__ & ~new_new_n7424__;
  assign new_new_n7427__ = ~new_new_n7425__ & ~new_new_n7426__;
  assign new_new_n7428__ = new_new_n7391__ & new_new_n7427__;
  assign new_new_n7429__ = ~new_new_n7391__ & ~new_new_n7427__;
  assign new_new_n7430__ = ~new_new_n7428__ & ~new_new_n7429__;
  assign new_new_n7431__ = ~new_new_n7284__ & ~new_new_n7287__;
  assign new_new_n7432__ = ~new_new_n7283__ & ~new_new_n7431__;
  assign new_new_n7433__ = new_new_n7430__ & ~new_new_n7432__;
  assign new_new_n7434__ = ~new_new_n7430__ & new_new_n7432__;
  assign new_new_n7435__ = ~new_new_n7433__ & ~new_new_n7434__;
  assign new_new_n7436__ = ~new_new_n7320__ & ~new_new_n7326__;
  assign new_new_n7437__ = ~new_new_n7321__ & ~new_new_n7436__;
  assign new_new_n7438__ = ~new_new_n7292__ & ~new_new_n7329__;
  assign new_new_n7439__ = ~new_new_n7291__ & ~new_new_n7438__;
  assign new_new_n7440__ = ~new_new_n7437__ & new_new_n7439__;
  assign new_new_n7441__ = new_new_n7437__ & ~new_new_n7439__;
  assign new_new_n7442__ = ~new_new_n7440__ & ~new_new_n7441__;
  assign new_new_n7443__ = ~new_new_n7118__ & ~new_new_n7153__;
  assign new_new_n7444__ = ~new_new_n7119__ & ~new_new_n7443__;
  assign new_new_n7445__ = ~new_new_n7234__ & ~new_new_n7240__;
  assign new_new_n7446__ = ~new_new_n7239__ & ~new_new_n7445__;
  assign new_new_n7447__ = ~new_new_n7253__ & ~new_new_n7258__;
  assign new_new_n7448__ = ~new_new_n7266__ & ~new_new_n7272__;
  assign new_new_n7449__ = ~new_new_n7271__ & ~new_new_n7448__;
  assign new_new_n7450__ = ~new_new_n7447__ & ~new_new_n7449__;
  assign new_new_n7451__ = new_new_n7447__ & new_new_n7449__;
  assign new_new_n7452__ = ~new_new_n7450__ & ~new_new_n7451__;
  assign new_new_n7453__ = new_new_n7446__ & ~new_new_n7452__;
  assign new_new_n7454__ = ~new_new_n7446__ & new_new_n7452__;
  assign new_new_n7455__ = ~new_new_n7453__ & ~new_new_n7454__;
  assign new_new_n7456__ = ~new_new_n7444__ & ~new_new_n7455__;
  assign new_new_n7457__ = new_new_n7444__ & new_new_n7455__;
  assign new_new_n7458__ = ~new_new_n7456__ & ~new_new_n7457__;
  assign new_new_n7459__ = ~new_new_n7103__ & ~new_new_n7114__;
  assign new_new_n7460__ = ~new_new_n7104__ & ~new_new_n7459__;
  assign new_new_n7461__ = ~new_new_n7085__ & ~new_new_n7089__;
  assign new_new_n7462__ = ~new_new_n7088__ & ~new_new_n7461__;
  assign new_new_n7463__ = ~new_new_n7203__ & ~new_new_n7207__;
  assign new_new_n7464__ = ~new_new_n7206__ & ~new_new_n7463__;
  assign new_new_n7465__ = ~new_new_n7106__ & ~new_new_n7110__;
  assign new_new_n7466__ = ~new_new_n7109__ & ~new_new_n7465__;
  assign new_new_n7467__ = ~new_new_n7464__ & ~new_new_n7466__;
  assign new_new_n7468__ = new_new_n7464__ & new_new_n7466__;
  assign new_new_n7469__ = ~new_new_n7467__ & ~new_new_n7468__;
  assign new_new_n7470__ = new_new_n7462__ & ~new_new_n7469__;
  assign new_new_n7471__ = ~new_new_n7462__ & new_new_n7469__;
  assign new_new_n7472__ = ~new_new_n7470__ & ~new_new_n7471__;
  assign new_new_n7473__ = new_new_n7460__ & new_new_n7472__;
  assign new_new_n7474__ = ~new_new_n7460__ & ~new_new_n7472__;
  assign new_new_n7475__ = ~new_new_n7473__ & ~new_new_n7474__;
  assign new_new_n7476__ = ~new_new_n7139__ & ~new_new_n7143__;
  assign new_new_n7477__ = ~new_new_n7142__ & ~new_new_n7476__;
  assign new_new_n7478__ = ~new_new_n7182__ & ~new_new_n7186__;
  assign new_new_n7479__ = ~new_new_n7185__ & ~new_new_n7478__;
  assign new_new_n7480__ = new_new_n7477__ & new_new_n7479__;
  assign new_new_n7481__ = ~new_new_n7477__ & ~new_new_n7479__;
  assign new_new_n7482__ = ~new_new_n7480__ & ~new_new_n7481__;
  assign new_new_n7483__ = ~new_new_n7121__ & ~new_new_n7125__;
  assign new_new_n7484__ = ~new_new_n7124__ & ~new_new_n7483__;
  assign new_new_n7485__ = ~new_new_n7482__ & new_new_n7484__;
  assign new_new_n7486__ = ~new_new_n7480__ & ~new_new_n7484__;
  assign new_new_n7487__ = ~new_new_n7481__ & new_new_n7486__;
  assign new_new_n7488__ = ~new_new_n7485__ & ~new_new_n7487__;
  assign new_new_n7489__ = ~new_new_n7475__ & new_new_n7488__;
  assign new_new_n7490__ = new_new_n7475__ & ~new_new_n7488__;
  assign new_new_n7491__ = ~new_new_n7489__ & ~new_new_n7490__;
  assign new_new_n7492__ = new_new_n7458__ & ~new_new_n7491__;
  assign new_new_n7493__ = ~new_new_n7458__ & new_new_n7491__;
  assign new_new_n7494__ = ~new_new_n7492__ & ~new_new_n7493__;
  assign new_new_n7495__ = ~new_new_n7165__ & new_new_n7217__;
  assign new_new_n7496__ = ~new_new_n7164__ & ~new_new_n7495__;
  assign new_new_n7497__ = new_new_n7494__ & new_new_n7496__;
  assign new_new_n7498__ = ~new_new_n7494__ & ~new_new_n7496__;
  assign new_new_n7499__ = ~new_new_n7497__ & ~new_new_n7498__;
  assign new_new_n7500__ = ~new_new_n7310__ & new_new_n7316__;
  assign new_new_n7501__ = ~new_new_n7311__ & ~new_new_n7500__;
  assign new_new_n7502__ = pi17 & pi37;
  assign new_new_n7503__ = pi16 & pi38;
  assign new_new_n7504__ = pi06 & pi48;
  assign new_new_n7505__ = ~new_new_n7503__ & ~new_new_n7504__;
  assign new_new_n7506__ = new_new_n7503__ & new_new_n7504__;
  assign new_new_n7507__ = ~new_new_n7505__ & ~new_new_n7506__;
  assign new_new_n7508__ = new_new_n7502__ & ~new_new_n7507__;
  assign new_new_n7509__ = ~new_new_n7502__ & new_new_n7507__;
  assign new_new_n7510__ = ~new_new_n7508__ & ~new_new_n7509__;
  assign new_new_n7511__ = pi20 & pi34;
  assign new_new_n7512__ = pi18 & pi36;
  assign new_new_n7513__ = pi05 & pi49;
  assign new_new_n7514__ = ~new_new_n7512__ & ~new_new_n7513__;
  assign new_new_n7515__ = new_new_n7512__ & new_new_n7513__;
  assign new_new_n7516__ = ~new_new_n7514__ & ~new_new_n7515__;
  assign new_new_n7517__ = new_new_n7511__ & ~new_new_n7516__;
  assign new_new_n7518__ = ~new_new_n7511__ & new_new_n7516__;
  assign new_new_n7519__ = ~new_new_n7517__ & ~new_new_n7518__;
  assign new_new_n7520__ = new_new_n7510__ & new_new_n7519__;
  assign new_new_n7521__ = ~new_new_n7510__ & ~new_new_n7519__;
  assign new_new_n7522__ = ~new_new_n7520__ & ~new_new_n7521__;
  assign new_new_n7523__ = pi13 & pi41;
  assign new_new_n7524__ = pi12 & pi42;
  assign new_new_n7525__ = pi11 & pi43;
  assign new_new_n7526__ = ~new_new_n7524__ & ~new_new_n7525__;
  assign new_new_n7527__ = new_new_n7524__ & new_new_n7525__;
  assign new_new_n7528__ = ~new_new_n7526__ & ~new_new_n7527__;
  assign new_new_n7529__ = new_new_n7523__ & ~new_new_n7528__;
  assign new_new_n7530__ = ~new_new_n7523__ & new_new_n7528__;
  assign new_new_n7531__ = ~new_new_n7529__ & ~new_new_n7530__;
  assign new_new_n7532__ = ~new_new_n7522__ & new_new_n7531__;
  assign new_new_n7533__ = new_new_n7522__ & ~new_new_n7531__;
  assign new_new_n7534__ = ~new_new_n7532__ & ~new_new_n7533__;
  assign new_new_n7535__ = ~new_new_n7501__ & new_new_n7534__;
  assign new_new_n7536__ = new_new_n7501__ & ~new_new_n7534__;
  assign new_new_n7537__ = ~new_new_n7535__ & ~new_new_n7536__;
  assign new_new_n7538__ = pi14 & pi40;
  assign new_new_n7539__ = pi09 & pi45;
  assign new_new_n7540__ = pi10 & pi44;
  assign new_new_n7541__ = ~new_new_n7539__ & ~new_new_n7540__;
  assign new_new_n7542__ = new_new_n7539__ & new_new_n7540__;
  assign new_new_n7543__ = ~new_new_n7541__ & ~new_new_n7542__;
  assign new_new_n7544__ = new_new_n7538__ & ~new_new_n7543__;
  assign new_new_n7545__ = ~new_new_n7538__ & new_new_n7543__;
  assign new_new_n7546__ = ~new_new_n7544__ & ~new_new_n7545__;
  assign new_new_n7547__ = pi04 & pi50;
  assign new_new_n7548__ = pi03 & pi51;
  assign new_new_n7549__ = pi02 & pi52;
  assign new_new_n7550__ = ~new_new_n7548__ & ~new_new_n7549__;
  assign new_new_n7551__ = new_new_n7548__ & new_new_n7549__;
  assign new_new_n7552__ = ~new_new_n7550__ & ~new_new_n7551__;
  assign new_new_n7553__ = new_new_n7547__ & ~new_new_n7552__;
  assign new_new_n7554__ = ~new_new_n7547__ & new_new_n7552__;
  assign new_new_n7555__ = ~new_new_n7553__ & ~new_new_n7554__;
  assign new_new_n7556__ = new_new_n7546__ & new_new_n7555__;
  assign new_new_n7557__ = ~new_new_n7546__ & ~new_new_n7555__;
  assign new_new_n7558__ = ~new_new_n7556__ & ~new_new_n7557__;
  assign new_new_n7559__ = pi15 & pi39;
  assign new_new_n7560__ = pi07 & pi47;
  assign new_new_n7561__ = pi08 & pi46;
  assign new_new_n7562__ = ~new_new_n7560__ & ~new_new_n7561__;
  assign new_new_n7563__ = new_new_n7560__ & new_new_n7561__;
  assign new_new_n7564__ = ~new_new_n7562__ & ~new_new_n7563__;
  assign new_new_n7565__ = new_new_n7559__ & ~new_new_n7564__;
  assign new_new_n7566__ = ~new_new_n7559__ & new_new_n7564__;
  assign new_new_n7567__ = ~new_new_n7565__ & ~new_new_n7566__;
  assign new_new_n7568__ = new_new_n7558__ & ~new_new_n7567__;
  assign new_new_n7569__ = ~new_new_n7558__ & new_new_n7567__;
  assign new_new_n7570__ = ~new_new_n7568__ & ~new_new_n7569__;
  assign new_new_n7571__ = new_new_n7537__ & ~new_new_n7570__;
  assign new_new_n7572__ = ~new_new_n7537__ & new_new_n7570__;
  assign new_new_n7573__ = ~new_new_n7571__ & ~new_new_n7572__;
  assign new_new_n7574__ = new_new_n7180__ & ~new_new_n7573__;
  assign new_new_n7575__ = new_new_n7179__ & new_new_n7573__;
  assign new_new_n7576__ = ~new_new_n7180__ & new_new_n7573__;
  assign new_new_n7577__ = new_new_n7211__ & ~new_new_n7576__;
  assign new_new_n7578__ = ~new_new_n7179__ & ~new_new_n7573__;
  assign new_new_n7579__ = ~new_new_n7211__ & ~new_new_n7578__;
  assign new_new_n7580__ = ~new_new_n7202__ & ~new_new_n7577__;
  assign new_new_n7581__ = ~new_new_n7579__ & new_new_n7580__;
  assign new_new_n7582__ = new_new_n7211__ & ~new_new_n7578__;
  assign new_new_n7583__ = ~new_new_n7211__ & ~new_new_n7576__;
  assign new_new_n7584__ = new_new_n7202__ & ~new_new_n7582__;
  assign new_new_n7585__ = ~new_new_n7583__ & new_new_n7584__;
  assign new_new_n7586__ = ~new_new_n7575__ & ~new_new_n7581__;
  assign new_new_n7587__ = ~new_new_n7585__ & new_new_n7586__;
  assign new_new_n7588__ = ~new_new_n7574__ & new_new_n7587__;
  assign new_new_n7589__ = ~new_new_n7200__ & ~new_new_n7211__;
  assign new_new_n7590__ = ~new_new_n7201__ & ~new_new_n7589__;
  assign new_new_n7591__ = ~new_new_n7129__ & ~new_new_n7148__;
  assign new_new_n7592__ = ~new_new_n7149__ & ~new_new_n7591__;
  assign new_new_n7593__ = ~new_new_n7590__ & ~new_new_n7592__;
  assign new_new_n7594__ = new_new_n7590__ & new_new_n7592__;
  assign new_new_n7595__ = ~new_new_n7593__ & ~new_new_n7594__;
  assign new_new_n7596__ = ~new_new_n7191__ & ~new_new_n7195__;
  assign new_new_n7597__ = ~new_new_n7194__ & ~new_new_n7596__;
  assign new_new_n7598__ = ~new_new_n7130__ & ~new_new_n7134__;
  assign new_new_n7599__ = new_new_n7133__ & ~new_new_n7598__;
  assign new_new_n7600__ = ~new_new_n7094__ & ~new_new_n7098__;
  assign new_new_n7601__ = ~new_new_n7097__ & ~new_new_n7600__;
  assign new_new_n7602__ = ~new_new_n7599__ & ~new_new_n7601__;
  assign new_new_n7603__ = new_new_n7599__ & new_new_n7601__;
  assign new_new_n7604__ = ~new_new_n7602__ & ~new_new_n7603__;
  assign new_new_n7605__ = new_new_n7597__ & ~new_new_n7604__;
  assign new_new_n7606__ = ~new_new_n7597__ & new_new_n7604__;
  assign new_new_n7607__ = ~new_new_n7605__ & ~new_new_n7606__;
  assign new_new_n7608__ = new_new_n7595__ & new_new_n7607__;
  assign new_new_n7609__ = ~new_new_n7595__ & ~new_new_n7607__;
  assign new_new_n7610__ = ~new_new_n7608__ & ~new_new_n7609__;
  assign new_new_n7611__ = new_new_n7588__ & ~new_new_n7610__;
  assign new_new_n7612__ = ~new_new_n7588__ & new_new_n7610__;
  assign new_new_n7613__ = ~new_new_n7611__ & ~new_new_n7612__;
  assign new_new_n7614__ = new_new_n7499__ & new_new_n7613__;
  assign new_new_n7615__ = ~new_new_n7499__ & ~new_new_n7613__;
  assign new_new_n7616__ = ~new_new_n7614__ & ~new_new_n7615__;
  assign new_new_n7617__ = new_new_n7442__ & ~new_new_n7616__;
  assign new_new_n7618__ = ~new_new_n7442__ & new_new_n7616__;
  assign new_new_n7619__ = ~new_new_n7617__ & ~new_new_n7618__;
  assign new_new_n7620__ = new_new_n7435__ & new_new_n7619__;
  assign new_new_n7621__ = ~new_new_n7435__ & ~new_new_n7619__;
  assign new_new_n7622__ = ~new_new_n7620__ & ~new_new_n7621__;
  assign new_new_n7623__ = new_new_n7384__ & new_new_n7622__;
  assign new_new_n7624__ = ~new_new_n7384__ & ~new_new_n7622__;
  assign po055 = ~new_new_n7623__ & ~new_new_n7624__;
  assign new_new_n7626__ = ~new_new_n7383__ & ~new_new_n7622__;
  assign new_new_n7627__ = ~new_new_n7382__ & ~new_new_n7626__;
  assign new_new_n7628__ = new_new_n7435__ & ~new_new_n7437__;
  assign new_new_n7629__ = ~new_new_n7435__ & new_new_n7437__;
  assign new_new_n7630__ = ~new_new_n7628__ & ~new_new_n7629__;
  assign new_new_n7631__ = ~new_new_n7616__ & new_new_n7630__;
  assign new_new_n7632__ = new_new_n7616__ & ~new_new_n7630__;
  assign new_new_n7633__ = ~new_new_n7439__ & ~new_new_n7632__;
  assign new_new_n7634__ = ~new_new_n7631__ & ~new_new_n7633__;
  assign new_new_n7635__ = new_new_n7627__ & new_new_n7634__;
  assign new_new_n7636__ = ~new_new_n7627__ & ~new_new_n7634__;
  assign new_new_n7637__ = ~new_new_n7635__ & ~new_new_n7636__;
  assign new_new_n7638__ = ~new_new_n7430__ & new_new_n7437__;
  assign new_new_n7639__ = new_new_n7432__ & ~new_new_n7638__;
  assign new_new_n7640__ = new_new_n7430__ & ~new_new_n7437__;
  assign new_new_n7641__ = ~new_new_n7639__ & ~new_new_n7640__;
  assign new_new_n7642__ = ~new_new_n7390__ & ~new_new_n7427__;
  assign new_new_n7643__ = ~new_new_n7389__ & ~new_new_n7642__;
  assign new_new_n7644__ = ~new_new_n7446__ & ~new_new_n7451__;
  assign new_new_n7645__ = ~new_new_n7450__ & ~new_new_n7644__;
  assign new_new_n7646__ = pi13 & pi42;
  assign new_new_n7647__ = pi10 & pi45;
  assign new_new_n7648__ = pi11 & pi44;
  assign new_new_n7649__ = ~new_new_n7647__ & ~new_new_n7648__;
  assign new_new_n7650__ = new_new_n7647__ & new_new_n7648__;
  assign new_new_n7651__ = ~new_new_n7649__ & ~new_new_n7650__;
  assign new_new_n7652__ = new_new_n7646__ & ~new_new_n7651__;
  assign new_new_n7653__ = ~new_new_n7646__ & new_new_n7651__;
  assign new_new_n7654__ = ~new_new_n7652__ & ~new_new_n7653__;
  assign new_new_n7655__ = pi27 & pi28;
  assign new_new_n7656__ = pi12 & pi43;
  assign new_new_n7657__ = pi26 & pi29;
  assign new_new_n7658__ = ~new_new_n7656__ & ~new_new_n7657__;
  assign new_new_n7659__ = new_new_n7656__ & new_new_n7657__;
  assign new_new_n7660__ = ~new_new_n7658__ & ~new_new_n7659__;
  assign new_new_n7661__ = new_new_n7655__ & ~new_new_n7660__;
  assign new_new_n7662__ = ~new_new_n7655__ & new_new_n7660__;
  assign new_new_n7663__ = ~new_new_n7661__ & ~new_new_n7662__;
  assign new_new_n7664__ = new_new_n7654__ & new_new_n7663__;
  assign new_new_n7665__ = ~new_new_n7654__ & ~new_new_n7663__;
  assign new_new_n7666__ = ~new_new_n7664__ & ~new_new_n7665__;
  assign new_new_n7667__ = pi16 & pi39;
  assign new_new_n7668__ = pi08 & pi47;
  assign new_new_n7669__ = pi07 & pi48;
  assign new_new_n7670__ = ~new_new_n7668__ & ~new_new_n7669__;
  assign new_new_n7671__ = new_new_n7668__ & new_new_n7669__;
  assign new_new_n7672__ = ~new_new_n7670__ & ~new_new_n7671__;
  assign new_new_n7673__ = new_new_n7667__ & ~new_new_n7672__;
  assign new_new_n7674__ = ~new_new_n7667__ & new_new_n7672__;
  assign new_new_n7675__ = ~new_new_n7673__ & ~new_new_n7674__;
  assign new_new_n7676__ = ~new_new_n7666__ & new_new_n7675__;
  assign new_new_n7677__ = new_new_n7666__ & ~new_new_n7675__;
  assign new_new_n7678__ = ~new_new_n7676__ & ~new_new_n7677__;
  assign new_new_n7679__ = ~new_new_n7645__ & ~new_new_n7678__;
  assign new_new_n7680__ = new_new_n7645__ & new_new_n7678__;
  assign new_new_n7681__ = ~new_new_n7679__ & ~new_new_n7680__;
  assign new_new_n7682__ = pi25 & pi30;
  assign new_new_n7683__ = pi24 & pi31;
  assign new_new_n7684__ = pi23 & pi32;
  assign new_new_n7685__ = ~new_new_n7683__ & ~new_new_n7684__;
  assign new_new_n7686__ = new_new_n7683__ & new_new_n7684__;
  assign new_new_n7687__ = ~new_new_n7685__ & ~new_new_n7686__;
  assign new_new_n7688__ = new_new_n7682__ & ~new_new_n7687__;
  assign new_new_n7689__ = ~new_new_n7682__ & new_new_n7687__;
  assign new_new_n7690__ = ~new_new_n7688__ & ~new_new_n7689__;
  assign new_new_n7691__ = pi04 & pi51;
  assign new_new_n7692__ = pi02 & pi53;
  assign new_new_n7693__ = pi00 & pi55;
  assign new_new_n7694__ = ~new_new_n7692__ & ~new_new_n7693__;
  assign new_new_n7695__ = new_new_n7692__ & new_new_n7693__;
  assign new_new_n7696__ = ~new_new_n7694__ & ~new_new_n7695__;
  assign new_new_n7697__ = new_new_n7691__ & ~new_new_n7696__;
  assign new_new_n7698__ = ~new_new_n7691__ & new_new_n7696__;
  assign new_new_n7699__ = ~new_new_n7697__ & ~new_new_n7698__;
  assign new_new_n7700__ = new_new_n7690__ & new_new_n7699__;
  assign new_new_n7701__ = ~new_new_n7690__ & ~new_new_n7699__;
  assign new_new_n7702__ = ~new_new_n7700__ & ~new_new_n7701__;
  assign new_new_n7703__ = pi22 & pi33;
  assign new_new_n7704__ = pi21 & pi34;
  assign new_new_n7705__ = pi20 & pi35;
  assign new_new_n7706__ = ~new_new_n7704__ & ~new_new_n7705__;
  assign new_new_n7707__ = new_new_n7704__ & new_new_n7705__;
  assign new_new_n7708__ = ~new_new_n7706__ & ~new_new_n7707__;
  assign new_new_n7709__ = new_new_n7703__ & ~new_new_n7708__;
  assign new_new_n7710__ = ~new_new_n7703__ & new_new_n7708__;
  assign new_new_n7711__ = ~new_new_n7709__ & ~new_new_n7710__;
  assign new_new_n7712__ = new_new_n7702__ & ~new_new_n7711__;
  assign new_new_n7713__ = ~new_new_n7702__ & new_new_n7711__;
  assign new_new_n7714__ = ~new_new_n7712__ & ~new_new_n7713__;
  assign new_new_n7715__ = new_new_n7681__ & ~new_new_n7714__;
  assign new_new_n7716__ = ~new_new_n7681__ & new_new_n7714__;
  assign new_new_n7717__ = ~new_new_n7715__ & ~new_new_n7716__;
  assign new_new_n7718__ = ~new_new_n7643__ & new_new_n7717__;
  assign new_new_n7719__ = new_new_n7643__ & ~new_new_n7717__;
  assign new_new_n7720__ = ~new_new_n7718__ & ~new_new_n7719__;
  assign new_new_n7721__ = ~new_new_n7556__ & ~new_new_n7567__;
  assign new_new_n7722__ = ~new_new_n7557__ & ~new_new_n7721__;
  assign new_new_n7723__ = ~new_new_n7520__ & ~new_new_n7531__;
  assign new_new_n7724__ = ~new_new_n7521__ & ~new_new_n7723__;
  assign new_new_n7725__ = ~new_new_n7416__ & ~new_new_n7420__;
  assign new_new_n7726__ = ~new_new_n7419__ & ~new_new_n7725__;
  assign new_new_n7727__ = ~new_new_n7502__ & ~new_new_n7506__;
  assign new_new_n7728__ = ~new_new_n7505__ & ~new_new_n7727__;
  assign new_new_n7729__ = ~new_new_n7392__ & ~new_new_n7396__;
  assign new_new_n7730__ = ~new_new_n7395__ & ~new_new_n7729__;
  assign new_new_n7731__ = ~new_new_n7728__ & ~new_new_n7730__;
  assign new_new_n7732__ = new_new_n7728__ & new_new_n7730__;
  assign new_new_n7733__ = ~new_new_n7731__ & ~new_new_n7732__;
  assign new_new_n7734__ = new_new_n7726__ & ~new_new_n7733__;
  assign new_new_n7735__ = ~new_new_n7726__ & new_new_n7733__;
  assign new_new_n7736__ = ~new_new_n7734__ & ~new_new_n7735__;
  assign new_new_n7737__ = ~new_new_n7724__ & ~new_new_n7736__;
  assign new_new_n7738__ = new_new_n7724__ & new_new_n7736__;
  assign new_new_n7739__ = ~new_new_n7737__ & ~new_new_n7738__;
  assign new_new_n7740__ = new_new_n7722__ & new_new_n7739__;
  assign new_new_n7741__ = ~new_new_n7722__ & ~new_new_n7739__;
  assign new_new_n7742__ = ~new_new_n7740__ & ~new_new_n7741__;
  assign new_new_n7743__ = new_new_n7720__ & ~new_new_n7742__;
  assign new_new_n7744__ = ~new_new_n7720__ & new_new_n7742__;
  assign new_new_n7745__ = ~new_new_n7743__ & ~new_new_n7744__;
  assign new_new_n7746__ = ~new_new_n7641__ & new_new_n7745__;
  assign new_new_n7747__ = new_new_n7641__ & ~new_new_n7745__;
  assign new_new_n7748__ = ~new_new_n7746__ & ~new_new_n7747__;
  assign new_new_n7749__ = ~new_new_n7536__ & new_new_n7570__;
  assign new_new_n7750__ = ~new_new_n7535__ & ~new_new_n7749__;
  assign new_new_n7751__ = ~new_new_n7597__ & ~new_new_n7603__;
  assign new_new_n7752__ = ~new_new_n7602__ & ~new_new_n7751__;
  assign new_new_n7753__ = ~new_new_n7462__ & ~new_new_n7468__;
  assign new_new_n7754__ = ~new_new_n7467__ & ~new_new_n7753__;
  assign new_new_n7755__ = pi26 & pi53;
  assign new_new_n7756__ = ~new_new_n7523__ & ~new_new_n7527__;
  assign new_new_n7757__ = ~new_new_n7526__ & ~new_new_n7756__;
  assign new_new_n7758__ = pi01 & ~pi54;
  assign new_new_n7759__ = ~new_new_n7757__ & ~new_new_n7758__;
  assign new_new_n7760__ = new_new_n7755__ & ~new_new_n7759__;
  assign new_new_n7761__ = pi28 & pi54;
  assign new_new_n7762__ = new_new_n7757__ & ~new_new_n7761__;
  assign new_new_n7763__ = new_new_n7760__ & ~new_new_n7762__;
  assign new_new_n7764__ = new_new_n7402__ & new_new_n7403__;
  assign new_new_n7765__ = pi01 & pi54;
  assign new_new_n7766__ = new_new_n7757__ & ~new_new_n7765__;
  assign new_new_n7767__ = ~new_new_n7757__ & new_new_n7765__;
  assign new_new_n7768__ = ~new_new_n7766__ & ~new_new_n7767__;
  assign new_new_n7769__ = pi28 & new_new_n7768__;
  assign new_new_n7770__ = ~pi28 & ~new_new_n7768__;
  assign new_new_n7771__ = ~new_new_n7764__ & ~new_new_n7769__;
  assign new_new_n7772__ = ~new_new_n7770__ & new_new_n7771__;
  assign new_new_n7773__ = ~new_new_n7763__ & ~new_new_n7772__;
  assign new_new_n7774__ = new_new_n7754__ & new_new_n7773__;
  assign new_new_n7775__ = ~new_new_n7754__ & ~new_new_n7773__;
  assign new_new_n7776__ = ~new_new_n7774__ & ~new_new_n7775__;
  assign new_new_n7777__ = new_new_n7752__ & ~new_new_n7776__;
  assign new_new_n7778__ = ~new_new_n7752__ & new_new_n7776__;
  assign new_new_n7779__ = ~new_new_n7777__ & ~new_new_n7778__;
  assign new_new_n7780__ = ~new_new_n7750__ & ~new_new_n7779__;
  assign new_new_n7781__ = new_new_n7750__ & new_new_n7779__;
  assign new_new_n7782__ = ~new_new_n7780__ & ~new_new_n7781__;
  assign new_new_n7783__ = ~new_new_n7511__ & ~new_new_n7515__;
  assign new_new_n7784__ = ~new_new_n7514__ & ~new_new_n7783__;
  assign new_new_n7785__ = ~new_new_n7538__ & ~new_new_n7542__;
  assign new_new_n7786__ = ~new_new_n7541__ & ~new_new_n7785__;
  assign new_new_n7787__ = ~new_new_n7784__ & ~new_new_n7786__;
  assign new_new_n7788__ = new_new_n7784__ & new_new_n7786__;
  assign new_new_n7789__ = ~new_new_n7787__ & ~new_new_n7788__;
  assign new_new_n7790__ = ~new_new_n7547__ & ~new_new_n7551__;
  assign new_new_n7791__ = ~new_new_n7550__ & ~new_new_n7790__;
  assign new_new_n7792__ = ~new_new_n7789__ & new_new_n7791__;
  assign new_new_n7793__ = ~new_new_n7788__ & ~new_new_n7791__;
  assign new_new_n7794__ = ~new_new_n7787__ & new_new_n7793__;
  assign new_new_n7795__ = ~new_new_n7792__ & ~new_new_n7794__;
  assign new_new_n7796__ = ~new_new_n7414__ & new_new_n7424__;
  assign new_new_n7797__ = ~new_new_n7413__ & ~new_new_n7796__;
  assign new_new_n7798__ = new_new_n7795__ & ~new_new_n7797__;
  assign new_new_n7799__ = ~new_new_n7795__ & new_new_n7797__;
  assign new_new_n7800__ = ~new_new_n7798__ & ~new_new_n7799__;
  assign new_new_n7801__ = ~new_new_n7559__ & ~new_new_n7563__;
  assign new_new_n7802__ = ~new_new_n7562__ & ~new_new_n7801__;
  assign new_new_n7803__ = ~new_new_n7401__ & ~new_new_n7407__;
  assign new_new_n7804__ = ~new_new_n7408__ & ~new_new_n7803__;
  assign new_new_n7805__ = new_new_n7802__ & new_new_n7804__;
  assign new_new_n7806__ = ~new_new_n7802__ & ~new_new_n7804__;
  assign new_new_n7807__ = ~new_new_n7805__ & ~new_new_n7806__;
  assign new_new_n7808__ = pi05 & pi50;
  assign new_new_n7809__ = ~new_new_n4095__ & ~new_new_n7808__;
  assign new_new_n7810__ = new_new_n4095__ & new_new_n7808__;
  assign new_new_n7811__ = ~new_new_n7809__ & ~new_new_n7810__;
  assign new_new_n7812__ = new_new_n3728__ & ~new_new_n7811__;
  assign new_new_n7813__ = ~new_new_n3728__ & new_new_n7811__;
  assign new_new_n7814__ = ~new_new_n7812__ & ~new_new_n7813__;
  assign new_new_n7815__ = new_new_n7807__ & ~new_new_n7814__;
  assign new_new_n7816__ = ~new_new_n7807__ & new_new_n7814__;
  assign new_new_n7817__ = ~new_new_n7815__ & ~new_new_n7816__;
  assign new_new_n7818__ = new_new_n7800__ & new_new_n7817__;
  assign new_new_n7819__ = ~new_new_n7800__ & ~new_new_n7817__;
  assign new_new_n7820__ = ~new_new_n7818__ & ~new_new_n7819__;
  assign new_new_n7821__ = new_new_n7782__ & new_new_n7820__;
  assign new_new_n7822__ = ~new_new_n7782__ & ~new_new_n7820__;
  assign new_new_n7823__ = ~new_new_n7821__ & ~new_new_n7822__;
  assign new_new_n7824__ = new_new_n7748__ & ~new_new_n7823__;
  assign new_new_n7825__ = ~new_new_n7748__ & new_new_n7823__;
  assign new_new_n7826__ = ~new_new_n7824__ & ~new_new_n7825__;
  assign new_new_n7827__ = ~new_new_n7498__ & ~new_new_n7613__;
  assign new_new_n7828__ = ~new_new_n7497__ & ~new_new_n7827__;
  assign new_new_n7829__ = new_new_n7588__ & new_new_n7610__;
  assign new_new_n7830__ = new_new_n7573__ & ~new_new_n7587__;
  assign new_new_n7831__ = ~new_new_n7829__ & ~new_new_n7830__;
  assign new_new_n7832__ = ~new_new_n7457__ & new_new_n7491__;
  assign new_new_n7833__ = ~new_new_n7456__ & ~new_new_n7832__;
  assign new_new_n7834__ = new_new_n7831__ & ~new_new_n7833__;
  assign new_new_n7835__ = ~new_new_n7831__ & new_new_n7833__;
  assign new_new_n7836__ = ~new_new_n7834__ & ~new_new_n7835__;
  assign new_new_n7837__ = ~new_new_n7594__ & ~new_new_n7607__;
  assign new_new_n7838__ = ~new_new_n7593__ & ~new_new_n7837__;
  assign new_new_n7839__ = pi15 & pi40;
  assign new_new_n7840__ = pi14 & pi41;
  assign new_new_n7841__ = pi09 & pi46;
  assign new_new_n7842__ = ~new_new_n7840__ & ~new_new_n7841__;
  assign new_new_n7843__ = new_new_n7840__ & new_new_n7841__;
  assign new_new_n7844__ = ~new_new_n7842__ & ~new_new_n7843__;
  assign new_new_n7845__ = new_new_n7839__ & ~new_new_n7844__;
  assign new_new_n7846__ = ~new_new_n7839__ & new_new_n7844__;
  assign new_new_n7847__ = ~new_new_n7845__ & ~new_new_n7846__;
  assign new_new_n7848__ = pi17 & pi38;
  assign new_new_n7849__ = pi06 & pi49;
  assign new_new_n7850__ = pi03 & pi52;
  assign new_new_n7851__ = ~new_new_n7849__ & ~new_new_n7850__;
  assign new_new_n7852__ = new_new_n7849__ & new_new_n7850__;
  assign new_new_n7853__ = ~new_new_n7851__ & ~new_new_n7852__;
  assign new_new_n7854__ = new_new_n7848__ & ~new_new_n7853__;
  assign new_new_n7855__ = ~new_new_n7848__ & new_new_n7853__;
  assign new_new_n7856__ = ~new_new_n7854__ & ~new_new_n7855__;
  assign new_new_n7857__ = new_new_n7847__ & new_new_n7856__;
  assign new_new_n7858__ = ~new_new_n7847__ & ~new_new_n7856__;
  assign new_new_n7859__ = ~new_new_n7857__ & ~new_new_n7858__;
  assign new_new_n7860__ = ~new_new_n7481__ & ~new_new_n7486__;
  assign new_new_n7861__ = new_new_n7859__ & ~new_new_n7860__;
  assign new_new_n7862__ = ~new_new_n7859__ & new_new_n7860__;
  assign new_new_n7863__ = ~new_new_n7861__ & ~new_new_n7862__;
  assign new_new_n7864__ = new_new_n7838__ & new_new_n7863__;
  assign new_new_n7865__ = ~new_new_n7838__ & ~new_new_n7863__;
  assign new_new_n7866__ = ~new_new_n7864__ & ~new_new_n7865__;
  assign new_new_n7867__ = ~new_new_n7473__ & ~new_new_n7488__;
  assign new_new_n7868__ = ~new_new_n7474__ & ~new_new_n7867__;
  assign new_new_n7869__ = new_new_n7866__ & ~new_new_n7868__;
  assign new_new_n7870__ = ~new_new_n7866__ & new_new_n7868__;
  assign new_new_n7871__ = ~new_new_n7869__ & ~new_new_n7870__;
  assign new_new_n7872__ = new_new_n7836__ & ~new_new_n7871__;
  assign new_new_n7873__ = ~new_new_n7836__ & new_new_n7871__;
  assign new_new_n7874__ = ~new_new_n7872__ & ~new_new_n7873__;
  assign new_new_n7875__ = new_new_n7828__ & ~new_new_n7874__;
  assign new_new_n7876__ = ~new_new_n7828__ & new_new_n7874__;
  assign new_new_n7877__ = ~new_new_n7875__ & ~new_new_n7876__;
  assign new_new_n7878__ = new_new_n7826__ & new_new_n7877__;
  assign new_new_n7879__ = ~new_new_n7826__ & ~new_new_n7877__;
  assign new_new_n7880__ = ~new_new_n7878__ & ~new_new_n7879__;
  assign new_new_n7881__ = new_new_n7637__ & new_new_n7880__;
  assign new_new_n7882__ = ~new_new_n7637__ & ~new_new_n7880__;
  assign po056 = new_new_n7881__ | new_new_n7882__;
  assign new_new_n7884__ = ~new_new_n7635__ & new_new_n7880__;
  assign new_new_n7885__ = ~new_new_n7636__ & ~new_new_n7884__;
  assign new_new_n7886__ = new_new_n7826__ & ~new_new_n7875__;
  assign new_new_n7887__ = ~new_new_n7876__ & ~new_new_n7886__;
  assign new_new_n7888__ = ~new_new_n7885__ & ~new_new_n7887__;
  assign new_new_n7889__ = new_new_n7885__ & new_new_n7887__;
  assign new_new_n7890__ = ~new_new_n7888__ & ~new_new_n7889__;
  assign new_new_n7891__ = ~new_new_n7746__ & ~new_new_n7823__;
  assign new_new_n7892__ = ~new_new_n7747__ & ~new_new_n7891__;
  assign new_new_n7893__ = pi16 & pi40;
  assign new_new_n7894__ = pi15 & pi41;
  assign new_new_n7895__ = pi08 & pi48;
  assign new_new_n7896__ = ~new_new_n7894__ & ~new_new_n7895__;
  assign new_new_n7897__ = new_new_n7894__ & new_new_n7895__;
  assign new_new_n7898__ = ~new_new_n7896__ & ~new_new_n7897__;
  assign new_new_n7899__ = new_new_n7893__ & ~new_new_n7898__;
  assign new_new_n7900__ = ~new_new_n7893__ & new_new_n7898__;
  assign new_new_n7901__ = ~new_new_n7899__ & ~new_new_n7900__;
  assign new_new_n7902__ = pi17 & pi39;
  assign new_new_n7903__ = pi07 & pi49;
  assign new_new_n7904__ = pi06 & pi50;
  assign new_new_n7905__ = ~new_new_n7903__ & ~new_new_n7904__;
  assign new_new_n7906__ = new_new_n7903__ & new_new_n7904__;
  assign new_new_n7907__ = ~new_new_n7905__ & ~new_new_n7906__;
  assign new_new_n7908__ = new_new_n7902__ & ~new_new_n7907__;
  assign new_new_n7909__ = ~new_new_n7902__ & new_new_n7907__;
  assign new_new_n7910__ = ~new_new_n7908__ & ~new_new_n7909__;
  assign new_new_n7911__ = new_new_n7901__ & new_new_n7910__;
  assign new_new_n7912__ = ~new_new_n7901__ & ~new_new_n7910__;
  assign new_new_n7913__ = ~new_new_n7911__ & ~new_new_n7912__;
  assign new_new_n7914__ = pi13 & pi43;
  assign new_new_n7915__ = pi11 & pi45;
  assign new_new_n7916__ = pi12 & pi44;
  assign new_new_n7917__ = ~new_new_n7915__ & ~new_new_n7916__;
  assign new_new_n7918__ = new_new_n7915__ & new_new_n7916__;
  assign new_new_n7919__ = ~new_new_n7917__ & ~new_new_n7918__;
  assign new_new_n7920__ = new_new_n7914__ & ~new_new_n7919__;
  assign new_new_n7921__ = ~new_new_n7914__ & new_new_n7919__;
  assign new_new_n7922__ = ~new_new_n7920__ & ~new_new_n7921__;
  assign new_new_n7923__ = new_new_n7913__ & ~new_new_n7922__;
  assign new_new_n7924__ = ~new_new_n7913__ & new_new_n7922__;
  assign new_new_n7925__ = ~new_new_n7923__ & ~new_new_n7924__;
  assign new_new_n7926__ = pi26 & pi30;
  assign new_new_n7927__ = pi24 & pi32;
  assign new_new_n7928__ = pi25 & pi31;
  assign new_new_n7929__ = ~new_new_n7927__ & ~new_new_n7928__;
  assign new_new_n7930__ = new_new_n7927__ & new_new_n7928__;
  assign new_new_n7931__ = ~new_new_n7929__ & ~new_new_n7930__;
  assign new_new_n7932__ = new_new_n7926__ & ~new_new_n7931__;
  assign new_new_n7933__ = ~new_new_n7926__ & new_new_n7931__;
  assign new_new_n7934__ = ~new_new_n7932__ & ~new_new_n7933__;
  assign new_new_n7935__ = pi23 & pi33;
  assign new_new_n7936__ = pi22 & pi34;
  assign new_new_n7937__ = pi20 & pi36;
  assign new_new_n7938__ = ~new_new_n7936__ & ~new_new_n7937__;
  assign new_new_n7939__ = new_new_n7936__ & new_new_n7937__;
  assign new_new_n7940__ = ~new_new_n7938__ & ~new_new_n7939__;
  assign new_new_n7941__ = new_new_n7935__ & ~new_new_n7940__;
  assign new_new_n7942__ = ~new_new_n7935__ & new_new_n7940__;
  assign new_new_n7943__ = ~new_new_n7941__ & ~new_new_n7942__;
  assign new_new_n7944__ = new_new_n7934__ & new_new_n7943__;
  assign new_new_n7945__ = ~new_new_n7934__ & ~new_new_n7943__;
  assign new_new_n7946__ = ~new_new_n7944__ & ~new_new_n7945__;
  assign new_new_n7947__ = pi14 & pi42;
  assign new_new_n7948__ = pi10 & pi46;
  assign new_new_n7949__ = pi09 & pi47;
  assign new_new_n7950__ = ~new_new_n7948__ & ~new_new_n7949__;
  assign new_new_n7951__ = new_new_n7948__ & new_new_n7949__;
  assign new_new_n7952__ = ~new_new_n7950__ & ~new_new_n7951__;
  assign new_new_n7953__ = new_new_n7947__ & ~new_new_n7952__;
  assign new_new_n7954__ = ~new_new_n7947__ & new_new_n7952__;
  assign new_new_n7955__ = ~new_new_n7953__ & ~new_new_n7954__;
  assign new_new_n7956__ = ~new_new_n7946__ & new_new_n7955__;
  assign new_new_n7957__ = new_new_n7946__ & ~new_new_n7955__;
  assign new_new_n7958__ = ~new_new_n7956__ & ~new_new_n7957__;
  assign new_new_n7959__ = ~new_new_n7925__ & ~new_new_n7958__;
  assign new_new_n7960__ = new_new_n7925__ & new_new_n7958__;
  assign new_new_n7961__ = ~new_new_n7959__ & ~new_new_n7960__;
  assign new_new_n7962__ = ~new_new_n7667__ & ~new_new_n7671__;
  assign new_new_n7963__ = ~new_new_n7670__ & ~new_new_n7962__;
  assign new_new_n7964__ = pi00 & pi56;
  assign new_new_n7965__ = pi02 & new_new_n2370__;
  assign new_new_n7966__ = ~pi02 & ~new_new_n2370__;
  assign new_new_n7967__ = pi54 & ~new_new_n7966__;
  assign new_new_n7968__ = ~new_new_n7965__ & new_new_n7967__;
  assign new_new_n7969__ = new_new_n7964__ & ~new_new_n7968__;
  assign new_new_n7970__ = ~new_new_n7964__ & new_new_n7968__;
  assign new_new_n7971__ = ~new_new_n7969__ & ~new_new_n7970__;
  assign new_new_n7972__ = new_new_n7963__ & ~new_new_n7971__;
  assign new_new_n7973__ = ~new_new_n7963__ & new_new_n7971__;
  assign new_new_n7974__ = ~new_new_n7972__ & ~new_new_n7973__;
  assign new_new_n7975__ = pi19 & pi37;
  assign new_new_n7976__ = pi04 & pi52;
  assign new_new_n7977__ = pi03 & pi53;
  assign new_new_n7978__ = ~new_new_n7976__ & ~new_new_n7977__;
  assign new_new_n7979__ = new_new_n7976__ & new_new_n7977__;
  assign new_new_n7980__ = ~new_new_n7978__ & ~new_new_n7979__;
  assign new_new_n7981__ = new_new_n7975__ & ~new_new_n7980__;
  assign new_new_n7982__ = ~new_new_n7975__ & new_new_n7980__;
  assign new_new_n7983__ = ~new_new_n7981__ & ~new_new_n7982__;
  assign new_new_n7984__ = ~new_new_n7974__ & new_new_n7983__;
  assign new_new_n7985__ = new_new_n7974__ & ~new_new_n7983__;
  assign new_new_n7986__ = ~new_new_n7984__ & ~new_new_n7985__;
  assign new_new_n7987__ = new_new_n7961__ & new_new_n7986__;
  assign new_new_n7988__ = ~new_new_n7961__ & ~new_new_n7986__;
  assign new_new_n7989__ = ~new_new_n7987__ & ~new_new_n7988__;
  assign new_new_n7990__ = ~new_new_n7664__ & ~new_new_n7675__;
  assign new_new_n7991__ = ~new_new_n7665__ & ~new_new_n7990__;
  assign new_new_n7992__ = pi01 & pi55;
  assign new_new_n7993__ = pi27 & pi29;
  assign new_new_n7994__ = new_new_n7992__ & ~new_new_n7993__;
  assign new_new_n7995__ = ~new_new_n7992__ & new_new_n7993__;
  assign new_new_n7996__ = ~new_new_n7994__ & ~new_new_n7995__;
  assign new_new_n7997__ = ~new_new_n7646__ & ~new_new_n7650__;
  assign new_new_n7998__ = ~new_new_n7649__ & ~new_new_n7997__;
  assign new_new_n7999__ = ~new_new_n7655__ & ~new_new_n7659__;
  assign new_new_n8000__ = ~new_new_n7658__ & ~new_new_n7999__;
  assign new_new_n8001__ = new_new_n7998__ & new_new_n8000__;
  assign new_new_n8002__ = ~new_new_n7998__ & ~new_new_n8000__;
  assign new_new_n8003__ = ~new_new_n8001__ & ~new_new_n8002__;
  assign new_new_n8004__ = new_new_n7996__ & new_new_n8003__;
  assign new_new_n8005__ = ~new_new_n7996__ & ~new_new_n8003__;
  assign new_new_n8006__ = ~new_new_n8004__ & ~new_new_n8005__;
  assign new_new_n8007__ = ~new_new_n7848__ & ~new_new_n7852__;
  assign new_new_n8008__ = ~new_new_n7851__ & ~new_new_n8007__;
  assign new_new_n8009__ = ~new_new_n7682__ & ~new_new_n7686__;
  assign new_new_n8010__ = ~new_new_n7685__ & ~new_new_n8009__;
  assign new_new_n8011__ = ~new_new_n7703__ & ~new_new_n7707__;
  assign new_new_n8012__ = ~new_new_n7706__ & ~new_new_n8011__;
  assign new_new_n8013__ = ~new_new_n8010__ & ~new_new_n8012__;
  assign new_new_n8014__ = new_new_n8010__ & new_new_n8012__;
  assign new_new_n8015__ = ~new_new_n8013__ & ~new_new_n8014__;
  assign new_new_n8016__ = new_new_n8008__ & ~new_new_n8015__;
  assign new_new_n8017__ = ~new_new_n8008__ & new_new_n8015__;
  assign new_new_n8018__ = ~new_new_n8016__ & ~new_new_n8017__;
  assign new_new_n8019__ = new_new_n8006__ & new_new_n8018__;
  assign new_new_n8020__ = ~new_new_n8006__ & ~new_new_n8018__;
  assign new_new_n8021__ = ~new_new_n8019__ & ~new_new_n8020__;
  assign new_new_n8022__ = new_new_n7991__ & ~new_new_n8021__;
  assign new_new_n8023__ = ~new_new_n7991__ & new_new_n8021__;
  assign new_new_n8024__ = ~new_new_n8022__ & ~new_new_n8023__;
  assign new_new_n8025__ = ~new_new_n7989__ & ~new_new_n8024__;
  assign new_new_n8026__ = new_new_n7989__ & new_new_n8024__;
  assign new_new_n8027__ = ~new_new_n8025__ & ~new_new_n8026__;
  assign new_new_n8028__ = ~new_new_n7864__ & ~new_new_n7868__;
  assign new_new_n8029__ = ~new_new_n7865__ & ~new_new_n8028__;
  assign new_new_n8030__ = new_new_n8027__ & ~new_new_n8029__;
  assign new_new_n8031__ = ~new_new_n8027__ & new_new_n8029__;
  assign new_new_n8032__ = ~new_new_n8030__ & ~new_new_n8031__;
  assign new_new_n8033__ = ~new_new_n7834__ & ~new_new_n7871__;
  assign new_new_n8034__ = ~new_new_n7835__ & ~new_new_n8033__;
  assign new_new_n8035__ = new_new_n8032__ & new_new_n8034__;
  assign new_new_n8036__ = ~new_new_n8032__ & ~new_new_n8034__;
  assign new_new_n8037__ = ~new_new_n8035__ & ~new_new_n8036__;
  assign new_new_n8038__ = ~new_new_n7700__ & ~new_new_n7711__;
  assign new_new_n8039__ = ~new_new_n7701__ & ~new_new_n8038__;
  assign new_new_n8040__ = ~new_new_n7726__ & ~new_new_n7732__;
  assign new_new_n8041__ = ~new_new_n7731__ & ~new_new_n8040__;
  assign new_new_n8042__ = new_new_n7807__ & new_new_n7814__;
  assign new_new_n8043__ = ~new_new_n7806__ & ~new_new_n8042__;
  assign new_new_n8044__ = new_new_n8041__ & new_new_n8043__;
  assign new_new_n8045__ = ~new_new_n8041__ & ~new_new_n8043__;
  assign new_new_n8046__ = ~new_new_n8044__ & ~new_new_n8045__;
  assign new_new_n8047__ = new_new_n8039__ & ~new_new_n8046__;
  assign new_new_n8048__ = ~new_new_n8039__ & new_new_n8046__;
  assign new_new_n8049__ = ~new_new_n8047__ & ~new_new_n8048__;
  assign new_new_n8050__ = ~new_new_n7752__ & ~new_new_n7774__;
  assign new_new_n8051__ = ~new_new_n7775__ & ~new_new_n8050__;
  assign new_new_n8052__ = ~new_new_n7857__ & new_new_n7860__;
  assign new_new_n8053__ = ~new_new_n7858__ & ~new_new_n8052__;
  assign new_new_n8054__ = new_new_n8051__ & ~new_new_n8053__;
  assign new_new_n8055__ = ~new_new_n8051__ & new_new_n8053__;
  assign new_new_n8056__ = ~new_new_n8054__ & ~new_new_n8055__;
  assign new_new_n8057__ = ~new_new_n3728__ & ~new_new_n7810__;
  assign new_new_n8058__ = ~new_new_n7809__ & ~new_new_n8057__;
  assign new_new_n8059__ = ~new_new_n7839__ & ~new_new_n7843__;
  assign new_new_n8060__ = ~new_new_n7842__ & ~new_new_n8059__;
  assign new_new_n8061__ = ~new_new_n8058__ & ~new_new_n8060__;
  assign new_new_n8062__ = new_new_n8058__ & new_new_n8060__;
  assign new_new_n8063__ = ~new_new_n7691__ & ~new_new_n7695__;
  assign new_new_n8064__ = ~new_new_n7694__ & ~new_new_n8063__;
  assign new_new_n8065__ = ~new_new_n8062__ & ~new_new_n8064__;
  assign new_new_n8066__ = ~new_new_n8061__ & new_new_n8065__;
  assign new_new_n8067__ = ~new_new_n8061__ & ~new_new_n8062__;
  assign new_new_n8068__ = new_new_n8064__ & ~new_new_n8067__;
  assign new_new_n8069__ = ~new_new_n8066__ & ~new_new_n8068__;
  assign new_new_n8070__ = new_new_n8056__ & new_new_n8069__;
  assign new_new_n8071__ = ~new_new_n8056__ & ~new_new_n8069__;
  assign new_new_n8072__ = ~new_new_n8070__ & ~new_new_n8071__;
  assign new_new_n8073__ = new_new_n8049__ & ~new_new_n8072__;
  assign new_new_n8074__ = ~new_new_n8049__ & new_new_n8072__;
  assign new_new_n8075__ = ~new_new_n7680__ & ~new_new_n7714__;
  assign new_new_n8076__ = ~new_new_n7679__ & ~new_new_n8075__;
  assign new_new_n8077__ = ~new_new_n8073__ & ~new_new_n8076__;
  assign new_new_n8078__ = ~new_new_n8074__ & ~new_new_n8077__;
  assign new_new_n8079__ = ~new_new_n8073__ & new_new_n8078__;
  assign new_new_n8080__ = ~new_new_n8074__ & new_new_n8077__;
  assign new_new_n8081__ = ~new_new_n8076__ & ~new_new_n8080__;
  assign new_new_n8082__ = ~new_new_n8079__ & ~new_new_n8081__;
  assign new_new_n8083__ = new_new_n8037__ & ~new_new_n8082__;
  assign new_new_n8084__ = ~new_new_n8037__ & new_new_n8082__;
  assign new_new_n8085__ = ~new_new_n8083__ & ~new_new_n8084__;
  assign new_new_n8086__ = new_new_n7892__ & ~new_new_n8085__;
  assign new_new_n8087__ = ~new_new_n7892__ & new_new_n8085__;
  assign new_new_n8088__ = ~new_new_n8086__ & ~new_new_n8087__;
  assign new_new_n8089__ = ~new_new_n7780__ & ~new_new_n7820__;
  assign new_new_n8090__ = ~new_new_n7781__ & ~new_new_n8089__;
  assign new_new_n8091__ = ~new_new_n7718__ & ~new_new_n7742__;
  assign new_new_n8092__ = ~new_new_n7719__ & ~new_new_n8091__;
  assign new_new_n8093__ = ~new_new_n8090__ & new_new_n8092__;
  assign new_new_n8094__ = new_new_n8090__ & ~new_new_n8092__;
  assign new_new_n8095__ = ~new_new_n8093__ & ~new_new_n8094__;
  assign new_new_n8096__ = ~new_new_n7722__ & ~new_new_n7738__;
  assign new_new_n8097__ = ~new_new_n7737__ & ~new_new_n8096__;
  assign new_new_n8098__ = ~new_new_n7799__ & ~new_new_n7817__;
  assign new_new_n8099__ = ~new_new_n7798__ & ~new_new_n8098__;
  assign new_new_n8100__ = new_new_n8097__ & ~new_new_n8099__;
  assign new_new_n8101__ = ~new_new_n8097__ & new_new_n8099__;
  assign new_new_n8102__ = ~new_new_n8100__ & ~new_new_n8101__;
  assign new_new_n8103__ = pi21 & pi35;
  assign new_new_n8104__ = pi18 & pi38;
  assign new_new_n8105__ = pi05 & pi51;
  assign new_new_n8106__ = ~new_new_n8104__ & ~new_new_n8105__;
  assign new_new_n8107__ = new_new_n8104__ & new_new_n8105__;
  assign new_new_n8108__ = ~new_new_n8106__ & ~new_new_n8107__;
  assign new_new_n8109__ = new_new_n8103__ & ~new_new_n8108__;
  assign new_new_n8110__ = ~new_new_n8103__ & new_new_n8108__;
  assign new_new_n8111__ = ~new_new_n8109__ & ~new_new_n8110__;
  assign new_new_n8112__ = ~new_new_n7760__ & ~new_new_n7766__;
  assign new_new_n8113__ = pi28 & ~new_new_n8112__;
  assign new_new_n8114__ = ~pi28 & new_new_n7765__;
  assign new_new_n8115__ = new_new_n7757__ & new_new_n8114__;
  assign new_new_n8116__ = ~new_new_n8113__ & ~new_new_n8115__;
  assign new_new_n8117__ = ~new_new_n8111__ & ~new_new_n8116__;
  assign new_new_n8118__ = new_new_n8111__ & new_new_n8116__;
  assign new_new_n8119__ = ~new_new_n8117__ & ~new_new_n8118__;
  assign new_new_n8120__ = ~new_new_n7787__ & ~new_new_n7793__;
  assign new_new_n8121__ = new_new_n8119__ & ~new_new_n8120__;
  assign new_new_n8122__ = ~new_new_n8119__ & new_new_n8120__;
  assign new_new_n8123__ = ~new_new_n8121__ & ~new_new_n8122__;
  assign new_new_n8124__ = new_new_n8102__ & ~new_new_n8123__;
  assign new_new_n8125__ = ~new_new_n8102__ & new_new_n8123__;
  assign new_new_n8126__ = ~new_new_n8124__ & ~new_new_n8125__;
  assign new_new_n8127__ = new_new_n8095__ & ~new_new_n8126__;
  assign new_new_n8128__ = ~new_new_n8095__ & new_new_n8126__;
  assign new_new_n8129__ = ~new_new_n8127__ & ~new_new_n8128__;
  assign new_new_n8130__ = new_new_n8088__ & new_new_n8129__;
  assign new_new_n8131__ = ~new_new_n8088__ & ~new_new_n8129__;
  assign new_new_n8132__ = ~new_new_n8130__ & ~new_new_n8131__;
  assign new_new_n8133__ = ~new_new_n7890__ & new_new_n8132__;
  assign new_new_n8134__ = new_new_n7890__ & ~new_new_n8132__;
  assign po057 = ~new_new_n8133__ & ~new_new_n8134__;
  assign new_new_n8136__ = ~new_new_n8035__ & ~new_new_n8082__;
  assign new_new_n8137__ = ~new_new_n8036__ & ~new_new_n8136__;
  assign new_new_n8138__ = ~new_new_n8093__ & ~new_new_n8127__;
  assign new_new_n8139__ = ~new_new_n7947__ & ~new_new_n7951__;
  assign new_new_n8140__ = ~new_new_n7950__ & ~new_new_n8139__;
  assign new_new_n8141__ = ~new_new_n8103__ & ~new_new_n8107__;
  assign new_new_n8142__ = ~new_new_n8106__ & ~new_new_n8141__;
  assign new_new_n8143__ = ~new_new_n8140__ & ~new_new_n8142__;
  assign new_new_n8144__ = new_new_n8140__ & new_new_n8142__;
  assign new_new_n8145__ = ~new_new_n8143__ & ~new_new_n8144__;
  assign new_new_n8146__ = ~new_new_n7914__ & ~new_new_n7918__;
  assign new_new_n8147__ = ~new_new_n7917__ & ~new_new_n8146__;
  assign new_new_n8148__ = ~new_new_n8145__ & new_new_n8147__;
  assign new_new_n8149__ = new_new_n8145__ & ~new_new_n8147__;
  assign new_new_n8150__ = ~new_new_n8148__ & ~new_new_n8149__;
  assign new_new_n8151__ = ~new_new_n8118__ & new_new_n8120__;
  assign new_new_n8152__ = ~new_new_n8117__ & ~new_new_n8151__;
  assign new_new_n8153__ = pi23 & pi34;
  assign new_new_n8154__ = pi22 & pi35;
  assign new_new_n8155__ = pi21 & pi36;
  assign new_new_n8156__ = ~new_new_n8154__ & ~new_new_n8155__;
  assign new_new_n8157__ = new_new_n8154__ & new_new_n8155__;
  assign new_new_n8158__ = ~new_new_n8156__ & ~new_new_n8157__;
  assign new_new_n8159__ = new_new_n8153__ & ~new_new_n8158__;
  assign new_new_n8160__ = ~new_new_n8153__ & new_new_n8158__;
  assign new_new_n8161__ = ~new_new_n8159__ & ~new_new_n8160__;
  assign new_new_n8162__ = pi26 & pi31;
  assign new_new_n8163__ = pi25 & pi32;
  assign new_new_n8164__ = pi24 & pi33;
  assign new_new_n8165__ = ~new_new_n8163__ & ~new_new_n8164__;
  assign new_new_n8166__ = new_new_n8163__ & new_new_n8164__;
  assign new_new_n8167__ = ~new_new_n8165__ & ~new_new_n8166__;
  assign new_new_n8168__ = new_new_n8162__ & ~new_new_n8167__;
  assign new_new_n8169__ = ~new_new_n8162__ & new_new_n8167__;
  assign new_new_n8170__ = ~new_new_n8168__ & ~new_new_n8169__;
  assign new_new_n8171__ = new_new_n8161__ & new_new_n8170__;
  assign new_new_n8172__ = ~new_new_n8161__ & ~new_new_n8170__;
  assign new_new_n8173__ = ~new_new_n8171__ & ~new_new_n8172__;
  assign new_new_n8174__ = pi16 & pi41;
  assign new_new_n8175__ = pi07 & pi50;
  assign new_new_n8176__ = pi08 & pi49;
  assign new_new_n8177__ = ~new_new_n8175__ & ~new_new_n8176__;
  assign new_new_n8178__ = new_new_n8175__ & new_new_n8176__;
  assign new_new_n8179__ = ~new_new_n8177__ & ~new_new_n8178__;
  assign new_new_n8180__ = new_new_n8174__ & ~new_new_n8179__;
  assign new_new_n8181__ = ~new_new_n8174__ & new_new_n8179__;
  assign new_new_n8182__ = ~new_new_n8180__ & ~new_new_n8181__;
  assign new_new_n8183__ = new_new_n8173__ & ~new_new_n8182__;
  assign new_new_n8184__ = ~new_new_n8173__ & new_new_n8182__;
  assign new_new_n8185__ = ~new_new_n8183__ & ~new_new_n8184__;
  assign new_new_n8186__ = new_new_n8152__ & ~new_new_n8185__;
  assign new_new_n8187__ = ~new_new_n8152__ & new_new_n8185__;
  assign new_new_n8188__ = ~new_new_n8186__ & ~new_new_n8187__;
  assign new_new_n8189__ = ~new_new_n8150__ & new_new_n8188__;
  assign new_new_n8190__ = new_new_n8150__ & ~new_new_n8188__;
  assign new_new_n8191__ = ~new_new_n8189__ & ~new_new_n8190__;
  assign new_new_n8192__ = new_new_n8039__ & ~new_new_n8044__;
  assign new_new_n8193__ = ~new_new_n8045__ & ~new_new_n8192__;
  assign new_new_n8194__ = pi18 & pi39;
  assign new_new_n8195__ = pi17 & pi40;
  assign new_new_n8196__ = pi06 & pi51;
  assign new_new_n8197__ = ~new_new_n8195__ & ~new_new_n8196__;
  assign new_new_n8198__ = new_new_n8195__ & new_new_n8196__;
  assign new_new_n8199__ = ~new_new_n8197__ & ~new_new_n8198__;
  assign new_new_n8200__ = new_new_n8194__ & ~new_new_n8199__;
  assign new_new_n8201__ = ~new_new_n8194__ & new_new_n8199__;
  assign new_new_n8202__ = ~new_new_n8200__ & ~new_new_n8201__;
  assign new_new_n8203__ = pi28 & pi29;
  assign new_new_n8204__ = pi12 & pi45;
  assign new_new_n8205__ = pi27 & pi30;
  assign new_new_n8206__ = ~new_new_n8204__ & ~new_new_n8205__;
  assign new_new_n8207__ = new_new_n8204__ & new_new_n8205__;
  assign new_new_n8208__ = ~new_new_n8206__ & ~new_new_n8207__;
  assign new_new_n8209__ = new_new_n8203__ & ~new_new_n8208__;
  assign new_new_n8210__ = ~new_new_n8203__ & new_new_n8208__;
  assign new_new_n8211__ = ~new_new_n8209__ & ~new_new_n8210__;
  assign new_new_n8212__ = new_new_n8202__ & new_new_n8211__;
  assign new_new_n8213__ = ~new_new_n8202__ & ~new_new_n8211__;
  assign new_new_n8214__ = ~new_new_n8212__ & ~new_new_n8213__;
  assign new_new_n8215__ = pi14 & pi43;
  assign new_new_n8216__ = pi13 & pi44;
  assign new_new_n8217__ = pi11 & pi46;
  assign new_new_n8218__ = ~new_new_n8216__ & ~new_new_n8217__;
  assign new_new_n8219__ = new_new_n8216__ & new_new_n8217__;
  assign new_new_n8220__ = ~new_new_n8218__ & ~new_new_n8219__;
  assign new_new_n8221__ = new_new_n8215__ & ~new_new_n8220__;
  assign new_new_n8222__ = ~new_new_n8215__ & new_new_n8220__;
  assign new_new_n8223__ = ~new_new_n8221__ & ~new_new_n8222__;
  assign new_new_n8224__ = ~new_new_n8214__ & new_new_n8223__;
  assign new_new_n8225__ = new_new_n8214__ & ~new_new_n8223__;
  assign new_new_n8226__ = ~new_new_n8224__ & ~new_new_n8225__;
  assign new_new_n8227__ = new_new_n8193__ & new_new_n8226__;
  assign new_new_n8228__ = ~new_new_n8193__ & ~new_new_n8226__;
  assign new_new_n8229__ = ~new_new_n8227__ & ~new_new_n8228__;
  assign new_new_n8230__ = pi04 & pi53;
  assign new_new_n8231__ = pi02 & pi55;
  assign new_new_n8232__ = pi03 & pi54;
  assign new_new_n8233__ = ~new_new_n8231__ & ~new_new_n8232__;
  assign new_new_n8234__ = new_new_n8231__ & new_new_n8232__;
  assign new_new_n8235__ = ~new_new_n8233__ & ~new_new_n8234__;
  assign new_new_n8236__ = new_new_n8230__ & ~new_new_n8235__;
  assign new_new_n8237__ = ~new_new_n8230__ & new_new_n8235__;
  assign new_new_n8238__ = ~new_new_n8236__ & ~new_new_n8237__;
  assign new_new_n8239__ = pi20 & pi37;
  assign new_new_n8240__ = pi19 & pi38;
  assign new_new_n8241__ = pi05 & pi52;
  assign new_new_n8242__ = ~new_new_n8240__ & ~new_new_n8241__;
  assign new_new_n8243__ = new_new_n8240__ & new_new_n8241__;
  assign new_new_n8244__ = ~new_new_n8242__ & ~new_new_n8243__;
  assign new_new_n8245__ = new_new_n8239__ & ~new_new_n8244__;
  assign new_new_n8246__ = ~new_new_n8239__ & new_new_n8244__;
  assign new_new_n8247__ = ~new_new_n8245__ & ~new_new_n8246__;
  assign new_new_n8248__ = pi15 & pi42;
  assign new_new_n8249__ = pi10 & pi47;
  assign new_new_n8250__ = pi09 & pi48;
  assign new_new_n8251__ = ~new_new_n8249__ & ~new_new_n8250__;
  assign new_new_n8252__ = new_new_n8249__ & new_new_n8250__;
  assign new_new_n8253__ = ~new_new_n8251__ & ~new_new_n8252__;
  assign new_new_n8254__ = new_new_n8248__ & ~new_new_n8253__;
  assign new_new_n8255__ = ~new_new_n8248__ & new_new_n8253__;
  assign new_new_n8256__ = ~new_new_n8254__ & ~new_new_n8255__;
  assign new_new_n8257__ = new_new_n8247__ & new_new_n8256__;
  assign new_new_n8258__ = ~new_new_n8247__ & ~new_new_n8256__;
  assign new_new_n8259__ = ~new_new_n8238__ & ~new_new_n8257__;
  assign new_new_n8260__ = ~new_new_n8258__ & ~new_new_n8259__;
  assign new_new_n8261__ = ~new_new_n8257__ & new_new_n8260__;
  assign new_new_n8262__ = new_new_n8238__ & ~new_new_n8261__;
  assign new_new_n8263__ = ~new_new_n8258__ & new_new_n8259__;
  assign new_new_n8264__ = ~new_new_n8262__ & ~new_new_n8263__;
  assign new_new_n8265__ = new_new_n8229__ & ~new_new_n8264__;
  assign new_new_n8266__ = ~new_new_n8229__ & new_new_n8264__;
  assign new_new_n8267__ = ~new_new_n8265__ & ~new_new_n8266__;
  assign new_new_n8268__ = ~new_new_n8191__ & new_new_n8267__;
  assign new_new_n8269__ = ~new_new_n8100__ & ~new_new_n8123__;
  assign new_new_n8270__ = new_new_n8191__ & ~new_new_n8267__;
  assign new_new_n8271__ = ~new_new_n8101__ & ~new_new_n8269__;
  assign new_new_n8272__ = ~new_new_n8270__ & new_new_n8271__;
  assign new_new_n8273__ = ~new_new_n8268__ & new_new_n8272__;
  assign new_new_n8274__ = ~new_new_n8097__ & new_new_n8270__;
  assign new_new_n8275__ = new_new_n8099__ & new_new_n8268__;
  assign new_new_n8276__ = ~new_new_n8274__ & ~new_new_n8275__;
  assign new_new_n8277__ = ~new_new_n8123__ & ~new_new_n8276__;
  assign new_new_n8278__ = ~new_new_n8097__ & new_new_n8268__;
  assign new_new_n8279__ = new_new_n8099__ & new_new_n8270__;
  assign new_new_n8280__ = ~new_new_n8278__ & ~new_new_n8279__;
  assign new_new_n8281__ = ~new_new_n8126__ & ~new_new_n8280__;
  assign new_new_n8282__ = ~new_new_n8273__ & ~new_new_n8277__;
  assign new_new_n8283__ = ~new_new_n8281__ & new_new_n8282__;
  assign new_new_n8284__ = ~new_new_n8138__ & new_new_n8283__;
  assign new_new_n8285__ = new_new_n8138__ & ~new_new_n8283__;
  assign new_new_n8286__ = ~new_new_n8284__ & ~new_new_n8285__;
  assign new_new_n8287__ = ~new_new_n7911__ & ~new_new_n7922__;
  assign new_new_n8288__ = ~new_new_n7912__ & ~new_new_n8287__;
  assign new_new_n8289__ = ~new_new_n7964__ & ~new_new_n7965__;
  assign new_new_n8290__ = new_new_n7967__ & ~new_new_n8289__;
  assign new_new_n8291__ = ~new_new_n7935__ & ~new_new_n7939__;
  assign new_new_n8292__ = ~new_new_n7938__ & ~new_new_n8291__;
  assign new_new_n8293__ = new_new_n8290__ & new_new_n8292__;
  assign new_new_n8294__ = ~new_new_n8290__ & ~new_new_n8292__;
  assign new_new_n8295__ = ~new_new_n8293__ & ~new_new_n8294__;
  assign new_new_n8296__ = ~new_new_n7975__ & ~new_new_n7979__;
  assign new_new_n8297__ = ~new_new_n7978__ & ~new_new_n8296__;
  assign new_new_n8298__ = ~new_new_n8295__ & new_new_n8297__;
  assign new_new_n8299__ = ~new_new_n8293__ & ~new_new_n8297__;
  assign new_new_n8300__ = ~new_new_n8294__ & new_new_n8299__;
  assign new_new_n8301__ = ~new_new_n8298__ & ~new_new_n8300__;
  assign new_new_n8302__ = new_new_n8288__ & ~new_new_n8301__;
  assign new_new_n8303__ = ~new_new_n8288__ & new_new_n8301__;
  assign new_new_n8304__ = ~new_new_n8302__ & ~new_new_n8303__;
  assign new_new_n8305__ = ~new_new_n7902__ & ~new_new_n7906__;
  assign new_new_n8306__ = ~new_new_n7905__ & ~new_new_n8305__;
  assign new_new_n8307__ = ~new_new_n7926__ & ~new_new_n7930__;
  assign new_new_n8308__ = ~new_new_n7929__ & ~new_new_n8307__;
  assign new_new_n8309__ = ~new_new_n7893__ & ~new_new_n7897__;
  assign new_new_n8310__ = ~new_new_n7896__ & ~new_new_n8309__;
  assign new_new_n8311__ = new_new_n8308__ & new_new_n8310__;
  assign new_new_n8312__ = ~new_new_n8308__ & ~new_new_n8310__;
  assign new_new_n8313__ = ~new_new_n8311__ & ~new_new_n8312__;
  assign new_new_n8314__ = new_new_n8306__ & ~new_new_n8313__;
  assign new_new_n8315__ = ~new_new_n8306__ & new_new_n8313__;
  assign new_new_n8316__ = ~new_new_n8314__ & ~new_new_n8315__;
  assign new_new_n8317__ = new_new_n8304__ & new_new_n8316__;
  assign new_new_n8318__ = ~new_new_n8304__ & ~new_new_n8316__;
  assign new_new_n8319__ = ~new_new_n8317__ & ~new_new_n8318__;
  assign new_new_n8320__ = new_new_n7996__ & ~new_new_n8001__;
  assign new_new_n8321__ = ~new_new_n8002__ & ~new_new_n8320__;
  assign new_new_n8322__ = ~new_new_n7972__ & new_new_n7983__;
  assign new_new_n8323__ = ~new_new_n7973__ & ~new_new_n8322__;
  assign new_new_n8324__ = new_new_n8321__ & new_new_n8323__;
  assign new_new_n8325__ = ~new_new_n8321__ & ~new_new_n8323__;
  assign new_new_n8326__ = ~new_new_n8324__ & ~new_new_n8325__;
  assign new_new_n8327__ = ~new_new_n7944__ & ~new_new_n7955__;
  assign new_new_n8328__ = ~new_new_n7945__ & ~new_new_n8327__;
  assign new_new_n8329__ = new_new_n8326__ & ~new_new_n8328__;
  assign new_new_n8330__ = ~new_new_n8326__ & new_new_n8328__;
  assign new_new_n8331__ = ~new_new_n8329__ & ~new_new_n8330__;
  assign new_new_n8332__ = ~new_new_n8319__ & ~new_new_n8331__;
  assign new_new_n8333__ = new_new_n8319__ & new_new_n8331__;
  assign new_new_n8334__ = ~new_new_n8332__ & ~new_new_n8333__;
  assign new_new_n8335__ = ~new_new_n7960__ & ~new_new_n7986__;
  assign new_new_n8336__ = ~new_new_n7959__ & ~new_new_n8335__;
  assign new_new_n8337__ = new_new_n8334__ & ~new_new_n8336__;
  assign new_new_n8338__ = ~new_new_n8334__ & new_new_n8336__;
  assign new_new_n8339__ = ~new_new_n8337__ & ~new_new_n8338__;
  assign new_new_n8340__ = new_new_n8286__ & ~new_new_n8339__;
  assign new_new_n8341__ = ~new_new_n8286__ & new_new_n8339__;
  assign new_new_n8342__ = ~new_new_n8340__ & ~new_new_n8341__;
  assign new_new_n8343__ = new_new_n8137__ & new_new_n8342__;
  assign new_new_n8344__ = ~new_new_n8137__ & ~new_new_n8342__;
  assign new_new_n8345__ = ~new_new_n8343__ & ~new_new_n8344__;
  assign new_new_n8346__ = ~new_new_n8087__ & ~new_new_n8129__;
  assign new_new_n8347__ = ~new_new_n8086__ & ~new_new_n8346__;
  assign new_new_n8348__ = ~new_new_n7889__ & new_new_n8132__;
  assign new_new_n8349__ = ~new_new_n7888__ & ~new_new_n8348__;
  assign new_new_n8350__ = new_new_n8347__ & ~new_new_n8349__;
  assign new_new_n8351__ = ~new_new_n8347__ & new_new_n8349__;
  assign new_new_n8352__ = ~new_new_n8350__ & ~new_new_n8351__;
  assign new_new_n8353__ = ~new_new_n8025__ & ~new_new_n8029__;
  assign new_new_n8354__ = ~new_new_n8026__ & ~new_new_n8353__;
  assign new_new_n8355__ = ~new_new_n8078__ & new_new_n8354__;
  assign new_new_n8356__ = new_new_n8078__ & ~new_new_n8354__;
  assign new_new_n8357__ = ~new_new_n8355__ & ~new_new_n8356__;
  assign new_new_n8358__ = ~new_new_n8055__ & ~new_new_n8069__;
  assign new_new_n8359__ = ~new_new_n8054__ & ~new_new_n8358__;
  assign new_new_n8360__ = ~new_new_n8008__ & ~new_new_n8014__;
  assign new_new_n8361__ = ~new_new_n8013__ & ~new_new_n8360__;
  assign new_new_n8362__ = ~new_new_n8061__ & ~new_new_n8065__;
  assign new_new_n8363__ = pi27 & pi55;
  assign new_new_n8364__ = pi01 & new_new_n8363__;
  assign new_new_n8365__ = pi29 & ~new_new_n8364__;
  assign new_new_n8366__ = pi00 & pi57;
  assign new_new_n8367__ = pi01 & pi56;
  assign new_new_n8368__ = new_new_n8366__ & ~new_new_n8367__;
  assign new_new_n8369__ = ~new_new_n8366__ & new_new_n8367__;
  assign new_new_n8370__ = ~new_new_n8368__ & ~new_new_n8369__;
  assign new_new_n8371__ = new_new_n8365__ & new_new_n8370__;
  assign new_new_n8372__ = ~new_new_n8365__ & ~new_new_n8370__;
  assign new_new_n8373__ = ~new_new_n8371__ & ~new_new_n8372__;
  assign new_new_n8374__ = new_new_n8362__ & ~new_new_n8373__;
  assign new_new_n8375__ = ~new_new_n8362__ & new_new_n8373__;
  assign new_new_n8376__ = ~new_new_n8374__ & ~new_new_n8375__;
  assign new_new_n8377__ = new_new_n8361__ & new_new_n8376__;
  assign new_new_n8378__ = ~new_new_n8361__ & ~new_new_n8376__;
  assign new_new_n8379__ = ~new_new_n8377__ & ~new_new_n8378__;
  assign new_new_n8380__ = new_new_n8359__ & ~new_new_n8379__;
  assign new_new_n8381__ = ~new_new_n8359__ & new_new_n8379__;
  assign new_new_n8382__ = ~new_new_n8380__ & ~new_new_n8381__;
  assign new_new_n8383__ = ~new_new_n7991__ & ~new_new_n8019__;
  assign new_new_n8384__ = ~new_new_n8020__ & ~new_new_n8383__;
  assign new_new_n8385__ = new_new_n8382__ & new_new_n8384__;
  assign new_new_n8386__ = ~new_new_n8382__ & ~new_new_n8384__;
  assign new_new_n8387__ = ~new_new_n8385__ & ~new_new_n8386__;
  assign new_new_n8388__ = new_new_n8357__ & ~new_new_n8387__;
  assign new_new_n8389__ = ~new_new_n8357__ & new_new_n8387__;
  assign new_new_n8390__ = ~new_new_n8388__ & ~new_new_n8389__;
  assign new_new_n8391__ = new_new_n8352__ & ~new_new_n8390__;
  assign new_new_n8392__ = ~new_new_n8352__ & new_new_n8390__;
  assign new_new_n8393__ = ~new_new_n8391__ & ~new_new_n8392__;
  assign new_new_n8394__ = new_new_n8345__ & new_new_n8393__;
  assign new_new_n8395__ = ~new_new_n8345__ & ~new_new_n8393__;
  assign po058 = new_new_n8394__ | new_new_n8395__;
  assign new_new_n8397__ = new_new_n8342__ & ~new_new_n8347__;
  assign new_new_n8398__ = new_new_n8349__ & new_new_n8397__;
  assign new_new_n8399__ = new_new_n8137__ & new_new_n8398__;
  assign new_new_n8400__ = ~new_new_n8342__ & ~new_new_n8351__;
  assign new_new_n8401__ = ~new_new_n8350__ & ~new_new_n8400__;
  assign new_new_n8402__ = ~new_new_n8137__ & ~new_new_n8401__;
  assign new_new_n8403__ = ~new_new_n8342__ & new_new_n8347__;
  assign new_new_n8404__ = ~new_new_n8349__ & new_new_n8403__;
  assign new_new_n8405__ = ~new_new_n8402__ & ~new_new_n8404__;
  assign new_new_n8406__ = ~new_new_n8390__ & ~new_new_n8405__;
  assign new_new_n8407__ = new_new_n8137__ & new_new_n8401__;
  assign new_new_n8408__ = ~new_new_n8398__ & ~new_new_n8407__;
  assign new_new_n8409__ = new_new_n8390__ & ~new_new_n8408__;
  assign new_new_n8410__ = ~new_new_n8137__ & ~new_new_n8349__;
  assign new_new_n8411__ = new_new_n8403__ & new_new_n8410__;
  assign new_new_n8412__ = ~new_new_n8285__ & new_new_n8339__;
  assign new_new_n8413__ = ~new_new_n8284__ & ~new_new_n8412__;
  assign new_new_n8414__ = ~new_new_n8355__ & ~new_new_n8387__;
  assign new_new_n8415__ = ~new_new_n8356__ & ~new_new_n8414__;
  assign new_new_n8416__ = ~new_new_n8227__ & ~new_new_n8264__;
  assign new_new_n8417__ = ~new_new_n8228__ & ~new_new_n8416__;
  assign new_new_n8418__ = ~new_new_n8215__ & ~new_new_n8219__;
  assign new_new_n8419__ = ~new_new_n8218__ & ~new_new_n8418__;
  assign new_new_n8420__ = ~new_new_n8248__ & ~new_new_n8252__;
  assign new_new_n8421__ = ~new_new_n8251__ & ~new_new_n8420__;
  assign new_new_n8422__ = ~new_new_n8162__ & ~new_new_n8166__;
  assign new_new_n8423__ = ~new_new_n8165__ & ~new_new_n8422__;
  assign new_new_n8424__ = new_new_n8421__ & new_new_n8423__;
  assign new_new_n8425__ = ~new_new_n8421__ & ~new_new_n8423__;
  assign new_new_n8426__ = ~new_new_n8424__ & ~new_new_n8425__;
  assign new_new_n8427__ = new_new_n8419__ & ~new_new_n8426__;
  assign new_new_n8428__ = ~new_new_n8419__ & new_new_n8426__;
  assign new_new_n8429__ = ~new_new_n8427__ & ~new_new_n8428__;
  assign new_new_n8430__ = ~new_new_n8171__ & ~new_new_n8182__;
  assign new_new_n8431__ = ~new_new_n8172__ & ~new_new_n8430__;
  assign new_new_n8432__ = ~new_new_n8153__ & ~new_new_n8157__;
  assign new_new_n8433__ = ~new_new_n8156__ & ~new_new_n8432__;
  assign new_new_n8434__ = ~new_new_n8239__ & ~new_new_n8243__;
  assign new_new_n8435__ = ~new_new_n8242__ & ~new_new_n8434__;
  assign new_new_n8436__ = ~new_new_n8230__ & ~new_new_n8234__;
  assign new_new_n8437__ = ~new_new_n8233__ & ~new_new_n8436__;
  assign new_new_n8438__ = new_new_n8435__ & ~new_new_n8437__;
  assign new_new_n8439__ = ~new_new_n8435__ & new_new_n8437__;
  assign new_new_n8440__ = ~new_new_n8438__ & ~new_new_n8439__;
  assign new_new_n8441__ = new_new_n8433__ & new_new_n8440__;
  assign new_new_n8442__ = ~new_new_n8433__ & ~new_new_n8440__;
  assign new_new_n8443__ = ~new_new_n8441__ & ~new_new_n8442__;
  assign new_new_n8444__ = new_new_n8431__ & ~new_new_n8443__;
  assign new_new_n8445__ = ~new_new_n8431__ & new_new_n8443__;
  assign new_new_n8446__ = ~new_new_n8444__ & ~new_new_n8445__;
  assign new_new_n8447__ = new_new_n8429__ & new_new_n8446__;
  assign new_new_n8448__ = ~new_new_n8429__ & ~new_new_n8446__;
  assign new_new_n8449__ = ~new_new_n8447__ & ~new_new_n8448__;
  assign new_new_n8450__ = new_new_n8417__ & new_new_n8449__;
  assign new_new_n8451__ = ~new_new_n8417__ & ~new_new_n8449__;
  assign new_new_n8452__ = ~new_new_n8450__ & ~new_new_n8451__;
  assign new_new_n8453__ = ~new_new_n8212__ & ~new_new_n8223__;
  assign new_new_n8454__ = ~new_new_n8213__ & ~new_new_n8453__;
  assign new_new_n8455__ = ~new_new_n8203__ & ~new_new_n8207__;
  assign new_new_n8456__ = ~new_new_n8206__ & ~new_new_n8455__;
  assign new_new_n8457__ = pi28 & pi30;
  assign new_new_n8458__ = pi29 & pi56;
  assign new_new_n8459__ = ~pi57 & ~new_new_n8458__;
  assign new_new_n8460__ = pi29 & pi57;
  assign new_new_n8461__ = pi56 & new_new_n8460__;
  assign new_new_n8462__ = pi01 & ~new_new_n8459__;
  assign new_new_n8463__ = ~new_new_n8461__ & new_new_n8462__;
  assign new_new_n8464__ = new_new_n8457__ & ~new_new_n8463__;
  assign new_new_n8465__ = ~new_new_n8457__ & new_new_n8463__;
  assign new_new_n8466__ = ~new_new_n8464__ & ~new_new_n8465__;
  assign new_new_n8467__ = new_new_n8456__ & new_new_n8466__;
  assign new_new_n8468__ = ~new_new_n8456__ & ~new_new_n8466__;
  assign new_new_n8469__ = ~new_new_n8467__ & ~new_new_n8468__;
  assign new_new_n8470__ = new_new_n8454__ & new_new_n8469__;
  assign new_new_n8471__ = ~new_new_n8454__ & ~new_new_n8469__;
  assign new_new_n8472__ = ~new_new_n8260__ & ~new_new_n8470__;
  assign new_new_n8473__ = ~new_new_n8471__ & ~new_new_n8472__;
  assign new_new_n8474__ = ~new_new_n8470__ & new_new_n8473__;
  assign new_new_n8475__ = ~new_new_n8471__ & new_new_n8472__;
  assign new_new_n8476__ = ~new_new_n8260__ & ~new_new_n8475__;
  assign new_new_n8477__ = ~new_new_n8474__ & ~new_new_n8476__;
  assign new_new_n8478__ = new_new_n8452__ & ~new_new_n8477__;
  assign new_new_n8479__ = ~new_new_n8452__ & new_new_n8477__;
  assign new_new_n8480__ = ~new_new_n8478__ & ~new_new_n8479__;
  assign new_new_n8481__ = ~new_new_n8415__ & new_new_n8480__;
  assign new_new_n8482__ = new_new_n8415__ & ~new_new_n8480__;
  assign new_new_n8483__ = ~new_new_n8481__ & ~new_new_n8482__;
  assign new_new_n8484__ = new_new_n8361__ & ~new_new_n8375__;
  assign new_new_n8485__ = ~new_new_n8374__ & ~new_new_n8484__;
  assign new_new_n8486__ = ~new_new_n8194__ & ~new_new_n8198__;
  assign new_new_n8487__ = ~new_new_n8197__ & ~new_new_n8486__;
  assign new_new_n8488__ = pi56 & ~new_new_n8366__;
  assign new_new_n8489__ = new_new_n8364__ & ~new_new_n8488__;
  assign new_new_n8490__ = ~new_new_n8368__ & ~new_new_n8489__;
  assign new_new_n8491__ = pi29 & ~new_new_n8490__;
  assign new_new_n8492__ = ~pi29 & new_new_n8366__;
  assign new_new_n8493__ = new_new_n8367__ & new_new_n8492__;
  assign new_new_n8494__ = ~new_new_n8491__ & ~new_new_n8493__;
  assign new_new_n8495__ = ~new_new_n8487__ & new_new_n8494__;
  assign new_new_n8496__ = new_new_n8487__ & ~new_new_n8494__;
  assign new_new_n8497__ = ~new_new_n8495__ & ~new_new_n8496__;
  assign new_new_n8498__ = ~new_new_n8174__ & ~new_new_n8178__;
  assign new_new_n8499__ = ~new_new_n8177__ & ~new_new_n8498__;
  assign new_new_n8500__ = pi15 & pi43;
  assign new_new_n8501__ = pi10 & pi48;
  assign new_new_n8502__ = pi11 & pi47;
  assign new_new_n8503__ = ~new_new_n8501__ & ~new_new_n8502__;
  assign new_new_n8504__ = new_new_n8501__ & new_new_n8502__;
  assign new_new_n8505__ = ~new_new_n8503__ & ~new_new_n8504__;
  assign new_new_n8506__ = new_new_n8500__ & ~new_new_n8505__;
  assign new_new_n8507__ = ~new_new_n8500__ & new_new_n8505__;
  assign new_new_n8508__ = ~new_new_n8506__ & ~new_new_n8507__;
  assign new_new_n8509__ = pi19 & pi39;
  assign new_new_n8510__ = pi06 & pi52;
  assign new_new_n8511__ = pi03 & pi55;
  assign new_new_n8512__ = ~new_new_n8510__ & ~new_new_n8511__;
  assign new_new_n8513__ = new_new_n8510__ & new_new_n8511__;
  assign new_new_n8514__ = ~new_new_n8512__ & ~new_new_n8513__;
  assign new_new_n8515__ = new_new_n8509__ & ~new_new_n8514__;
  assign new_new_n8516__ = ~new_new_n8509__ & new_new_n8514__;
  assign new_new_n8517__ = ~new_new_n8515__ & ~new_new_n8516__;
  assign new_new_n8518__ = new_new_n8508__ & new_new_n8517__;
  assign new_new_n8519__ = ~new_new_n8508__ & ~new_new_n8517__;
  assign new_new_n8520__ = ~new_new_n8518__ & ~new_new_n8519__;
  assign new_new_n8521__ = pi14 & pi44;
  assign new_new_n8522__ = pi13 & pi45;
  assign new_new_n8523__ = pi12 & pi46;
  assign new_new_n8524__ = ~new_new_n8522__ & ~new_new_n8523__;
  assign new_new_n8525__ = new_new_n8522__ & new_new_n8523__;
  assign new_new_n8526__ = ~new_new_n8524__ & ~new_new_n8525__;
  assign new_new_n8527__ = new_new_n8521__ & ~new_new_n8526__;
  assign new_new_n8528__ = ~new_new_n8521__ & new_new_n8526__;
  assign new_new_n8529__ = ~new_new_n8527__ & ~new_new_n8528__;
  assign new_new_n8530__ = ~new_new_n8520__ & new_new_n8529__;
  assign new_new_n8531__ = new_new_n8520__ & ~new_new_n8529__;
  assign new_new_n8532__ = ~new_new_n8530__ & ~new_new_n8531__;
  assign new_new_n8533__ = new_new_n8499__ & new_new_n8532__;
  assign new_new_n8534__ = ~new_new_n8499__ & ~new_new_n8532__;
  assign new_new_n8535__ = ~new_new_n8533__ & ~new_new_n8534__;
  assign new_new_n8536__ = new_new_n8497__ & ~new_new_n8535__;
  assign new_new_n8537__ = ~new_new_n8497__ & new_new_n8535__;
  assign new_new_n8538__ = ~new_new_n8536__ & ~new_new_n8537__;
  assign new_new_n8539__ = new_new_n8485__ & new_new_n8538__;
  assign new_new_n8540__ = ~new_new_n8485__ & ~new_new_n8538__;
  assign new_new_n8541__ = ~new_new_n8539__ & ~new_new_n8540__;
  assign new_new_n8542__ = ~new_new_n8324__ & new_new_n8328__;
  assign new_new_n8543__ = ~new_new_n8325__ & ~new_new_n8542__;
  assign new_new_n8544__ = pi27 & pi31;
  assign new_new_n8545__ = pi25 & pi33;
  assign new_new_n8546__ = pi26 & pi32;
  assign new_new_n8547__ = ~new_new_n8545__ & ~new_new_n8546__;
  assign new_new_n8548__ = new_new_n8545__ & new_new_n8546__;
  assign new_new_n8549__ = ~new_new_n8547__ & ~new_new_n8548__;
  assign new_new_n8550__ = new_new_n8544__ & ~new_new_n8549__;
  assign new_new_n8551__ = ~new_new_n8544__ & new_new_n8549__;
  assign new_new_n8552__ = ~new_new_n8550__ & ~new_new_n8551__;
  assign new_new_n8553__ = pi24 & pi34;
  assign new_new_n8554__ = pi22 & pi36;
  assign new_new_n8555__ = pi23 & pi35;
  assign new_new_n8556__ = ~new_new_n8554__ & ~new_new_n8555__;
  assign new_new_n8557__ = new_new_n8554__ & new_new_n8555__;
  assign new_new_n8558__ = ~new_new_n8556__ & ~new_new_n8557__;
  assign new_new_n8559__ = new_new_n8553__ & ~new_new_n8558__;
  assign new_new_n8560__ = ~new_new_n8553__ & new_new_n8558__;
  assign new_new_n8561__ = ~new_new_n8559__ & ~new_new_n8560__;
  assign new_new_n8562__ = new_new_n8552__ & new_new_n8561__;
  assign new_new_n8563__ = ~new_new_n8552__ & ~new_new_n8561__;
  assign new_new_n8564__ = ~new_new_n8562__ & ~new_new_n8563__;
  assign new_new_n8565__ = pi18 & pi40;
  assign new_new_n8566__ = pi08 & pi50;
  assign new_new_n8567__ = pi07 & pi51;
  assign new_new_n8568__ = ~new_new_n8566__ & ~new_new_n8567__;
  assign new_new_n8569__ = new_new_n8566__ & new_new_n8567__;
  assign new_new_n8570__ = ~new_new_n8568__ & ~new_new_n8569__;
  assign new_new_n8571__ = new_new_n8565__ & ~new_new_n8570__;
  assign new_new_n8572__ = ~new_new_n8565__ & new_new_n8570__;
  assign new_new_n8573__ = ~new_new_n8571__ & ~new_new_n8572__;
  assign new_new_n8574__ = new_new_n8564__ & ~new_new_n8573__;
  assign new_new_n8575__ = ~new_new_n8564__ & new_new_n8573__;
  assign new_new_n8576__ = ~new_new_n8574__ & ~new_new_n8575__;
  assign new_new_n8577__ = ~new_new_n8543__ & ~new_new_n8576__;
  assign new_new_n8578__ = new_new_n8543__ & new_new_n8576__;
  assign new_new_n8579__ = ~new_new_n8577__ & ~new_new_n8578__;
  assign new_new_n8580__ = pi21 & pi37;
  assign new_new_n8581__ = pi05 & pi53;
  assign new_new_n8582__ = ~new_new_n4093__ & ~new_new_n8581__;
  assign new_new_n8583__ = new_new_n4093__ & new_new_n8581__;
  assign new_new_n8584__ = ~new_new_n8582__ & ~new_new_n8583__;
  assign new_new_n8585__ = new_new_n8580__ & ~new_new_n8584__;
  assign new_new_n8586__ = ~new_new_n8580__ & new_new_n8584__;
  assign new_new_n8587__ = ~new_new_n8585__ & ~new_new_n8586__;
  assign new_new_n8588__ = pi04 & pi54;
  assign new_new_n8589__ = pi02 & pi56;
  assign new_new_n8590__ = pi00 & pi58;
  assign new_new_n8591__ = ~new_new_n8589__ & ~new_new_n8590__;
  assign new_new_n8592__ = new_new_n8589__ & new_new_n8590__;
  assign new_new_n8593__ = ~new_new_n8591__ & ~new_new_n8592__;
  assign new_new_n8594__ = new_new_n8588__ & ~new_new_n8593__;
  assign new_new_n8595__ = ~new_new_n8588__ & new_new_n8593__;
  assign new_new_n8596__ = ~new_new_n8594__ & ~new_new_n8595__;
  assign new_new_n8597__ = new_new_n8587__ & new_new_n8596__;
  assign new_new_n8598__ = ~new_new_n8587__ & ~new_new_n8596__;
  assign new_new_n8599__ = ~new_new_n8597__ & ~new_new_n8598__;
  assign new_new_n8600__ = pi17 & pi41;
  assign new_new_n8601__ = pi16 & pi42;
  assign new_new_n8602__ = pi09 & pi49;
  assign new_new_n8603__ = ~new_new_n8601__ & ~new_new_n8602__;
  assign new_new_n8604__ = new_new_n8601__ & new_new_n8602__;
  assign new_new_n8605__ = ~new_new_n8603__ & ~new_new_n8604__;
  assign new_new_n8606__ = new_new_n8600__ & ~new_new_n8605__;
  assign new_new_n8607__ = ~new_new_n8600__ & new_new_n8605__;
  assign new_new_n8608__ = ~new_new_n8606__ & ~new_new_n8607__;
  assign new_new_n8609__ = ~new_new_n8599__ & new_new_n8608__;
  assign new_new_n8610__ = new_new_n8599__ & ~new_new_n8608__;
  assign new_new_n8611__ = ~new_new_n8609__ & ~new_new_n8610__;
  assign new_new_n8612__ = new_new_n8579__ & new_new_n8611__;
  assign new_new_n8613__ = ~new_new_n8579__ & ~new_new_n8611__;
  assign new_new_n8614__ = ~new_new_n8612__ & ~new_new_n8613__;
  assign new_new_n8615__ = ~new_new_n8541__ & ~new_new_n8614__;
  assign new_new_n8616__ = new_new_n8541__ & new_new_n8614__;
  assign new_new_n8617__ = ~new_new_n8615__ & ~new_new_n8616__;
  assign new_new_n8618__ = ~new_new_n8380__ & ~new_new_n8384__;
  assign new_new_n8619__ = ~new_new_n8381__ & ~new_new_n8618__;
  assign new_new_n8620__ = new_new_n8617__ & new_new_n8619__;
  assign new_new_n8621__ = ~new_new_n8617__ & ~new_new_n8619__;
  assign new_new_n8622__ = ~new_new_n8620__ & ~new_new_n8621__;
  assign new_new_n8623__ = new_new_n8483__ & new_new_n8622__;
  assign new_new_n8624__ = ~new_new_n8483__ & ~new_new_n8622__;
  assign new_new_n8625__ = ~new_new_n8623__ & ~new_new_n8624__;
  assign new_new_n8626__ = new_new_n8413__ & ~new_new_n8625__;
  assign new_new_n8627__ = ~new_new_n8413__ & new_new_n8625__;
  assign new_new_n8628__ = ~new_new_n8626__ & ~new_new_n8627__;
  assign new_new_n8629__ = ~new_new_n8268__ & ~new_new_n8272__;
  assign new_new_n8630__ = ~new_new_n8333__ & ~new_new_n8336__;
  assign new_new_n8631__ = ~new_new_n8332__ & ~new_new_n8630__;
  assign new_new_n8632__ = new_new_n8629__ & new_new_n8631__;
  assign new_new_n8633__ = ~new_new_n8629__ & ~new_new_n8631__;
  assign new_new_n8634__ = ~new_new_n8632__ & ~new_new_n8633__;
  assign new_new_n8635__ = new_new_n8150__ & ~new_new_n8187__;
  assign new_new_n8636__ = ~new_new_n8186__ & ~new_new_n8635__;
  assign new_new_n8637__ = ~new_new_n8144__ & ~new_new_n8147__;
  assign new_new_n8638__ = ~new_new_n8143__ & ~new_new_n8637__;
  assign new_new_n8639__ = ~new_new_n8294__ & ~new_new_n8299__;
  assign new_new_n8640__ = ~new_new_n8306__ & ~new_new_n8311__;
  assign new_new_n8641__ = ~new_new_n8312__ & ~new_new_n8640__;
  assign new_new_n8642__ = new_new_n8639__ & new_new_n8641__;
  assign new_new_n8643__ = ~new_new_n8639__ & ~new_new_n8641__;
  assign new_new_n8644__ = ~new_new_n8642__ & ~new_new_n8643__;
  assign new_new_n8645__ = new_new_n8638__ & ~new_new_n8644__;
  assign new_new_n8646__ = ~new_new_n8638__ & new_new_n8644__;
  assign new_new_n8647__ = ~new_new_n8645__ & ~new_new_n8646__;
  assign new_new_n8648__ = ~new_new_n8636__ & new_new_n8647__;
  assign new_new_n8649__ = new_new_n8636__ & ~new_new_n8647__;
  assign new_new_n8650__ = ~new_new_n8648__ & ~new_new_n8649__;
  assign new_new_n8651__ = ~new_new_n8288__ & ~new_new_n8301__;
  assign new_new_n8652__ = new_new_n8288__ & new_new_n8301__;
  assign new_new_n8653__ = ~new_new_n8316__ & ~new_new_n8652__;
  assign new_new_n8654__ = ~new_new_n8651__ & ~new_new_n8653__;
  assign new_new_n8655__ = new_new_n8650__ & ~new_new_n8654__;
  assign new_new_n8656__ = ~new_new_n8650__ & new_new_n8654__;
  assign new_new_n8657__ = ~new_new_n8655__ & ~new_new_n8656__;
  assign new_new_n8658__ = new_new_n8634__ & new_new_n8657__;
  assign new_new_n8659__ = ~new_new_n8634__ & ~new_new_n8657__;
  assign new_new_n8660__ = ~new_new_n8658__ & ~new_new_n8659__;
  assign new_new_n8661__ = new_new_n8628__ & ~new_new_n8660__;
  assign new_new_n8662__ = ~new_new_n8628__ & new_new_n8660__;
  assign new_new_n8663__ = ~new_new_n8661__ & ~new_new_n8662__;
  assign new_new_n8664__ = ~new_new_n8399__ & ~new_new_n8663__;
  assign new_new_n8665__ = ~new_new_n8411__ & new_new_n8664__;
  assign new_new_n8666__ = ~new_new_n8406__ & new_new_n8665__;
  assign new_new_n8667__ = ~new_new_n8409__ & new_new_n8666__;
  assign new_new_n8668__ = ~new_new_n8343__ & ~new_new_n8390__;
  assign new_new_n8669__ = ~new_new_n8344__ & ~new_new_n8668__;
  assign new_new_n8670__ = new_new_n8350__ & new_new_n8669__;
  assign new_new_n8671__ = new_new_n8343__ & new_new_n8390__;
  assign new_new_n8672__ = new_new_n8344__ & ~new_new_n8390__;
  assign new_new_n8673__ = ~new_new_n8671__ & ~new_new_n8672__;
  assign new_new_n8674__ = new_new_n8352__ & new_new_n8673__;
  assign new_new_n8675__ = new_new_n8351__ & ~new_new_n8669__;
  assign new_new_n8676__ = new_new_n8663__ & ~new_new_n8670__;
  assign new_new_n8677__ = ~new_new_n8675__ & new_new_n8676__;
  assign new_new_n8678__ = ~new_new_n8674__ & new_new_n8677__;
  assign po059 = ~new_new_n8667__ & ~new_new_n8678__;
  assign new_new_n8680__ = ~new_new_n8410__ & ~new_new_n8663__;
  assign new_new_n8681__ = ~new_new_n8390__ & ~new_new_n8680__;
  assign new_new_n8682__ = new_new_n8137__ & new_new_n8349__;
  assign new_new_n8683__ = new_new_n8663__ & ~new_new_n8682__;
  assign new_new_n8684__ = ~new_new_n8403__ & ~new_new_n8683__;
  assign new_new_n8685__ = ~new_new_n8681__ & new_new_n8684__;
  assign new_new_n8686__ = new_new_n8397__ & ~new_new_n8663__;
  assign new_new_n8687__ = ~new_new_n8390__ & ~new_new_n8682__;
  assign new_new_n8688__ = ~new_new_n8397__ & new_new_n8663__;
  assign new_new_n8689__ = ~new_new_n8410__ & ~new_new_n8688__;
  assign new_new_n8690__ = ~new_new_n8687__ & new_new_n8689__;
  assign new_new_n8691__ = ~new_new_n8686__ & ~new_new_n8690__;
  assign new_new_n8692__ = ~new_new_n8685__ & new_new_n8691__;
  assign new_new_n8693__ = ~new_new_n8482__ & ~new_new_n8622__;
  assign new_new_n8694__ = ~new_new_n8481__ & ~new_new_n8693__;
  assign new_new_n8695__ = pi29 & pi30;
  assign new_new_n8696__ = pi13 & pi46;
  assign new_new_n8697__ = pi17 & pi42;
  assign new_new_n8698__ = pi08 & pi51;
  assign new_new_n8699__ = pi16 & pi43;
  assign new_new_n8700__ = ~new_new_n8698__ & ~new_new_n8699__;
  assign new_new_n8701__ = new_new_n8698__ & new_new_n8699__;
  assign new_new_n8702__ = ~new_new_n8700__ & ~new_new_n8701__;
  assign new_new_n8703__ = new_new_n8697__ & ~new_new_n8702__;
  assign new_new_n8704__ = ~new_new_n8697__ & new_new_n8702__;
  assign new_new_n8705__ = ~new_new_n8703__ & ~new_new_n8704__;
  assign new_new_n8706__ = pi28 & pi31;
  assign new_new_n8707__ = pi14 & pi45;
  assign new_new_n8708__ = pi11 & pi48;
  assign new_new_n8709__ = pi12 & pi47;
  assign new_new_n8710__ = ~new_new_n8708__ & ~new_new_n8709__;
  assign new_new_n8711__ = new_new_n8708__ & new_new_n8709__;
  assign new_new_n8712__ = ~new_new_n8710__ & ~new_new_n8711__;
  assign new_new_n8713__ = new_new_n8707__ & ~new_new_n8712__;
  assign new_new_n8714__ = ~new_new_n8707__ & new_new_n8712__;
  assign new_new_n8715__ = ~new_new_n8713__ & ~new_new_n8714__;
  assign new_new_n8716__ = new_new_n8706__ & ~new_new_n8715__;
  assign new_new_n8717__ = ~new_new_n8706__ & new_new_n8715__;
  assign new_new_n8718__ = ~new_new_n8716__ & ~new_new_n8717__;
  assign new_new_n8719__ = new_new_n8705__ & new_new_n8718__;
  assign new_new_n8720__ = ~new_new_n8705__ & ~new_new_n8718__;
  assign new_new_n8721__ = ~new_new_n8719__ & ~new_new_n8720__;
  assign new_new_n8722__ = new_new_n8696__ & ~new_new_n8721__;
  assign new_new_n8723__ = ~new_new_n8696__ & new_new_n8721__;
  assign new_new_n8724__ = ~new_new_n8722__ & ~new_new_n8723__;
  assign new_new_n8725__ = new_new_n8695__ & new_new_n8724__;
  assign new_new_n8726__ = ~new_new_n8695__ & ~new_new_n8724__;
  assign new_new_n8727__ = ~new_new_n8725__ & ~new_new_n8726__;
  assign new_new_n8728__ = ~new_new_n8473__ & new_new_n8727__;
  assign new_new_n8729__ = new_new_n8473__ & ~new_new_n8727__;
  assign new_new_n8730__ = ~new_new_n8728__ & ~new_new_n8729__;
  assign new_new_n8731__ = pi19 & pi40;
  assign new_new_n8732__ = pi05 & pi54;
  assign new_new_n8733__ = pi04 & pi55;
  assign new_new_n8734__ = ~new_new_n8732__ & ~new_new_n8733__;
  assign new_new_n8735__ = new_new_n8732__ & new_new_n8733__;
  assign new_new_n8736__ = ~new_new_n8734__ & ~new_new_n8735__;
  assign new_new_n8737__ = new_new_n8731__ & ~new_new_n8736__;
  assign new_new_n8738__ = ~new_new_n8731__ & new_new_n8736__;
  assign new_new_n8739__ = ~new_new_n8737__ & ~new_new_n8738__;
  assign new_new_n8740__ = pi03 & pi56;
  assign new_new_n8741__ = pi30 & new_new_n2370__;
  assign new_new_n8742__ = ~pi02 & ~new_new_n8741__;
  assign new_new_n8743__ = pi57 & ~new_new_n8742__;
  assign new_new_n8744__ = pi30 & new_new_n7965__;
  assign new_new_n8745__ = new_new_n8743__ & ~new_new_n8744__;
  assign new_new_n8746__ = new_new_n8740__ & ~new_new_n8745__;
  assign new_new_n8747__ = ~new_new_n8740__ & new_new_n8745__;
  assign new_new_n8748__ = ~new_new_n8746__ & ~new_new_n8747__;
  assign new_new_n8749__ = new_new_n8739__ & new_new_n8748__;
  assign new_new_n8750__ = ~new_new_n8739__ & ~new_new_n8748__;
  assign new_new_n8751__ = ~new_new_n8749__ & ~new_new_n8750__;
  assign new_new_n8752__ = ~new_new_n8544__ & ~new_new_n8548__;
  assign new_new_n8753__ = ~new_new_n8547__ & ~new_new_n8752__;
  assign new_new_n8754__ = new_new_n8751__ & new_new_n8753__;
  assign new_new_n8755__ = ~new_new_n8751__ & ~new_new_n8753__;
  assign new_new_n8756__ = ~new_new_n8754__ & ~new_new_n8755__;
  assign new_new_n8757__ = new_new_n8730__ & ~new_new_n8756__;
  assign new_new_n8758__ = ~new_new_n8730__ & new_new_n8756__;
  assign new_new_n8759__ = ~new_new_n8757__ & ~new_new_n8758__;
  assign new_new_n8760__ = pi15 & pi44;
  assign new_new_n8761__ = pi10 & pi49;
  assign new_new_n8762__ = pi09 & pi50;
  assign new_new_n8763__ = ~new_new_n8761__ & ~new_new_n8762__;
  assign new_new_n8764__ = new_new_n8761__ & new_new_n8762__;
  assign new_new_n8765__ = ~new_new_n8763__ & ~new_new_n8764__;
  assign new_new_n8766__ = new_new_n8760__ & ~new_new_n8765__;
  assign new_new_n8767__ = ~new_new_n8760__ & new_new_n8765__;
  assign new_new_n8768__ = ~new_new_n8766__ & ~new_new_n8767__;
  assign new_new_n8769__ = ~new_new_n8456__ & ~new_new_n8458__;
  assign new_new_n8770__ = pi57 & ~new_new_n8457__;
  assign new_new_n8771__ = ~new_new_n8769__ & new_new_n8770__;
  assign new_new_n8772__ = ~pi57 & new_new_n8457__;
  assign new_new_n8773__ = ~new_new_n8456__ & ~new_new_n8772__;
  assign new_new_n8774__ = new_new_n8458__ & ~new_new_n8773__;
  assign new_new_n8775__ = ~new_new_n8771__ & ~new_new_n8774__;
  assign new_new_n8776__ = pi01 & ~new_new_n8775__;
  assign new_new_n8777__ = pi01 & pi57;
  assign new_new_n8778__ = new_new_n8457__ & ~new_new_n8777__;
  assign new_new_n8779__ = new_new_n8456__ & new_new_n8778__;
  assign new_new_n8780__ = ~new_new_n8776__ & ~new_new_n8779__;
  assign new_new_n8781__ = new_new_n8768__ & new_new_n8780__;
  assign new_new_n8782__ = ~new_new_n8768__ & ~new_new_n8780__;
  assign new_new_n8783__ = ~new_new_n8781__ & ~new_new_n8782__;
  assign new_new_n8784__ = pi18 & pi41;
  assign new_new_n8785__ = pi07 & pi52;
  assign new_new_n8786__ = pi06 & pi53;
  assign new_new_n8787__ = ~new_new_n8785__ & ~new_new_n8786__;
  assign new_new_n8788__ = new_new_n8785__ & new_new_n8786__;
  assign new_new_n8789__ = ~new_new_n8787__ & ~new_new_n8788__;
  assign new_new_n8790__ = new_new_n8784__ & ~new_new_n8789__;
  assign new_new_n8791__ = ~new_new_n8784__ & new_new_n8789__;
  assign new_new_n8792__ = ~new_new_n8790__ & ~new_new_n8791__;
  assign new_new_n8793__ = ~new_new_n8783__ & new_new_n8792__;
  assign new_new_n8794__ = new_new_n8783__ & ~new_new_n8792__;
  assign new_new_n8795__ = ~new_new_n8793__ & ~new_new_n8794__;
  assign new_new_n8796__ = new_new_n8759__ & ~new_new_n8795__;
  assign new_new_n8797__ = ~new_new_n8759__ & new_new_n8795__;
  assign new_new_n8798__ = ~new_new_n8796__ & ~new_new_n8797__;
  assign new_new_n8799__ = ~new_new_n8632__ & ~new_new_n8657__;
  assign new_new_n8800__ = ~new_new_n8633__ & ~new_new_n8799__;
  assign new_new_n8801__ = ~new_new_n8562__ & ~new_new_n8573__;
  assign new_new_n8802__ = ~new_new_n8563__ & ~new_new_n8801__;
  assign new_new_n8803__ = ~new_new_n8518__ & ~new_new_n8529__;
  assign new_new_n8804__ = ~new_new_n8519__ & ~new_new_n8803__;
  assign new_new_n8805__ = ~new_new_n8597__ & ~new_new_n8608__;
  assign new_new_n8806__ = ~new_new_n8598__ & ~new_new_n8805__;
  assign new_new_n8807__ = new_new_n8804__ & new_new_n8806__;
  assign new_new_n8808__ = ~new_new_n8804__ & ~new_new_n8806__;
  assign new_new_n8809__ = ~new_new_n8807__ & ~new_new_n8808__;
  assign new_new_n8810__ = new_new_n8802__ & new_new_n8809__;
  assign new_new_n8811__ = ~new_new_n8802__ & ~new_new_n8809__;
  assign new_new_n8812__ = ~new_new_n8810__ & ~new_new_n8811__;
  assign new_new_n8813__ = ~new_new_n8578__ & ~new_new_n8611__;
  assign new_new_n8814__ = ~new_new_n8577__ & ~new_new_n8813__;
  assign new_new_n8815__ = ~new_new_n8588__ & ~new_new_n8592__;
  assign new_new_n8816__ = ~new_new_n8591__ & ~new_new_n8815__;
  assign new_new_n8817__ = ~new_new_n8509__ & ~new_new_n8513__;
  assign new_new_n8818__ = ~new_new_n8512__ & ~new_new_n8817__;
  assign new_new_n8819__ = ~new_new_n8816__ & ~new_new_n8818__;
  assign new_new_n8820__ = new_new_n8816__ & new_new_n8818__;
  assign new_new_n8821__ = ~new_new_n8819__ & ~new_new_n8820__;
  assign new_new_n8822__ = ~new_new_n8600__ & ~new_new_n8604__;
  assign new_new_n8823__ = ~new_new_n8603__ & ~new_new_n8822__;
  assign new_new_n8824__ = ~new_new_n8821__ & new_new_n8823__;
  assign new_new_n8825__ = new_new_n8821__ & ~new_new_n8823__;
  assign new_new_n8826__ = ~new_new_n8824__ & ~new_new_n8825__;
  assign new_new_n8827__ = pi30 & pi58;
  assign new_new_n8828__ = pi01 & new_new_n8827__;
  assign new_new_n8829__ = pi01 & pi58;
  assign new_new_n8830__ = ~pi30 & ~new_new_n8829__;
  assign new_new_n8831__ = ~new_new_n8828__ & ~new_new_n8830__;
  assign new_new_n8832__ = ~new_new_n8500__ & ~new_new_n8504__;
  assign new_new_n8833__ = ~new_new_n8503__ & ~new_new_n8832__;
  assign new_new_n8834__ = ~new_new_n8521__ & ~new_new_n8525__;
  assign new_new_n8835__ = ~new_new_n8524__ & ~new_new_n8834__;
  assign new_new_n8836__ = new_new_n8833__ & new_new_n8835__;
  assign new_new_n8837__ = ~new_new_n8833__ & ~new_new_n8835__;
  assign new_new_n8838__ = ~new_new_n8836__ & ~new_new_n8837__;
  assign new_new_n8839__ = new_new_n8831__ & ~new_new_n8838__;
  assign new_new_n8840__ = ~new_new_n8831__ & new_new_n8838__;
  assign new_new_n8841__ = ~new_new_n8839__ & ~new_new_n8840__;
  assign new_new_n8842__ = new_new_n8826__ & new_new_n8841__;
  assign new_new_n8843__ = ~new_new_n8826__ & ~new_new_n8841__;
  assign new_new_n8844__ = ~new_new_n8842__ & ~new_new_n8843__;
  assign new_new_n8845__ = ~new_new_n8580__ & ~new_new_n8583__;
  assign new_new_n8846__ = ~new_new_n8582__ & ~new_new_n8845__;
  assign new_new_n8847__ = ~new_new_n8553__ & ~new_new_n8557__;
  assign new_new_n8848__ = ~new_new_n8556__ & ~new_new_n8847__;
  assign new_new_n8849__ = ~new_new_n8565__ & ~new_new_n8569__;
  assign new_new_n8850__ = ~new_new_n8568__ & ~new_new_n8849__;
  assign new_new_n8851__ = new_new_n8848__ & new_new_n8850__;
  assign new_new_n8852__ = ~new_new_n8848__ & ~new_new_n8850__;
  assign new_new_n8853__ = ~new_new_n8851__ & ~new_new_n8852__;
  assign new_new_n8854__ = new_new_n8846__ & ~new_new_n8853__;
  assign new_new_n8855__ = ~new_new_n8846__ & new_new_n8853__;
  assign new_new_n8856__ = ~new_new_n8854__ & ~new_new_n8855__;
  assign new_new_n8857__ = new_new_n8844__ & ~new_new_n8856__;
  assign new_new_n8858__ = ~new_new_n8844__ & new_new_n8856__;
  assign new_new_n8859__ = ~new_new_n8857__ & ~new_new_n8858__;
  assign new_new_n8860__ = ~new_new_n8814__ & ~new_new_n8859__;
  assign new_new_n8861__ = new_new_n8814__ & new_new_n8859__;
  assign new_new_n8862__ = ~new_new_n8860__ & ~new_new_n8861__;
  assign new_new_n8863__ = new_new_n8812__ & new_new_n8862__;
  assign new_new_n8864__ = ~new_new_n8812__ & ~new_new_n8862__;
  assign new_new_n8865__ = ~new_new_n8863__ & ~new_new_n8864__;
  assign new_new_n8866__ = ~new_new_n8800__ & new_new_n8865__;
  assign new_new_n8867__ = new_new_n8800__ & ~new_new_n8865__;
  assign new_new_n8868__ = ~new_new_n8866__ & ~new_new_n8867__;
  assign new_new_n8869__ = ~new_new_n8638__ & ~new_new_n8642__;
  assign new_new_n8870__ = ~new_new_n8643__ & ~new_new_n8869__;
  assign new_new_n8871__ = pi27 & pi32;
  assign new_new_n8872__ = pi26 & pi33;
  assign new_new_n8873__ = pi00 & pi59;
  assign new_new_n8874__ = ~new_new_n8872__ & ~new_new_n8873__;
  assign new_new_n8875__ = new_new_n8872__ & new_new_n8873__;
  assign new_new_n8876__ = ~new_new_n8874__ & ~new_new_n8875__;
  assign new_new_n8877__ = new_new_n8871__ & ~new_new_n8876__;
  assign new_new_n8878__ = ~new_new_n8871__ & new_new_n8876__;
  assign new_new_n8879__ = ~new_new_n8877__ & ~new_new_n8878__;
  assign new_new_n8880__ = pi25 & pi34;
  assign new_new_n8881__ = pi23 & pi36;
  assign new_new_n8882__ = pi24 & pi35;
  assign new_new_n8883__ = ~new_new_n8881__ & ~new_new_n8882__;
  assign new_new_n8884__ = new_new_n8881__ & new_new_n8882__;
  assign new_new_n8885__ = ~new_new_n8883__ & ~new_new_n8884__;
  assign new_new_n8886__ = new_new_n8880__ & ~new_new_n8885__;
  assign new_new_n8887__ = ~new_new_n8880__ & new_new_n8885__;
  assign new_new_n8888__ = ~new_new_n8886__ & ~new_new_n8887__;
  assign new_new_n8889__ = new_new_n8879__ & new_new_n8888__;
  assign new_new_n8890__ = ~new_new_n8879__ & ~new_new_n8888__;
  assign new_new_n8891__ = ~new_new_n8889__ & ~new_new_n8890__;
  assign new_new_n8892__ = pi22 & pi37;
  assign new_new_n8893__ = pi21 & pi38;
  assign new_new_n8894__ = ~new_new_n4298__ & ~new_new_n8893__;
  assign new_new_n8895__ = new_new_n4298__ & new_new_n8893__;
  assign new_new_n8896__ = ~new_new_n8894__ & ~new_new_n8895__;
  assign new_new_n8897__ = new_new_n8892__ & ~new_new_n8896__;
  assign new_new_n8898__ = ~new_new_n8892__ & new_new_n8896__;
  assign new_new_n8899__ = ~new_new_n8897__ & ~new_new_n8898__;
  assign new_new_n8900__ = new_new_n8891__ & ~new_new_n8899__;
  assign new_new_n8901__ = ~new_new_n8891__ & new_new_n8899__;
  assign new_new_n8902__ = ~new_new_n8900__ & ~new_new_n8901__;
  assign new_new_n8903__ = new_new_n8870__ & new_new_n8902__;
  assign new_new_n8904__ = ~new_new_n8870__ & ~new_new_n8902__;
  assign new_new_n8905__ = ~new_new_n8903__ & ~new_new_n8904__;
  assign new_new_n8906__ = ~new_new_n8648__ & ~new_new_n8654__;
  assign new_new_n8907__ = ~new_new_n8649__ & ~new_new_n8906__;
  assign new_new_n8908__ = new_new_n8905__ & ~new_new_n8907__;
  assign new_new_n8909__ = ~new_new_n8905__ & new_new_n8907__;
  assign new_new_n8910__ = ~new_new_n8908__ & ~new_new_n8909__;
  assign new_new_n8911__ = new_new_n8868__ & ~new_new_n8910__;
  assign new_new_n8912__ = ~new_new_n8868__ & new_new_n8910__;
  assign new_new_n8913__ = ~new_new_n8911__ & ~new_new_n8912__;
  assign new_new_n8914__ = new_new_n8798__ & new_new_n8913__;
  assign new_new_n8915__ = ~new_new_n8798__ & ~new_new_n8913__;
  assign new_new_n8916__ = ~new_new_n8914__ & ~new_new_n8915__;
  assign new_new_n8917__ = ~new_new_n8694__ & ~new_new_n8916__;
  assign new_new_n8918__ = new_new_n8694__ & new_new_n8916__;
  assign new_new_n8919__ = ~new_new_n8917__ & ~new_new_n8918__;
  assign new_new_n8920__ = ~new_new_n8615__ & ~new_new_n8620__;
  assign new_new_n8921__ = ~new_new_n8485__ & new_new_n8532__;
  assign new_new_n8922__ = new_new_n8485__ & ~new_new_n8532__;
  assign new_new_n8923__ = ~new_new_n8497__ & new_new_n8499__;
  assign new_new_n8924__ = new_new_n8497__ & ~new_new_n8499__;
  assign new_new_n8925__ = ~new_new_n8923__ & ~new_new_n8924__;
  assign new_new_n8926__ = ~new_new_n8922__ & ~new_new_n8925__;
  assign new_new_n8927__ = ~new_new_n8921__ & ~new_new_n8926__;
  assign new_new_n8928__ = ~new_new_n8424__ & ~new_new_n8433__;
  assign new_new_n8929__ = ~new_new_n8425__ & ~new_new_n8928__;
  assign new_new_n8930__ = ~new_new_n8495__ & new_new_n8499__;
  assign new_new_n8931__ = ~new_new_n8496__ & ~new_new_n8930__;
  assign new_new_n8932__ = new_new_n8929__ & ~new_new_n8931__;
  assign new_new_n8933__ = ~new_new_n8929__ & new_new_n8931__;
  assign new_new_n8934__ = ~new_new_n8932__ & ~new_new_n8933__;
  assign new_new_n8935__ = ~new_new_n8419__ & ~new_new_n8437__;
  assign new_new_n8936__ = new_new_n8419__ & new_new_n8437__;
  assign new_new_n8937__ = ~new_new_n8435__ & ~new_new_n8936__;
  assign new_new_n8938__ = ~new_new_n8935__ & ~new_new_n8937__;
  assign new_new_n8939__ = new_new_n8934__ & ~new_new_n8938__;
  assign new_new_n8940__ = ~new_new_n8934__ & new_new_n8938__;
  assign new_new_n8941__ = ~new_new_n8939__ & ~new_new_n8940__;
  assign new_new_n8942__ = ~new_new_n8927__ & ~new_new_n8941__;
  assign new_new_n8943__ = new_new_n8927__ & new_new_n8941__;
  assign new_new_n8944__ = ~new_new_n8942__ & ~new_new_n8943__;
  assign new_new_n8945__ = new_new_n8426__ & ~new_new_n8433__;
  assign new_new_n8946__ = ~new_new_n8426__ & new_new_n8433__;
  assign new_new_n8947__ = ~new_new_n8945__ & ~new_new_n8946__;
  assign new_new_n8948__ = new_new_n8431__ & new_new_n8947__;
  assign new_new_n8949__ = ~new_new_n8431__ & ~new_new_n8947__;
  assign new_new_n8950__ = new_new_n8419__ & new_new_n8440__;
  assign new_new_n8951__ = ~new_new_n8419__ & ~new_new_n8440__;
  assign new_new_n8952__ = ~new_new_n8950__ & ~new_new_n8951__;
  assign new_new_n8953__ = ~new_new_n8949__ & new_new_n8952__;
  assign new_new_n8954__ = ~new_new_n8948__ & ~new_new_n8953__;
  assign new_new_n8955__ = ~new_new_n8944__ & new_new_n8954__;
  assign new_new_n8956__ = new_new_n8944__ & ~new_new_n8954__;
  assign new_new_n8957__ = ~new_new_n8955__ & ~new_new_n8956__;
  assign new_new_n8958__ = ~new_new_n8920__ & new_new_n8957__;
  assign new_new_n8959__ = new_new_n8920__ & ~new_new_n8957__;
  assign new_new_n8960__ = ~new_new_n8958__ & ~new_new_n8959__;
  assign new_new_n8961__ = ~new_new_n8451__ & ~new_new_n8477__;
  assign new_new_n8962__ = ~new_new_n8450__ & ~new_new_n8961__;
  assign new_new_n8963__ = new_new_n8960__ & ~new_new_n8962__;
  assign new_new_n8964__ = ~new_new_n8960__ & new_new_n8962__;
  assign new_new_n8965__ = ~new_new_n8963__ & ~new_new_n8964__;
  assign new_new_n8966__ = new_new_n8919__ & ~new_new_n8965__;
  assign new_new_n8967__ = ~new_new_n8919__ & new_new_n8965__;
  assign new_new_n8968__ = ~new_new_n8966__ & ~new_new_n8967__;
  assign new_new_n8969__ = new_new_n8692__ & new_new_n8968__;
  assign new_new_n8970__ = ~new_new_n8692__ & ~new_new_n8968__;
  assign new_new_n8971__ = ~new_new_n8969__ & ~new_new_n8970__;
  assign new_new_n8972__ = ~new_new_n8627__ & new_new_n8660__;
  assign new_new_n8973__ = ~new_new_n8626__ & ~new_new_n8972__;
  assign new_new_n8974__ = new_new_n8971__ & new_new_n8973__;
  assign new_new_n8975__ = ~new_new_n8971__ & ~new_new_n8973__;
  assign po060 = new_new_n8974__ | new_new_n8975__;
  assign new_new_n8977__ = ~new_new_n8958__ & ~new_new_n8962__;
  assign new_new_n8978__ = ~new_new_n8959__ & ~new_new_n8977__;
  assign new_new_n8979__ = ~new_new_n8781__ & ~new_new_n8792__;
  assign new_new_n8980__ = ~new_new_n8782__ & ~new_new_n8979__;
  assign new_new_n8981__ = ~new_new_n8740__ & ~new_new_n8744__;
  assign new_new_n8982__ = new_new_n8743__ & ~new_new_n8981__;
  assign new_new_n8983__ = ~new_new_n8871__ & ~new_new_n8875__;
  assign new_new_n8984__ = ~new_new_n8874__ & ~new_new_n8983__;
  assign new_new_n8985__ = ~new_new_n8760__ & ~new_new_n8764__;
  assign new_new_n8986__ = ~new_new_n8763__ & ~new_new_n8985__;
  assign new_new_n8987__ = new_new_n8984__ & ~new_new_n8986__;
  assign new_new_n8988__ = ~new_new_n8984__ & new_new_n8986__;
  assign new_new_n8989__ = ~new_new_n8987__ & ~new_new_n8988__;
  assign new_new_n8990__ = new_new_n8982__ & new_new_n8989__;
  assign new_new_n8991__ = ~new_new_n8982__ & ~new_new_n8989__;
  assign new_new_n8992__ = ~new_new_n8990__ & ~new_new_n8991__;
  assign new_new_n8993__ = new_new_n8980__ & ~new_new_n8992__;
  assign new_new_n8994__ = ~new_new_n8980__ & new_new_n8992__;
  assign new_new_n8995__ = ~new_new_n8993__ & ~new_new_n8994__;
  assign new_new_n8996__ = ~new_new_n8892__ & ~new_new_n8895__;
  assign new_new_n8997__ = ~new_new_n8894__ & ~new_new_n8996__;
  assign new_new_n8998__ = ~new_new_n8731__ & ~new_new_n8735__;
  assign new_new_n8999__ = ~new_new_n8734__ & ~new_new_n8998__;
  assign new_new_n9000__ = ~new_new_n8880__ & ~new_new_n8884__;
  assign new_new_n9001__ = ~new_new_n8883__ & ~new_new_n9000__;
  assign new_new_n9002__ = new_new_n8999__ & new_new_n9001__;
  assign new_new_n9003__ = ~new_new_n8999__ & ~new_new_n9001__;
  assign new_new_n9004__ = ~new_new_n9002__ & ~new_new_n9003__;
  assign new_new_n9005__ = new_new_n8997__ & ~new_new_n9004__;
  assign new_new_n9006__ = ~new_new_n8997__ & new_new_n9004__;
  assign new_new_n9007__ = ~new_new_n9005__ & ~new_new_n9006__;
  assign new_new_n9008__ = ~new_new_n8728__ & ~new_new_n8756__;
  assign new_new_n9009__ = ~new_new_n8729__ & ~new_new_n9008__;
  assign new_new_n9010__ = new_new_n9007__ & ~new_new_n9009__;
  assign new_new_n9011__ = ~new_new_n9007__ & new_new_n9009__;
  assign new_new_n9012__ = ~new_new_n9010__ & ~new_new_n9011__;
  assign new_new_n9013__ = new_new_n8995__ & new_new_n9012__;
  assign new_new_n9014__ = ~new_new_n8995__ & ~new_new_n9012__;
  assign new_new_n9015__ = ~new_new_n9013__ & ~new_new_n9014__;
  assign new_new_n9016__ = new_new_n8978__ & ~new_new_n9015__;
  assign new_new_n9017__ = ~new_new_n8978__ & new_new_n9015__;
  assign new_new_n9018__ = ~new_new_n9016__ & ~new_new_n9017__;
  assign new_new_n9019__ = ~new_new_n8933__ & new_new_n8938__;
  assign new_new_n9020__ = ~new_new_n8932__ & ~new_new_n9019__;
  assign new_new_n9021__ = ~new_new_n8707__ & ~new_new_n8711__;
  assign new_new_n9022__ = ~new_new_n8710__ & ~new_new_n9021__;
  assign new_new_n9023__ = pi15 & pi45;
  assign new_new_n9024__ = pi10 & pi50;
  assign new_new_n9025__ = pi11 & pi49;
  assign new_new_n9026__ = ~new_new_n9024__ & ~new_new_n9025__;
  assign new_new_n9027__ = new_new_n9024__ & new_new_n9025__;
  assign new_new_n9028__ = ~new_new_n9026__ & ~new_new_n9027__;
  assign new_new_n9029__ = new_new_n9023__ & ~new_new_n9028__;
  assign new_new_n9030__ = ~new_new_n9023__ & new_new_n9028__;
  assign new_new_n9031__ = ~new_new_n9029__ & ~new_new_n9030__;
  assign new_new_n9032__ = ~new_new_n9022__ & new_new_n9031__;
  assign new_new_n9033__ = new_new_n9022__ & ~new_new_n9031__;
  assign new_new_n9034__ = ~new_new_n9032__ & ~new_new_n9033__;
  assign new_new_n9035__ = pi17 & pi43;
  assign new_new_n9036__ = pi16 & pi44;
  assign new_new_n9037__ = pi09 & pi51;
  assign new_new_n9038__ = ~new_new_n9036__ & ~new_new_n9037__;
  assign new_new_n9039__ = new_new_n9036__ & new_new_n9037__;
  assign new_new_n9040__ = ~new_new_n9038__ & ~new_new_n9039__;
  assign new_new_n9041__ = new_new_n9035__ & ~new_new_n9040__;
  assign new_new_n9042__ = ~new_new_n9035__ & new_new_n9040__;
  assign new_new_n9043__ = ~new_new_n9041__ & ~new_new_n9042__;
  assign new_new_n9044__ = ~new_new_n9034__ & new_new_n9043__;
  assign new_new_n9045__ = new_new_n9034__ & ~new_new_n9043__;
  assign new_new_n9046__ = ~new_new_n9044__ & ~new_new_n9045__;
  assign new_new_n9047__ = ~new_new_n9020__ & new_new_n9046__;
  assign new_new_n9048__ = new_new_n9020__ & ~new_new_n9046__;
  assign new_new_n9049__ = ~new_new_n9047__ & ~new_new_n9048__;
  assign new_new_n9050__ = pi22 & pi38;
  assign new_new_n9051__ = pi21 & pi39;
  assign new_new_n9052__ = pi20 & pi40;
  assign new_new_n9053__ = ~new_new_n9051__ & ~new_new_n9052__;
  assign new_new_n9054__ = new_new_n9051__ & new_new_n9052__;
  assign new_new_n9055__ = ~new_new_n9053__ & ~new_new_n9054__;
  assign new_new_n9056__ = new_new_n9050__ & ~new_new_n9055__;
  assign new_new_n9057__ = ~new_new_n9050__ & new_new_n9055__;
  assign new_new_n9058__ = ~new_new_n9056__ & ~new_new_n9057__;
  assign new_new_n9059__ = pi26 & pi34;
  assign new_new_n9060__ = pi24 & pi36;
  assign new_new_n9061__ = pi25 & pi35;
  assign new_new_n9062__ = ~new_new_n9060__ & ~new_new_n9061__;
  assign new_new_n9063__ = new_new_n9060__ & new_new_n9061__;
  assign new_new_n9064__ = ~new_new_n9062__ & ~new_new_n9063__;
  assign new_new_n9065__ = new_new_n9059__ & ~new_new_n9064__;
  assign new_new_n9066__ = ~new_new_n9059__ & new_new_n9064__;
  assign new_new_n9067__ = ~new_new_n9065__ & ~new_new_n9066__;
  assign new_new_n9068__ = ~new_new_n9058__ & ~new_new_n9067__;
  assign new_new_n9069__ = new_new_n9058__ & new_new_n9067__;
  assign new_new_n9070__ = ~new_new_n9068__ & ~new_new_n9069__;
  assign new_new_n9071__ = pi04 & pi56;
  assign new_new_n9072__ = pi02 & pi58;
  assign new_new_n9073__ = pi03 & pi57;
  assign new_new_n9074__ = ~new_new_n9072__ & ~new_new_n9073__;
  assign new_new_n9075__ = new_new_n9072__ & new_new_n9073__;
  assign new_new_n9076__ = ~new_new_n9074__ & ~new_new_n9075__;
  assign new_new_n9077__ = new_new_n9071__ & ~new_new_n9076__;
  assign new_new_n9078__ = ~new_new_n9071__ & new_new_n9076__;
  assign new_new_n9079__ = ~new_new_n9077__ & ~new_new_n9078__;
  assign new_new_n9080__ = ~new_new_n9070__ & new_new_n9079__;
  assign new_new_n9081__ = new_new_n9070__ & ~new_new_n9079__;
  assign new_new_n9082__ = ~new_new_n9080__ & ~new_new_n9081__;
  assign new_new_n9083__ = new_new_n9049__ & ~new_new_n9082__;
  assign new_new_n9084__ = ~new_new_n9049__ & new_new_n9082__;
  assign new_new_n9085__ = ~new_new_n9083__ & ~new_new_n9084__;
  assign new_new_n9086__ = ~new_new_n8843__ & new_new_n8856__;
  assign new_new_n9087__ = ~new_new_n8842__ & ~new_new_n9086__;
  assign new_new_n9088__ = pi19 & pi41;
  assign new_new_n9089__ = pi05 & pi55;
  assign new_new_n9090__ = pi06 & pi54;
  assign new_new_n9091__ = ~new_new_n9089__ & ~new_new_n9090__;
  assign new_new_n9092__ = new_new_n9089__ & new_new_n9090__;
  assign new_new_n9093__ = ~new_new_n9091__ & ~new_new_n9092__;
  assign new_new_n9094__ = new_new_n9088__ & ~new_new_n9093__;
  assign new_new_n9095__ = ~new_new_n9088__ & new_new_n9093__;
  assign new_new_n9096__ = ~new_new_n9094__ & ~new_new_n9095__;
  assign new_new_n9097__ = pi18 & pi42;
  assign new_new_n9098__ = pi07 & pi53;
  assign new_new_n9099__ = pi08 & pi52;
  assign new_new_n9100__ = ~new_new_n9098__ & ~new_new_n9099__;
  assign new_new_n9101__ = new_new_n9098__ & new_new_n9099__;
  assign new_new_n9102__ = ~new_new_n9100__ & ~new_new_n9101__;
  assign new_new_n9103__ = new_new_n9097__ & ~new_new_n9102__;
  assign new_new_n9104__ = ~new_new_n9097__ & new_new_n9102__;
  assign new_new_n9105__ = ~new_new_n9103__ & ~new_new_n9104__;
  assign new_new_n9106__ = new_new_n9096__ & new_new_n9105__;
  assign new_new_n9107__ = ~new_new_n9096__ & ~new_new_n9105__;
  assign new_new_n9108__ = ~new_new_n9106__ & ~new_new_n9107__;
  assign new_new_n9109__ = pi14 & pi46;
  assign new_new_n9110__ = pi12 & pi48;
  assign new_new_n9111__ = pi13 & pi47;
  assign new_new_n9112__ = ~new_new_n9110__ & ~new_new_n9111__;
  assign new_new_n9113__ = new_new_n9110__ & new_new_n9111__;
  assign new_new_n9114__ = ~new_new_n9112__ & ~new_new_n9113__;
  assign new_new_n9115__ = new_new_n9109__ & ~new_new_n9114__;
  assign new_new_n9116__ = ~new_new_n9109__ & new_new_n9114__;
  assign new_new_n9117__ = ~new_new_n9115__ & ~new_new_n9116__;
  assign new_new_n9118__ = ~new_new_n9108__ & new_new_n9117__;
  assign new_new_n9119__ = new_new_n9108__ & ~new_new_n9117__;
  assign new_new_n9120__ = ~new_new_n9118__ & ~new_new_n9119__;
  assign new_new_n9121__ = ~new_new_n9087__ & ~new_new_n9120__;
  assign new_new_n9122__ = new_new_n9087__ & new_new_n9120__;
  assign new_new_n9123__ = ~new_new_n9121__ & ~new_new_n9122__;
  assign new_new_n9124__ = ~new_new_n8831__ & ~new_new_n8836__;
  assign new_new_n9125__ = ~new_new_n8837__ & ~new_new_n9124__;
  assign new_new_n9126__ = pi00 & pi60;
  assign new_new_n9127__ = pi29 & pi31;
  assign new_new_n9128__ = pi01 & pi59;
  assign new_new_n9129__ = ~new_new_n9127__ & new_new_n9128__;
  assign new_new_n9130__ = new_new_n9127__ & ~new_new_n9128__;
  assign new_new_n9131__ = ~new_new_n9129__ & ~new_new_n9130__;
  assign new_new_n9132__ = ~new_new_n9126__ & new_new_n9131__;
  assign new_new_n9133__ = new_new_n9126__ & ~new_new_n9131__;
  assign new_new_n9134__ = ~new_new_n9132__ & ~new_new_n9133__;
  assign new_new_n9135__ = new_new_n8828__ & new_new_n9134__;
  assign new_new_n9136__ = ~new_new_n8828__ & ~new_new_n9134__;
  assign new_new_n9137__ = ~new_new_n9135__ & ~new_new_n9136__;
  assign new_new_n9138__ = ~new_new_n9125__ & ~new_new_n9137__;
  assign new_new_n9139__ = new_new_n9125__ & new_new_n9137__;
  assign new_new_n9140__ = ~new_new_n9138__ & ~new_new_n9139__;
  assign new_new_n9141__ = pi28 & pi32;
  assign new_new_n9142__ = pi27 & pi33;
  assign new_new_n9143__ = pi23 & pi37;
  assign new_new_n9144__ = ~new_new_n9142__ & ~new_new_n9143__;
  assign new_new_n9145__ = new_new_n9142__ & new_new_n9143__;
  assign new_new_n9146__ = ~new_new_n9144__ & ~new_new_n9145__;
  assign new_new_n9147__ = new_new_n9141__ & ~new_new_n9146__;
  assign new_new_n9148__ = ~new_new_n9141__ & new_new_n9146__;
  assign new_new_n9149__ = ~new_new_n9147__ & ~new_new_n9148__;
  assign new_new_n9150__ = new_new_n9140__ & ~new_new_n9149__;
  assign new_new_n9151__ = ~new_new_n9140__ & new_new_n9149__;
  assign new_new_n9152__ = ~new_new_n9150__ & ~new_new_n9151__;
  assign new_new_n9153__ = new_new_n9123__ & new_new_n9152__;
  assign new_new_n9154__ = ~new_new_n9123__ & ~new_new_n9152__;
  assign new_new_n9155__ = ~new_new_n9153__ & ~new_new_n9154__;
  assign new_new_n9156__ = new_new_n9085__ & ~new_new_n9155__;
  assign new_new_n9157__ = ~new_new_n9085__ & new_new_n9155__;
  assign new_new_n9158__ = ~new_new_n9156__ & ~new_new_n9157__;
  assign new_new_n9159__ = ~new_new_n8943__ & new_new_n8954__;
  assign new_new_n9160__ = ~new_new_n8942__ & ~new_new_n9159__;
  assign new_new_n9161__ = new_new_n9158__ & new_new_n9160__;
  assign new_new_n9162__ = ~new_new_n9158__ & ~new_new_n9160__;
  assign new_new_n9163__ = ~new_new_n9161__ & ~new_new_n9162__;
  assign new_new_n9164__ = ~new_new_n8889__ & ~new_new_n8899__;
  assign new_new_n9165__ = ~new_new_n8890__ & ~new_new_n9164__;
  assign new_new_n9166__ = ~new_new_n8697__ & ~new_new_n8701__;
  assign new_new_n9167__ = ~new_new_n8700__ & ~new_new_n9166__;
  assign new_new_n9168__ = ~new_new_n8784__ & ~new_new_n8788__;
  assign new_new_n9169__ = ~new_new_n8787__ & ~new_new_n9168__;
  assign new_new_n9170__ = ~new_new_n9167__ & ~new_new_n9169__;
  assign new_new_n9171__ = new_new_n9167__ & new_new_n9169__;
  assign new_new_n9172__ = ~new_new_n9170__ & ~new_new_n9171__;
  assign new_new_n9173__ = ~new_new_n8695__ & ~new_new_n8706__;
  assign new_new_n9174__ = new_new_n8695__ & new_new_n8706__;
  assign new_new_n9175__ = ~new_new_n8696__ & ~new_new_n9174__;
  assign new_new_n9176__ = ~new_new_n9173__ & ~new_new_n9175__;
  assign new_new_n9177__ = ~new_new_n9172__ & new_new_n9176__;
  assign new_new_n9178__ = new_new_n9172__ & ~new_new_n9176__;
  assign new_new_n9179__ = ~new_new_n9177__ & ~new_new_n9178__;
  assign new_new_n9180__ = new_new_n8705__ & new_new_n8715__;
  assign new_new_n9181__ = ~new_new_n8705__ & ~new_new_n8715__;
  assign new_new_n9182__ = ~new_new_n9173__ & ~new_new_n9174__;
  assign new_new_n9183__ = new_new_n8696__ & ~new_new_n9182__;
  assign new_new_n9184__ = ~new_new_n8696__ & new_new_n9182__;
  assign new_new_n9185__ = ~new_new_n9183__ & ~new_new_n9184__;
  assign new_new_n9186__ = ~new_new_n9181__ & new_new_n9185__;
  assign new_new_n9187__ = ~new_new_n9180__ & ~new_new_n9186__;
  assign new_new_n9188__ = ~new_new_n9179__ & new_new_n9187__;
  assign new_new_n9189__ = new_new_n9179__ & ~new_new_n9187__;
  assign new_new_n9190__ = ~new_new_n9188__ & ~new_new_n9189__;
  assign new_new_n9191__ = new_new_n9165__ & new_new_n9190__;
  assign new_new_n9192__ = ~new_new_n9165__ & ~new_new_n9190__;
  assign new_new_n9193__ = ~new_new_n9191__ & ~new_new_n9192__;
  assign new_new_n9194__ = new_new_n9163__ & ~new_new_n9193__;
  assign new_new_n9195__ = ~new_new_n9163__ & new_new_n9193__;
  assign new_new_n9196__ = ~new_new_n9194__ & ~new_new_n9195__;
  assign new_new_n9197__ = new_new_n9018__ & new_new_n9196__;
  assign new_new_n9198__ = ~new_new_n9018__ & ~new_new_n9196__;
  assign new_new_n9199__ = ~new_new_n9197__ & ~new_new_n9198__;
  assign new_new_n9200__ = new_new_n8759__ & new_new_n8907__;
  assign new_new_n9201__ = ~new_new_n8759__ & ~new_new_n8907__;
  assign new_new_n9202__ = ~new_new_n9200__ & ~new_new_n9201__;
  assign new_new_n9203__ = ~new_new_n8795__ & new_new_n8905__;
  assign new_new_n9204__ = new_new_n8795__ & ~new_new_n8905__;
  assign new_new_n9205__ = ~new_new_n9203__ & ~new_new_n9204__;
  assign new_new_n9206__ = ~new_new_n9202__ & ~new_new_n9205__;
  assign new_new_n9207__ = new_new_n9202__ & new_new_n9205__;
  assign new_new_n9208__ = ~new_new_n9206__ & ~new_new_n9207__;
  assign new_new_n9209__ = ~new_new_n8867__ & new_new_n9208__;
  assign new_new_n9210__ = ~new_new_n8866__ & ~new_new_n9209__;
  assign new_new_n9211__ = ~new_new_n9199__ & ~new_new_n9210__;
  assign new_new_n9212__ = new_new_n9199__ & new_new_n9210__;
  assign new_new_n9213__ = ~new_new_n9211__ & ~new_new_n9212__;
  assign new_new_n9214__ = ~new_new_n8918__ & new_new_n8965__;
  assign new_new_n9215__ = ~new_new_n8917__ & ~new_new_n9214__;
  assign new_new_n9216__ = ~new_new_n8969__ & ~new_new_n8973__;
  assign new_new_n9217__ = ~new_new_n8970__ & ~new_new_n9216__;
  assign new_new_n9218__ = ~new_new_n9215__ & ~new_new_n9217__;
  assign new_new_n9219__ = new_new_n9215__ & new_new_n9217__;
  assign new_new_n9220__ = ~new_new_n9218__ & ~new_new_n9219__;
  assign new_new_n9221__ = new_new_n9213__ & ~new_new_n9220__;
  assign new_new_n9222__ = ~new_new_n9213__ & new_new_n9220__;
  assign new_new_n9223__ = ~new_new_n9221__ & ~new_new_n9222__;
  assign new_new_n9224__ = new_new_n8812__ & ~new_new_n8861__;
  assign new_new_n9225__ = ~new_new_n8860__ & ~new_new_n9224__;
  assign new_new_n9226__ = ~new_new_n8807__ & ~new_new_n8810__;
  assign new_new_n9227__ = ~new_new_n8749__ & new_new_n8753__;
  assign new_new_n9228__ = ~new_new_n8750__ & ~new_new_n9227__;
  assign new_new_n9229__ = ~new_new_n8846__ & ~new_new_n8851__;
  assign new_new_n9230__ = ~new_new_n8852__ & ~new_new_n9229__;
  assign new_new_n9231__ = ~new_new_n8820__ & ~new_new_n8823__;
  assign new_new_n9232__ = ~new_new_n8819__ & ~new_new_n9231__;
  assign new_new_n9233__ = new_new_n9230__ & new_new_n9232__;
  assign new_new_n9234__ = ~new_new_n9230__ & ~new_new_n9232__;
  assign new_new_n9235__ = ~new_new_n9233__ & ~new_new_n9234__;
  assign new_new_n9236__ = new_new_n9228__ & ~new_new_n9235__;
  assign new_new_n9237__ = ~new_new_n9228__ & new_new_n9235__;
  assign new_new_n9238__ = ~new_new_n9236__ & ~new_new_n9237__;
  assign new_new_n9239__ = ~new_new_n9226__ & ~new_new_n9238__;
  assign new_new_n9240__ = new_new_n9226__ & new_new_n9238__;
  assign new_new_n9241__ = ~new_new_n9239__ & ~new_new_n9240__;
  assign new_new_n9242__ = new_new_n8795__ & ~new_new_n8904__;
  assign new_new_n9243__ = ~new_new_n8903__ & ~new_new_n9242__;
  assign new_new_n9244__ = new_new_n9241__ & ~new_new_n9243__;
  assign new_new_n9245__ = ~new_new_n9241__ & new_new_n9243__;
  assign new_new_n9246__ = ~new_new_n9244__ & ~new_new_n9245__;
  assign new_new_n9247__ = new_new_n9225__ & new_new_n9246__;
  assign new_new_n9248__ = ~new_new_n9225__ & ~new_new_n9246__;
  assign new_new_n9249__ = ~new_new_n9247__ & ~new_new_n9248__;
  assign new_new_n9250__ = ~new_new_n9200__ & ~new_new_n9205__;
  assign new_new_n9251__ = ~new_new_n9201__ & ~new_new_n9250__;
  assign new_new_n9252__ = new_new_n9249__ & ~new_new_n9251__;
  assign new_new_n9253__ = ~new_new_n9249__ & new_new_n9251__;
  assign new_new_n9254__ = ~new_new_n9252__ & ~new_new_n9253__;
  assign new_new_n9255__ = new_new_n9223__ & new_new_n9254__;
  assign new_new_n9256__ = ~new_new_n9223__ & ~new_new_n9254__;
  assign po061 = new_new_n9255__ | new_new_n9256__;
  assign new_new_n9258__ = pi19 & pi42;
  assign new_new_n9259__ = pi08 & pi53;
  assign new_new_n9260__ = pi07 & pi54;
  assign new_new_n9261__ = ~new_new_n9259__ & ~new_new_n9260__;
  assign new_new_n9262__ = new_new_n9259__ & new_new_n9260__;
  assign new_new_n9263__ = ~new_new_n9261__ & ~new_new_n9262__;
  assign new_new_n9264__ = new_new_n9258__ & ~new_new_n9263__;
  assign new_new_n9265__ = ~new_new_n9258__ & new_new_n9263__;
  assign new_new_n9266__ = ~new_new_n9264__ & ~new_new_n9265__;
  assign new_new_n9267__ = pi18 & pi43;
  assign new_new_n9268__ = pi17 & pi44;
  assign new_new_n9269__ = pi09 & pi52;
  assign new_new_n9270__ = ~new_new_n9268__ & ~new_new_n9269__;
  assign new_new_n9271__ = new_new_n9268__ & new_new_n9269__;
  assign new_new_n9272__ = ~new_new_n9270__ & ~new_new_n9271__;
  assign new_new_n9273__ = new_new_n9267__ & ~new_new_n9272__;
  assign new_new_n9274__ = ~new_new_n9267__ & new_new_n9272__;
  assign new_new_n9275__ = ~new_new_n9273__ & ~new_new_n9274__;
  assign new_new_n9276__ = new_new_n9266__ & new_new_n9275__;
  assign new_new_n9277__ = ~new_new_n9266__ & ~new_new_n9275__;
  assign new_new_n9278__ = ~new_new_n9276__ & ~new_new_n9277__;
  assign new_new_n9279__ = pi28 & pi33;
  assign new_new_n9280__ = pi27 & pi34;
  assign new_new_n9281__ = pi26 & pi35;
  assign new_new_n9282__ = ~new_new_n9280__ & ~new_new_n9281__;
  assign new_new_n9283__ = new_new_n9280__ & new_new_n9281__;
  assign new_new_n9284__ = ~new_new_n9282__ & ~new_new_n9283__;
  assign new_new_n9285__ = new_new_n9279__ & ~new_new_n9284__;
  assign new_new_n9286__ = ~new_new_n9279__ & new_new_n9284__;
  assign new_new_n9287__ = ~new_new_n9285__ & ~new_new_n9286__;
  assign new_new_n9288__ = ~new_new_n9278__ & new_new_n9287__;
  assign new_new_n9289__ = new_new_n9278__ & ~new_new_n9287__;
  assign new_new_n9290__ = ~new_new_n9288__ & ~new_new_n9289__;
  assign new_new_n9291__ = ~new_new_n8980__ & ~new_new_n9007__;
  assign new_new_n9292__ = new_new_n8980__ & new_new_n9007__;
  assign new_new_n9293__ = ~new_new_n8992__ & ~new_new_n9292__;
  assign new_new_n9294__ = ~new_new_n9291__ & ~new_new_n9293__;
  assign new_new_n9295__ = ~new_new_n9290__ & new_new_n9294__;
  assign new_new_n9296__ = new_new_n9290__ & ~new_new_n9294__;
  assign new_new_n9297__ = ~new_new_n9295__ & ~new_new_n9296__;
  assign new_new_n9298__ = new_new_n9165__ & ~new_new_n9188__;
  assign new_new_n9299__ = ~new_new_n9189__ & ~new_new_n9298__;
  assign new_new_n9300__ = new_new_n9297__ & ~new_new_n9299__;
  assign new_new_n9301__ = ~new_new_n9297__ & new_new_n9299__;
  assign new_new_n9302__ = ~new_new_n9300__ & ~new_new_n9301__;
  assign new_new_n9303__ = ~new_new_n9156__ & ~new_new_n9160__;
  assign new_new_n9304__ = ~new_new_n9157__ & ~new_new_n9303__;
  assign new_new_n9305__ = ~new_new_n9302__ & ~new_new_n9304__;
  assign new_new_n9306__ = new_new_n9302__ & new_new_n9304__;
  assign new_new_n9307__ = ~new_new_n9305__ & ~new_new_n9306__;
  assign new_new_n9308__ = ~new_new_n9171__ & ~new_new_n9176__;
  assign new_new_n9309__ = ~new_new_n9170__ & ~new_new_n9308__;
  assign new_new_n9310__ = pi23 & pi38;
  assign new_new_n9311__ = pi04 & pi57;
  assign new_new_n9312__ = pi03 & pi58;
  assign new_new_n9313__ = ~new_new_n9311__ & ~new_new_n9312__;
  assign new_new_n9314__ = new_new_n9311__ & new_new_n9312__;
  assign new_new_n9315__ = ~new_new_n9313__ & ~new_new_n9314__;
  assign new_new_n9316__ = new_new_n9310__ & ~new_new_n9315__;
  assign new_new_n9317__ = ~new_new_n9310__ & new_new_n9315__;
  assign new_new_n9318__ = ~new_new_n9316__ & ~new_new_n9317__;
  assign new_new_n9319__ = ~new_new_n9309__ & new_new_n9318__;
  assign new_new_n9320__ = new_new_n9309__ & ~new_new_n9318__;
  assign new_new_n9321__ = ~new_new_n9319__ & ~new_new_n9320__;
  assign new_new_n9322__ = ~new_new_n8982__ & ~new_new_n8984__;
  assign new_new_n9323__ = new_new_n8982__ & new_new_n8984__;
  assign new_new_n9324__ = ~new_new_n8986__ & ~new_new_n9323__;
  assign new_new_n9325__ = ~new_new_n9322__ & ~new_new_n9324__;
  assign new_new_n9326__ = ~new_new_n9321__ & new_new_n9325__;
  assign new_new_n9327__ = new_new_n9321__ & ~new_new_n9325__;
  assign new_new_n9328__ = ~new_new_n9326__ & ~new_new_n9327__;
  assign new_new_n9329__ = ~new_new_n9048__ & new_new_n9082__;
  assign new_new_n9330__ = ~new_new_n9047__ & ~new_new_n9329__;
  assign new_new_n9331__ = ~new_new_n8997__ & ~new_new_n9002__;
  assign new_new_n9332__ = ~new_new_n9003__ & ~new_new_n9331__;
  assign new_new_n9333__ = pi29 & pi59;
  assign new_new_n9334__ = ~new_new_n9109__ & ~new_new_n9113__;
  assign new_new_n9335__ = ~new_new_n9112__ & ~new_new_n9334__;
  assign new_new_n9336__ = pi01 & ~pi60;
  assign new_new_n9337__ = ~new_new_n9335__ & ~new_new_n9336__;
  assign new_new_n9338__ = new_new_n9333__ & ~new_new_n9337__;
  assign new_new_n9339__ = pi31 & pi60;
  assign new_new_n9340__ = new_new_n9335__ & ~new_new_n9339__;
  assign new_new_n9341__ = new_new_n9338__ & ~new_new_n9340__;
  assign new_new_n9342__ = new_new_n9127__ & new_new_n9128__;
  assign new_new_n9343__ = pi01 & pi60;
  assign new_new_n9344__ = new_new_n9335__ & ~new_new_n9343__;
  assign new_new_n9345__ = ~new_new_n9335__ & new_new_n9343__;
  assign new_new_n9346__ = ~new_new_n9344__ & ~new_new_n9345__;
  assign new_new_n9347__ = pi31 & new_new_n9346__;
  assign new_new_n9348__ = ~pi31 & ~new_new_n9346__;
  assign new_new_n9349__ = ~new_new_n9342__ & ~new_new_n9347__;
  assign new_new_n9350__ = ~new_new_n9348__ & new_new_n9349__;
  assign new_new_n9351__ = ~new_new_n9341__ & ~new_new_n9350__;
  assign new_new_n9352__ = new_new_n9332__ & new_new_n9351__;
  assign new_new_n9353__ = ~new_new_n9332__ & ~new_new_n9351__;
  assign new_new_n9354__ = ~new_new_n9352__ & ~new_new_n9353__;
  assign new_new_n9355__ = ~new_new_n9033__ & new_new_n9043__;
  assign new_new_n9356__ = ~new_new_n9032__ & ~new_new_n9355__;
  assign new_new_n9357__ = new_new_n9354__ & ~new_new_n9356__;
  assign new_new_n9358__ = ~new_new_n9354__ & new_new_n9356__;
  assign new_new_n9359__ = ~new_new_n9357__ & ~new_new_n9358__;
  assign new_new_n9360__ = new_new_n9330__ & ~new_new_n9359__;
  assign new_new_n9361__ = ~new_new_n9330__ & new_new_n9359__;
  assign new_new_n9362__ = ~new_new_n9360__ & ~new_new_n9361__;
  assign new_new_n9363__ = new_new_n9328__ & new_new_n9362__;
  assign new_new_n9364__ = ~new_new_n9328__ & ~new_new_n9362__;
  assign new_new_n9365__ = ~new_new_n9363__ & ~new_new_n9364__;
  assign new_new_n9366__ = new_new_n9307__ & ~new_new_n9365__;
  assign new_new_n9367__ = ~new_new_n9307__ & new_new_n9365__;
  assign new_new_n9368__ = ~new_new_n9366__ & ~new_new_n9367__;
  assign new_new_n9369__ = ~new_new_n9015__ & ~new_new_n9193__;
  assign new_new_n9370__ = new_new_n9015__ & new_new_n9193__;
  assign new_new_n9371__ = ~new_new_n9369__ & ~new_new_n9370__;
  assign new_new_n9372__ = ~new_new_n8978__ & new_new_n9371__;
  assign new_new_n9373__ = new_new_n9163__ & ~new_new_n9372__;
  assign new_new_n9374__ = new_new_n8978__ & ~new_new_n9371__;
  assign new_new_n9375__ = ~new_new_n9373__ & ~new_new_n9374__;
  assign new_new_n9376__ = new_new_n9368__ & ~new_new_n9375__;
  assign new_new_n9377__ = ~new_new_n9368__ & new_new_n9375__;
  assign new_new_n9378__ = ~new_new_n9376__ & ~new_new_n9377__;
  assign new_new_n9379__ = new_new_n9009__ & new_new_n9015__;
  assign new_new_n9380__ = ~new_new_n9369__ & ~new_new_n9379__;
  assign new_new_n9381__ = ~new_new_n9239__ & ~new_new_n9243__;
  assign new_new_n9382__ = ~new_new_n9240__ & ~new_new_n9381__;
  assign new_new_n9383__ = new_new_n9380__ & new_new_n9382__;
  assign new_new_n9384__ = ~new_new_n9380__ & ~new_new_n9382__;
  assign new_new_n9385__ = ~new_new_n9383__ & ~new_new_n9384__;
  assign new_new_n9386__ = ~new_new_n9228__ & ~new_new_n9234__;
  assign new_new_n9387__ = ~new_new_n9233__ & ~new_new_n9386__;
  assign new_new_n9388__ = pi14 & pi47;
  assign new_new_n9389__ = pi11 & pi50;
  assign new_new_n9390__ = pi12 & pi49;
  assign new_new_n9391__ = ~new_new_n9389__ & ~new_new_n9390__;
  assign new_new_n9392__ = new_new_n9389__ & new_new_n9390__;
  assign new_new_n9393__ = ~new_new_n9391__ & ~new_new_n9392__;
  assign new_new_n9394__ = new_new_n9388__ & ~new_new_n9393__;
  assign new_new_n9395__ = ~new_new_n9388__ & new_new_n9393__;
  assign new_new_n9396__ = ~new_new_n9394__ & ~new_new_n9395__;
  assign new_new_n9397__ = pi30 & pi31;
  assign new_new_n9398__ = pi13 & pi48;
  assign new_new_n9399__ = pi29 & pi32;
  assign new_new_n9400__ = ~new_new_n9398__ & ~new_new_n9399__;
  assign new_new_n9401__ = new_new_n9398__ & new_new_n9399__;
  assign new_new_n9402__ = ~new_new_n9400__ & ~new_new_n9401__;
  assign new_new_n9403__ = new_new_n9397__ & ~new_new_n9402__;
  assign new_new_n9404__ = ~new_new_n9397__ & new_new_n9402__;
  assign new_new_n9405__ = ~new_new_n9403__ & ~new_new_n9404__;
  assign new_new_n9406__ = new_new_n9396__ & new_new_n9405__;
  assign new_new_n9407__ = ~new_new_n9396__ & ~new_new_n9405__;
  assign new_new_n9408__ = ~new_new_n9406__ & ~new_new_n9407__;
  assign new_new_n9409__ = pi16 & pi45;
  assign new_new_n9410__ = pi15 & pi46;
  assign new_new_n9411__ = pi10 & pi51;
  assign new_new_n9412__ = ~new_new_n9410__ & ~new_new_n9411__;
  assign new_new_n9413__ = new_new_n9410__ & new_new_n9411__;
  assign new_new_n9414__ = ~new_new_n9412__ & ~new_new_n9413__;
  assign new_new_n9415__ = new_new_n9409__ & ~new_new_n9414__;
  assign new_new_n9416__ = ~new_new_n9409__ & new_new_n9414__;
  assign new_new_n9417__ = ~new_new_n9415__ & ~new_new_n9416__;
  assign new_new_n9418__ = new_new_n9408__ & ~new_new_n9417__;
  assign new_new_n9419__ = ~new_new_n9408__ & new_new_n9417__;
  assign new_new_n9420__ = ~new_new_n9418__ & ~new_new_n9419__;
  assign new_new_n9421__ = new_new_n9387__ & ~new_new_n9420__;
  assign new_new_n9422__ = ~new_new_n9387__ & new_new_n9420__;
  assign new_new_n9423__ = ~new_new_n9421__ & ~new_new_n9422__;
  assign new_new_n9424__ = pi05 & pi56;
  assign new_new_n9425__ = pi02 & pi59;
  assign new_new_n9426__ = pi00 & pi61;
  assign new_new_n9427__ = ~new_new_n9425__ & ~new_new_n9426__;
  assign new_new_n9428__ = new_new_n9425__ & new_new_n9426__;
  assign new_new_n9429__ = ~new_new_n9427__ & ~new_new_n9428__;
  assign new_new_n9430__ = new_new_n9424__ & ~new_new_n9429__;
  assign new_new_n9431__ = ~new_new_n9424__ & new_new_n9429__;
  assign new_new_n9432__ = ~new_new_n9430__ & ~new_new_n9431__;
  assign new_new_n9433__ = pi25 & pi36;
  assign new_new_n9434__ = pi24 & pi37;
  assign new_new_n9435__ = pi22 & pi39;
  assign new_new_n9436__ = ~new_new_n9434__ & ~new_new_n9435__;
  assign new_new_n9437__ = new_new_n9434__ & new_new_n9435__;
  assign new_new_n9438__ = ~new_new_n9436__ & ~new_new_n9437__;
  assign new_new_n9439__ = new_new_n9433__ & ~new_new_n9438__;
  assign new_new_n9440__ = ~new_new_n9433__ & new_new_n9438__;
  assign new_new_n9441__ = ~new_new_n9439__ & ~new_new_n9440__;
  assign new_new_n9442__ = new_new_n9432__ & new_new_n9441__;
  assign new_new_n9443__ = ~new_new_n9432__ & ~new_new_n9441__;
  assign new_new_n9444__ = ~new_new_n9442__ & ~new_new_n9443__;
  assign new_new_n9445__ = pi06 & pi55;
  assign new_new_n9446__ = ~new_new_n4946__ & ~new_new_n9445__;
  assign new_new_n9447__ = new_new_n4946__ & new_new_n9445__;
  assign new_new_n9448__ = ~new_new_n9446__ & ~new_new_n9447__;
  assign new_new_n9449__ = new_new_n4701__ & ~new_new_n9448__;
  assign new_new_n9450__ = ~new_new_n4701__ & new_new_n9448__;
  assign new_new_n9451__ = ~new_new_n9449__ & ~new_new_n9450__;
  assign new_new_n9452__ = ~new_new_n9444__ & new_new_n9451__;
  assign new_new_n9453__ = new_new_n9444__ & ~new_new_n9451__;
  assign new_new_n9454__ = ~new_new_n9452__ & ~new_new_n9453__;
  assign new_new_n9455__ = new_new_n9423__ & new_new_n9454__;
  assign new_new_n9456__ = ~new_new_n9423__ & ~new_new_n9454__;
  assign new_new_n9457__ = ~new_new_n9455__ & ~new_new_n9456__;
  assign new_new_n9458__ = new_new_n9385__ & ~new_new_n9457__;
  assign new_new_n9459__ = ~new_new_n9385__ & new_new_n9457__;
  assign new_new_n9460__ = ~new_new_n9458__ & ~new_new_n9459__;
  assign new_new_n9461__ = ~new_new_n9247__ & new_new_n9251__;
  assign new_new_n9462__ = ~new_new_n9248__ & ~new_new_n9461__;
  assign new_new_n9463__ = new_new_n9460__ & ~new_new_n9462__;
  assign new_new_n9464__ = ~new_new_n9460__ & new_new_n9462__;
  assign new_new_n9465__ = ~new_new_n9463__ & ~new_new_n9464__;
  assign new_new_n9466__ = ~new_new_n9069__ & ~new_new_n9079__;
  assign new_new_n9467__ = ~new_new_n9068__ & ~new_new_n9466__;
  assign new_new_n9468__ = ~new_new_n9059__ & ~new_new_n9063__;
  assign new_new_n9469__ = ~new_new_n9062__ & ~new_new_n9468__;
  assign new_new_n9470__ = ~new_new_n9050__ & ~new_new_n9054__;
  assign new_new_n9471__ = ~new_new_n9053__ & ~new_new_n9470__;
  assign new_new_n9472__ = ~new_new_n9141__ & ~new_new_n9145__;
  assign new_new_n9473__ = ~new_new_n9144__ & ~new_new_n9472__;
  assign new_new_n9474__ = ~new_new_n9471__ & ~new_new_n9473__;
  assign new_new_n9475__ = new_new_n9471__ & new_new_n9473__;
  assign new_new_n9476__ = ~new_new_n9474__ & ~new_new_n9475__;
  assign new_new_n9477__ = new_new_n9469__ & ~new_new_n9476__;
  assign new_new_n9478__ = ~new_new_n9469__ & new_new_n9476__;
  assign new_new_n9479__ = ~new_new_n9477__ & ~new_new_n9478__;
  assign new_new_n9480__ = ~new_new_n9467__ & ~new_new_n9479__;
  assign new_new_n9481__ = new_new_n9467__ & new_new_n9479__;
  assign new_new_n9482__ = ~new_new_n9480__ & ~new_new_n9481__;
  assign new_new_n9483__ = ~new_new_n9088__ & ~new_new_n9092__;
  assign new_new_n9484__ = ~new_new_n9091__ & ~new_new_n9483__;
  assign new_new_n9485__ = ~new_new_n9023__ & ~new_new_n9027__;
  assign new_new_n9486__ = ~new_new_n9026__ & ~new_new_n9485__;
  assign new_new_n9487__ = ~new_new_n9071__ & ~new_new_n9075__;
  assign new_new_n9488__ = ~new_new_n9074__ & ~new_new_n9487__;
  assign new_new_n9489__ = ~new_new_n9486__ & ~new_new_n9488__;
  assign new_new_n9490__ = new_new_n9486__ & new_new_n9488__;
  assign new_new_n9491__ = ~new_new_n9489__ & ~new_new_n9490__;
  assign new_new_n9492__ = new_new_n9484__ & ~new_new_n9491__;
  assign new_new_n9493__ = ~new_new_n9484__ & new_new_n9491__;
  assign new_new_n9494__ = ~new_new_n9492__ & ~new_new_n9493__;
  assign new_new_n9495__ = new_new_n9482__ & new_new_n9494__;
  assign new_new_n9496__ = ~new_new_n9482__ & ~new_new_n9494__;
  assign new_new_n9497__ = ~new_new_n9495__ & ~new_new_n9496__;
  assign new_new_n9498__ = ~new_new_n9122__ & ~new_new_n9152__;
  assign new_new_n9499__ = ~new_new_n9121__ & ~new_new_n9498__;
  assign new_new_n9500__ = new_new_n9497__ & ~new_new_n9499__;
  assign new_new_n9501__ = ~new_new_n9497__ & new_new_n9499__;
  assign new_new_n9502__ = ~new_new_n9500__ & ~new_new_n9501__;
  assign new_new_n9503__ = ~new_new_n9035__ & ~new_new_n9039__;
  assign new_new_n9504__ = ~new_new_n9038__ & ~new_new_n9503__;
  assign new_new_n9505__ = ~new_new_n9097__ & ~new_new_n9101__;
  assign new_new_n9506__ = ~new_new_n9100__ & ~new_new_n9505__;
  assign new_new_n9507__ = ~new_new_n9504__ & ~new_new_n9506__;
  assign new_new_n9508__ = new_new_n9504__ & new_new_n9506__;
  assign new_new_n9509__ = ~new_new_n9507__ & ~new_new_n9508__;
  assign new_new_n9510__ = new_new_n8828__ & ~new_new_n9132__;
  assign new_new_n9511__ = ~new_new_n9133__ & ~new_new_n9510__;
  assign new_new_n9512__ = new_new_n9509__ & ~new_new_n9511__;
  assign new_new_n9513__ = ~new_new_n9509__ & new_new_n9511__;
  assign new_new_n9514__ = ~new_new_n9512__ & ~new_new_n9513__;
  assign new_new_n9515__ = ~new_new_n9106__ & ~new_new_n9117__;
  assign new_new_n9516__ = ~new_new_n9107__ & ~new_new_n9515__;
  assign new_new_n9517__ = ~new_new_n9139__ & new_new_n9149__;
  assign new_new_n9518__ = ~new_new_n9138__ & ~new_new_n9517__;
  assign new_new_n9519__ = ~new_new_n9516__ & new_new_n9518__;
  assign new_new_n9520__ = new_new_n9516__ & ~new_new_n9518__;
  assign new_new_n9521__ = ~new_new_n9519__ & ~new_new_n9520__;
  assign new_new_n9522__ = ~new_new_n9514__ & new_new_n9521__;
  assign new_new_n9523__ = new_new_n9514__ & ~new_new_n9521__;
  assign new_new_n9524__ = ~new_new_n9522__ & ~new_new_n9523__;
  assign new_new_n9525__ = new_new_n9502__ & new_new_n9524__;
  assign new_new_n9526__ = ~new_new_n9502__ & ~new_new_n9524__;
  assign new_new_n9527__ = ~new_new_n9525__ & ~new_new_n9526__;
  assign new_new_n9528__ = new_new_n9465__ & new_new_n9527__;
  assign new_new_n9529__ = ~new_new_n9465__ & ~new_new_n9527__;
  assign new_new_n9530__ = ~new_new_n9528__ & ~new_new_n9529__;
  assign new_new_n9531__ = new_new_n9378__ & ~new_new_n9530__;
  assign new_new_n9532__ = ~new_new_n9378__ & new_new_n9530__;
  assign new_new_n9533__ = ~new_new_n9531__ & ~new_new_n9532__;
  assign new_new_n9534__ = ~new_new_n9212__ & ~new_new_n9254__;
  assign new_new_n9535__ = ~new_new_n9211__ & ~new_new_n9534__;
  assign new_new_n9536__ = new_new_n9219__ & new_new_n9535__;
  assign new_new_n9537__ = new_new_n9212__ & new_new_n9254__;
  assign new_new_n9538__ = new_new_n9211__ & ~new_new_n9254__;
  assign new_new_n9539__ = ~new_new_n9537__ & ~new_new_n9538__;
  assign new_new_n9540__ = new_new_n9220__ & new_new_n9539__;
  assign new_new_n9541__ = new_new_n9218__ & ~new_new_n9535__;
  assign new_new_n9542__ = ~new_new_n9536__ & ~new_new_n9541__;
  assign new_new_n9543__ = ~new_new_n9540__ & new_new_n9542__;
  assign new_new_n9544__ = ~new_new_n9533__ & ~new_new_n9543__;
  assign new_new_n9545__ = new_new_n9199__ & new_new_n9218__;
  assign new_new_n9546__ = new_new_n9210__ & new_new_n9545__;
  assign new_new_n9547__ = ~new_new_n9199__ & ~new_new_n9218__;
  assign new_new_n9548__ = new_new_n9210__ & ~new_new_n9219__;
  assign new_new_n9549__ = ~new_new_n9547__ & new_new_n9548__;
  assign new_new_n9550__ = ~new_new_n9545__ & ~new_new_n9549__;
  assign new_new_n9551__ = new_new_n9254__ & ~new_new_n9550__;
  assign new_new_n9552__ = ~new_new_n9212__ & new_new_n9219__;
  assign new_new_n9553__ = ~new_new_n9210__ & new_new_n9547__;
  assign new_new_n9554__ = ~new_new_n9552__ & ~new_new_n9553__;
  assign new_new_n9555__ = ~new_new_n9254__ & ~new_new_n9554__;
  assign new_new_n9556__ = new_new_n9211__ & new_new_n9219__;
  assign new_new_n9557__ = ~new_new_n9546__ & ~new_new_n9556__;
  assign new_new_n9558__ = ~new_new_n9551__ & new_new_n9557__;
  assign new_new_n9559__ = ~new_new_n9555__ & new_new_n9558__;
  assign new_new_n9560__ = new_new_n9533__ & ~new_new_n9559__;
  assign po062 = new_new_n9544__ | new_new_n9560__;
  assign new_new_n9562__ = ~new_new_n9218__ & ~new_new_n9535__;
  assign new_new_n9563__ = new_new_n9533__ & ~new_new_n9562__;
  assign new_new_n9564__ = new_new_n9533__ & ~new_new_n9538__;
  assign new_new_n9565__ = ~new_new_n9537__ & ~new_new_n9564__;
  assign new_new_n9566__ = ~new_new_n9219__ & ~new_new_n9565__;
  assign new_new_n9567__ = new_new_n9218__ & new_new_n9535__;
  assign new_new_n9568__ = ~new_new_n9566__ & ~new_new_n9567__;
  assign new_new_n9569__ = ~new_new_n9563__ & new_new_n9568__;
  assign new_new_n9570__ = ~new_new_n9463__ & ~new_new_n9527__;
  assign new_new_n9571__ = ~new_new_n9464__ & ~new_new_n9570__;
  assign new_new_n9572__ = ~new_new_n9352__ & ~new_new_n9356__;
  assign new_new_n9573__ = ~new_new_n9353__ & ~new_new_n9572__;
  assign new_new_n9574__ = ~new_new_n9481__ & ~new_new_n9494__;
  assign new_new_n9575__ = ~new_new_n9480__ & ~new_new_n9574__;
  assign new_new_n9576__ = new_new_n9573__ & ~new_new_n9575__;
  assign new_new_n9577__ = ~new_new_n9573__ & new_new_n9575__;
  assign new_new_n9578__ = ~new_new_n9576__ & ~new_new_n9577__;
  assign new_new_n9579__ = new_new_n9514__ & ~new_new_n9520__;
  assign new_new_n9580__ = ~new_new_n9519__ & ~new_new_n9579__;
  assign new_new_n9581__ = new_new_n9578__ & ~new_new_n9580__;
  assign new_new_n9582__ = ~new_new_n9578__ & new_new_n9580__;
  assign new_new_n9583__ = ~new_new_n9581__ & ~new_new_n9582__;
  assign new_new_n9584__ = ~new_new_n9484__ & ~new_new_n9490__;
  assign new_new_n9585__ = ~new_new_n9489__ & ~new_new_n9584__;
  assign new_new_n9586__ = ~new_new_n9442__ & ~new_new_n9451__;
  assign new_new_n9587__ = ~new_new_n9443__ & ~new_new_n9586__;
  assign new_new_n9588__ = ~new_new_n9585__ & new_new_n9587__;
  assign new_new_n9589__ = new_new_n9585__ & ~new_new_n9587__;
  assign new_new_n9590__ = ~new_new_n9588__ & ~new_new_n9589__;
  assign new_new_n9591__ = ~new_new_n9406__ & ~new_new_n9417__;
  assign new_new_n9592__ = ~new_new_n9407__ & ~new_new_n9591__;
  assign new_new_n9593__ = new_new_n9590__ & new_new_n9592__;
  assign new_new_n9594__ = ~new_new_n9590__ & ~new_new_n9592__;
  assign new_new_n9595__ = ~new_new_n9593__ & ~new_new_n9594__;
  assign new_new_n9596__ = ~new_new_n9295__ & ~new_new_n9300__;
  assign new_new_n9597__ = ~new_new_n9424__ & ~new_new_n9428__;
  assign new_new_n9598__ = ~new_new_n9427__ & ~new_new_n9597__;
  assign new_new_n9599__ = ~new_new_n9258__ & ~new_new_n9262__;
  assign new_new_n9600__ = ~new_new_n9261__ & ~new_new_n9599__;
  assign new_new_n9601__ = ~new_new_n9598__ & ~new_new_n9600__;
  assign new_new_n9602__ = new_new_n9598__ & new_new_n9600__;
  assign new_new_n9603__ = ~new_new_n9601__ & ~new_new_n9602__;
  assign new_new_n9604__ = ~new_new_n4701__ & ~new_new_n9447__;
  assign new_new_n9605__ = ~new_new_n9446__ & ~new_new_n9604__;
  assign new_new_n9606__ = ~new_new_n9603__ & new_new_n9605__;
  assign new_new_n9607__ = new_new_n9603__ & ~new_new_n9605__;
  assign new_new_n9608__ = ~new_new_n9606__ & ~new_new_n9607__;
  assign new_new_n9609__ = pi01 & pi61;
  assign new_new_n9610__ = pi30 & pi32;
  assign new_new_n9611__ = new_new_n9609__ & ~new_new_n9610__;
  assign new_new_n9612__ = ~new_new_n9609__ & new_new_n9610__;
  assign new_new_n9613__ = ~new_new_n9611__ & ~new_new_n9612__;
  assign new_new_n9614__ = ~new_new_n9397__ & ~new_new_n9401__;
  assign new_new_n9615__ = ~new_new_n9400__ & ~new_new_n9614__;
  assign new_new_n9616__ = ~new_new_n9388__ & ~new_new_n9392__;
  assign new_new_n9617__ = ~new_new_n9391__ & ~new_new_n9616__;
  assign new_new_n9618__ = new_new_n9615__ & new_new_n9617__;
  assign new_new_n9619__ = ~new_new_n9615__ & ~new_new_n9617__;
  assign new_new_n9620__ = ~new_new_n9618__ & ~new_new_n9619__;
  assign new_new_n9621__ = new_new_n9613__ & new_new_n9620__;
  assign new_new_n9622__ = ~new_new_n9613__ & ~new_new_n9620__;
  assign new_new_n9623__ = ~new_new_n9621__ & ~new_new_n9622__;
  assign new_new_n9624__ = ~new_new_n9608__ & ~new_new_n9623__;
  assign new_new_n9625__ = new_new_n9608__ & new_new_n9623__;
  assign new_new_n9626__ = ~new_new_n9624__ & ~new_new_n9625__;
  assign new_new_n9627__ = ~new_new_n9433__ & ~new_new_n9437__;
  assign new_new_n9628__ = ~new_new_n9436__ & ~new_new_n9627__;
  assign new_new_n9629__ = ~new_new_n9310__ & ~new_new_n9314__;
  assign new_new_n9630__ = ~new_new_n9313__ & ~new_new_n9629__;
  assign new_new_n9631__ = ~new_new_n9279__ & ~new_new_n9283__;
  assign new_new_n9632__ = ~new_new_n9282__ & ~new_new_n9631__;
  assign new_new_n9633__ = ~new_new_n9630__ & ~new_new_n9632__;
  assign new_new_n9634__ = new_new_n9630__ & new_new_n9632__;
  assign new_new_n9635__ = ~new_new_n9633__ & ~new_new_n9634__;
  assign new_new_n9636__ = new_new_n9628__ & ~new_new_n9635__;
  assign new_new_n9637__ = ~new_new_n9628__ & new_new_n9635__;
  assign new_new_n9638__ = ~new_new_n9636__ & ~new_new_n9637__;
  assign new_new_n9639__ = new_new_n9626__ & new_new_n9638__;
  assign new_new_n9640__ = ~new_new_n9626__ & ~new_new_n9638__;
  assign new_new_n9641__ = ~new_new_n9639__ & ~new_new_n9640__;
  assign new_new_n9642__ = ~new_new_n9596__ & new_new_n9641__;
  assign new_new_n9643__ = new_new_n9596__ & ~new_new_n9641__;
  assign new_new_n9644__ = ~new_new_n9642__ & ~new_new_n9643__;
  assign new_new_n9645__ = ~new_new_n9384__ & ~new_new_n9457__;
  assign new_new_n9646__ = ~new_new_n9383__ & ~new_new_n9645__;
  assign new_new_n9647__ = new_new_n9644__ & new_new_n9646__;
  assign new_new_n9648__ = ~new_new_n9644__ & ~new_new_n9646__;
  assign new_new_n9649__ = ~new_new_n9647__ & ~new_new_n9648__;
  assign new_new_n9650__ = new_new_n9595__ & ~new_new_n9649__;
  assign new_new_n9651__ = ~new_new_n9595__ & new_new_n9649__;
  assign new_new_n9652__ = ~new_new_n9650__ & ~new_new_n9651__;
  assign new_new_n9653__ = new_new_n9583__ & new_new_n9652__;
  assign new_new_n9654__ = ~new_new_n9583__ & ~new_new_n9652__;
  assign new_new_n9655__ = ~new_new_n9653__ & ~new_new_n9654__;
  assign new_new_n9656__ = new_new_n9571__ & ~new_new_n9655__;
  assign new_new_n9657__ = ~new_new_n9571__ & new_new_n9655__;
  assign new_new_n9658__ = ~new_new_n9656__ & ~new_new_n9657__;
  assign new_new_n9659__ = pi29 & pi33;
  assign new_new_n9660__ = pi27 & pi35;
  assign new_new_n9661__ = pi28 & pi34;
  assign new_new_n9662__ = ~new_new_n9660__ & ~new_new_n9661__;
  assign new_new_n9663__ = new_new_n9660__ & new_new_n9661__;
  assign new_new_n9664__ = ~new_new_n9662__ & ~new_new_n9663__;
  assign new_new_n9665__ = new_new_n9659__ & ~new_new_n9664__;
  assign new_new_n9666__ = ~new_new_n9659__ & new_new_n9664__;
  assign new_new_n9667__ = ~new_new_n9665__ & ~new_new_n9666__;
  assign new_new_n9668__ = pi19 & pi43;
  assign new_new_n9669__ = pi08 & pi54;
  assign new_new_n9670__ = pi18 & pi44;
  assign new_new_n9671__ = ~new_new_n9669__ & ~new_new_n9670__;
  assign new_new_n9672__ = new_new_n9669__ & new_new_n9670__;
  assign new_new_n9673__ = ~new_new_n9671__ & ~new_new_n9672__;
  assign new_new_n9674__ = new_new_n9668__ & ~new_new_n9673__;
  assign new_new_n9675__ = ~new_new_n9668__ & new_new_n9673__;
  assign new_new_n9676__ = ~new_new_n9674__ & ~new_new_n9675__;
  assign new_new_n9677__ = ~new_new_n9667__ & ~new_new_n9676__;
  assign new_new_n9678__ = new_new_n9667__ & new_new_n9676__;
  assign new_new_n9679__ = ~new_new_n9677__ & ~new_new_n9678__;
  assign new_new_n9680__ = pi24 & pi38;
  assign new_new_n9681__ = pi23 & pi39;
  assign new_new_n9682__ = pi22 & pi40;
  assign new_new_n9683__ = ~new_new_n9681__ & ~new_new_n9682__;
  assign new_new_n9684__ = new_new_n9681__ & new_new_n9682__;
  assign new_new_n9685__ = ~new_new_n9683__ & ~new_new_n9684__;
  assign new_new_n9686__ = new_new_n9680__ & ~new_new_n9685__;
  assign new_new_n9687__ = ~new_new_n9680__ & new_new_n9685__;
  assign new_new_n9688__ = ~new_new_n9686__ & ~new_new_n9687__;
  assign new_new_n9689__ = new_new_n9679__ & ~new_new_n9688__;
  assign new_new_n9690__ = ~new_new_n9679__ & new_new_n9688__;
  assign new_new_n9691__ = ~new_new_n9689__ & ~new_new_n9690__;
  assign new_new_n9692__ = pi17 & pi45;
  assign new_new_n9693__ = pi10 & pi52;
  assign new_new_n9694__ = pi09 & pi53;
  assign new_new_n9695__ = ~new_new_n9693__ & ~new_new_n9694__;
  assign new_new_n9696__ = new_new_n9693__ & new_new_n9694__;
  assign new_new_n9697__ = ~new_new_n9695__ & ~new_new_n9696__;
  assign new_new_n9698__ = new_new_n9692__ & ~new_new_n9697__;
  assign new_new_n9699__ = ~new_new_n9692__ & new_new_n9697__;
  assign new_new_n9700__ = ~new_new_n9698__ & ~new_new_n9699__;
  assign new_new_n9701__ = pi00 & pi62;
  assign new_new_n9702__ = pi02 & new_new_n2803__;
  assign new_new_n9703__ = ~pi02 & ~new_new_n2803__;
  assign new_new_n9704__ = pi60 & ~new_new_n9703__;
  assign new_new_n9705__ = ~new_new_n9702__ & new_new_n9704__;
  assign new_new_n9706__ = new_new_n9701__ & ~new_new_n9705__;
  assign new_new_n9707__ = ~new_new_n9701__ & new_new_n9705__;
  assign new_new_n9708__ = ~new_new_n9706__ & ~new_new_n9707__;
  assign new_new_n9709__ = new_new_n9700__ & new_new_n9708__;
  assign new_new_n9710__ = ~new_new_n9700__ & ~new_new_n9708__;
  assign new_new_n9711__ = ~new_new_n9709__ & ~new_new_n9710__;
  assign new_new_n9712__ = pi26 & pi36;
  assign new_new_n9713__ = pi25 & pi37;
  assign new_new_n9714__ = pi21 & pi41;
  assign new_new_n9715__ = ~new_new_n9713__ & ~new_new_n9714__;
  assign new_new_n9716__ = new_new_n9713__ & new_new_n9714__;
  assign new_new_n9717__ = ~new_new_n9715__ & ~new_new_n9716__;
  assign new_new_n9718__ = new_new_n9712__ & ~new_new_n9717__;
  assign new_new_n9719__ = ~new_new_n9712__ & new_new_n9717__;
  assign new_new_n9720__ = ~new_new_n9718__ & ~new_new_n9719__;
  assign new_new_n9721__ = ~new_new_n9711__ & new_new_n9720__;
  assign new_new_n9722__ = new_new_n9711__ & ~new_new_n9720__;
  assign new_new_n9723__ = ~new_new_n9721__ & ~new_new_n9722__;
  assign new_new_n9724__ = ~new_new_n9691__ & ~new_new_n9723__;
  assign new_new_n9725__ = new_new_n9691__ & new_new_n9723__;
  assign new_new_n9726__ = ~new_new_n9724__ & ~new_new_n9725__;
  assign new_new_n9727__ = pi07 & pi55;
  assign new_new_n9728__ = pi06 & pi56;
  assign new_new_n9729__ = ~new_new_n9727__ & ~new_new_n9728__;
  assign new_new_n9730__ = new_new_n9727__ & new_new_n9728__;
  assign new_new_n9731__ = ~new_new_n9729__ & ~new_new_n9730__;
  assign new_new_n9732__ = new_new_n4882__ & ~new_new_n9731__;
  assign new_new_n9733__ = ~new_new_n4882__ & new_new_n9731__;
  assign new_new_n9734__ = ~new_new_n9732__ & ~new_new_n9733__;
  assign new_new_n9735__ = pi16 & pi46;
  assign new_new_n9736__ = pi15 & pi47;
  assign new_new_n9737__ = pi11 & pi51;
  assign new_new_n9738__ = ~new_new_n9736__ & ~new_new_n9737__;
  assign new_new_n9739__ = new_new_n9736__ & new_new_n9737__;
  assign new_new_n9740__ = ~new_new_n9738__ & ~new_new_n9739__;
  assign new_new_n9741__ = new_new_n9735__ & ~new_new_n9740__;
  assign new_new_n9742__ = ~new_new_n9735__ & new_new_n9740__;
  assign new_new_n9743__ = ~new_new_n9741__ & ~new_new_n9742__;
  assign new_new_n9744__ = new_new_n9734__ & new_new_n9743__;
  assign new_new_n9745__ = ~new_new_n9734__ & ~new_new_n9743__;
  assign new_new_n9746__ = ~new_new_n9744__ & ~new_new_n9745__;
  assign new_new_n9747__ = pi14 & pi48;
  assign new_new_n9748__ = pi12 & pi50;
  assign new_new_n9749__ = pi13 & pi49;
  assign new_new_n9750__ = ~new_new_n9748__ & ~new_new_n9749__;
  assign new_new_n9751__ = new_new_n9748__ & new_new_n9749__;
  assign new_new_n9752__ = ~new_new_n9750__ & ~new_new_n9751__;
  assign new_new_n9753__ = new_new_n9747__ & ~new_new_n9752__;
  assign new_new_n9754__ = ~new_new_n9747__ & new_new_n9752__;
  assign new_new_n9755__ = ~new_new_n9753__ & ~new_new_n9754__;
  assign new_new_n9756__ = new_new_n9746__ & new_new_n9755__;
  assign new_new_n9757__ = ~new_new_n9746__ & ~new_new_n9755__;
  assign new_new_n9758__ = ~new_new_n9756__ & ~new_new_n9757__;
  assign new_new_n9759__ = new_new_n9726__ & ~new_new_n9758__;
  assign new_new_n9760__ = ~new_new_n9726__ & new_new_n9758__;
  assign new_new_n9761__ = ~new_new_n9759__ & ~new_new_n9760__;
  assign new_new_n9762__ = ~new_new_n9500__ & ~new_new_n9524__;
  assign new_new_n9763__ = ~new_new_n9501__ & ~new_new_n9762__;
  assign new_new_n9764__ = ~new_new_n9761__ & new_new_n9763__;
  assign new_new_n9765__ = new_new_n9761__ & ~new_new_n9763__;
  assign new_new_n9766__ = ~new_new_n9764__ & ~new_new_n9765__;
  assign new_new_n9767__ = ~new_new_n9330__ & ~new_new_n9359__;
  assign new_new_n9768__ = new_new_n9330__ & new_new_n9359__;
  assign new_new_n9769__ = ~new_new_n9328__ & ~new_new_n9768__;
  assign new_new_n9770__ = ~new_new_n9767__ & ~new_new_n9769__;
  assign new_new_n9771__ = new_new_n9766__ & ~new_new_n9770__;
  assign new_new_n9772__ = ~new_new_n9766__ & new_new_n9770__;
  assign new_new_n9773__ = ~new_new_n9771__ & ~new_new_n9772__;
  assign new_new_n9774__ = ~new_new_n9306__ & new_new_n9365__;
  assign new_new_n9775__ = ~new_new_n9305__ & ~new_new_n9774__;
  assign new_new_n9776__ = ~new_new_n9773__ & new_new_n9775__;
  assign new_new_n9777__ = new_new_n9773__ & ~new_new_n9775__;
  assign new_new_n9778__ = ~new_new_n9776__ & ~new_new_n9777__;
  assign new_new_n9779__ = ~new_new_n9469__ & ~new_new_n9475__;
  assign new_new_n9780__ = ~new_new_n9474__ & ~new_new_n9779__;
  assign new_new_n9781__ = ~new_new_n9507__ & ~new_new_n9511__;
  assign new_new_n9782__ = ~new_new_n9508__ & ~new_new_n9781__;
  assign new_new_n9783__ = ~new_new_n9338__ & ~new_new_n9344__;
  assign new_new_n9784__ = pi31 & ~new_new_n9783__;
  assign new_new_n9785__ = ~pi31 & new_new_n9343__;
  assign new_new_n9786__ = new_new_n9335__ & new_new_n9785__;
  assign new_new_n9787__ = ~new_new_n9784__ & ~new_new_n9786__;
  assign new_new_n9788__ = ~new_new_n9782__ & ~new_new_n9787__;
  assign new_new_n9789__ = new_new_n9782__ & new_new_n9787__;
  assign new_new_n9790__ = ~new_new_n9788__ & ~new_new_n9789__;
  assign new_new_n9791__ = new_new_n9780__ & ~new_new_n9790__;
  assign new_new_n9792__ = ~new_new_n9780__ & new_new_n9790__;
  assign new_new_n9793__ = ~new_new_n9791__ & ~new_new_n9792__;
  assign new_new_n9794__ = ~new_new_n9276__ & ~new_new_n9287__;
  assign new_new_n9795__ = ~new_new_n9277__ & ~new_new_n9794__;
  assign new_new_n9796__ = ~new_new_n9319__ & new_new_n9325__;
  assign new_new_n9797__ = ~new_new_n9320__ & ~new_new_n9796__;
  assign new_new_n9798__ = ~new_new_n9409__ & ~new_new_n9413__;
  assign new_new_n9799__ = ~new_new_n9412__ & ~new_new_n9798__;
  assign new_new_n9800__ = ~new_new_n9267__ & ~new_new_n9271__;
  assign new_new_n9801__ = ~new_new_n9270__ & ~new_new_n9800__;
  assign new_new_n9802__ = pi05 & pi57;
  assign new_new_n9803__ = pi04 & pi58;
  assign new_new_n9804__ = pi03 & pi59;
  assign new_new_n9805__ = ~new_new_n9803__ & ~new_new_n9804__;
  assign new_new_n9806__ = new_new_n9803__ & new_new_n9804__;
  assign new_new_n9807__ = ~new_new_n9805__ & ~new_new_n9806__;
  assign new_new_n9808__ = new_new_n9802__ & ~new_new_n9807__;
  assign new_new_n9809__ = ~new_new_n9802__ & new_new_n9807__;
  assign new_new_n9810__ = ~new_new_n9808__ & ~new_new_n9809__;
  assign new_new_n9811__ = new_new_n9801__ & ~new_new_n9810__;
  assign new_new_n9812__ = ~new_new_n9801__ & new_new_n9810__;
  assign new_new_n9813__ = ~new_new_n9811__ & ~new_new_n9812__;
  assign new_new_n9814__ = new_new_n9799__ & ~new_new_n9813__;
  assign new_new_n9815__ = ~new_new_n9799__ & new_new_n9813__;
  assign new_new_n9816__ = ~new_new_n9814__ & ~new_new_n9815__;
  assign new_new_n9817__ = new_new_n9797__ & new_new_n9816__;
  assign new_new_n9818__ = ~new_new_n9797__ & ~new_new_n9816__;
  assign new_new_n9819__ = ~new_new_n9817__ & ~new_new_n9818__;
  assign new_new_n9820__ = new_new_n9795__ & new_new_n9819__;
  assign new_new_n9821__ = ~new_new_n9795__ & ~new_new_n9819__;
  assign new_new_n9822__ = ~new_new_n9820__ & ~new_new_n9821__;
  assign new_new_n9823__ = new_new_n9793__ & new_new_n9822__;
  assign new_new_n9824__ = ~new_new_n9793__ & ~new_new_n9822__;
  assign new_new_n9825__ = ~new_new_n9823__ & ~new_new_n9824__;
  assign new_new_n9826__ = ~new_new_n9421__ & new_new_n9454__;
  assign new_new_n9827__ = ~new_new_n9422__ & ~new_new_n9826__;
  assign new_new_n9828__ = new_new_n9825__ & new_new_n9827__;
  assign new_new_n9829__ = ~new_new_n9825__ & ~new_new_n9827__;
  assign new_new_n9830__ = ~new_new_n9828__ & ~new_new_n9829__;
  assign new_new_n9831__ = new_new_n9778__ & ~new_new_n9830__;
  assign new_new_n9832__ = ~new_new_n9778__ & new_new_n9830__;
  assign new_new_n9833__ = ~new_new_n9831__ & ~new_new_n9832__;
  assign new_new_n9834__ = new_new_n9658__ & new_new_n9833__;
  assign new_new_n9835__ = ~new_new_n9658__ & ~new_new_n9833__;
  assign new_new_n9836__ = ~new_new_n9834__ & ~new_new_n9835__;
  assign new_new_n9837__ = ~new_new_n9569__ & new_new_n9836__;
  assign new_new_n9838__ = new_new_n9569__ & ~new_new_n9836__;
  assign new_new_n9839__ = ~new_new_n9837__ & ~new_new_n9838__;
  assign new_new_n9840__ = ~new_new_n9377__ & new_new_n9530__;
  assign new_new_n9841__ = ~new_new_n9376__ & ~new_new_n9840__;
  assign new_new_n9842__ = new_new_n9839__ & ~new_new_n9841__;
  assign new_new_n9843__ = ~new_new_n9839__ & new_new_n9841__;
  assign po063 = new_new_n9842__ | new_new_n9843__;
  assign new_new_n9845__ = ~new_new_n9657__ & ~new_new_n9833__;
  assign new_new_n9846__ = ~new_new_n9656__ & ~new_new_n9845__;
  assign new_new_n9847__ = ~new_new_n9837__ & ~new_new_n9841__;
  assign new_new_n9848__ = ~new_new_n9838__ & ~new_new_n9847__;
  assign new_new_n9849__ = ~new_new_n9846__ & ~new_new_n9848__;
  assign new_new_n9850__ = new_new_n9846__ & new_new_n9848__;
  assign new_new_n9851__ = ~new_new_n9849__ & ~new_new_n9850__;
  assign new_new_n9852__ = ~new_new_n9776__ & ~new_new_n9830__;
  assign new_new_n9853__ = ~new_new_n9777__ & ~new_new_n9852__;
  assign new_new_n9854__ = ~new_new_n9668__ & ~new_new_n9672__;
  assign new_new_n9855__ = ~new_new_n9671__ & ~new_new_n9854__;
  assign new_new_n9856__ = ~new_new_n9678__ & ~new_new_n9688__;
  assign new_new_n9857__ = ~new_new_n9677__ & ~new_new_n9856__;
  assign new_new_n9858__ = ~new_new_n9744__ & ~new_new_n9755__;
  assign new_new_n9859__ = ~new_new_n9745__ & ~new_new_n9858__;
  assign new_new_n9860__ = new_new_n9857__ & new_new_n9859__;
  assign new_new_n9861__ = ~new_new_n9857__ & ~new_new_n9859__;
  assign new_new_n9862__ = ~new_new_n9860__ & ~new_new_n9861__;
  assign new_new_n9863__ = new_new_n9855__ & ~new_new_n9862__;
  assign new_new_n9864__ = ~new_new_n9855__ & new_new_n9862__;
  assign new_new_n9865__ = ~new_new_n9863__ & ~new_new_n9864__;
  assign new_new_n9866__ = new_new_n9780__ & ~new_new_n9789__;
  assign new_new_n9867__ = ~new_new_n9788__ & ~new_new_n9866__;
  assign new_new_n9868__ = new_new_n9865__ & ~new_new_n9867__;
  assign new_new_n9869__ = ~new_new_n9865__ & new_new_n9867__;
  assign new_new_n9870__ = ~new_new_n9868__ & ~new_new_n9869__;
  assign new_new_n9871__ = ~new_new_n9709__ & ~new_new_n9720__;
  assign new_new_n9872__ = ~new_new_n9710__ & ~new_new_n9871__;
  assign new_new_n9873__ = ~new_new_n9692__ & ~new_new_n9696__;
  assign new_new_n9874__ = ~new_new_n9695__ & ~new_new_n9873__;
  assign new_new_n9875__ = ~new_new_n9659__ & ~new_new_n9663__;
  assign new_new_n9876__ = ~new_new_n9662__ & ~new_new_n9875__;
  assign new_new_n9877__ = ~new_new_n9874__ & ~new_new_n9876__;
  assign new_new_n9878__ = new_new_n9874__ & new_new_n9876__;
  assign new_new_n9879__ = ~new_new_n9877__ & ~new_new_n9878__;
  assign new_new_n9880__ = pi00 & pi63;
  assign new_new_n9881__ = pi30 & pi61;
  assign new_new_n9882__ = ~pi62 & ~new_new_n9881__;
  assign new_new_n9883__ = pi32 & ~new_new_n9881__;
  assign new_new_n9884__ = pi62 & ~new_new_n9883__;
  assign new_new_n9885__ = pi01 & ~new_new_n9882__;
  assign new_new_n9886__ = ~new_new_n9884__ & new_new_n9885__;
  assign new_new_n9887__ = pi32 & ~new_new_n9886__;
  assign new_new_n9888__ = pi01 & new_new_n9884__;
  assign new_new_n9889__ = ~new_new_n9887__ & ~new_new_n9888__;
  assign new_new_n9890__ = new_new_n9880__ & ~new_new_n9889__;
  assign new_new_n9891__ = ~new_new_n9880__ & new_new_n9889__;
  assign new_new_n9892__ = ~new_new_n9890__ & ~new_new_n9891__;
  assign new_new_n9893__ = pi29 & pi34;
  assign new_new_n9894__ = pi28 & pi35;
  assign new_new_n9895__ = pi27 & pi36;
  assign new_new_n9896__ = ~new_new_n9894__ & ~new_new_n9895__;
  assign new_new_n9897__ = new_new_n9894__ & new_new_n9895__;
  assign new_new_n9898__ = ~new_new_n9896__ & ~new_new_n9897__;
  assign new_new_n9899__ = new_new_n9893__ & ~new_new_n9898__;
  assign new_new_n9900__ = ~new_new_n9893__ & new_new_n9898__;
  assign new_new_n9901__ = ~new_new_n9899__ & ~new_new_n9900__;
  assign new_new_n9902__ = ~new_new_n9892__ & new_new_n9901__;
  assign new_new_n9903__ = new_new_n9892__ & ~new_new_n9901__;
  assign new_new_n9904__ = ~new_new_n9902__ & ~new_new_n9903__;
  assign new_new_n9905__ = pi26 & pi37;
  assign new_new_n9906__ = pi24 & pi39;
  assign new_new_n9907__ = pi25 & pi38;
  assign new_new_n9908__ = ~new_new_n9906__ & ~new_new_n9907__;
  assign new_new_n9909__ = new_new_n9906__ & new_new_n9907__;
  assign new_new_n9910__ = ~new_new_n9908__ & ~new_new_n9909__;
  assign new_new_n9911__ = new_new_n9905__ & ~new_new_n9910__;
  assign new_new_n9912__ = ~new_new_n9905__ & new_new_n9910__;
  assign new_new_n9913__ = ~new_new_n9911__ & ~new_new_n9912__;
  assign new_new_n9914__ = new_new_n9904__ & new_new_n9913__;
  assign new_new_n9915__ = ~new_new_n9904__ & ~new_new_n9913__;
  assign new_new_n9916__ = ~new_new_n9914__ & ~new_new_n9915__;
  assign new_new_n9917__ = new_new_n9879__ & ~new_new_n9916__;
  assign new_new_n9918__ = ~new_new_n9879__ & new_new_n9916__;
  assign new_new_n9919__ = ~new_new_n9917__ & ~new_new_n9918__;
  assign new_new_n9920__ = new_new_n9872__ & new_new_n9919__;
  assign new_new_n9921__ = ~new_new_n9872__ & ~new_new_n9919__;
  assign new_new_n9922__ = ~new_new_n9920__ & ~new_new_n9921__;
  assign new_new_n9923__ = ~new_new_n9577__ & ~new_new_n9580__;
  assign new_new_n9924__ = ~new_new_n9576__ & ~new_new_n9923__;
  assign new_new_n9925__ = new_new_n9922__ & ~new_new_n9924__;
  assign new_new_n9926__ = ~new_new_n9922__ & new_new_n9924__;
  assign new_new_n9927__ = ~new_new_n9925__ & ~new_new_n9926__;
  assign new_new_n9928__ = new_new_n9870__ & new_new_n9927__;
  assign new_new_n9929__ = ~new_new_n9870__ & ~new_new_n9927__;
  assign new_new_n9930__ = ~new_new_n9928__ & ~new_new_n9929__;
  assign new_new_n9931__ = ~new_new_n9583__ & ~new_new_n9646__;
  assign new_new_n9932__ = new_new_n9583__ & new_new_n9646__;
  assign new_new_n9933__ = new_new_n9595__ & ~new_new_n9644__;
  assign new_new_n9934__ = ~new_new_n9595__ & new_new_n9644__;
  assign new_new_n9935__ = ~new_new_n9933__ & ~new_new_n9934__;
  assign new_new_n9936__ = ~new_new_n9932__ & ~new_new_n9935__;
  assign new_new_n9937__ = ~new_new_n9931__ & ~new_new_n9936__;
  assign new_new_n9938__ = new_new_n9930__ & new_new_n9937__;
  assign new_new_n9939__ = ~new_new_n9930__ & ~new_new_n9937__;
  assign new_new_n9940__ = ~new_new_n9938__ & ~new_new_n9939__;
  assign new_new_n9941__ = ~new_new_n9823__ & ~new_new_n9827__;
  assign new_new_n9942__ = ~new_new_n9824__ & ~new_new_n9941__;
  assign new_new_n9943__ = ~new_new_n9595__ & ~new_new_n9642__;
  assign new_new_n9944__ = ~new_new_n9643__ & ~new_new_n9943__;
  assign new_new_n9945__ = new_new_n9942__ & new_new_n9944__;
  assign new_new_n9946__ = ~new_new_n9942__ & ~new_new_n9944__;
  assign new_new_n9947__ = ~new_new_n9945__ & ~new_new_n9946__;
  assign new_new_n9948__ = pi31 & pi32;
  assign new_new_n9949__ = pi30 & pi33;
  assign new_new_n9950__ = pi14 & pi49;
  assign new_new_n9951__ = ~new_new_n9949__ & ~new_new_n9950__;
  assign new_new_n9952__ = new_new_n9949__ & new_new_n9950__;
  assign new_new_n9953__ = ~new_new_n9951__ & ~new_new_n9952__;
  assign new_new_n9954__ = new_new_n9948__ & ~new_new_n9953__;
  assign new_new_n9955__ = ~new_new_n9948__ & new_new_n9953__;
  assign new_new_n9956__ = ~new_new_n9954__ & ~new_new_n9955__;
  assign new_new_n9957__ = pi19 & pi44;
  assign new_new_n9958__ = pi07 & pi56;
  assign new_new_n9959__ = pi08 & pi55;
  assign new_new_n9960__ = ~new_new_n9958__ & ~new_new_n9959__;
  assign new_new_n9961__ = new_new_n9958__ & new_new_n9959__;
  assign new_new_n9962__ = ~new_new_n9960__ & ~new_new_n9961__;
  assign new_new_n9963__ = new_new_n9957__ & ~new_new_n9962__;
  assign new_new_n9964__ = ~new_new_n9957__ & new_new_n9962__;
  assign new_new_n9965__ = ~new_new_n9963__ & ~new_new_n9964__;
  assign new_new_n9966__ = new_new_n9956__ & new_new_n9965__;
  assign new_new_n9967__ = ~new_new_n9956__ & ~new_new_n9965__;
  assign new_new_n9968__ = ~new_new_n9966__ & ~new_new_n9967__;
  assign new_new_n9969__ = pi23 & pi40;
  assign new_new_n9970__ = pi20 & pi43;
  assign new_new_n9971__ = pi06 & pi57;
  assign new_new_n9972__ = ~new_new_n9970__ & ~new_new_n9971__;
  assign new_new_n9973__ = new_new_n9970__ & new_new_n9971__;
  assign new_new_n9974__ = ~new_new_n9972__ & ~new_new_n9973__;
  assign new_new_n9975__ = new_new_n9969__ & ~new_new_n9974__;
  assign new_new_n9976__ = ~new_new_n9969__ & new_new_n9974__;
  assign new_new_n9977__ = ~new_new_n9975__ & ~new_new_n9976__;
  assign new_new_n9978__ = ~new_new_n9968__ & new_new_n9977__;
  assign new_new_n9979__ = new_new_n9968__ & ~new_new_n9977__;
  assign new_new_n9980__ = ~new_new_n9978__ & ~new_new_n9979__;
  assign new_new_n9981__ = ~new_new_n9735__ & ~new_new_n9739__;
  assign new_new_n9982__ = ~new_new_n9738__ & ~new_new_n9981__;
  assign new_new_n9983__ = pi04 & pi59;
  assign new_new_n9984__ = pi02 & pi61;
  assign new_new_n9985__ = pi03 & pi60;
  assign new_new_n9986__ = ~new_new_n9984__ & ~new_new_n9985__;
  assign new_new_n9987__ = new_new_n9984__ & new_new_n9985__;
  assign new_new_n9988__ = ~new_new_n9986__ & ~new_new_n9987__;
  assign new_new_n9989__ = new_new_n9983__ & ~new_new_n9988__;
  assign new_new_n9990__ = ~new_new_n9983__ & new_new_n9988__;
  assign new_new_n9991__ = ~new_new_n9989__ & ~new_new_n9990__;
  assign new_new_n9992__ = new_new_n9982__ & ~new_new_n9991__;
  assign new_new_n9993__ = ~new_new_n9982__ & new_new_n9991__;
  assign new_new_n9994__ = ~new_new_n9992__ & ~new_new_n9993__;
  assign new_new_n9995__ = pi22 & pi41;
  assign new_new_n9996__ = pi21 & pi42;
  assign new_new_n9997__ = pi05 & pi58;
  assign new_new_n9998__ = ~new_new_n9996__ & ~new_new_n9997__;
  assign new_new_n9999__ = new_new_n9996__ & new_new_n9997__;
  assign new_new_n10000__ = ~new_new_n9998__ & ~new_new_n9999__;
  assign new_new_n10001__ = new_new_n9995__ & ~new_new_n10000__;
  assign new_new_n10002__ = ~new_new_n9995__ & new_new_n10000__;
  assign new_new_n10003__ = ~new_new_n10001__ & ~new_new_n10002__;
  assign new_new_n10004__ = new_new_n9994__ & ~new_new_n10003__;
  assign new_new_n10005__ = ~new_new_n9994__ & new_new_n10003__;
  assign new_new_n10006__ = ~new_new_n10004__ & ~new_new_n10005__;
  assign new_new_n10007__ = ~new_new_n9980__ & ~new_new_n10006__;
  assign new_new_n10008__ = new_new_n9980__ & new_new_n10006__;
  assign new_new_n10009__ = ~new_new_n10007__ & ~new_new_n10008__;
  assign new_new_n10010__ = pi18 & pi45;
  assign new_new_n10011__ = pi17 & pi46;
  assign new_new_n10012__ = pi09 & pi54;
  assign new_new_n10013__ = ~new_new_n10011__ & ~new_new_n10012__;
  assign new_new_n10014__ = new_new_n10011__ & new_new_n10012__;
  assign new_new_n10015__ = ~new_new_n10013__ & ~new_new_n10014__;
  assign new_new_n10016__ = new_new_n10010__ & ~new_new_n10015__;
  assign new_new_n10017__ = ~new_new_n10010__ & new_new_n10015__;
  assign new_new_n10018__ = ~new_new_n10016__ & ~new_new_n10017__;
  assign new_new_n10019__ = pi15 & pi48;
  assign new_new_n10020__ = pi13 & pi50;
  assign new_new_n10021__ = pi12 & pi51;
  assign new_new_n10022__ = ~new_new_n10020__ & ~new_new_n10021__;
  assign new_new_n10023__ = new_new_n10020__ & new_new_n10021__;
  assign new_new_n10024__ = ~new_new_n10022__ & ~new_new_n10023__;
  assign new_new_n10025__ = new_new_n10019__ & ~new_new_n10024__;
  assign new_new_n10026__ = ~new_new_n10019__ & new_new_n10024__;
  assign new_new_n10027__ = ~new_new_n10025__ & ~new_new_n10026__;
  assign new_new_n10028__ = new_new_n10018__ & new_new_n10027__;
  assign new_new_n10029__ = ~new_new_n10018__ & ~new_new_n10027__;
  assign new_new_n10030__ = ~new_new_n10028__ & ~new_new_n10029__;
  assign new_new_n10031__ = pi16 & pi47;
  assign new_new_n10032__ = pi10 & pi53;
  assign new_new_n10033__ = pi11 & pi52;
  assign new_new_n10034__ = ~new_new_n10032__ & ~new_new_n10033__;
  assign new_new_n10035__ = new_new_n10032__ & new_new_n10033__;
  assign new_new_n10036__ = ~new_new_n10034__ & ~new_new_n10035__;
  assign new_new_n10037__ = new_new_n10031__ & ~new_new_n10036__;
  assign new_new_n10038__ = ~new_new_n10031__ & new_new_n10036__;
  assign new_new_n10039__ = ~new_new_n10037__ & ~new_new_n10038__;
  assign new_new_n10040__ = ~new_new_n10030__ & new_new_n10039__;
  assign new_new_n10041__ = new_new_n10030__ & ~new_new_n10039__;
  assign new_new_n10042__ = ~new_new_n10040__ & ~new_new_n10041__;
  assign new_new_n10043__ = new_new_n10009__ & ~new_new_n10042__;
  assign new_new_n10044__ = ~new_new_n10009__ & new_new_n10042__;
  assign new_new_n10045__ = ~new_new_n10043__ & ~new_new_n10044__;
  assign new_new_n10046__ = new_new_n9947__ & ~new_new_n10045__;
  assign new_new_n10047__ = ~new_new_n9947__ & new_new_n10045__;
  assign new_new_n10048__ = ~new_new_n10046__ & ~new_new_n10047__;
  assign new_new_n10049__ = new_new_n9940__ & new_new_n10048__;
  assign new_new_n10050__ = ~new_new_n9940__ & ~new_new_n10048__;
  assign new_new_n10051__ = ~new_new_n10049__ & ~new_new_n10050__;
  assign new_new_n10052__ = ~new_new_n9853__ & new_new_n10051__;
  assign new_new_n10053__ = new_new_n9853__ & ~new_new_n10051__;
  assign new_new_n10054__ = ~new_new_n10052__ & ~new_new_n10053__;
  assign new_new_n10055__ = ~new_new_n9628__ & ~new_new_n9634__;
  assign new_new_n10056__ = ~new_new_n9633__ & ~new_new_n10055__;
  assign new_new_n10057__ = new_new_n9613__ & ~new_new_n9618__;
  assign new_new_n10058__ = ~new_new_n9619__ & ~new_new_n10057__;
  assign new_new_n10059__ = new_new_n9799__ & ~new_new_n9812__;
  assign new_new_n10060__ = ~new_new_n9811__ & ~new_new_n10059__;
  assign new_new_n10061__ = new_new_n10058__ & ~new_new_n10060__;
  assign new_new_n10062__ = ~new_new_n10058__ & new_new_n10060__;
  assign new_new_n10063__ = ~new_new_n10061__ & ~new_new_n10062__;
  assign new_new_n10064__ = new_new_n10056__ & new_new_n10063__;
  assign new_new_n10065__ = ~new_new_n10056__ & ~new_new_n10063__;
  assign new_new_n10066__ = ~new_new_n10064__ & ~new_new_n10065__;
  assign new_new_n10067__ = ~new_new_n9724__ & ~new_new_n9758__;
  assign new_new_n10068__ = ~new_new_n9725__ & ~new_new_n10067__;
  assign new_new_n10069__ = new_new_n10066__ & ~new_new_n10068__;
  assign new_new_n10070__ = ~new_new_n10066__ & new_new_n10068__;
  assign new_new_n10071__ = ~new_new_n10069__ & ~new_new_n10070__;
  assign new_new_n10072__ = ~new_new_n9602__ & ~new_new_n9605__;
  assign new_new_n10073__ = ~new_new_n9601__ & ~new_new_n10072__;
  assign new_new_n10074__ = ~new_new_n9701__ & ~new_new_n9702__;
  assign new_new_n10075__ = new_new_n9704__ & ~new_new_n10074__;
  assign new_new_n10076__ = ~new_new_n9802__ & ~new_new_n9806__;
  assign new_new_n10077__ = ~new_new_n9805__ & ~new_new_n10076__;
  assign new_new_n10078__ = new_new_n10075__ & new_new_n10077__;
  assign new_new_n10079__ = ~new_new_n10075__ & ~new_new_n10077__;
  assign new_new_n10080__ = ~new_new_n10078__ & ~new_new_n10079__;
  assign new_new_n10081__ = ~new_new_n9712__ & ~new_new_n9716__;
  assign new_new_n10082__ = ~new_new_n9715__ & ~new_new_n10081__;
  assign new_new_n10083__ = ~new_new_n10080__ & new_new_n10082__;
  assign new_new_n10084__ = new_new_n10080__ & ~new_new_n10082__;
  assign new_new_n10085__ = ~new_new_n10083__ & ~new_new_n10084__;
  assign new_new_n10086__ = ~new_new_n9747__ & ~new_new_n9751__;
  assign new_new_n10087__ = ~new_new_n9750__ & ~new_new_n10086__;
  assign new_new_n10088__ = ~new_new_n9680__ & ~new_new_n9684__;
  assign new_new_n10089__ = ~new_new_n9683__ & ~new_new_n10088__;
  assign new_new_n10090__ = ~new_new_n4882__ & ~new_new_n9730__;
  assign new_new_n10091__ = ~new_new_n9729__ & ~new_new_n10090__;
  assign new_new_n10092__ = new_new_n10089__ & new_new_n10091__;
  assign new_new_n10093__ = ~new_new_n10089__ & ~new_new_n10091__;
  assign new_new_n10094__ = ~new_new_n10092__ & ~new_new_n10093__;
  assign new_new_n10095__ = new_new_n10087__ & ~new_new_n10094__;
  assign new_new_n10096__ = ~new_new_n10087__ & new_new_n10094__;
  assign new_new_n10097__ = ~new_new_n10095__ & ~new_new_n10096__;
  assign new_new_n10098__ = ~new_new_n10085__ & ~new_new_n10097__;
  assign new_new_n10099__ = new_new_n10085__ & new_new_n10097__;
  assign new_new_n10100__ = ~new_new_n10098__ & ~new_new_n10099__;
  assign new_new_n10101__ = new_new_n10073__ & ~new_new_n10100__;
  assign new_new_n10102__ = ~new_new_n10073__ & new_new_n10100__;
  assign new_new_n10103__ = ~new_new_n10101__ & ~new_new_n10102__;
  assign new_new_n10104__ = new_new_n10071__ & ~new_new_n10103__;
  assign new_new_n10105__ = ~new_new_n10071__ & new_new_n10103__;
  assign new_new_n10106__ = ~new_new_n10104__ & ~new_new_n10105__;
  assign new_new_n10107__ = ~new_new_n9764__ & ~new_new_n9770__;
  assign new_new_n10108__ = ~new_new_n9765__ & ~new_new_n10107__;
  assign new_new_n10109__ = ~new_new_n9588__ & ~new_new_n9593__;
  assign new_new_n10110__ = ~new_new_n9795__ & ~new_new_n9817__;
  assign new_new_n10111__ = ~new_new_n9818__ & ~new_new_n10110__;
  assign new_new_n10112__ = ~new_new_n10109__ & new_new_n10111__;
  assign new_new_n10113__ = new_new_n10109__ & ~new_new_n10111__;
  assign new_new_n10114__ = ~new_new_n10112__ & ~new_new_n10113__;
  assign new_new_n10115__ = ~new_new_n9625__ & ~new_new_n9638__;
  assign new_new_n10116__ = ~new_new_n9624__ & ~new_new_n10115__;
  assign new_new_n10117__ = new_new_n10114__ & ~new_new_n10116__;
  assign new_new_n10118__ = ~new_new_n10114__ & new_new_n10116__;
  assign new_new_n10119__ = ~new_new_n10117__ & ~new_new_n10118__;
  assign new_new_n10120__ = ~new_new_n10108__ & new_new_n10119__;
  assign new_new_n10121__ = new_new_n10108__ & ~new_new_n10119__;
  assign new_new_n10122__ = ~new_new_n10120__ & ~new_new_n10121__;
  assign new_new_n10123__ = new_new_n10106__ & new_new_n10122__;
  assign new_new_n10124__ = ~new_new_n10106__ & ~new_new_n10122__;
  assign new_new_n10125__ = ~new_new_n10123__ & ~new_new_n10124__;
  assign new_new_n10126__ = new_new_n10054__ & ~new_new_n10125__;
  assign new_new_n10127__ = ~new_new_n10054__ & new_new_n10125__;
  assign new_new_n10128__ = ~new_new_n10126__ & ~new_new_n10127__;
  assign new_new_n10129__ = new_new_n9851__ & new_new_n10128__;
  assign new_new_n10130__ = ~new_new_n9851__ & ~new_new_n10128__;
  assign po064 = new_new_n10129__ | new_new_n10130__;
  assign new_new_n10132__ = ~new_new_n10052__ & ~new_new_n10125__;
  assign new_new_n10133__ = ~new_new_n10053__ & ~new_new_n10132__;
  assign new_new_n10134__ = ~new_new_n9849__ & new_new_n10133__;
  assign new_new_n10135__ = ~new_new_n9850__ & ~new_new_n10133__;
  assign new_new_n10136__ = ~new_new_n10134__ & ~new_new_n10135__;
  assign new_new_n10137__ = ~new_new_n9938__ & ~new_new_n10048__;
  assign new_new_n10138__ = ~new_new_n9939__ & ~new_new_n10137__;
  assign new_new_n10139__ = ~new_new_n10069__ & ~new_new_n10104__;
  assign new_new_n10140__ = pi29 & pi35;
  assign new_new_n10141__ = pi27 & pi37;
  assign new_new_n10142__ = pi28 & pi36;
  assign new_new_n10143__ = ~new_new_n10141__ & ~new_new_n10142__;
  assign new_new_n10144__ = new_new_n10141__ & new_new_n10142__;
  assign new_new_n10145__ = ~new_new_n10143__ & ~new_new_n10144__;
  assign new_new_n10146__ = new_new_n10140__ & ~new_new_n10145__;
  assign new_new_n10147__ = ~new_new_n10140__ & new_new_n10145__;
  assign new_new_n10148__ = ~new_new_n10146__ & ~new_new_n10147__;
  assign new_new_n10149__ = pi26 & pi38;
  assign new_new_n10150__ = pi16 & pi48;
  assign new_new_n10151__ = pi08 & pi56;
  assign new_new_n10152__ = ~new_new_n10150__ & ~new_new_n10151__;
  assign new_new_n10153__ = new_new_n10150__ & new_new_n10151__;
  assign new_new_n10154__ = ~new_new_n10152__ & ~new_new_n10153__;
  assign new_new_n10155__ = new_new_n10149__ & ~new_new_n10154__;
  assign new_new_n10156__ = ~new_new_n10149__ & new_new_n10154__;
  assign new_new_n10157__ = ~new_new_n10155__ & ~new_new_n10156__;
  assign new_new_n10158__ = ~new_new_n10148__ & ~new_new_n10157__;
  assign new_new_n10159__ = new_new_n10148__ & new_new_n10157__;
  assign new_new_n10160__ = ~new_new_n10158__ & ~new_new_n10159__;
  assign new_new_n10161__ = pi31 & pi33;
  assign new_new_n10162__ = pi30 & pi34;
  assign new_new_n10163__ = pi14 & pi50;
  assign new_new_n10164__ = ~new_new_n10162__ & ~new_new_n10163__;
  assign new_new_n10165__ = new_new_n10162__ & new_new_n10163__;
  assign new_new_n10166__ = ~new_new_n10164__ & ~new_new_n10165__;
  assign new_new_n10167__ = new_new_n10161__ & ~new_new_n10166__;
  assign new_new_n10168__ = ~new_new_n10161__ & new_new_n10166__;
  assign new_new_n10169__ = ~new_new_n10167__ & ~new_new_n10168__;
  assign new_new_n10170__ = ~new_new_n10160__ & new_new_n10169__;
  assign new_new_n10171__ = new_new_n10160__ & ~new_new_n10169__;
  assign new_new_n10172__ = ~new_new_n10170__ & ~new_new_n10171__;
  assign new_new_n10173__ = pi20 & pi44;
  assign new_new_n10174__ = pi25 & pi39;
  assign new_new_n10175__ = pi24 & pi40;
  assign new_new_n10176__ = pi23 & pi41;
  assign new_new_n10177__ = ~new_new_n10175__ & ~new_new_n10176__;
  assign new_new_n10178__ = new_new_n10175__ & new_new_n10176__;
  assign new_new_n10179__ = ~new_new_n10177__ & ~new_new_n10178__;
  assign new_new_n10180__ = new_new_n10174__ & ~new_new_n10179__;
  assign new_new_n10181__ = ~new_new_n10174__ & new_new_n10179__;
  assign new_new_n10182__ = ~new_new_n10180__ & ~new_new_n10181__;
  assign new_new_n10183__ = pi17 & pi47;
  assign new_new_n10184__ = pi07 & pi57;
  assign new_new_n10185__ = pi06 & pi58;
  assign new_new_n10186__ = ~new_new_n10184__ & ~new_new_n10185__;
  assign new_new_n10187__ = new_new_n10184__ & new_new_n10185__;
  assign new_new_n10188__ = ~new_new_n10186__ & ~new_new_n10187__;
  assign new_new_n10189__ = new_new_n10183__ & ~new_new_n10188__;
  assign new_new_n10190__ = ~new_new_n10183__ & new_new_n10188__;
  assign new_new_n10191__ = ~new_new_n10189__ & ~new_new_n10190__;
  assign new_new_n10192__ = new_new_n4944__ & ~new_new_n10191__;
  assign new_new_n10193__ = ~new_new_n4944__ & new_new_n10191__;
  assign new_new_n10194__ = ~new_new_n10192__ & ~new_new_n10193__;
  assign new_new_n10195__ = new_new_n10182__ & new_new_n10194__;
  assign new_new_n10196__ = ~new_new_n10182__ & ~new_new_n10194__;
  assign new_new_n10197__ = ~new_new_n10195__ & ~new_new_n10196__;
  assign new_new_n10198__ = new_new_n5236__ & ~new_new_n10197__;
  assign new_new_n10199__ = ~new_new_n5236__ & new_new_n10197__;
  assign new_new_n10200__ = ~new_new_n10198__ & ~new_new_n10199__;
  assign new_new_n10201__ = new_new_n10173__ & new_new_n10200__;
  assign new_new_n10202__ = ~new_new_n10173__ & ~new_new_n10200__;
  assign new_new_n10203__ = ~new_new_n10201__ & ~new_new_n10202__;
  assign new_new_n10204__ = ~new_new_n10172__ & ~new_new_n10203__;
  assign new_new_n10205__ = new_new_n10172__ & new_new_n10203__;
  assign new_new_n10206__ = ~new_new_n10204__ & ~new_new_n10205__;
  assign new_new_n10207__ = pi04 & pi60;
  assign new_new_n10208__ = pi03 & pi61;
  assign new_new_n10209__ = pi02 & pi62;
  assign new_new_n10210__ = ~new_new_n10208__ & ~new_new_n10209__;
  assign new_new_n10211__ = new_new_n10208__ & new_new_n10209__;
  assign new_new_n10212__ = ~new_new_n10210__ & ~new_new_n10211__;
  assign new_new_n10213__ = new_new_n10207__ & ~new_new_n10212__;
  assign new_new_n10214__ = ~new_new_n10207__ & new_new_n10212__;
  assign new_new_n10215__ = ~new_new_n10213__ & ~new_new_n10214__;
  assign new_new_n10216__ = pi01 & pi62;
  assign new_new_n10217__ = ~new_new_n9881__ & new_new_n10216__;
  assign new_new_n10218__ = new_new_n9880__ & ~new_new_n10217__;
  assign new_new_n10219__ = pi01 & ~pi62;
  assign new_new_n10220__ = new_new_n9881__ & new_new_n10219__;
  assign new_new_n10221__ = ~new_new_n10218__ & ~new_new_n10220__;
  assign new_new_n10222__ = pi32 & ~new_new_n10221__;
  assign new_new_n10223__ = ~pi32 & new_new_n9880__;
  assign new_new_n10224__ = new_new_n10216__ & new_new_n10223__;
  assign new_new_n10225__ = ~new_new_n10222__ & ~new_new_n10224__;
  assign new_new_n10226__ = new_new_n10215__ & new_new_n10225__;
  assign new_new_n10227__ = ~new_new_n10215__ & ~new_new_n10225__;
  assign new_new_n10228__ = ~new_new_n10226__ & ~new_new_n10227__;
  assign new_new_n10229__ = pi19 & pi45;
  assign new_new_n10230__ = pi18 & pi46;
  assign new_new_n10231__ = pi05 & pi59;
  assign new_new_n10232__ = ~new_new_n10230__ & ~new_new_n10231__;
  assign new_new_n10233__ = new_new_n10230__ & new_new_n10231__;
  assign new_new_n10234__ = ~new_new_n10232__ & ~new_new_n10233__;
  assign new_new_n10235__ = new_new_n10229__ & ~new_new_n10234__;
  assign new_new_n10236__ = ~new_new_n10229__ & new_new_n10234__;
  assign new_new_n10237__ = ~new_new_n10235__ & ~new_new_n10236__;
  assign new_new_n10238__ = new_new_n10228__ & ~new_new_n10237__;
  assign new_new_n10239__ = ~new_new_n10228__ & new_new_n10237__;
  assign new_new_n10240__ = ~new_new_n10238__ & ~new_new_n10239__;
  assign new_new_n10241__ = new_new_n10206__ & ~new_new_n10240__;
  assign new_new_n10242__ = ~new_new_n10206__ & new_new_n10240__;
  assign new_new_n10243__ = ~new_new_n10241__ & ~new_new_n10242__;
  assign new_new_n10244__ = new_new_n10139__ & new_new_n10243__;
  assign new_new_n10245__ = ~new_new_n10139__ & ~new_new_n10243__;
  assign new_new_n10246__ = ~new_new_n10244__ & ~new_new_n10245__;
  assign new_new_n10247__ = new_new_n9865__ & new_new_n9879__;
  assign new_new_n10248__ = ~new_new_n9865__ & ~new_new_n9879__;
  assign new_new_n10249__ = ~new_new_n10247__ & ~new_new_n10248__;
  assign new_new_n10250__ = ~new_new_n9860__ & new_new_n10249__;
  assign new_new_n10251__ = ~new_new_n9861__ & ~new_new_n10250__;
  assign new_new_n10252__ = ~new_new_n9855__ & ~new_new_n9878__;
  assign new_new_n10253__ = ~new_new_n9877__ & ~new_new_n10252__;
  assign new_new_n10254__ = ~new_new_n10087__ & ~new_new_n10092__;
  assign new_new_n10255__ = ~new_new_n10093__ & ~new_new_n10254__;
  assign new_new_n10256__ = new_new_n10253__ & new_new_n10255__;
  assign new_new_n10257__ = ~new_new_n10253__ & ~new_new_n10255__;
  assign new_new_n10258__ = ~new_new_n10256__ & ~new_new_n10257__;
  assign new_new_n10259__ = ~new_new_n10078__ & ~new_new_n10082__;
  assign new_new_n10260__ = ~new_new_n10079__ & ~new_new_n10259__;
  assign new_new_n10261__ = ~new_new_n10258__ & new_new_n10260__;
  assign new_new_n10262__ = new_new_n10258__ & ~new_new_n10260__;
  assign new_new_n10263__ = ~new_new_n10261__ & ~new_new_n10262__;
  assign new_new_n10264__ = ~new_new_n10251__ & ~new_new_n10263__;
  assign new_new_n10265__ = new_new_n10251__ & new_new_n10263__;
  assign new_new_n10266__ = new_new_n10073__ & ~new_new_n10099__;
  assign new_new_n10267__ = ~new_new_n10098__ & ~new_new_n10266__;
  assign new_new_n10268__ = ~new_new_n10264__ & new_new_n10267__;
  assign new_new_n10269__ = ~new_new_n10265__ & ~new_new_n10268__;
  assign new_new_n10270__ = ~new_new_n10264__ & new_new_n10269__;
  assign new_new_n10271__ = ~new_new_n10265__ & new_new_n10268__;
  assign new_new_n10272__ = new_new_n10267__ & ~new_new_n10271__;
  assign new_new_n10273__ = ~new_new_n10270__ & ~new_new_n10272__;
  assign new_new_n10274__ = new_new_n10246__ & ~new_new_n10273__;
  assign new_new_n10275__ = ~new_new_n10246__ & new_new_n10273__;
  assign new_new_n10276__ = ~new_new_n10274__ & ~new_new_n10275__;
  assign new_new_n10277__ = new_new_n10106__ & ~new_new_n10121__;
  assign new_new_n10278__ = ~new_new_n10120__ & ~new_new_n10277__;
  assign new_new_n10279__ = ~new_new_n10276__ & ~new_new_n10278__;
  assign new_new_n10280__ = new_new_n10276__ & new_new_n10278__;
  assign new_new_n10281__ = ~new_new_n10279__ & ~new_new_n10280__;
  assign new_new_n10282__ = ~new_new_n10112__ & ~new_new_n10116__;
  assign new_new_n10283__ = ~new_new_n10113__ & ~new_new_n10282__;
  assign new_new_n10284__ = new_new_n10056__ & ~new_new_n10062__;
  assign new_new_n10285__ = ~new_new_n10061__ & ~new_new_n10284__;
  assign new_new_n10286__ = ~new_new_n9948__ & ~new_new_n9952__;
  assign new_new_n10287__ = ~new_new_n9951__ & ~new_new_n10286__;
  assign new_new_n10288__ = pi15 & pi49;
  assign new_new_n10289__ = pi10 & pi54;
  assign new_new_n10290__ = pi09 & pi55;
  assign new_new_n10291__ = ~new_new_n10289__ & ~new_new_n10290__;
  assign new_new_n10292__ = new_new_n10289__ & new_new_n10290__;
  assign new_new_n10293__ = ~new_new_n10291__ & ~new_new_n10292__;
  assign new_new_n10294__ = new_new_n10288__ & ~new_new_n10293__;
  assign new_new_n10295__ = ~new_new_n10288__ & new_new_n10293__;
  assign new_new_n10296__ = ~new_new_n10294__ & ~new_new_n10295__;
  assign new_new_n10297__ = new_new_n10287__ & ~new_new_n10296__;
  assign new_new_n10298__ = ~new_new_n10287__ & new_new_n10296__;
  assign new_new_n10299__ = ~new_new_n10297__ & ~new_new_n10298__;
  assign new_new_n10300__ = pi32 & pi62;
  assign new_new_n10301__ = pi63 & new_new_n10300__;
  assign new_new_n10302__ = ~pi63 & ~new_new_n10300__;
  assign new_new_n10303__ = pi01 & ~new_new_n10302__;
  assign new_new_n10304__ = ~new_new_n10301__ & new_new_n10303__;
  assign new_new_n10305__ = pi13 & pi51;
  assign new_new_n10306__ = pi11 & pi53;
  assign new_new_n10307__ = pi12 & pi52;
  assign new_new_n10308__ = ~new_new_n10306__ & ~new_new_n10307__;
  assign new_new_n10309__ = new_new_n10306__ & new_new_n10307__;
  assign new_new_n10310__ = ~new_new_n10308__ & ~new_new_n10309__;
  assign new_new_n10311__ = new_new_n10305__ & ~new_new_n10310__;
  assign new_new_n10312__ = ~new_new_n10305__ & new_new_n10310__;
  assign new_new_n10313__ = ~new_new_n10311__ & ~new_new_n10312__;
  assign new_new_n10314__ = new_new_n10304__ & ~new_new_n10313__;
  assign new_new_n10315__ = ~new_new_n10304__ & new_new_n10313__;
  assign new_new_n10316__ = ~new_new_n10314__ & ~new_new_n10315__;
  assign new_new_n10317__ = new_new_n10299__ & new_new_n10316__;
  assign new_new_n10318__ = ~new_new_n10299__ & ~new_new_n10316__;
  assign new_new_n10319__ = ~new_new_n10317__ & ~new_new_n10318__;
  assign new_new_n10320__ = new_new_n10285__ & ~new_new_n10319__;
  assign new_new_n10321__ = ~new_new_n10285__ & new_new_n10319__;
  assign new_new_n10322__ = ~new_new_n10320__ & ~new_new_n10321__;
  assign new_new_n10323__ = ~new_new_n9993__ & ~new_new_n10003__;
  assign new_new_n10324__ = ~new_new_n9992__ & ~new_new_n10323__;
  assign new_new_n10325__ = new_new_n10322__ & ~new_new_n10324__;
  assign new_new_n10326__ = ~new_new_n10322__ & new_new_n10324__;
  assign new_new_n10327__ = ~new_new_n10325__ & ~new_new_n10326__;
  assign new_new_n10328__ = ~new_new_n10283__ & new_new_n10327__;
  assign new_new_n10329__ = new_new_n10283__ & ~new_new_n10327__;
  assign new_new_n10330__ = ~new_new_n10328__ & ~new_new_n10329__;
  assign new_new_n10331__ = ~new_new_n10019__ & ~new_new_n10023__;
  assign new_new_n10332__ = ~new_new_n10022__ & ~new_new_n10331__;
  assign new_new_n10333__ = ~new_new_n9905__ & ~new_new_n9909__;
  assign new_new_n10334__ = ~new_new_n9908__ & ~new_new_n10333__;
  assign new_new_n10335__ = ~new_new_n10332__ & ~new_new_n10334__;
  assign new_new_n10336__ = new_new_n10332__ & new_new_n10334__;
  assign new_new_n10337__ = ~new_new_n10335__ & ~new_new_n10336__;
  assign new_new_n10338__ = ~new_new_n10031__ & ~new_new_n10035__;
  assign new_new_n10339__ = ~new_new_n10034__ & ~new_new_n10338__;
  assign new_new_n10340__ = ~new_new_n10337__ & new_new_n10339__;
  assign new_new_n10341__ = new_new_n10337__ & ~new_new_n10339__;
  assign new_new_n10342__ = ~new_new_n10340__ & ~new_new_n10341__;
  assign new_new_n10343__ = ~new_new_n10028__ & ~new_new_n10039__;
  assign new_new_n10344__ = ~new_new_n10029__ & ~new_new_n10343__;
  assign new_new_n10345__ = ~new_new_n9966__ & ~new_new_n9977__;
  assign new_new_n10346__ = ~new_new_n9967__ & ~new_new_n10345__;
  assign new_new_n10347__ = ~new_new_n10344__ & ~new_new_n10346__;
  assign new_new_n10348__ = new_new_n10344__ & new_new_n10346__;
  assign new_new_n10349__ = ~new_new_n10347__ & ~new_new_n10348__;
  assign new_new_n10350__ = new_new_n10342__ & new_new_n10349__;
  assign new_new_n10351__ = ~new_new_n10342__ & ~new_new_n10349__;
  assign new_new_n10352__ = ~new_new_n10350__ & ~new_new_n10351__;
  assign new_new_n10353__ = new_new_n10330__ & ~new_new_n10352__;
  assign new_new_n10354__ = ~new_new_n10330__ & new_new_n10352__;
  assign new_new_n10355__ = ~new_new_n10353__ & ~new_new_n10354__;
  assign new_new_n10356__ = new_new_n10281__ & ~new_new_n10355__;
  assign new_new_n10357__ = ~new_new_n10281__ & new_new_n10355__;
  assign new_new_n10358__ = ~new_new_n10356__ & ~new_new_n10357__;
  assign new_new_n10359__ = ~new_new_n10138__ & new_new_n10358__;
  assign new_new_n10360__ = new_new_n10138__ & ~new_new_n10358__;
  assign new_new_n10361__ = ~new_new_n10359__ & ~new_new_n10360__;
  assign new_new_n10362__ = ~new_new_n9945__ & ~new_new_n10045__;
  assign new_new_n10363__ = ~new_new_n9946__ & ~new_new_n10362__;
  assign new_new_n10364__ = ~new_new_n9902__ & ~new_new_n9913__;
  assign new_new_n10365__ = ~new_new_n9903__ & ~new_new_n10364__;
  assign new_new_n10366__ = ~new_new_n9957__ & ~new_new_n9961__;
  assign new_new_n10367__ = ~new_new_n9960__ & ~new_new_n10366__;
  assign new_new_n10368__ = ~new_new_n9995__ & ~new_new_n9999__;
  assign new_new_n10369__ = ~new_new_n9998__ & ~new_new_n10368__;
  assign new_new_n10370__ = ~new_new_n10367__ & ~new_new_n10369__;
  assign new_new_n10371__ = new_new_n10367__ & new_new_n10369__;
  assign new_new_n10372__ = ~new_new_n10370__ & ~new_new_n10371__;
  assign new_new_n10373__ = ~new_new_n9983__ & ~new_new_n9987__;
  assign new_new_n10374__ = ~new_new_n9986__ & ~new_new_n10373__;
  assign new_new_n10375__ = ~new_new_n10372__ & new_new_n10374__;
  assign new_new_n10376__ = new_new_n10372__ & ~new_new_n10374__;
  assign new_new_n10377__ = ~new_new_n10375__ & ~new_new_n10376__;
  assign new_new_n10378__ = ~new_new_n10010__ & ~new_new_n10014__;
  assign new_new_n10379__ = ~new_new_n10013__ & ~new_new_n10378__;
  assign new_new_n10380__ = ~new_new_n9893__ & ~new_new_n9897__;
  assign new_new_n10381__ = ~new_new_n9896__ & ~new_new_n10380__;
  assign new_new_n10382__ = ~new_new_n10379__ & ~new_new_n10381__;
  assign new_new_n10383__ = new_new_n10379__ & new_new_n10381__;
  assign new_new_n10384__ = ~new_new_n10382__ & ~new_new_n10383__;
  assign new_new_n10385__ = ~new_new_n9969__ & ~new_new_n9973__;
  assign new_new_n10386__ = ~new_new_n9972__ & ~new_new_n10385__;
  assign new_new_n10387__ = ~new_new_n10384__ & new_new_n10386__;
  assign new_new_n10388__ = ~new_new_n10383__ & ~new_new_n10386__;
  assign new_new_n10389__ = ~new_new_n10382__ & new_new_n10388__;
  assign new_new_n10390__ = ~new_new_n10387__ & ~new_new_n10389__;
  assign new_new_n10391__ = new_new_n10377__ & ~new_new_n10390__;
  assign new_new_n10392__ = ~new_new_n10377__ & new_new_n10390__;
  assign new_new_n10393__ = ~new_new_n10391__ & ~new_new_n10392__;
  assign new_new_n10394__ = new_new_n10365__ & new_new_n10393__;
  assign new_new_n10395__ = ~new_new_n10365__ & ~new_new_n10393__;
  assign new_new_n10396__ = ~new_new_n10394__ & ~new_new_n10395__;
  assign new_new_n10397__ = ~new_new_n10008__ & ~new_new_n10042__;
  assign new_new_n10398__ = ~new_new_n10007__ & ~new_new_n10397__;
  assign new_new_n10399__ = new_new_n10396__ & new_new_n10398__;
  assign new_new_n10400__ = ~new_new_n10396__ & ~new_new_n10398__;
  assign new_new_n10401__ = ~new_new_n10399__ & ~new_new_n10400__;
  assign new_new_n10402__ = ~new_new_n9867__ & ~new_new_n9916__;
  assign new_new_n10403__ = new_new_n9867__ & new_new_n9916__;
  assign new_new_n10404__ = ~new_new_n9872__ & ~new_new_n10403__;
  assign new_new_n10405__ = ~new_new_n10402__ & ~new_new_n10404__;
  assign new_new_n10406__ = new_new_n10401__ & ~new_new_n10405__;
  assign new_new_n10407__ = ~new_new_n10401__ & new_new_n10405__;
  assign new_new_n10408__ = ~new_new_n10406__ & ~new_new_n10407__;
  assign new_new_n10409__ = new_new_n10363__ & ~new_new_n10408__;
  assign new_new_n10410__ = ~new_new_n10363__ & new_new_n10408__;
  assign new_new_n10411__ = ~new_new_n10409__ & ~new_new_n10410__;
  assign new_new_n10412__ = ~new_new_n9924__ & ~new_new_n10249__;
  assign new_new_n10413__ = new_new_n9924__ & new_new_n10249__;
  assign new_new_n10414__ = ~new_new_n10402__ & ~new_new_n10403__;
  assign new_new_n10415__ = ~new_new_n9872__ & ~new_new_n10414__;
  assign new_new_n10416__ = new_new_n9872__ & new_new_n10414__;
  assign new_new_n10417__ = ~new_new_n10415__ & ~new_new_n10416__;
  assign new_new_n10418__ = ~new_new_n10413__ & ~new_new_n10417__;
  assign new_new_n10419__ = ~new_new_n10412__ & ~new_new_n10418__;
  assign new_new_n10420__ = new_new_n10411__ & new_new_n10419__;
  assign new_new_n10421__ = ~new_new_n10411__ & ~new_new_n10419__;
  assign new_new_n10422__ = ~new_new_n10420__ & ~new_new_n10421__;
  assign new_new_n10423__ = new_new_n10361__ & ~new_new_n10422__;
  assign new_new_n10424__ = ~new_new_n10361__ & new_new_n10422__;
  assign new_new_n10425__ = ~new_new_n10423__ & ~new_new_n10424__;
  assign new_new_n10426__ = new_new_n10052__ & new_new_n10125__;
  assign new_new_n10427__ = new_new_n10053__ & ~new_new_n10125__;
  assign new_new_n10428__ = ~new_new_n10426__ & ~new_new_n10427__;
  assign new_new_n10429__ = new_new_n9851__ & new_new_n10428__;
  assign new_new_n10430__ = ~new_new_n10136__ & ~new_new_n10425__;
  assign new_new_n10431__ = ~new_new_n10429__ & new_new_n10430__;
  assign new_new_n10432__ = new_new_n9850__ & new_new_n10052__;
  assign new_new_n10433__ = new_new_n9849__ & ~new_new_n10051__;
  assign new_new_n10434__ = new_new_n9853__ & new_new_n10433__;
  assign new_new_n10435__ = ~new_new_n9849__ & new_new_n10051__;
  assign new_new_n10436__ = ~new_new_n9853__ & new_new_n10435__;
  assign new_new_n10437__ = new_new_n9850__ & ~new_new_n10053__;
  assign new_new_n10438__ = new_new_n10125__ & ~new_new_n10437__;
  assign new_new_n10439__ = ~new_new_n10436__ & new_new_n10438__;
  assign new_new_n10440__ = ~new_new_n9850__ & new_new_n9853__;
  assign new_new_n10441__ = ~new_new_n10435__ & new_new_n10440__;
  assign new_new_n10442__ = ~new_new_n10125__ & ~new_new_n10433__;
  assign new_new_n10443__ = ~new_new_n10441__ & new_new_n10442__;
  assign new_new_n10444__ = ~new_new_n10439__ & ~new_new_n10443__;
  assign new_new_n10445__ = new_new_n10425__ & ~new_new_n10432__;
  assign new_new_n10446__ = ~new_new_n10434__ & new_new_n10445__;
  assign new_new_n10447__ = ~new_new_n10444__ & new_new_n10446__;
  assign po065 = ~new_new_n10431__ & ~new_new_n10447__;
  assign new_new_n10449__ = ~new_new_n10359__ & ~new_new_n10422__;
  assign new_new_n10450__ = ~new_new_n10360__ & ~new_new_n10449__;
  assign new_new_n10451__ = ~new_new_n10244__ & new_new_n10273__;
  assign new_new_n10452__ = ~new_new_n10245__ & ~new_new_n10451__;
  assign new_new_n10453__ = ~new_new_n10183__ & ~new_new_n10187__;
  assign new_new_n10454__ = ~new_new_n10186__ & ~new_new_n10453__;
  assign new_new_n10455__ = ~new_new_n10207__ & ~new_new_n10211__;
  assign new_new_n10456__ = ~new_new_n10210__ & ~new_new_n10455__;
  assign new_new_n10457__ = ~new_new_n10149__ & ~new_new_n10153__;
  assign new_new_n10458__ = ~new_new_n10152__ & ~new_new_n10457__;
  assign new_new_n10459__ = ~new_new_n10456__ & ~new_new_n10458__;
  assign new_new_n10460__ = new_new_n10456__ & new_new_n10458__;
  assign new_new_n10461__ = ~new_new_n10459__ & ~new_new_n10460__;
  assign new_new_n10462__ = new_new_n10454__ & ~new_new_n10461__;
  assign new_new_n10463__ = ~new_new_n10454__ & new_new_n10461__;
  assign new_new_n10464__ = ~new_new_n10462__ & ~new_new_n10463__;
  assign new_new_n10465__ = ~new_new_n10229__ & ~new_new_n10233__;
  assign new_new_n10466__ = ~new_new_n10232__ & ~new_new_n10465__;
  assign new_new_n10467__ = ~new_new_n10174__ & ~new_new_n10178__;
  assign new_new_n10468__ = ~new_new_n10177__ & ~new_new_n10467__;
  assign new_new_n10469__ = ~new_new_n10288__ & ~new_new_n10292__;
  assign new_new_n10470__ = ~new_new_n10291__ & ~new_new_n10469__;
  assign new_new_n10471__ = new_new_n10468__ & new_new_n10470__;
  assign new_new_n10472__ = ~new_new_n10468__ & ~new_new_n10470__;
  assign new_new_n10473__ = ~new_new_n10471__ & ~new_new_n10472__;
  assign new_new_n10474__ = new_new_n10466__ & ~new_new_n10473__;
  assign new_new_n10475__ = ~new_new_n10466__ & new_new_n10473__;
  assign new_new_n10476__ = ~new_new_n10474__ & ~new_new_n10475__;
  assign new_new_n10477__ = ~new_new_n10313__ & ~new_new_n10319__;
  assign new_new_n10478__ = new_new_n10313__ & new_new_n10319__;
  assign new_new_n10479__ = ~new_new_n10296__ & ~new_new_n10478__;
  assign new_new_n10480__ = ~new_new_n10477__ & ~new_new_n10479__;
  assign new_new_n10481__ = new_new_n10476__ & ~new_new_n10480__;
  assign new_new_n10482__ = ~new_new_n10476__ & new_new_n10480__;
  assign new_new_n10483__ = ~new_new_n10481__ & ~new_new_n10482__;
  assign new_new_n10484__ = new_new_n10464__ & new_new_n10483__;
  assign new_new_n10485__ = ~new_new_n10464__ & ~new_new_n10483__;
  assign new_new_n10486__ = ~new_new_n10484__ & ~new_new_n10485__;
  assign new_new_n10487__ = ~new_new_n10205__ & ~new_new_n10240__;
  assign new_new_n10488__ = ~new_new_n10204__ & ~new_new_n10487__;
  assign new_new_n10489__ = ~new_new_n10486__ & ~new_new_n10488__;
  assign new_new_n10490__ = new_new_n10486__ & new_new_n10488__;
  assign new_new_n10491__ = ~new_new_n10489__ & ~new_new_n10490__;
  assign new_new_n10492__ = ~new_new_n10321__ & new_new_n10324__;
  assign new_new_n10493__ = ~new_new_n10320__ & ~new_new_n10492__;
  assign new_new_n10494__ = new_new_n10491__ & ~new_new_n10493__;
  assign new_new_n10495__ = ~new_new_n10491__ & new_new_n10493__;
  assign new_new_n10496__ = ~new_new_n10494__ & ~new_new_n10495__;
  assign new_new_n10497__ = new_new_n10452__ & new_new_n10496__;
  assign new_new_n10498__ = ~new_new_n10452__ & ~new_new_n10496__;
  assign new_new_n10499__ = ~new_new_n10497__ & ~new_new_n10498__;
  assign new_new_n10500__ = ~new_new_n10329__ & ~new_new_n10352__;
  assign new_new_n10501__ = ~new_new_n10328__ & ~new_new_n10500__;
  assign new_new_n10502__ = new_new_n10499__ & new_new_n10501__;
  assign new_new_n10503__ = ~new_new_n10499__ & ~new_new_n10501__;
  assign new_new_n10504__ = ~new_new_n10502__ & ~new_new_n10503__;
  assign new_new_n10505__ = new_new_n10450__ & new_new_n10504__;
  assign new_new_n10506__ = ~new_new_n10450__ & ~new_new_n10504__;
  assign new_new_n10507__ = ~new_new_n10505__ & ~new_new_n10506__;
  assign new_new_n10508__ = ~new_new_n10134__ & ~new_new_n10425__;
  assign new_new_n10509__ = new_new_n10425__ & ~new_new_n10427__;
  assign new_new_n10510__ = ~new_new_n10426__ & ~new_new_n10509__;
  assign new_new_n10511__ = ~new_new_n9850__ & new_new_n10510__;
  assign new_new_n10512__ = new_new_n9849__ & ~new_new_n10133__;
  assign new_new_n10513__ = ~new_new_n10511__ & ~new_new_n10512__;
  assign new_new_n10514__ = ~new_new_n10508__ & new_new_n10513__;
  assign new_new_n10515__ = ~new_new_n10409__ & ~new_new_n10419__;
  assign new_new_n10516__ = ~new_new_n10410__ & ~new_new_n10515__;
  assign new_new_n10517__ = ~new_new_n10399__ & new_new_n10405__;
  assign new_new_n10518__ = ~new_new_n10400__ & ~new_new_n10517__;
  assign new_new_n10519__ = pi07 & pi58;
  assign new_new_n10520__ = pi06 & pi59;
  assign new_new_n10521__ = pi05 & pi60;
  assign new_new_n10522__ = ~new_new_n10520__ & ~new_new_n10521__;
  assign new_new_n10523__ = new_new_n10520__ & new_new_n10521__;
  assign new_new_n10524__ = ~new_new_n10522__ & ~new_new_n10523__;
  assign new_new_n10525__ = new_new_n10519__ & ~new_new_n10524__;
  assign new_new_n10526__ = ~new_new_n10519__ & new_new_n10524__;
  assign new_new_n10527__ = ~new_new_n10525__ & ~new_new_n10526__;
  assign new_new_n10528__ = pi22 & pi43;
  assign new_new_n10529__ = pi21 & pi44;
  assign new_new_n10530__ = pi08 & pi57;
  assign new_new_n10531__ = ~new_new_n10529__ & ~new_new_n10530__;
  assign new_new_n10532__ = new_new_n10529__ & new_new_n10530__;
  assign new_new_n10533__ = ~new_new_n10531__ & ~new_new_n10532__;
  assign new_new_n10534__ = new_new_n10528__ & ~new_new_n10533__;
  assign new_new_n10535__ = ~new_new_n10528__ & new_new_n10533__;
  assign new_new_n10536__ = ~new_new_n10534__ & ~new_new_n10535__;
  assign new_new_n10537__ = new_new_n10527__ & new_new_n10536__;
  assign new_new_n10538__ = ~new_new_n10527__ & ~new_new_n10536__;
  assign new_new_n10539__ = ~new_new_n10537__ & ~new_new_n10538__;
  assign new_new_n10540__ = ~new_new_n10287__ & ~new_new_n10301__;
  assign new_new_n10541__ = new_new_n10303__ & ~new_new_n10540__;
  assign new_new_n10542__ = ~new_new_n10539__ & new_new_n10541__;
  assign new_new_n10543__ = new_new_n10539__ & ~new_new_n10541__;
  assign new_new_n10544__ = ~new_new_n10542__ & ~new_new_n10543__;
  assign new_new_n10545__ = pi17 & pi48;
  assign new_new_n10546__ = pi03 & pi62;
  assign new_new_n10547__ = ~pi33 & ~new_new_n10546__;
  assign new_new_n10548__ = pi33 & new_new_n10546__;
  assign new_new_n10549__ = ~new_new_n10547__ & ~new_new_n10548__;
  assign new_new_n10550__ = new_new_n10545__ & ~new_new_n10549__;
  assign new_new_n10551__ = ~new_new_n10545__ & new_new_n10549__;
  assign new_new_n10552__ = ~new_new_n10550__ & ~new_new_n10551__;
  assign new_new_n10553__ = pi31 & pi34;
  assign new_new_n10554__ = pi30 & pi35;
  assign new_new_n10555__ = ~new_new_n10553__ & ~new_new_n10554__;
  assign new_new_n10556__ = new_new_n10553__ & new_new_n10554__;
  assign new_new_n10557__ = ~new_new_n10555__ & ~new_new_n10556__;
  assign new_new_n10558__ = new_new_n6289__ & ~new_new_n10557__;
  assign new_new_n10559__ = ~new_new_n6289__ & new_new_n10557__;
  assign new_new_n10560__ = ~new_new_n10558__ & ~new_new_n10559__;
  assign new_new_n10561__ = ~new_new_n10552__ & ~new_new_n10560__;
  assign new_new_n10562__ = new_new_n10552__ & new_new_n10560__;
  assign new_new_n10563__ = ~new_new_n10561__ & ~new_new_n10562__;
  assign new_new_n10564__ = pi29 & pi36;
  assign new_new_n10565__ = pi19 & pi46;
  assign new_new_n10566__ = pi11 & pi54;
  assign new_new_n10567__ = ~new_new_n10565__ & ~new_new_n10566__;
  assign new_new_n10568__ = new_new_n10565__ & new_new_n10566__;
  assign new_new_n10569__ = ~new_new_n10567__ & ~new_new_n10568__;
  assign new_new_n10570__ = new_new_n10564__ & ~new_new_n10569__;
  assign new_new_n10571__ = ~new_new_n10564__ & new_new_n10569__;
  assign new_new_n10572__ = ~new_new_n10570__ & ~new_new_n10571__;
  assign new_new_n10573__ = ~new_new_n10563__ & new_new_n10572__;
  assign new_new_n10574__ = new_new_n10563__ & ~new_new_n10572__;
  assign new_new_n10575__ = ~new_new_n10573__ & ~new_new_n10574__;
  assign new_new_n10576__ = ~new_new_n10544__ & new_new_n10575__;
  assign new_new_n10577__ = new_new_n10544__ & ~new_new_n10575__;
  assign new_new_n10578__ = ~new_new_n10576__ & ~new_new_n10577__;
  assign new_new_n10579__ = pi25 & pi40;
  assign new_new_n10580__ = pi24 & pi41;
  assign new_new_n10581__ = pi23 & pi42;
  assign new_new_n10582__ = ~new_new_n10580__ & ~new_new_n10581__;
  assign new_new_n10583__ = new_new_n10580__ & new_new_n10581__;
  assign new_new_n10584__ = ~new_new_n10582__ & ~new_new_n10583__;
  assign new_new_n10585__ = new_new_n10579__ & ~new_new_n10584__;
  assign new_new_n10586__ = ~new_new_n10579__ & new_new_n10584__;
  assign new_new_n10587__ = ~new_new_n10585__ & ~new_new_n10586__;
  assign new_new_n10588__ = pi28 & pi37;
  assign new_new_n10589__ = pi27 & pi38;
  assign new_new_n10590__ = pi26 & pi39;
  assign new_new_n10591__ = ~new_new_n10589__ & ~new_new_n10590__;
  assign new_new_n10592__ = new_new_n10589__ & new_new_n10590__;
  assign new_new_n10593__ = ~new_new_n10591__ & ~new_new_n10592__;
  assign new_new_n10594__ = new_new_n10588__ & ~new_new_n10593__;
  assign new_new_n10595__ = ~new_new_n10588__ & new_new_n10593__;
  assign new_new_n10596__ = ~new_new_n10594__ & ~new_new_n10595__;
  assign new_new_n10597__ = pi20 & pi45;
  assign new_new_n10598__ = pi10 & pi55;
  assign new_new_n10599__ = pi09 & pi56;
  assign new_new_n10600__ = ~new_new_n10598__ & ~new_new_n10599__;
  assign new_new_n10601__ = new_new_n10598__ & new_new_n10599__;
  assign new_new_n10602__ = ~new_new_n10600__ & ~new_new_n10601__;
  assign new_new_n10603__ = new_new_n10597__ & ~new_new_n10602__;
  assign new_new_n10604__ = ~new_new_n10597__ & new_new_n10602__;
  assign new_new_n10605__ = ~new_new_n10603__ & ~new_new_n10604__;
  assign new_new_n10606__ = new_new_n10596__ & new_new_n10605__;
  assign new_new_n10607__ = ~new_new_n10596__ & ~new_new_n10605__;
  assign new_new_n10608__ = ~new_new_n10606__ & ~new_new_n10607__;
  assign new_new_n10609__ = ~new_new_n10587__ & new_new_n10608__;
  assign new_new_n10610__ = new_new_n10587__ & ~new_new_n10608__;
  assign new_new_n10611__ = ~new_new_n10609__ & ~new_new_n10610__;
  assign new_new_n10612__ = new_new_n10578__ & ~new_new_n10611__;
  assign new_new_n10613__ = ~new_new_n10578__ & new_new_n10611__;
  assign new_new_n10614__ = ~new_new_n10612__ & ~new_new_n10613__;
  assign new_new_n10615__ = new_new_n10518__ & ~new_new_n10614__;
  assign new_new_n10616__ = ~new_new_n10518__ & new_new_n10614__;
  assign new_new_n10617__ = ~new_new_n10615__ & ~new_new_n10616__;
  assign new_new_n10618__ = ~new_new_n10342__ & ~new_new_n10348__;
  assign new_new_n10619__ = ~new_new_n10347__ & ~new_new_n10618__;
  assign new_new_n10620__ = new_new_n10377__ & new_new_n10390__;
  assign new_new_n10621__ = ~new_new_n10365__ & ~new_new_n10620__;
  assign new_new_n10622__ = ~new_new_n10377__ & ~new_new_n10390__;
  assign new_new_n10623__ = ~new_new_n10621__ & ~new_new_n10622__;
  assign new_new_n10624__ = ~new_new_n10619__ & ~new_new_n10623__;
  assign new_new_n10625__ = new_new_n10619__ & new_new_n10623__;
  assign new_new_n10626__ = ~new_new_n10624__ & ~new_new_n10625__;
  assign new_new_n10627__ = ~new_new_n10382__ & ~new_new_n10388__;
  assign new_new_n10628__ = ~new_new_n10336__ & ~new_new_n10339__;
  assign new_new_n10629__ = ~new_new_n10335__ & ~new_new_n10628__;
  assign new_new_n10630__ = new_new_n10627__ & new_new_n10629__;
  assign new_new_n10631__ = ~new_new_n10371__ & ~new_new_n10374__;
  assign new_new_n10632__ = ~new_new_n10627__ & ~new_new_n10629__;
  assign new_new_n10633__ = ~new_new_n10370__ & ~new_new_n10631__;
  assign new_new_n10634__ = ~new_new_n10632__ & new_new_n10633__;
  assign new_new_n10635__ = ~new_new_n10630__ & new_new_n10634__;
  assign new_new_n10636__ = ~new_new_n10367__ & new_new_n10630__;
  assign new_new_n10637__ = ~new_new_n10374__ & new_new_n10632__;
  assign new_new_n10638__ = ~new_new_n10636__ & ~new_new_n10637__;
  assign new_new_n10639__ = ~new_new_n10369__ & ~new_new_n10638__;
  assign new_new_n10640__ = ~new_new_n10374__ & new_new_n10630__;
  assign new_new_n10641__ = ~new_new_n10367__ & new_new_n10632__;
  assign new_new_n10642__ = ~new_new_n10640__ & ~new_new_n10641__;
  assign new_new_n10643__ = ~new_new_n10377__ & ~new_new_n10642__;
  assign new_new_n10644__ = ~new_new_n10635__ & ~new_new_n10639__;
  assign new_new_n10645__ = ~new_new_n10643__ & new_new_n10644__;
  assign new_new_n10646__ = ~new_new_n10626__ & new_new_n10645__;
  assign new_new_n10647__ = new_new_n10626__ & ~new_new_n10645__;
  assign new_new_n10648__ = ~new_new_n10646__ & ~new_new_n10647__;
  assign new_new_n10649__ = new_new_n10617__ & new_new_n10648__;
  assign new_new_n10650__ = ~new_new_n10617__ & ~new_new_n10648__;
  assign new_new_n10651__ = ~new_new_n10649__ & ~new_new_n10650__;
  assign new_new_n10652__ = new_new_n10516__ & new_new_n10651__;
  assign new_new_n10653__ = ~new_new_n10516__ & ~new_new_n10651__;
  assign new_new_n10654__ = ~new_new_n10652__ & ~new_new_n10653__;
  assign new_new_n10655__ = ~new_new_n10226__ & ~new_new_n10237__;
  assign new_new_n10656__ = ~new_new_n10227__ & ~new_new_n10655__;
  assign new_new_n10657__ = ~new_new_n10256__ & ~new_new_n10260__;
  assign new_new_n10658__ = ~new_new_n10257__ & ~new_new_n10657__;
  assign new_new_n10659__ = new_new_n10656__ & ~new_new_n10658__;
  assign new_new_n10660__ = ~new_new_n10656__ & new_new_n10658__;
  assign new_new_n10661__ = ~new_new_n10659__ & ~new_new_n10660__;
  assign new_new_n10662__ = ~new_new_n10161__ & ~new_new_n10165__;
  assign new_new_n10663__ = ~new_new_n10164__ & ~new_new_n10662__;
  assign new_new_n10664__ = pi04 & pi61;
  assign new_new_n10665__ = pi02 & pi63;
  assign new_new_n10666__ = ~new_new_n10664__ & ~new_new_n10665__;
  assign new_new_n10667__ = new_new_n10664__ & new_new_n10665__;
  assign new_new_n10668__ = ~new_new_n10666__ & ~new_new_n10667__;
  assign new_new_n10669__ = new_new_n10663__ & ~new_new_n10668__;
  assign new_new_n10670__ = ~new_new_n10663__ & new_new_n10668__;
  assign new_new_n10671__ = ~new_new_n10669__ & ~new_new_n10670__;
  assign new_new_n10672__ = pi18 & pi47;
  assign new_new_n10673__ = pi12 & pi53;
  assign new_new_n10674__ = pi13 & pi52;
  assign new_new_n10675__ = ~new_new_n10673__ & ~new_new_n10674__;
  assign new_new_n10676__ = new_new_n10673__ & new_new_n10674__;
  assign new_new_n10677__ = ~new_new_n10675__ & ~new_new_n10676__;
  assign new_new_n10678__ = new_new_n10672__ & ~new_new_n10677__;
  assign new_new_n10679__ = ~new_new_n10672__ & new_new_n10677__;
  assign new_new_n10680__ = ~new_new_n10678__ & ~new_new_n10679__;
  assign new_new_n10681__ = new_new_n10671__ & new_new_n10680__;
  assign new_new_n10682__ = ~new_new_n10671__ & ~new_new_n10680__;
  assign new_new_n10683__ = ~new_new_n10681__ & ~new_new_n10682__;
  assign new_new_n10684__ = pi16 & pi49;
  assign new_new_n10685__ = pi15 & pi50;
  assign new_new_n10686__ = pi14 & pi51;
  assign new_new_n10687__ = ~new_new_n10685__ & ~new_new_n10686__;
  assign new_new_n10688__ = new_new_n10685__ & new_new_n10686__;
  assign new_new_n10689__ = ~new_new_n10687__ & ~new_new_n10688__;
  assign new_new_n10690__ = new_new_n10684__ & ~new_new_n10689__;
  assign new_new_n10691__ = ~new_new_n10684__ & new_new_n10689__;
  assign new_new_n10692__ = ~new_new_n10690__ & ~new_new_n10691__;
  assign new_new_n10693__ = new_new_n10683__ & new_new_n10692__;
  assign new_new_n10694__ = ~new_new_n10683__ & ~new_new_n10692__;
  assign new_new_n10695__ = ~new_new_n10693__ & ~new_new_n10694__;
  assign new_new_n10696__ = new_new_n10661__ & ~new_new_n10695__;
  assign new_new_n10697__ = ~new_new_n10661__ & new_new_n10695__;
  assign new_new_n10698__ = ~new_new_n10696__ & ~new_new_n10697__;
  assign new_new_n10699__ = ~new_new_n10269__ & ~new_new_n10698__;
  assign new_new_n10700__ = new_new_n10269__ & new_new_n10698__;
  assign new_new_n10701__ = ~new_new_n10699__ & ~new_new_n10700__;
  assign new_new_n10702__ = ~new_new_n10159__ & ~new_new_n10169__;
  assign new_new_n10703__ = ~new_new_n10158__ & ~new_new_n10702__;
  assign new_new_n10704__ = ~new_new_n10305__ & ~new_new_n10309__;
  assign new_new_n10705__ = ~new_new_n10308__ & ~new_new_n10704__;
  assign new_new_n10706__ = ~new_new_n10140__ & ~new_new_n10144__;
  assign new_new_n10707__ = ~new_new_n10143__ & ~new_new_n10706__;
  assign new_new_n10708__ = ~new_new_n10705__ & ~new_new_n10707__;
  assign new_new_n10709__ = new_new_n10705__ & new_new_n10707__;
  assign new_new_n10710__ = ~new_new_n10708__ & ~new_new_n10709__;
  assign new_new_n10711__ = ~new_new_n4944__ & ~new_new_n5236__;
  assign new_new_n10712__ = new_new_n4944__ & new_new_n5236__;
  assign new_new_n10713__ = ~new_new_n10173__ & ~new_new_n10712__;
  assign new_new_n10714__ = ~new_new_n10711__ & ~new_new_n10713__;
  assign new_new_n10715__ = ~new_new_n10710__ & new_new_n10714__;
  assign new_new_n10716__ = ~new_new_n10709__ & ~new_new_n10714__;
  assign new_new_n10717__ = ~new_new_n10708__ & new_new_n10716__;
  assign new_new_n10718__ = ~new_new_n10715__ & ~new_new_n10717__;
  assign new_new_n10719__ = new_new_n10182__ & new_new_n10191__;
  assign new_new_n10720__ = ~new_new_n10182__ & ~new_new_n10191__;
  assign new_new_n10721__ = ~new_new_n10711__ & ~new_new_n10712__;
  assign new_new_n10722__ = new_new_n10173__ & ~new_new_n10721__;
  assign new_new_n10723__ = ~new_new_n10173__ & new_new_n10721__;
  assign new_new_n10724__ = ~new_new_n10722__ & ~new_new_n10723__;
  assign new_new_n10725__ = ~new_new_n10720__ & new_new_n10724__;
  assign new_new_n10726__ = ~new_new_n10719__ & ~new_new_n10725__;
  assign new_new_n10727__ = new_new_n10718__ & ~new_new_n10726__;
  assign new_new_n10728__ = ~new_new_n10718__ & new_new_n10726__;
  assign new_new_n10729__ = ~new_new_n10727__ & ~new_new_n10728__;
  assign new_new_n10730__ = new_new_n10703__ & ~new_new_n10729__;
  assign new_new_n10731__ = ~new_new_n10703__ & new_new_n10729__;
  assign new_new_n10732__ = ~new_new_n10730__ & ~new_new_n10731__;
  assign new_new_n10733__ = new_new_n10701__ & ~new_new_n10732__;
  assign new_new_n10734__ = ~new_new_n10701__ & new_new_n10732__;
  assign new_new_n10735__ = ~new_new_n10733__ & ~new_new_n10734__;
  assign new_new_n10736__ = new_new_n10654__ & ~new_new_n10735__;
  assign new_new_n10737__ = ~new_new_n10654__ & new_new_n10735__;
  assign new_new_n10738__ = ~new_new_n10736__ & ~new_new_n10737__;
  assign new_new_n10739__ = ~new_new_n10514__ & ~new_new_n10738__;
  assign new_new_n10740__ = new_new_n10514__ & new_new_n10738__;
  assign new_new_n10741__ = ~new_new_n10739__ & ~new_new_n10740__;
  assign new_new_n10742__ = ~new_new_n10280__ & new_new_n10355__;
  assign new_new_n10743__ = ~new_new_n10279__ & ~new_new_n10742__;
  assign new_new_n10744__ = new_new_n10741__ & ~new_new_n10743__;
  assign new_new_n10745__ = ~new_new_n10741__ & new_new_n10743__;
  assign new_new_n10746__ = ~new_new_n10744__ & ~new_new_n10745__;
  assign new_new_n10747__ = new_new_n10507__ & new_new_n10746__;
  assign new_new_n10748__ = ~new_new_n10507__ & ~new_new_n10746__;
  assign po066 = ~new_new_n10747__ & ~new_new_n10748__;
  assign new_new_n10750__ = ~new_new_n10652__ & ~new_new_n10735__;
  assign new_new_n10751__ = ~new_new_n10653__ & ~new_new_n10750__;
  assign new_new_n10752__ = ~new_new_n10577__ & new_new_n10611__;
  assign new_new_n10753__ = ~new_new_n10576__ & ~new_new_n10752__;
  assign new_new_n10754__ = ~new_new_n10659__ & ~new_new_n10695__;
  assign new_new_n10755__ = ~new_new_n10660__ & ~new_new_n10754__;
  assign new_new_n10756__ = ~new_new_n10753__ & ~new_new_n10755__;
  assign new_new_n10757__ = new_new_n10753__ & new_new_n10755__;
  assign new_new_n10758__ = ~new_new_n10756__ & ~new_new_n10757__;
  assign new_new_n10759__ = ~new_new_n10587__ & ~new_new_n10606__;
  assign new_new_n10760__ = ~new_new_n10607__ & ~new_new_n10759__;
  assign new_new_n10761__ = ~new_new_n10672__ & ~new_new_n10676__;
  assign new_new_n10762__ = ~new_new_n10675__ & ~new_new_n10761__;
  assign new_new_n10763__ = ~new_new_n10579__ & ~new_new_n10583__;
  assign new_new_n10764__ = ~new_new_n10582__ & ~new_new_n10763__;
  assign new_new_n10765__ = ~new_new_n10762__ & ~new_new_n10764__;
  assign new_new_n10766__ = new_new_n10762__ & new_new_n10764__;
  assign new_new_n10767__ = ~new_new_n10765__ & ~new_new_n10766__;
  assign new_new_n10768__ = ~new_new_n10597__ & ~new_new_n10601__;
  assign new_new_n10769__ = ~new_new_n10600__ & ~new_new_n10768__;
  assign new_new_n10770__ = ~new_new_n10767__ & new_new_n10769__;
  assign new_new_n10771__ = ~new_new_n10766__ & ~new_new_n10769__;
  assign new_new_n10772__ = ~new_new_n10765__ & new_new_n10771__;
  assign new_new_n10773__ = ~new_new_n10770__ & ~new_new_n10772__;
  assign new_new_n10774__ = ~new_new_n10537__ & new_new_n10541__;
  assign new_new_n10775__ = ~new_new_n10538__ & ~new_new_n10774__;
  assign new_new_n10776__ = ~new_new_n10773__ & ~new_new_n10775__;
  assign new_new_n10777__ = new_new_n10773__ & new_new_n10775__;
  assign new_new_n10778__ = ~new_new_n10776__ & ~new_new_n10777__;
  assign new_new_n10779__ = new_new_n10760__ & ~new_new_n10778__;
  assign new_new_n10780__ = ~new_new_n10760__ & new_new_n10778__;
  assign new_new_n10781__ = ~new_new_n10779__ & ~new_new_n10780__;
  assign new_new_n10782__ = new_new_n10758__ & ~new_new_n10781__;
  assign new_new_n10783__ = ~new_new_n10758__ & new_new_n10781__;
  assign new_new_n10784__ = ~new_new_n10782__ & ~new_new_n10783__;
  assign new_new_n10785__ = ~new_new_n10630__ & ~new_new_n10634__;
  assign new_new_n10786__ = ~new_new_n10681__ & ~new_new_n10692__;
  assign new_new_n10787__ = ~new_new_n10682__ & ~new_new_n10786__;
  assign new_new_n10788__ = ~new_new_n10785__ & ~new_new_n10787__;
  assign new_new_n10789__ = new_new_n10785__ & new_new_n10787__;
  assign new_new_n10790__ = ~new_new_n10788__ & ~new_new_n10789__;
  assign new_new_n10791__ = ~new_new_n10663__ & ~new_new_n10667__;
  assign new_new_n10792__ = ~new_new_n10666__ & ~new_new_n10791__;
  assign new_new_n10793__ = pi08 & pi58;
  assign new_new_n10794__ = pi06 & pi60;
  assign new_new_n10795__ = pi07 & pi59;
  assign new_new_n10796__ = ~new_new_n10794__ & ~new_new_n10795__;
  assign new_new_n10797__ = new_new_n10794__ & new_new_n10795__;
  assign new_new_n10798__ = ~new_new_n10796__ & ~new_new_n10797__;
  assign new_new_n10799__ = new_new_n10793__ & ~new_new_n10798__;
  assign new_new_n10800__ = ~new_new_n10793__ & new_new_n10798__;
  assign new_new_n10801__ = ~new_new_n10799__ & ~new_new_n10800__;
  assign new_new_n10802__ = ~new_new_n10792__ & new_new_n10801__;
  assign new_new_n10803__ = new_new_n10792__ & ~new_new_n10801__;
  assign new_new_n10804__ = ~new_new_n10588__ & ~new_new_n10592__;
  assign new_new_n10805__ = ~new_new_n10591__ & ~new_new_n10804__;
  assign new_new_n10806__ = ~new_new_n10802__ & new_new_n10805__;
  assign new_new_n10807__ = ~new_new_n10803__ & ~new_new_n10806__;
  assign new_new_n10808__ = ~new_new_n10802__ & new_new_n10807__;
  assign new_new_n10809__ = ~new_new_n10803__ & new_new_n10806__;
  assign new_new_n10810__ = new_new_n10805__ & ~new_new_n10809__;
  assign new_new_n10811__ = ~new_new_n10808__ & ~new_new_n10810__;
  assign new_new_n10812__ = new_new_n10790__ & ~new_new_n10811__;
  assign new_new_n10813__ = ~new_new_n10790__ & new_new_n10811__;
  assign new_new_n10814__ = ~new_new_n10812__ & ~new_new_n10813__;
  assign new_new_n10815__ = ~new_new_n10684__ & ~new_new_n10688__;
  assign new_new_n10816__ = ~new_new_n10687__ & ~new_new_n10815__;
  assign new_new_n10817__ = ~new_new_n6289__ & ~new_new_n10556__;
  assign new_new_n10818__ = ~new_new_n10555__ & ~new_new_n10817__;
  assign new_new_n10819__ = new_new_n10816__ & new_new_n10818__;
  assign new_new_n10820__ = ~new_new_n10816__ & ~new_new_n10818__;
  assign new_new_n10821__ = ~new_new_n10819__ & ~new_new_n10820__;
  assign new_new_n10822__ = ~new_new_n10545__ & ~new_new_n10548__;
  assign new_new_n10823__ = ~new_new_n10547__ & ~new_new_n10822__;
  assign new_new_n10824__ = ~new_new_n10821__ & new_new_n10823__;
  assign new_new_n10825__ = ~new_new_n10819__ & ~new_new_n10823__;
  assign new_new_n10826__ = ~new_new_n10820__ & new_new_n10825__;
  assign new_new_n10827__ = ~new_new_n10824__ & ~new_new_n10826__;
  assign new_new_n10828__ = ~new_new_n10519__ & ~new_new_n10523__;
  assign new_new_n10829__ = ~new_new_n10522__ & ~new_new_n10828__;
  assign new_new_n10830__ = ~new_new_n10528__ & ~new_new_n10532__;
  assign new_new_n10831__ = ~new_new_n10531__ & ~new_new_n10830__;
  assign new_new_n10832__ = ~new_new_n10829__ & ~new_new_n10831__;
  assign new_new_n10833__ = new_new_n10829__ & new_new_n10831__;
  assign new_new_n10834__ = ~new_new_n10832__ & ~new_new_n10833__;
  assign new_new_n10835__ = ~new_new_n10564__ & ~new_new_n10568__;
  assign new_new_n10836__ = ~new_new_n10567__ & ~new_new_n10835__;
  assign new_new_n10837__ = ~new_new_n10834__ & new_new_n10836__;
  assign new_new_n10838__ = new_new_n10834__ & ~new_new_n10836__;
  assign new_new_n10839__ = ~new_new_n10837__ & ~new_new_n10838__;
  assign new_new_n10840__ = ~new_new_n10827__ & ~new_new_n10839__;
  assign new_new_n10841__ = new_new_n10827__ & new_new_n10839__;
  assign new_new_n10842__ = ~new_new_n10840__ & ~new_new_n10841__;
  assign new_new_n10843__ = ~new_new_n10561__ & new_new_n10572__;
  assign new_new_n10844__ = ~new_new_n10562__ & ~new_new_n10843__;
  assign new_new_n10845__ = new_new_n10842__ & ~new_new_n10844__;
  assign new_new_n10846__ = ~new_new_n10842__ & new_new_n10844__;
  assign new_new_n10847__ = ~new_new_n10845__ & ~new_new_n10846__;
  assign new_new_n10848__ = new_new_n10814__ & ~new_new_n10847__;
  assign new_new_n10849__ = ~new_new_n10814__ & new_new_n10847__;
  assign new_new_n10850__ = ~new_new_n10848__ & ~new_new_n10849__;
  assign new_new_n10851__ = ~new_new_n10625__ & new_new_n10645__;
  assign new_new_n10852__ = ~new_new_n10624__ & ~new_new_n10851__;
  assign new_new_n10853__ = new_new_n10850__ & new_new_n10852__;
  assign new_new_n10854__ = ~new_new_n10850__ & ~new_new_n10852__;
  assign new_new_n10855__ = ~new_new_n10853__ & ~new_new_n10854__;
  assign new_new_n10856__ = ~new_new_n10784__ & ~new_new_n10855__;
  assign new_new_n10857__ = new_new_n10784__ & new_new_n10855__;
  assign new_new_n10858__ = ~new_new_n10856__ & ~new_new_n10857__;
  assign new_new_n10859__ = ~new_new_n10700__ & ~new_new_n10732__;
  assign new_new_n10860__ = ~new_new_n10699__ & ~new_new_n10859__;
  assign new_new_n10861__ = new_new_n10858__ & new_new_n10860__;
  assign new_new_n10862__ = ~new_new_n10858__ & ~new_new_n10860__;
  assign new_new_n10863__ = ~new_new_n10861__ & ~new_new_n10862__;
  assign new_new_n10864__ = new_new_n10751__ & ~new_new_n10863__;
  assign new_new_n10865__ = ~new_new_n10751__ & new_new_n10863__;
  assign new_new_n10866__ = ~new_new_n10864__ & ~new_new_n10865__;
  assign new_new_n10867__ = ~new_new_n10497__ & ~new_new_n10501__;
  assign new_new_n10868__ = ~new_new_n10498__ & ~new_new_n10867__;
  assign new_new_n10869__ = ~new_new_n10490__ & ~new_new_n10493__;
  assign new_new_n10870__ = ~new_new_n10489__ & ~new_new_n10869__;
  assign new_new_n10871__ = pi26 & pi40;
  assign new_new_n10872__ = pi25 & pi41;
  assign new_new_n10873__ = pi10 & pi56;
  assign new_new_n10874__ = ~new_new_n10872__ & ~new_new_n10873__;
  assign new_new_n10875__ = new_new_n10872__ & new_new_n10873__;
  assign new_new_n10876__ = ~new_new_n10874__ & ~new_new_n10875__;
  assign new_new_n10877__ = new_new_n10871__ & ~new_new_n10876__;
  assign new_new_n10878__ = ~new_new_n10871__ & new_new_n10876__;
  assign new_new_n10879__ = ~new_new_n10877__ & ~new_new_n10878__;
  assign new_new_n10880__ = pi22 & pi44;
  assign new_new_n10881__ = pi21 & pi45;
  assign new_new_n10882__ = pi20 & pi46;
  assign new_new_n10883__ = ~new_new_n10881__ & ~new_new_n10882__;
  assign new_new_n10884__ = new_new_n10881__ & new_new_n10882__;
  assign new_new_n10885__ = ~new_new_n10883__ & ~new_new_n10884__;
  assign new_new_n10886__ = new_new_n10880__ & ~new_new_n10885__;
  assign new_new_n10887__ = ~new_new_n10880__ & new_new_n10885__;
  assign new_new_n10888__ = ~new_new_n10886__ & ~new_new_n10887__;
  assign new_new_n10889__ = new_new_n10879__ & new_new_n10888__;
  assign new_new_n10890__ = ~new_new_n10879__ & ~new_new_n10888__;
  assign new_new_n10891__ = ~new_new_n10889__ & ~new_new_n10890__;
  assign new_new_n10892__ = pi24 & pi42;
  assign new_new_n10893__ = pi23 & pi43;
  assign new_new_n10894__ = pi09 & pi57;
  assign new_new_n10895__ = ~new_new_n10893__ & ~new_new_n10894__;
  assign new_new_n10896__ = new_new_n10893__ & new_new_n10894__;
  assign new_new_n10897__ = ~new_new_n10895__ & ~new_new_n10896__;
  assign new_new_n10898__ = new_new_n10892__ & ~new_new_n10897__;
  assign new_new_n10899__ = ~new_new_n10892__ & new_new_n10897__;
  assign new_new_n10900__ = ~new_new_n10898__ & ~new_new_n10899__;
  assign new_new_n10901__ = new_new_n10891__ & ~new_new_n10900__;
  assign new_new_n10902__ = ~new_new_n10891__ & new_new_n10900__;
  assign new_new_n10903__ = ~new_new_n10901__ & ~new_new_n10902__;
  assign new_new_n10904__ = pi18 & pi48;
  assign new_new_n10905__ = pi15 & pi51;
  assign new_new_n10906__ = pi13 & pi53;
  assign new_new_n10907__ = ~new_new_n10905__ & ~new_new_n10906__;
  assign new_new_n10908__ = new_new_n10905__ & new_new_n10906__;
  assign new_new_n10909__ = ~new_new_n10907__ & ~new_new_n10908__;
  assign new_new_n10910__ = new_new_n10904__ & ~new_new_n10909__;
  assign new_new_n10911__ = ~new_new_n10904__ & new_new_n10909__;
  assign new_new_n10912__ = ~new_new_n10910__ & ~new_new_n10911__;
  assign new_new_n10913__ = pi32 & pi34;
  assign new_new_n10914__ = pi17 & pi49;
  assign new_new_n10915__ = pi16 & pi50;
  assign new_new_n10916__ = ~new_new_n10914__ & ~new_new_n10915__;
  assign new_new_n10917__ = new_new_n10914__ & new_new_n10915__;
  assign new_new_n10918__ = ~new_new_n10916__ & ~new_new_n10917__;
  assign new_new_n10919__ = new_new_n10913__ & ~new_new_n10918__;
  assign new_new_n10920__ = ~new_new_n10913__ & new_new_n10918__;
  assign new_new_n10921__ = ~new_new_n10919__ & ~new_new_n10920__;
  assign new_new_n10922__ = ~new_new_n10912__ & ~new_new_n10921__;
  assign new_new_n10923__ = new_new_n10912__ & new_new_n10921__;
  assign new_new_n10924__ = ~new_new_n10922__ & ~new_new_n10923__;
  assign new_new_n10925__ = pi31 & pi35;
  assign new_new_n10926__ = pi30 & pi36;
  assign new_new_n10927__ = pi14 & pi52;
  assign new_new_n10928__ = ~new_new_n10926__ & ~new_new_n10927__;
  assign new_new_n10929__ = new_new_n10926__ & new_new_n10927__;
  assign new_new_n10930__ = ~new_new_n10928__ & ~new_new_n10929__;
  assign new_new_n10931__ = new_new_n10925__ & ~new_new_n10930__;
  assign new_new_n10932__ = ~new_new_n10925__ & new_new_n10930__;
  assign new_new_n10933__ = ~new_new_n10931__ & ~new_new_n10932__;
  assign new_new_n10934__ = ~new_new_n10924__ & new_new_n10933__;
  assign new_new_n10935__ = new_new_n10924__ & ~new_new_n10933__;
  assign new_new_n10936__ = ~new_new_n10934__ & ~new_new_n10935__;
  assign new_new_n10937__ = pi19 & pi47;
  assign new_new_n10938__ = pi12 & pi54;
  assign new_new_n10939__ = pi11 & pi55;
  assign new_new_n10940__ = ~new_new_n10938__ & ~new_new_n10939__;
  assign new_new_n10941__ = new_new_n10938__ & new_new_n10939__;
  assign new_new_n10942__ = ~new_new_n10940__ & ~new_new_n10941__;
  assign new_new_n10943__ = new_new_n10937__ & ~new_new_n10942__;
  assign new_new_n10944__ = ~new_new_n10937__ & new_new_n10942__;
  assign new_new_n10945__ = ~new_new_n10943__ & ~new_new_n10944__;
  assign new_new_n10946__ = pi05 & pi61;
  assign new_new_n10947__ = pi04 & pi62;
  assign new_new_n10948__ = pi03 & pi63;
  assign new_new_n10949__ = ~new_new_n10947__ & ~new_new_n10948__;
  assign new_new_n10950__ = new_new_n10947__ & new_new_n10948__;
  assign new_new_n10951__ = ~new_new_n10949__ & ~new_new_n10950__;
  assign new_new_n10952__ = new_new_n10946__ & ~new_new_n10951__;
  assign new_new_n10953__ = ~new_new_n10946__ & new_new_n10951__;
  assign new_new_n10954__ = ~new_new_n10952__ & ~new_new_n10953__;
  assign new_new_n10955__ = new_new_n10945__ & new_new_n10954__;
  assign new_new_n10956__ = ~new_new_n10945__ & ~new_new_n10954__;
  assign new_new_n10957__ = ~new_new_n10955__ & ~new_new_n10956__;
  assign new_new_n10958__ = pi29 & pi37;
  assign new_new_n10959__ = pi27 & pi39;
  assign new_new_n10960__ = pi28 & pi38;
  assign new_new_n10961__ = ~new_new_n10959__ & ~new_new_n10960__;
  assign new_new_n10962__ = new_new_n10959__ & new_new_n10960__;
  assign new_new_n10963__ = ~new_new_n10961__ & ~new_new_n10962__;
  assign new_new_n10964__ = new_new_n10958__ & ~new_new_n10963__;
  assign new_new_n10965__ = ~new_new_n10958__ & new_new_n10963__;
  assign new_new_n10966__ = ~new_new_n10964__ & ~new_new_n10965__;
  assign new_new_n10967__ = new_new_n10957__ & ~new_new_n10966__;
  assign new_new_n10968__ = ~new_new_n10957__ & new_new_n10966__;
  assign new_new_n10969__ = ~new_new_n10967__ & ~new_new_n10968__;
  assign new_new_n10970__ = ~new_new_n10936__ & ~new_new_n10969__;
  assign new_new_n10971__ = new_new_n10936__ & new_new_n10969__;
  assign new_new_n10972__ = ~new_new_n10970__ & ~new_new_n10971__;
  assign new_new_n10973__ = new_new_n10903__ & new_new_n10972__;
  assign new_new_n10974__ = ~new_new_n10903__ & ~new_new_n10972__;
  assign new_new_n10975__ = ~new_new_n10973__ & ~new_new_n10974__;
  assign new_new_n10976__ = new_new_n10870__ & new_new_n10975__;
  assign new_new_n10977__ = ~new_new_n10870__ & ~new_new_n10975__;
  assign new_new_n10978__ = ~new_new_n10976__ & ~new_new_n10977__;
  assign new_new_n10979__ = new_new_n10461__ & ~new_new_n10466__;
  assign new_new_n10980__ = ~new_new_n10461__ & new_new_n10466__;
  assign new_new_n10981__ = ~new_new_n10979__ & ~new_new_n10980__;
  assign new_new_n10982__ = new_new_n10480__ & new_new_n10981__;
  assign new_new_n10983__ = ~new_new_n10480__ & ~new_new_n10981__;
  assign new_new_n10984__ = new_new_n10454__ & ~new_new_n10473__;
  assign new_new_n10985__ = ~new_new_n10454__ & new_new_n10473__;
  assign new_new_n10986__ = ~new_new_n10984__ & ~new_new_n10985__;
  assign new_new_n10987__ = ~new_new_n10983__ & new_new_n10986__;
  assign new_new_n10988__ = ~new_new_n10982__ & ~new_new_n10987__;
  assign new_new_n10989__ = ~new_new_n10454__ & ~new_new_n10471__;
  assign new_new_n10990__ = ~new_new_n10472__ & ~new_new_n10989__;
  assign new_new_n10991__ = ~new_new_n10460__ & ~new_new_n10466__;
  assign new_new_n10992__ = ~new_new_n10459__ & ~new_new_n10991__;
  assign new_new_n10993__ = ~new_new_n10708__ & ~new_new_n10716__;
  assign new_new_n10994__ = new_new_n10992__ & new_new_n10993__;
  assign new_new_n10995__ = ~new_new_n10992__ & ~new_new_n10993__;
  assign new_new_n10996__ = ~new_new_n10994__ & ~new_new_n10995__;
  assign new_new_n10997__ = new_new_n10990__ & ~new_new_n10996__;
  assign new_new_n10998__ = ~new_new_n10990__ & new_new_n10996__;
  assign new_new_n10999__ = ~new_new_n10997__ & ~new_new_n10998__;
  assign new_new_n11000__ = ~new_new_n10988__ & new_new_n10999__;
  assign new_new_n11001__ = new_new_n10988__ & ~new_new_n10999__;
  assign new_new_n11002__ = ~new_new_n11000__ & ~new_new_n11001__;
  assign new_new_n11003__ = new_new_n10703__ & ~new_new_n10728__;
  assign new_new_n11004__ = ~new_new_n10727__ & ~new_new_n11003__;
  assign new_new_n11005__ = new_new_n11002__ & ~new_new_n11004__;
  assign new_new_n11006__ = ~new_new_n11002__ & new_new_n11004__;
  assign new_new_n11007__ = ~new_new_n11005__ & ~new_new_n11006__;
  assign new_new_n11008__ = new_new_n10978__ & ~new_new_n11007__;
  assign new_new_n11009__ = ~new_new_n10978__ & new_new_n11007__;
  assign new_new_n11010__ = ~new_new_n11008__ & ~new_new_n11009__;
  assign new_new_n11011__ = new_new_n10868__ & ~new_new_n11010__;
  assign new_new_n11012__ = ~new_new_n10868__ & new_new_n11010__;
  assign new_new_n11013__ = ~new_new_n10615__ & new_new_n10648__;
  assign new_new_n11014__ = ~new_new_n10616__ & ~new_new_n11013__;
  assign new_new_n11015__ = ~new_new_n11011__ & new_new_n11014__;
  assign new_new_n11016__ = ~new_new_n11012__ & ~new_new_n11015__;
  assign new_new_n11017__ = ~new_new_n11011__ & new_new_n11016__;
  assign new_new_n11018__ = ~new_new_n11012__ & new_new_n11015__;
  assign new_new_n11019__ = new_new_n11014__ & ~new_new_n11018__;
  assign new_new_n11020__ = ~new_new_n11017__ & ~new_new_n11019__;
  assign new_new_n11021__ = new_new_n10866__ & ~new_new_n11020__;
  assign new_new_n11022__ = ~new_new_n10866__ & new_new_n11020__;
  assign new_new_n11023__ = ~new_new_n11021__ & ~new_new_n11022__;
  assign new_new_n11024__ = ~new_new_n10505__ & ~new_new_n10743__;
  assign new_new_n11025__ = ~new_new_n10506__ & ~new_new_n11024__;
  assign new_new_n11026__ = ~new_new_n10739__ & ~new_new_n11025__;
  assign new_new_n11027__ = ~new_new_n10740__ & new_new_n11025__;
  assign new_new_n11028__ = ~new_new_n11026__ & ~new_new_n11027__;
  assign new_new_n11029__ = new_new_n10506__ & ~new_new_n10743__;
  assign new_new_n11030__ = new_new_n10505__ & new_new_n10743__;
  assign new_new_n11031__ = ~new_new_n11029__ & ~new_new_n11030__;
  assign new_new_n11032__ = new_new_n10741__ & new_new_n11031__;
  assign new_new_n11033__ = ~new_new_n11028__ & ~new_new_n11032__;
  assign new_new_n11034__ = ~new_new_n11023__ & ~new_new_n11033__;
  assign new_new_n11035__ = new_new_n10505__ & new_new_n10739__;
  assign new_new_n11036__ = new_new_n10450__ & new_new_n10739__;
  assign new_new_n11037__ = ~new_new_n10450__ & ~new_new_n10739__;
  assign new_new_n11038__ = new_new_n10504__ & ~new_new_n10740__;
  assign new_new_n11039__ = ~new_new_n11037__ & new_new_n11038__;
  assign new_new_n11040__ = ~new_new_n11036__ & ~new_new_n11039__;
  assign new_new_n11041__ = new_new_n10743__ & ~new_new_n11040__;
  assign new_new_n11042__ = new_new_n10506__ & new_new_n10740__;
  assign new_new_n11043__ = ~new_new_n10505__ & new_new_n10740__;
  assign new_new_n11044__ = new_new_n10506__ & ~new_new_n10739__;
  assign new_new_n11045__ = ~new_new_n11043__ & ~new_new_n11044__;
  assign new_new_n11046__ = ~new_new_n10743__ & ~new_new_n11045__;
  assign new_new_n11047__ = ~new_new_n11035__ & ~new_new_n11042__;
  assign new_new_n11048__ = ~new_new_n11046__ & new_new_n11047__;
  assign new_new_n11049__ = ~new_new_n11041__ & new_new_n11048__;
  assign new_new_n11050__ = new_new_n11023__ & ~new_new_n11049__;
  assign po067 = new_new_n11034__ | new_new_n11050__;
  assign new_new_n11052__ = ~new_new_n11023__ & ~new_new_n11026__;
  assign new_new_n11053__ = new_new_n10739__ & new_new_n11025__;
  assign new_new_n11054__ = ~new_new_n11023__ & ~new_new_n11029__;
  assign new_new_n11055__ = ~new_new_n11030__ & ~new_new_n11054__;
  assign new_new_n11056__ = ~new_new_n10740__ & ~new_new_n11055__;
  assign new_new_n11057__ = ~new_new_n11053__ & ~new_new_n11056__;
  assign new_new_n11058__ = ~new_new_n11052__ & new_new_n11057__;
  assign new_new_n11059__ = ~new_new_n10865__ & new_new_n11020__;
  assign new_new_n11060__ = ~new_new_n10864__ & ~new_new_n11059__;
  assign new_new_n11061__ = ~new_new_n11058__ & ~new_new_n11060__;
  assign new_new_n11062__ = new_new_n11058__ & new_new_n11060__;
  assign new_new_n11063__ = ~new_new_n11061__ & ~new_new_n11062__;
  assign new_new_n11064__ = ~new_new_n10857__ & new_new_n10860__;
  assign new_new_n11065__ = ~new_new_n10856__ & ~new_new_n11064__;
  assign new_new_n11066__ = pi24 & pi43;
  assign new_new_n11067__ = ~pi22 & ~new_new_n5601__;
  assign new_new_n11068__ = ~new_new_n5602__ & ~new_new_n11067__;
  assign new_new_n11069__ = pi22 & new_new_n5604__;
  assign new_new_n11070__ = new_new_n11068__ & ~new_new_n11069__;
  assign new_new_n11071__ = new_new_n11066__ & ~new_new_n11070__;
  assign new_new_n11072__ = ~new_new_n11066__ & new_new_n11070__;
  assign new_new_n11073__ = ~new_new_n11071__ & ~new_new_n11072__;
  assign new_new_n11074__ = pi30 & pi37;
  assign new_new_n11075__ = pi16 & pi51;
  assign new_new_n11076__ = pi15 & pi52;
  assign new_new_n11077__ = ~new_new_n11075__ & ~new_new_n11076__;
  assign new_new_n11078__ = new_new_n11075__ & new_new_n11076__;
  assign new_new_n11079__ = ~new_new_n11077__ & ~new_new_n11078__;
  assign new_new_n11080__ = new_new_n11074__ & ~new_new_n11079__;
  assign new_new_n11081__ = ~new_new_n11074__ & new_new_n11079__;
  assign new_new_n11082__ = ~new_new_n11080__ & ~new_new_n11081__;
  assign new_new_n11083__ = new_new_n11073__ & new_new_n11082__;
  assign new_new_n11084__ = ~new_new_n11073__ & ~new_new_n11082__;
  assign new_new_n11085__ = ~new_new_n11083__ & ~new_new_n11084__;
  assign new_new_n11086__ = pi26 & pi41;
  assign new_new_n11087__ = pi25 & pi42;
  assign new_new_n11088__ = pi21 & pi46;
  assign new_new_n11089__ = ~new_new_n11087__ & ~new_new_n11088__;
  assign new_new_n11090__ = new_new_n11087__ & new_new_n11088__;
  assign new_new_n11091__ = ~new_new_n11089__ & ~new_new_n11090__;
  assign new_new_n11092__ = new_new_n11086__ & ~new_new_n11091__;
  assign new_new_n11093__ = ~new_new_n11086__ & new_new_n11091__;
  assign new_new_n11094__ = ~new_new_n11092__ & ~new_new_n11093__;
  assign new_new_n11095__ = pi28 & pi39;
  assign new_new_n11096__ = pi04 & pi63;
  assign new_new_n11097__ = pi27 & pi40;
  assign new_new_n11098__ = ~new_new_n11096__ & ~new_new_n11097__;
  assign new_new_n11099__ = new_new_n11096__ & new_new_n11097__;
  assign new_new_n11100__ = ~new_new_n11098__ & ~new_new_n11099__;
  assign new_new_n11101__ = new_new_n11095__ & ~new_new_n11100__;
  assign new_new_n11102__ = ~new_new_n11095__ & new_new_n11100__;
  assign new_new_n11103__ = ~new_new_n11101__ & ~new_new_n11102__;
  assign new_new_n11104__ = new_new_n11094__ & new_new_n11103__;
  assign new_new_n11105__ = ~new_new_n11094__ & ~new_new_n11103__;
  assign new_new_n11106__ = ~new_new_n11104__ & ~new_new_n11105__;
  assign new_new_n11107__ = pi19 & pi48;
  assign new_new_n11108__ = pi17 & pi50;
  assign new_new_n11109__ = pi14 & pi53;
  assign new_new_n11110__ = ~new_new_n11108__ & ~new_new_n11109__;
  assign new_new_n11111__ = new_new_n11108__ & new_new_n11109__;
  assign new_new_n11112__ = ~new_new_n11110__ & ~new_new_n11111__;
  assign new_new_n11113__ = new_new_n11107__ & ~new_new_n11112__;
  assign new_new_n11114__ = ~new_new_n11107__ & new_new_n11112__;
  assign new_new_n11115__ = ~new_new_n11113__ & ~new_new_n11114__;
  assign new_new_n11116__ = new_new_n11106__ & ~new_new_n11115__;
  assign new_new_n11117__ = ~new_new_n11106__ & new_new_n11115__;
  assign new_new_n11118__ = ~new_new_n11116__ & ~new_new_n11117__;
  assign new_new_n11119__ = new_new_n11085__ & ~new_new_n11118__;
  assign new_new_n11120__ = ~new_new_n11085__ & new_new_n11118__;
  assign new_new_n11121__ = ~new_new_n11119__ & ~new_new_n11120__;
  assign new_new_n11122__ = pi18 & pi49;
  assign new_new_n11123__ = pi05 & pi62;
  assign new_new_n11124__ = ~new_new_n11122__ & ~new_new_n11123__;
  assign new_new_n11125__ = new_new_n11122__ & new_new_n11123__;
  assign new_new_n11126__ = ~new_new_n11124__ & ~new_new_n11125__;
  assign new_new_n11127__ = pi34 & ~new_new_n11126__;
  assign new_new_n11128__ = ~pi34 & ~new_new_n11125__;
  assign new_new_n11129__ = ~new_new_n11124__ & new_new_n11128__;
  assign new_new_n11130__ = ~new_new_n11127__ & ~new_new_n11129__;
  assign new_new_n11131__ = pi29 & pi38;
  assign new_new_n11132__ = pi12 & pi55;
  assign new_new_n11133__ = pi13 & pi54;
  assign new_new_n11134__ = ~new_new_n11132__ & ~new_new_n11133__;
  assign new_new_n11135__ = new_new_n11132__ & new_new_n11133__;
  assign new_new_n11136__ = ~new_new_n11134__ & ~new_new_n11135__;
  assign new_new_n11137__ = new_new_n11131__ & ~new_new_n11136__;
  assign new_new_n11138__ = ~new_new_n11131__ & new_new_n11136__;
  assign new_new_n11139__ = ~new_new_n11137__ & ~new_new_n11138__;
  assign new_new_n11140__ = pi33 & pi34;
  assign new_new_n11141__ = pi32 & pi35;
  assign new_new_n11142__ = pi31 & pi36;
  assign new_new_n11143__ = ~new_new_n11141__ & ~new_new_n11142__;
  assign new_new_n11144__ = new_new_n11141__ & new_new_n11142__;
  assign new_new_n11145__ = ~new_new_n11143__ & ~new_new_n11144__;
  assign new_new_n11146__ = new_new_n11140__ & ~new_new_n11145__;
  assign new_new_n11147__ = ~new_new_n11140__ & new_new_n11145__;
  assign new_new_n11148__ = ~new_new_n11146__ & ~new_new_n11147__;
  assign new_new_n11149__ = pi09 & pi58;
  assign new_new_n11150__ = pi07 & pi60;
  assign new_new_n11151__ = pi08 & pi59;
  assign new_new_n11152__ = ~new_new_n11150__ & ~new_new_n11151__;
  assign new_new_n11153__ = new_new_n11150__ & new_new_n11151__;
  assign new_new_n11154__ = ~new_new_n11152__ & ~new_new_n11153__;
  assign new_new_n11155__ = new_new_n11149__ & ~new_new_n11154__;
  assign new_new_n11156__ = ~new_new_n11149__ & new_new_n11154__;
  assign new_new_n11157__ = ~new_new_n11155__ & ~new_new_n11156__;
  assign new_new_n11158__ = new_new_n11148__ & ~new_new_n11157__;
  assign new_new_n11159__ = ~new_new_n11148__ & new_new_n11157__;
  assign new_new_n11160__ = ~new_new_n11158__ & ~new_new_n11159__;
  assign new_new_n11161__ = new_new_n11139__ & new_new_n11160__;
  assign new_new_n11162__ = ~new_new_n11139__ & ~new_new_n11160__;
  assign new_new_n11163__ = ~new_new_n11161__ & ~new_new_n11162__;
  assign new_new_n11164__ = new_new_n11130__ & ~new_new_n11163__;
  assign new_new_n11165__ = ~new_new_n11130__ & new_new_n11163__;
  assign new_new_n11166__ = ~new_new_n11164__ & ~new_new_n11165__;
  assign new_new_n11167__ = new_new_n11121__ & new_new_n11166__;
  assign new_new_n11168__ = ~new_new_n11121__ & ~new_new_n11166__;
  assign new_new_n11169__ = ~new_new_n11167__ & ~new_new_n11168__;
  assign new_new_n11170__ = ~new_new_n10757__ & new_new_n10781__;
  assign new_new_n11171__ = ~new_new_n10756__ & ~new_new_n11170__;
  assign new_new_n11172__ = ~new_new_n10833__ & ~new_new_n10836__;
  assign new_new_n11173__ = ~new_new_n10832__ & ~new_new_n11172__;
  assign new_new_n11174__ = ~new_new_n10765__ & ~new_new_n10771__;
  assign new_new_n11175__ = ~new_new_n11173__ & ~new_new_n11174__;
  assign new_new_n11176__ = new_new_n11173__ & new_new_n11174__;
  assign new_new_n11177__ = ~new_new_n11175__ & ~new_new_n11176__;
  assign new_new_n11178__ = ~new_new_n10820__ & ~new_new_n10825__;
  assign new_new_n11179__ = new_new_n11177__ & ~new_new_n11178__;
  assign new_new_n11180__ = ~new_new_n11177__ & new_new_n11178__;
  assign new_new_n11181__ = ~new_new_n11179__ & ~new_new_n11180__;
  assign new_new_n11182__ = ~new_new_n10840__ & ~new_new_n10844__;
  assign new_new_n11183__ = ~new_new_n10841__ & ~new_new_n11182__;
  assign new_new_n11184__ = ~new_new_n11181__ & new_new_n11183__;
  assign new_new_n11185__ = new_new_n11181__ & ~new_new_n11183__;
  assign new_new_n11186__ = ~new_new_n11184__ & ~new_new_n11185__;
  assign new_new_n11187__ = ~new_new_n10760__ & ~new_new_n10777__;
  assign new_new_n11188__ = ~new_new_n10776__ & ~new_new_n11187__;
  assign new_new_n11189__ = new_new_n11186__ & new_new_n11188__;
  assign new_new_n11190__ = ~new_new_n11186__ & ~new_new_n11188__;
  assign new_new_n11191__ = ~new_new_n11189__ & ~new_new_n11190__;
  assign new_new_n11192__ = ~new_new_n11171__ & ~new_new_n11191__;
  assign new_new_n11193__ = new_new_n11171__ & new_new_n11191__;
  assign new_new_n11194__ = ~new_new_n11192__ & ~new_new_n11193__;
  assign new_new_n11195__ = ~new_new_n10976__ & new_new_n11007__;
  assign new_new_n11196__ = ~new_new_n10977__ & ~new_new_n11195__;
  assign new_new_n11197__ = new_new_n11194__ & ~new_new_n11196__;
  assign new_new_n11198__ = ~new_new_n11194__ & new_new_n11196__;
  assign new_new_n11199__ = ~new_new_n11197__ & ~new_new_n11198__;
  assign new_new_n11200__ = new_new_n11169__ & new_new_n11199__;
  assign new_new_n11201__ = ~new_new_n11169__ & ~new_new_n11199__;
  assign new_new_n11202__ = ~new_new_n11200__ & ~new_new_n11201__;
  assign new_new_n11203__ = new_new_n11065__ & new_new_n11202__;
  assign new_new_n11204__ = ~new_new_n11065__ & ~new_new_n11202__;
  assign new_new_n11205__ = ~new_new_n11203__ & ~new_new_n11204__;
  assign new_new_n11206__ = ~new_new_n10849__ & ~new_new_n10852__;
  assign new_new_n11207__ = ~new_new_n10848__ & ~new_new_n11206__;
  assign new_new_n11208__ = ~new_new_n10955__ & ~new_new_n10966__;
  assign new_new_n11209__ = ~new_new_n10956__ & ~new_new_n11208__;
  assign new_new_n11210__ = ~new_new_n10807__ & ~new_new_n11209__;
  assign new_new_n11211__ = new_new_n10807__ & new_new_n11209__;
  assign new_new_n11212__ = ~new_new_n11210__ & ~new_new_n11211__;
  assign new_new_n11213__ = ~new_new_n10889__ & ~new_new_n10900__;
  assign new_new_n11214__ = ~new_new_n10890__ & ~new_new_n11213__;
  assign new_new_n11215__ = ~new_new_n11212__ & new_new_n11214__;
  assign new_new_n11216__ = ~new_new_n11211__ & ~new_new_n11214__;
  assign new_new_n11217__ = ~new_new_n11210__ & new_new_n11216__;
  assign new_new_n11218__ = ~new_new_n11215__ & ~new_new_n11217__;
  assign new_new_n11219__ = ~new_new_n10958__ & ~new_new_n10962__;
  assign new_new_n11220__ = ~new_new_n10961__ & ~new_new_n11219__;
  assign new_new_n11221__ = ~new_new_n10946__ & ~new_new_n10950__;
  assign new_new_n11222__ = ~new_new_n10949__ & ~new_new_n11221__;
  assign new_new_n11223__ = ~new_new_n10793__ & ~new_new_n10797__;
  assign new_new_n11224__ = ~new_new_n10796__ & ~new_new_n11223__;
  assign new_new_n11225__ = ~new_new_n11222__ & ~new_new_n11224__;
  assign new_new_n11226__ = new_new_n11222__ & new_new_n11224__;
  assign new_new_n11227__ = ~new_new_n11225__ & ~new_new_n11226__;
  assign new_new_n11228__ = new_new_n11220__ & ~new_new_n11227__;
  assign new_new_n11229__ = ~new_new_n11220__ & new_new_n11227__;
  assign new_new_n11230__ = ~new_new_n11228__ & ~new_new_n11229__;
  assign new_new_n11231__ = ~new_new_n10925__ & ~new_new_n10929__;
  assign new_new_n11232__ = ~new_new_n10928__ & ~new_new_n11231__;
  assign new_new_n11233__ = ~new_new_n10913__ & ~new_new_n10917__;
  assign new_new_n11234__ = ~new_new_n10916__ & ~new_new_n11233__;
  assign new_new_n11235__ = pi06 & pi61;
  assign new_new_n11236__ = new_new_n11234__ & ~new_new_n11235__;
  assign new_new_n11237__ = ~new_new_n11234__ & new_new_n11235__;
  assign new_new_n11238__ = ~new_new_n11236__ & ~new_new_n11237__;
  assign new_new_n11239__ = new_new_n11232__ & new_new_n11238__;
  assign new_new_n11240__ = ~new_new_n11232__ & ~new_new_n11238__;
  assign new_new_n11241__ = ~new_new_n11239__ & ~new_new_n11240__;
  assign new_new_n11242__ = new_new_n11230__ & new_new_n11241__;
  assign new_new_n11243__ = ~new_new_n11230__ & ~new_new_n11241__;
  assign new_new_n11244__ = ~new_new_n11242__ & ~new_new_n11243__;
  assign new_new_n11245__ = ~new_new_n10892__ & ~new_new_n10896__;
  assign new_new_n11246__ = ~new_new_n10895__ & ~new_new_n11245__;
  assign new_new_n11247__ = ~new_new_n10871__ & ~new_new_n10875__;
  assign new_new_n11248__ = ~new_new_n10874__ & ~new_new_n11247__;
  assign new_new_n11249__ = ~new_new_n10880__ & ~new_new_n10884__;
  assign new_new_n11250__ = ~new_new_n10883__ & ~new_new_n11249__;
  assign new_new_n11251__ = ~new_new_n11248__ & ~new_new_n11250__;
  assign new_new_n11252__ = new_new_n11248__ & new_new_n11250__;
  assign new_new_n11253__ = ~new_new_n11251__ & ~new_new_n11252__;
  assign new_new_n11254__ = new_new_n11246__ & ~new_new_n11253__;
  assign new_new_n11255__ = ~new_new_n11246__ & new_new_n11253__;
  assign new_new_n11256__ = ~new_new_n11254__ & ~new_new_n11255__;
  assign new_new_n11257__ = new_new_n11244__ & ~new_new_n11256__;
  assign new_new_n11258__ = ~new_new_n11244__ & new_new_n11256__;
  assign new_new_n11259__ = ~new_new_n11257__ & ~new_new_n11258__;
  assign new_new_n11260__ = ~new_new_n11218__ & ~new_new_n11259__;
  assign new_new_n11261__ = new_new_n11218__ & new_new_n11259__;
  assign new_new_n11262__ = ~new_new_n11260__ & ~new_new_n11261__;
  assign new_new_n11263__ = ~new_new_n11000__ & new_new_n11004__;
  assign new_new_n11264__ = ~new_new_n11001__ & ~new_new_n11263__;
  assign new_new_n11265__ = new_new_n11262__ & ~new_new_n11264__;
  assign new_new_n11266__ = ~new_new_n11262__ & new_new_n11264__;
  assign new_new_n11267__ = ~new_new_n11265__ & ~new_new_n11266__;
  assign new_new_n11268__ = ~new_new_n11207__ & new_new_n11267__;
  assign new_new_n11269__ = new_new_n11207__ & ~new_new_n11267__;
  assign new_new_n11270__ = ~new_new_n11268__ & ~new_new_n11269__;
  assign new_new_n11271__ = ~new_new_n10789__ & ~new_new_n10811__;
  assign new_new_n11272__ = ~new_new_n10788__ & ~new_new_n11271__;
  assign new_new_n11273__ = ~new_new_n10990__ & ~new_new_n10994__;
  assign new_new_n11274__ = ~new_new_n10995__ & ~new_new_n11273__;
  assign new_new_n11275__ = ~new_new_n10923__ & ~new_new_n10933__;
  assign new_new_n11276__ = ~new_new_n10922__ & ~new_new_n11275__;
  assign new_new_n11277__ = ~new_new_n11274__ & new_new_n11276__;
  assign new_new_n11278__ = new_new_n11274__ & ~new_new_n11276__;
  assign new_new_n11279__ = ~new_new_n11277__ & ~new_new_n11278__;
  assign new_new_n11280__ = ~new_new_n10937__ & ~new_new_n10941__;
  assign new_new_n11281__ = ~new_new_n10940__ & ~new_new_n11280__;
  assign new_new_n11282__ = ~new_new_n10904__ & ~new_new_n10908__;
  assign new_new_n11283__ = ~new_new_n10907__ & ~new_new_n11282__;
  assign new_new_n11284__ = ~new_new_n11281__ & ~new_new_n11283__;
  assign new_new_n11285__ = new_new_n11281__ & new_new_n11283__;
  assign new_new_n11286__ = pi20 & pi47;
  assign new_new_n11287__ = pi11 & pi56;
  assign new_new_n11288__ = pi10 & pi57;
  assign new_new_n11289__ = ~new_new_n11287__ & ~new_new_n11288__;
  assign new_new_n11290__ = new_new_n11287__ & new_new_n11288__;
  assign new_new_n11291__ = ~new_new_n11289__ & ~new_new_n11290__;
  assign new_new_n11292__ = new_new_n11286__ & ~new_new_n11291__;
  assign new_new_n11293__ = ~new_new_n11286__ & new_new_n11291__;
  assign new_new_n11294__ = ~new_new_n11292__ & ~new_new_n11293__;
  assign new_new_n11295__ = ~new_new_n11284__ & ~new_new_n11294__;
  assign new_new_n11296__ = ~new_new_n11285__ & ~new_new_n11295__;
  assign new_new_n11297__ = ~new_new_n11284__ & new_new_n11296__;
  assign new_new_n11298__ = ~new_new_n11285__ & new_new_n11295__;
  assign new_new_n11299__ = ~new_new_n11294__ & ~new_new_n11298__;
  assign new_new_n11300__ = ~new_new_n11297__ & ~new_new_n11299__;
  assign new_new_n11301__ = new_new_n11279__ & ~new_new_n11300__;
  assign new_new_n11302__ = ~new_new_n11279__ & new_new_n11300__;
  assign new_new_n11303__ = ~new_new_n11301__ & ~new_new_n11302__;
  assign new_new_n11304__ = ~new_new_n11272__ & new_new_n11303__;
  assign new_new_n11305__ = new_new_n11272__ & ~new_new_n11303__;
  assign new_new_n11306__ = ~new_new_n11304__ & ~new_new_n11305__;
  assign new_new_n11307__ = ~new_new_n10903__ & ~new_new_n10971__;
  assign new_new_n11308__ = ~new_new_n10970__ & ~new_new_n11307__;
  assign new_new_n11309__ = ~new_new_n11306__ & new_new_n11308__;
  assign new_new_n11310__ = new_new_n11306__ & ~new_new_n11308__;
  assign new_new_n11311__ = ~new_new_n11309__ & ~new_new_n11310__;
  assign new_new_n11312__ = new_new_n11270__ & new_new_n11311__;
  assign new_new_n11313__ = ~new_new_n11270__ & ~new_new_n11311__;
  assign new_new_n11314__ = ~new_new_n11312__ & ~new_new_n11313__;
  assign new_new_n11315__ = new_new_n11205__ & new_new_n11314__;
  assign new_new_n11316__ = ~new_new_n11205__ & ~new_new_n11314__;
  assign new_new_n11317__ = ~new_new_n11315__ & ~new_new_n11316__;
  assign new_new_n11318__ = new_new_n11016__ & ~new_new_n11317__;
  assign new_new_n11319__ = ~new_new_n11016__ & new_new_n11317__;
  assign new_new_n11320__ = ~new_new_n11318__ & ~new_new_n11319__;
  assign new_new_n11321__ = new_new_n11063__ & ~new_new_n11320__;
  assign new_new_n11322__ = ~new_new_n11063__ & new_new_n11320__;
  assign po068 = new_new_n11321__ | new_new_n11322__;
  assign new_new_n11324__ = ~new_new_n11196__ & ~new_new_n11202__;
  assign new_new_n11325__ = ~new_new_n11203__ & ~new_new_n11324__;
  assign new_new_n11326__ = ~new_new_n11016__ & ~new_new_n11315__;
  assign new_new_n11327__ = ~new_new_n11316__ & ~new_new_n11326__;
  assign new_new_n11328__ = ~new_new_n11325__ & new_new_n11327__;
  assign new_new_n11329__ = new_new_n11325__ & ~new_new_n11327__;
  assign new_new_n11330__ = ~new_new_n11328__ & ~new_new_n11329__;
  assign new_new_n11331__ = ~new_new_n11269__ & ~new_new_n11311__;
  assign new_new_n11332__ = ~new_new_n11268__ & ~new_new_n11331__;
  assign new_new_n11333__ = ~new_new_n11242__ & ~new_new_n11256__;
  assign new_new_n11334__ = ~new_new_n11243__ & ~new_new_n11333__;
  assign new_new_n11335__ = ~new_new_n11277__ & ~new_new_n11300__;
  assign new_new_n11336__ = ~new_new_n11278__ & ~new_new_n11335__;
  assign new_new_n11337__ = new_new_n11334__ & new_new_n11336__;
  assign new_new_n11338__ = ~new_new_n11334__ & ~new_new_n11336__;
  assign new_new_n11339__ = ~new_new_n11337__ & ~new_new_n11338__;
  assign new_new_n11340__ = ~new_new_n11210__ & ~new_new_n11216__;
  assign new_new_n11341__ = ~new_new_n11339__ & new_new_n11340__;
  assign new_new_n11342__ = ~new_new_n11337__ & ~new_new_n11340__;
  assign new_new_n11343__ = ~new_new_n11338__ & new_new_n11342__;
  assign new_new_n11344__ = ~new_new_n11341__ & ~new_new_n11343__;
  assign new_new_n11345__ = pi26 & pi42;
  assign new_new_n11346__ = pi25 & pi43;
  assign new_new_n11347__ = pi24 & pi44;
  assign new_new_n11348__ = ~new_new_n11346__ & ~new_new_n11347__;
  assign new_new_n11349__ = new_new_n11346__ & new_new_n11347__;
  assign new_new_n11350__ = ~new_new_n11348__ & ~new_new_n11349__;
  assign new_new_n11351__ = new_new_n11345__ & ~new_new_n11350__;
  assign new_new_n11352__ = ~new_new_n11345__ & new_new_n11350__;
  assign new_new_n11353__ = ~new_new_n11351__ & ~new_new_n11352__;
  assign new_new_n11354__ = pi16 & pi52;
  assign new_new_n11355__ = pi15 & pi53;
  assign new_new_n11356__ = pi14 & pi54;
  assign new_new_n11357__ = ~new_new_n11355__ & ~new_new_n11356__;
  assign new_new_n11358__ = new_new_n11355__ & new_new_n11356__;
  assign new_new_n11359__ = ~new_new_n11357__ & ~new_new_n11358__;
  assign new_new_n11360__ = new_new_n11354__ & ~new_new_n11359__;
  assign new_new_n11361__ = ~new_new_n11354__ & new_new_n11359__;
  assign new_new_n11362__ = ~new_new_n11360__ & ~new_new_n11361__;
  assign new_new_n11363__ = new_new_n11353__ & new_new_n11362__;
  assign new_new_n11364__ = ~new_new_n11353__ & ~new_new_n11362__;
  assign new_new_n11365__ = ~new_new_n11363__ & ~new_new_n11364__;
  assign new_new_n11366__ = pi22 & pi46;
  assign new_new_n11367__ = pi20 & pi48;
  assign new_new_n11368__ = ~new_new_n11366__ & ~new_new_n11367__;
  assign new_new_n11369__ = new_new_n11366__ & new_new_n11367__;
  assign new_new_n11370__ = ~new_new_n11368__ & ~new_new_n11369__;
  assign new_new_n11371__ = new_new_n5603__ & ~new_new_n11370__;
  assign new_new_n11372__ = ~new_new_n5603__ & new_new_n11370__;
  assign new_new_n11373__ = ~new_new_n11371__ & ~new_new_n11372__;
  assign new_new_n11374__ = new_new_n11365__ & ~new_new_n11373__;
  assign new_new_n11375__ = ~new_new_n11365__ & new_new_n11373__;
  assign new_new_n11376__ = ~new_new_n11374__ & ~new_new_n11375__;
  assign new_new_n11377__ = pi17 & pi51;
  assign new_new_n11378__ = pi13 & pi55;
  assign new_new_n11379__ = pi12 & pi56;
  assign new_new_n11380__ = ~new_new_n11378__ & ~new_new_n11379__;
  assign new_new_n11381__ = new_new_n11378__ & new_new_n11379__;
  assign new_new_n11382__ = ~new_new_n11380__ & ~new_new_n11381__;
  assign new_new_n11383__ = new_new_n11377__ & ~new_new_n11382__;
  assign new_new_n11384__ = ~new_new_n11377__ & new_new_n11382__;
  assign new_new_n11385__ = ~new_new_n11383__ & ~new_new_n11384__;
  assign new_new_n11386__ = pi32 & pi36;
  assign new_new_n11387__ = pi31 & pi37;
  assign new_new_n11388__ = pi30 & pi38;
  assign new_new_n11389__ = ~new_new_n11387__ & ~new_new_n11388__;
  assign new_new_n11390__ = new_new_n11387__ & new_new_n11388__;
  assign new_new_n11391__ = ~new_new_n11389__ & ~new_new_n11390__;
  assign new_new_n11392__ = new_new_n11386__ & ~new_new_n11391__;
  assign new_new_n11393__ = ~new_new_n11386__ & new_new_n11391__;
  assign new_new_n11394__ = ~new_new_n11392__ & ~new_new_n11393__;
  assign new_new_n11395__ = new_new_n11385__ & new_new_n11394__;
  assign new_new_n11396__ = ~new_new_n11385__ & ~new_new_n11394__;
  assign new_new_n11397__ = ~new_new_n11395__ & ~new_new_n11396__;
  assign new_new_n11398__ = pi33 & pi35;
  assign new_new_n11399__ = pi18 & pi50;
  assign new_new_n11400__ = pi19 & pi49;
  assign new_new_n11401__ = ~new_new_n11399__ & ~new_new_n11400__;
  assign new_new_n11402__ = new_new_n11399__ & new_new_n11400__;
  assign new_new_n11403__ = ~new_new_n11401__ & ~new_new_n11402__;
  assign new_new_n11404__ = new_new_n11398__ & ~new_new_n11403__;
  assign new_new_n11405__ = ~new_new_n11398__ & new_new_n11403__;
  assign new_new_n11406__ = ~new_new_n11404__ & ~new_new_n11405__;
  assign new_new_n11407__ = new_new_n11397__ & ~new_new_n11406__;
  assign new_new_n11408__ = ~new_new_n11397__ & new_new_n11406__;
  assign new_new_n11409__ = ~new_new_n11407__ & ~new_new_n11408__;
  assign new_new_n11410__ = ~new_new_n11376__ & ~new_new_n11409__;
  assign new_new_n11411__ = new_new_n11376__ & new_new_n11409__;
  assign new_new_n11412__ = ~new_new_n11410__ & ~new_new_n11411__;
  assign new_new_n11413__ = pi29 & pi39;
  assign new_new_n11414__ = pi28 & pi40;
  assign new_new_n11415__ = pi27 & pi41;
  assign new_new_n11416__ = ~new_new_n11414__ & ~new_new_n11415__;
  assign new_new_n11417__ = new_new_n11414__ & new_new_n11415__;
  assign new_new_n11418__ = ~new_new_n11416__ & ~new_new_n11417__;
  assign new_new_n11419__ = new_new_n11413__ & ~new_new_n11418__;
  assign new_new_n11420__ = ~new_new_n11413__ & new_new_n11418__;
  assign new_new_n11421__ = ~new_new_n11419__ & ~new_new_n11420__;
  assign new_new_n11422__ = pi21 & pi47;
  assign new_new_n11423__ = pi06 & pi62;
  assign new_new_n11424__ = pi05 & pi63;
  assign new_new_n11425__ = ~new_new_n11423__ & ~new_new_n11424__;
  assign new_new_n11426__ = new_new_n11423__ & new_new_n11424__;
  assign new_new_n11427__ = ~new_new_n11425__ & ~new_new_n11426__;
  assign new_new_n11428__ = new_new_n11422__ & ~new_new_n11427__;
  assign new_new_n11429__ = ~new_new_n11422__ & new_new_n11427__;
  assign new_new_n11430__ = ~new_new_n11428__ & ~new_new_n11429__;
  assign new_new_n11431__ = ~new_new_n11421__ & ~new_new_n11430__;
  assign new_new_n11432__ = new_new_n11421__ & new_new_n11430__;
  assign new_new_n11433__ = ~new_new_n11431__ & ~new_new_n11432__;
  assign new_new_n11434__ = pi11 & pi57;
  assign new_new_n11435__ = pi10 & pi58;
  assign new_new_n11436__ = pi09 & pi59;
  assign new_new_n11437__ = ~new_new_n11435__ & ~new_new_n11436__;
  assign new_new_n11438__ = new_new_n11435__ & new_new_n11436__;
  assign new_new_n11439__ = ~new_new_n11437__ & ~new_new_n11438__;
  assign new_new_n11440__ = new_new_n11434__ & ~new_new_n11439__;
  assign new_new_n11441__ = ~new_new_n11434__ & new_new_n11439__;
  assign new_new_n11442__ = ~new_new_n11440__ & ~new_new_n11441__;
  assign new_new_n11443__ = new_new_n11433__ & ~new_new_n11442__;
  assign new_new_n11444__ = ~new_new_n11433__ & new_new_n11442__;
  assign new_new_n11445__ = ~new_new_n11443__ & ~new_new_n11444__;
  assign new_new_n11446__ = new_new_n11412__ & new_new_n11445__;
  assign new_new_n11447__ = ~new_new_n11412__ & ~new_new_n11445__;
  assign new_new_n11448__ = ~new_new_n11446__ & ~new_new_n11447__;
  assign new_new_n11449__ = new_new_n11344__ & new_new_n11448__;
  assign new_new_n11450__ = ~new_new_n11344__ & ~new_new_n11448__;
  assign new_new_n11451__ = ~new_new_n11449__ & ~new_new_n11450__;
  assign new_new_n11452__ = ~new_new_n11304__ & ~new_new_n11308__;
  assign new_new_n11453__ = ~new_new_n11305__ & ~new_new_n11452__;
  assign new_new_n11454__ = new_new_n11451__ & ~new_new_n11453__;
  assign new_new_n11455__ = ~new_new_n11451__ & new_new_n11453__;
  assign new_new_n11456__ = ~new_new_n11454__ & ~new_new_n11455__;
  assign new_new_n11457__ = new_new_n11332__ & new_new_n11456__;
  assign new_new_n11458__ = ~new_new_n11332__ & ~new_new_n11456__;
  assign new_new_n11459__ = ~new_new_n11457__ & ~new_new_n11458__;
  assign new_new_n11460__ = ~new_new_n11169__ & ~new_new_n11193__;
  assign new_new_n11461__ = ~new_new_n11192__ & ~new_new_n11460__;
  assign new_new_n11462__ = new_new_n11459__ & ~new_new_n11461__;
  assign new_new_n11463__ = ~new_new_n11459__ & new_new_n11461__;
  assign new_new_n11464__ = ~new_new_n11462__ & ~new_new_n11463__;
  assign new_new_n11465__ = ~new_new_n11062__ & ~new_new_n11320__;
  assign new_new_n11466__ = ~new_new_n11061__ & ~new_new_n11465__;
  assign new_new_n11467__ = ~new_new_n11464__ & ~new_new_n11466__;
  assign new_new_n11468__ = new_new_n11464__ & new_new_n11466__;
  assign new_new_n11469__ = ~new_new_n11467__ & ~new_new_n11468__;
  assign new_new_n11470__ = ~new_new_n11260__ & ~new_new_n11264__;
  assign new_new_n11471__ = ~new_new_n11261__ & ~new_new_n11470__;
  assign new_new_n11472__ = ~new_new_n11246__ & ~new_new_n11252__;
  assign new_new_n11473__ = ~new_new_n11251__ & ~new_new_n11472__;
  assign new_new_n11474__ = ~new_new_n11083__ & ~new_new_n11157__;
  assign new_new_n11475__ = ~new_new_n11084__ & ~new_new_n11474__;
  assign new_new_n11476__ = new_new_n11296__ & new_new_n11475__;
  assign new_new_n11477__ = ~new_new_n11296__ & ~new_new_n11475__;
  assign new_new_n11478__ = ~new_new_n11476__ & ~new_new_n11477__;
  assign new_new_n11479__ = new_new_n11473__ & ~new_new_n11478__;
  assign new_new_n11480__ = ~new_new_n11473__ & new_new_n11478__;
  assign new_new_n11481__ = ~new_new_n11479__ & ~new_new_n11480__;
  assign new_new_n11482__ = new_new_n11085__ & new_new_n11157__;
  assign new_new_n11483__ = ~new_new_n11085__ & ~new_new_n11157__;
  assign new_new_n11484__ = ~new_new_n11482__ & ~new_new_n11483__;
  assign new_new_n11485__ = new_new_n11118__ & ~new_new_n11484__;
  assign new_new_n11486__ = ~new_new_n11118__ & new_new_n11484__;
  assign new_new_n11487__ = ~new_new_n11130__ & ~new_new_n11148__;
  assign new_new_n11488__ = new_new_n11130__ & new_new_n11148__;
  assign new_new_n11489__ = ~new_new_n11487__ & ~new_new_n11488__;
  assign new_new_n11490__ = new_new_n11139__ & new_new_n11489__;
  assign new_new_n11491__ = ~new_new_n11139__ & ~new_new_n11489__;
  assign new_new_n11492__ = ~new_new_n11490__ & ~new_new_n11491__;
  assign new_new_n11493__ = ~new_new_n11486__ & ~new_new_n11492__;
  assign new_new_n11494__ = ~new_new_n11485__ & ~new_new_n11493__;
  assign new_new_n11495__ = new_new_n11481__ & new_new_n11494__;
  assign new_new_n11496__ = ~new_new_n11481__ & ~new_new_n11494__;
  assign new_new_n11497__ = ~new_new_n11495__ & ~new_new_n11496__;
  assign new_new_n11498__ = ~new_new_n11220__ & ~new_new_n11226__;
  assign new_new_n11499__ = ~new_new_n11225__ & ~new_new_n11498__;
  assign new_new_n11500__ = pi08 & pi60;
  assign new_new_n11501__ = pi07 & pi61;
  assign new_new_n11502__ = ~new_new_n11500__ & ~new_new_n11501__;
  assign new_new_n11503__ = new_new_n11500__ & new_new_n11501__;
  assign new_new_n11504__ = ~new_new_n11502__ & ~new_new_n11503__;
  assign new_new_n11505__ = ~new_new_n11124__ & ~new_new_n11128__;
  assign new_new_n11506__ = ~new_new_n11504__ & new_new_n11505__;
  assign new_new_n11507__ = new_new_n11504__ & ~new_new_n11505__;
  assign new_new_n11508__ = ~new_new_n11506__ & ~new_new_n11507__;
  assign new_new_n11509__ = ~new_new_n11234__ & ~new_new_n11235__;
  assign new_new_n11510__ = new_new_n11234__ & new_new_n11235__;
  assign new_new_n11511__ = ~new_new_n11232__ & ~new_new_n11510__;
  assign new_new_n11512__ = ~new_new_n11509__ & ~new_new_n11511__;
  assign new_new_n11513__ = ~new_new_n11508__ & new_new_n11512__;
  assign new_new_n11514__ = new_new_n11508__ & ~new_new_n11512__;
  assign new_new_n11515__ = ~new_new_n11513__ & ~new_new_n11514__;
  assign new_new_n11516__ = new_new_n11499__ & ~new_new_n11515__;
  assign new_new_n11517__ = ~new_new_n11499__ & new_new_n11515__;
  assign new_new_n11518__ = ~new_new_n11516__ & ~new_new_n11517__;
  assign new_new_n11519__ = new_new_n11497__ & ~new_new_n11518__;
  assign new_new_n11520__ = ~new_new_n11497__ & new_new_n11518__;
  assign new_new_n11521__ = ~new_new_n11519__ & ~new_new_n11520__;
  assign new_new_n11522__ = ~new_new_n11471__ & new_new_n11521__;
  assign new_new_n11523__ = new_new_n11471__ & ~new_new_n11521__;
  assign new_new_n11524__ = ~new_new_n11522__ & ~new_new_n11523__;
  assign new_new_n11525__ = ~new_new_n11104__ & ~new_new_n11115__;
  assign new_new_n11526__ = ~new_new_n11105__ & ~new_new_n11525__;
  assign new_new_n11527__ = ~new_new_n11139__ & ~new_new_n11488__;
  assign new_new_n11528__ = ~new_new_n11487__ & ~new_new_n11527__;
  assign new_new_n11529__ = new_new_n11526__ & ~new_new_n11528__;
  assign new_new_n11530__ = ~new_new_n11526__ & new_new_n11528__;
  assign new_new_n11531__ = ~new_new_n11529__ & ~new_new_n11530__;
  assign new_new_n11532__ = ~new_new_n11131__ & ~new_new_n11135__;
  assign new_new_n11533__ = ~new_new_n11134__ & ~new_new_n11532__;
  assign new_new_n11534__ = ~new_new_n11086__ & ~new_new_n11090__;
  assign new_new_n11535__ = ~new_new_n11089__ & ~new_new_n11534__;
  assign new_new_n11536__ = ~new_new_n11107__ & ~new_new_n11111__;
  assign new_new_n11537__ = ~new_new_n11110__ & ~new_new_n11536__;
  assign new_new_n11538__ = ~new_new_n11535__ & ~new_new_n11537__;
  assign new_new_n11539__ = new_new_n11535__ & new_new_n11537__;
  assign new_new_n11540__ = ~new_new_n11538__ & ~new_new_n11539__;
  assign new_new_n11541__ = new_new_n11533__ & ~new_new_n11540__;
  assign new_new_n11542__ = ~new_new_n11533__ & new_new_n11540__;
  assign new_new_n11543__ = ~new_new_n11541__ & ~new_new_n11542__;
  assign new_new_n11544__ = new_new_n11531__ & ~new_new_n11543__;
  assign new_new_n11545__ = ~new_new_n11531__ & new_new_n11543__;
  assign new_new_n11546__ = ~new_new_n11544__ & ~new_new_n11545__;
  assign new_new_n11547__ = ~new_new_n11185__ & ~new_new_n11188__;
  assign new_new_n11548__ = ~new_new_n11184__ & ~new_new_n11547__;
  assign new_new_n11549__ = ~new_new_n11175__ & ~new_new_n11179__;
  assign new_new_n11550__ = ~new_new_n11095__ & ~new_new_n11099__;
  assign new_new_n11551__ = ~new_new_n11098__ & ~new_new_n11550__;
  assign new_new_n11552__ = ~new_new_n11140__ & ~new_new_n11144__;
  assign new_new_n11553__ = ~new_new_n11143__ & ~new_new_n11552__;
  assign new_new_n11554__ = ~new_new_n11074__ & ~new_new_n11078__;
  assign new_new_n11555__ = ~new_new_n11077__ & ~new_new_n11554__;
  assign new_new_n11556__ = new_new_n11553__ & new_new_n11555__;
  assign new_new_n11557__ = ~new_new_n11553__ & ~new_new_n11555__;
  assign new_new_n11558__ = ~new_new_n11556__ & ~new_new_n11557__;
  assign new_new_n11559__ = new_new_n11551__ & ~new_new_n11558__;
  assign new_new_n11560__ = ~new_new_n11551__ & new_new_n11558__;
  assign new_new_n11561__ = ~new_new_n11559__ & ~new_new_n11560__;
  assign new_new_n11562__ = new_new_n11549__ & ~new_new_n11561__;
  assign new_new_n11563__ = ~new_new_n11549__ & new_new_n11561__;
  assign new_new_n11564__ = ~new_new_n11562__ & ~new_new_n11563__;
  assign new_new_n11565__ = ~new_new_n11149__ & ~new_new_n11153__;
  assign new_new_n11566__ = ~new_new_n11152__ & ~new_new_n11565__;
  assign new_new_n11567__ = ~new_new_n11066__ & ~new_new_n11069__;
  assign new_new_n11568__ = new_new_n11068__ & ~new_new_n11567__;
  assign new_new_n11569__ = ~new_new_n11566__ & ~new_new_n11568__;
  assign new_new_n11570__ = new_new_n11566__ & new_new_n11568__;
  assign new_new_n11571__ = ~new_new_n11569__ & ~new_new_n11570__;
  assign new_new_n11572__ = ~new_new_n11286__ & ~new_new_n11290__;
  assign new_new_n11573__ = ~new_new_n11289__ & ~new_new_n11572__;
  assign new_new_n11574__ = new_new_n11571__ & ~new_new_n11573__;
  assign new_new_n11575__ = ~new_new_n11571__ & new_new_n11573__;
  assign new_new_n11576__ = ~new_new_n11574__ & ~new_new_n11575__;
  assign new_new_n11577__ = new_new_n11564__ & new_new_n11576__;
  assign new_new_n11578__ = ~new_new_n11564__ & ~new_new_n11576__;
  assign new_new_n11579__ = ~new_new_n11577__ & ~new_new_n11578__;
  assign new_new_n11580__ = ~new_new_n11548__ & new_new_n11579__;
  assign new_new_n11581__ = new_new_n11548__ & ~new_new_n11579__;
  assign new_new_n11582__ = ~new_new_n11580__ & ~new_new_n11581__;
  assign new_new_n11583__ = new_new_n11546__ & new_new_n11582__;
  assign new_new_n11584__ = ~new_new_n11546__ & ~new_new_n11582__;
  assign new_new_n11585__ = ~new_new_n11583__ & ~new_new_n11584__;
  assign new_new_n11586__ = new_new_n11524__ & ~new_new_n11585__;
  assign new_new_n11587__ = ~new_new_n11524__ & new_new_n11585__;
  assign new_new_n11588__ = ~new_new_n11586__ & ~new_new_n11587__;
  assign new_new_n11589__ = new_new_n11469__ & ~new_new_n11588__;
  assign new_new_n11590__ = ~new_new_n11469__ & new_new_n11588__;
  assign new_new_n11591__ = ~new_new_n11589__ & ~new_new_n11590__;
  assign new_new_n11592__ = new_new_n11330__ & new_new_n11591__;
  assign new_new_n11593__ = ~new_new_n11330__ & ~new_new_n11591__;
  assign po069 = ~new_new_n11592__ & ~new_new_n11593__;
  assign new_new_n11595__ = ~new_new_n11329__ & new_new_n11588__;
  assign new_new_n11596__ = ~new_new_n11328__ & ~new_new_n11595__;
  assign new_new_n11597__ = new_new_n11467__ & new_new_n11596__;
  assign new_new_n11598__ = new_new_n11329__ & ~new_new_n11588__;
  assign new_new_n11599__ = new_new_n11328__ & new_new_n11588__;
  assign new_new_n11600__ = ~new_new_n11598__ & ~new_new_n11599__;
  assign new_new_n11601__ = new_new_n11469__ & new_new_n11600__;
  assign new_new_n11602__ = ~new_new_n11457__ & ~new_new_n11461__;
  assign new_new_n11603__ = ~new_new_n11458__ & ~new_new_n11602__;
  assign new_new_n11604__ = ~new_new_n11363__ & ~new_new_n11373__;
  assign new_new_n11605__ = ~new_new_n11364__ & ~new_new_n11604__;
  assign new_new_n11606__ = ~new_new_n11395__ & ~new_new_n11406__;
  assign new_new_n11607__ = ~new_new_n11396__ & ~new_new_n11606__;
  assign new_new_n11608__ = new_new_n11605__ & new_new_n11607__;
  assign new_new_n11609__ = ~new_new_n11605__ & ~new_new_n11607__;
  assign new_new_n11610__ = ~new_new_n11608__ & ~new_new_n11609__;
  assign new_new_n11611__ = new_new_n11499__ & ~new_new_n11514__;
  assign new_new_n11612__ = ~new_new_n11513__ & ~new_new_n11611__;
  assign new_new_n11613__ = new_new_n11610__ & ~new_new_n11612__;
  assign new_new_n11614__ = ~new_new_n11610__ & new_new_n11612__;
  assign new_new_n11615__ = ~new_new_n11613__ & ~new_new_n11614__;
  assign new_new_n11616__ = ~new_new_n11432__ & ~new_new_n11442__;
  assign new_new_n11617__ = ~new_new_n11431__ & ~new_new_n11616__;
  assign new_new_n11618__ = ~new_new_n11434__ & ~new_new_n11438__;
  assign new_new_n11619__ = ~new_new_n11437__ & ~new_new_n11618__;
  assign new_new_n11620__ = ~new_new_n5603__ & ~new_new_n11369__;
  assign new_new_n11621__ = ~new_new_n11368__ & ~new_new_n11620__;
  assign new_new_n11622__ = ~new_new_n11619__ & ~new_new_n11621__;
  assign new_new_n11623__ = new_new_n11619__ & new_new_n11621__;
  assign new_new_n11624__ = ~new_new_n11622__ & ~new_new_n11623__;
  assign new_new_n11625__ = new_new_n11617__ & ~new_new_n11624__;
  assign new_new_n11626__ = ~new_new_n11617__ & new_new_n11624__;
  assign new_new_n11627__ = ~new_new_n11625__ & ~new_new_n11626__;
  assign new_new_n11628__ = ~new_new_n11422__ & ~new_new_n11426__;
  assign new_new_n11629__ = ~new_new_n11425__ & ~new_new_n11628__;
  assign new_new_n11630__ = ~new_new_n11398__ & ~new_new_n11402__;
  assign new_new_n11631__ = ~new_new_n11401__ & ~new_new_n11630__;
  assign new_new_n11632__ = ~new_new_n11354__ & ~new_new_n11358__;
  assign new_new_n11633__ = ~new_new_n11357__ & ~new_new_n11632__;
  assign new_new_n11634__ = ~new_new_n11631__ & ~new_new_n11633__;
  assign new_new_n11635__ = new_new_n11631__ & new_new_n11633__;
  assign new_new_n11636__ = ~new_new_n11634__ & ~new_new_n11635__;
  assign new_new_n11637__ = ~new_new_n11386__ & ~new_new_n11390__;
  assign new_new_n11638__ = ~new_new_n11389__ & ~new_new_n11637__;
  assign new_new_n11639__ = ~new_new_n11636__ & new_new_n11638__;
  assign new_new_n11640__ = ~new_new_n11635__ & ~new_new_n11638__;
  assign new_new_n11641__ = ~new_new_n11634__ & new_new_n11640__;
  assign new_new_n11642__ = ~new_new_n11639__ & ~new_new_n11641__;
  assign new_new_n11643__ = new_new_n11629__ & ~new_new_n11642__;
  assign new_new_n11644__ = ~new_new_n11629__ & new_new_n11642__;
  assign new_new_n11645__ = ~new_new_n11643__ & ~new_new_n11644__;
  assign new_new_n11646__ = new_new_n11627__ & new_new_n11645__;
  assign new_new_n11647__ = ~new_new_n11627__ & ~new_new_n11645__;
  assign new_new_n11648__ = ~new_new_n11646__ & ~new_new_n11647__;
  assign new_new_n11649__ = ~new_new_n11615__ & ~new_new_n11648__;
  assign new_new_n11650__ = new_new_n11615__ & new_new_n11648__;
  assign new_new_n11651__ = ~new_new_n11649__ & ~new_new_n11650__;
  assign new_new_n11652__ = ~new_new_n11338__ & ~new_new_n11342__;
  assign new_new_n11653__ = new_new_n11651__ & new_new_n11652__;
  assign new_new_n11654__ = ~new_new_n11651__ & ~new_new_n11652__;
  assign new_new_n11655__ = ~new_new_n11653__ & ~new_new_n11654__;
  assign new_new_n11656__ = new_new_n11548__ & new_new_n11579__;
  assign new_new_n11657__ = ~new_new_n11546__ & ~new_new_n11656__;
  assign new_new_n11658__ = ~new_new_n11548__ & ~new_new_n11579__;
  assign new_new_n11659__ = ~new_new_n11657__ & ~new_new_n11658__;
  assign new_new_n11660__ = new_new_n11655__ & new_new_n11659__;
  assign new_new_n11661__ = ~new_new_n11655__ & ~new_new_n11659__;
  assign new_new_n11662__ = ~new_new_n11660__ & ~new_new_n11661__;
  assign new_new_n11663__ = ~new_new_n11533__ & ~new_new_n11539__;
  assign new_new_n11664__ = ~new_new_n11538__ & ~new_new_n11663__;
  assign new_new_n11665__ = ~new_new_n11551__ & ~new_new_n11556__;
  assign new_new_n11666__ = ~new_new_n11557__ & ~new_new_n11665__;
  assign new_new_n11667__ = new_new_n11664__ & new_new_n11666__;
  assign new_new_n11668__ = ~new_new_n11664__ & ~new_new_n11666__;
  assign new_new_n11669__ = ~new_new_n11667__ & ~new_new_n11668__;
  assign new_new_n11670__ = ~new_new_n11377__ & ~new_new_n11381__;
  assign new_new_n11671__ = ~new_new_n11380__ & ~new_new_n11670__;
  assign new_new_n11672__ = ~new_new_n11413__ & ~new_new_n11417__;
  assign new_new_n11673__ = ~new_new_n11416__ & ~new_new_n11672__;
  assign new_new_n11674__ = ~new_new_n11345__ & ~new_new_n11349__;
  assign new_new_n11675__ = ~new_new_n11348__ & ~new_new_n11674__;
  assign new_new_n11676__ = ~new_new_n11673__ & ~new_new_n11675__;
  assign new_new_n11677__ = new_new_n11673__ & new_new_n11675__;
  assign new_new_n11678__ = ~new_new_n11676__ & ~new_new_n11677__;
  assign new_new_n11679__ = new_new_n11671__ & ~new_new_n11678__;
  assign new_new_n11680__ = ~new_new_n11671__ & new_new_n11678__;
  assign new_new_n11681__ = ~new_new_n11679__ & ~new_new_n11680__;
  assign new_new_n11682__ = new_new_n11669__ & new_new_n11681__;
  assign new_new_n11683__ = ~new_new_n11669__ & ~new_new_n11681__;
  assign new_new_n11684__ = ~new_new_n11682__ & ~new_new_n11683__;
  assign new_new_n11685__ = ~new_new_n11571__ & ~new_new_n11573__;
  assign new_new_n11686__ = new_new_n11571__ & new_new_n11573__;
  assign new_new_n11687__ = ~new_new_n11685__ & ~new_new_n11686__;
  assign new_new_n11688__ = ~new_new_n11563__ & new_new_n11687__;
  assign new_new_n11689__ = ~new_new_n11562__ & ~new_new_n11688__;
  assign new_new_n11690__ = new_new_n11684__ & new_new_n11689__;
  assign new_new_n11691__ = ~new_new_n11684__ & ~new_new_n11689__;
  assign new_new_n11692__ = ~new_new_n11690__ & ~new_new_n11691__;
  assign new_new_n11693__ = ~new_new_n11411__ & ~new_new_n11445__;
  assign new_new_n11694__ = ~new_new_n11410__ & ~new_new_n11693__;
  assign new_new_n11695__ = new_new_n11692__ & ~new_new_n11694__;
  assign new_new_n11696__ = ~new_new_n11692__ & new_new_n11694__;
  assign new_new_n11697__ = ~new_new_n11695__ & ~new_new_n11696__;
  assign new_new_n11698__ = new_new_n11662__ & ~new_new_n11697__;
  assign new_new_n11699__ = ~new_new_n11662__ & new_new_n11697__;
  assign new_new_n11700__ = ~new_new_n11698__ & ~new_new_n11699__;
  assign new_new_n11701__ = new_new_n11603__ & ~new_new_n11700__;
  assign new_new_n11702__ = ~new_new_n11603__ & new_new_n11700__;
  assign new_new_n11703__ = ~new_new_n11701__ & ~new_new_n11702__;
  assign new_new_n11704__ = ~new_new_n11495__ & ~new_new_n11518__;
  assign new_new_n11705__ = ~new_new_n11496__ & ~new_new_n11704__;
  assign new_new_n11706__ = ~new_new_n11473__ & ~new_new_n11477__;
  assign new_new_n11707__ = ~new_new_n11476__ & ~new_new_n11706__;
  assign new_new_n11708__ = pi10 & pi59;
  assign new_new_n11709__ = pi08 & pi61;
  assign new_new_n11710__ = pi09 & pi60;
  assign new_new_n11711__ = ~new_new_n11709__ & ~new_new_n11710__;
  assign new_new_n11712__ = new_new_n11709__ & new_new_n11710__;
  assign new_new_n11713__ = ~new_new_n11711__ & ~new_new_n11712__;
  assign new_new_n11714__ = new_new_n11708__ & ~new_new_n11713__;
  assign new_new_n11715__ = ~new_new_n11708__ & new_new_n11713__;
  assign new_new_n11716__ = ~new_new_n11714__ & ~new_new_n11715__;
  assign new_new_n11717__ = pi27 & pi42;
  assign new_new_n11718__ = pi26 & pi43;
  assign new_new_n11719__ = pi06 & pi63;
  assign new_new_n11720__ = ~new_new_n11718__ & ~new_new_n11719__;
  assign new_new_n11721__ = new_new_n11718__ & new_new_n11719__;
  assign new_new_n11722__ = ~new_new_n11720__ & ~new_new_n11721__;
  assign new_new_n11723__ = new_new_n11717__ & ~new_new_n11722__;
  assign new_new_n11724__ = ~new_new_n11717__ & new_new_n11722__;
  assign new_new_n11725__ = ~new_new_n11723__ & ~new_new_n11724__;
  assign new_new_n11726__ = new_new_n11716__ & new_new_n11725__;
  assign new_new_n11727__ = ~new_new_n11716__ & ~new_new_n11725__;
  assign new_new_n11728__ = ~new_new_n11726__ & ~new_new_n11727__;
  assign new_new_n11729__ = pi25 & pi44;
  assign new_new_n11730__ = pi24 & pi45;
  assign new_new_n11731__ = pi23 & pi46;
  assign new_new_n11732__ = ~new_new_n11730__ & ~new_new_n11731__;
  assign new_new_n11733__ = new_new_n11730__ & new_new_n11731__;
  assign new_new_n11734__ = ~new_new_n11732__ & ~new_new_n11733__;
  assign new_new_n11735__ = new_new_n11729__ & ~new_new_n11734__;
  assign new_new_n11736__ = ~new_new_n11729__ & new_new_n11734__;
  assign new_new_n11737__ = ~new_new_n11735__ & ~new_new_n11736__;
  assign new_new_n11738__ = ~new_new_n11728__ & new_new_n11737__;
  assign new_new_n11739__ = new_new_n11728__ & ~new_new_n11737__;
  assign new_new_n11740__ = ~new_new_n11738__ & ~new_new_n11739__;
  assign new_new_n11741__ = new_new_n11707__ & new_new_n11740__;
  assign new_new_n11742__ = ~new_new_n11707__ & ~new_new_n11740__;
  assign new_new_n11743__ = ~new_new_n11741__ & ~new_new_n11742__;
  assign new_new_n11744__ = ~new_new_n11503__ & ~new_new_n11505__;
  assign new_new_n11745__ = ~new_new_n11502__ & ~new_new_n11744__;
  assign new_new_n11746__ = pi22 & pi47;
  assign new_new_n11747__ = pi21 & pi48;
  assign new_new_n11748__ = pi14 & pi55;
  assign new_new_n11749__ = ~new_new_n11747__ & ~new_new_n11748__;
  assign new_new_n11750__ = new_new_n11747__ & new_new_n11748__;
  assign new_new_n11751__ = ~new_new_n11749__ & ~new_new_n11750__;
  assign new_new_n11752__ = new_new_n11746__ & ~new_new_n11751__;
  assign new_new_n11753__ = ~new_new_n11746__ & new_new_n11751__;
  assign new_new_n11754__ = ~new_new_n11752__ & ~new_new_n11753__;
  assign new_new_n11755__ = ~new_new_n11745__ & new_new_n11754__;
  assign new_new_n11756__ = new_new_n11745__ & ~new_new_n11754__;
  assign new_new_n11757__ = ~new_new_n11755__ & ~new_new_n11756__;
  assign new_new_n11758__ = pi13 & pi56;
  assign new_new_n11759__ = pi12 & pi57;
  assign new_new_n11760__ = pi11 & pi58;
  assign new_new_n11761__ = ~new_new_n11759__ & ~new_new_n11760__;
  assign new_new_n11762__ = new_new_n11759__ & new_new_n11760__;
  assign new_new_n11763__ = ~new_new_n11761__ & ~new_new_n11762__;
  assign new_new_n11764__ = new_new_n11758__ & ~new_new_n11763__;
  assign new_new_n11765__ = ~new_new_n11758__ & new_new_n11763__;
  assign new_new_n11766__ = ~new_new_n11764__ & ~new_new_n11765__;
  assign new_new_n11767__ = new_new_n11757__ & ~new_new_n11766__;
  assign new_new_n11768__ = ~new_new_n11757__ & new_new_n11766__;
  assign new_new_n11769__ = ~new_new_n11767__ & ~new_new_n11768__;
  assign new_new_n11770__ = new_new_n11743__ & ~new_new_n11769__;
  assign new_new_n11771__ = ~new_new_n11743__ & new_new_n11769__;
  assign new_new_n11772__ = ~new_new_n11770__ & ~new_new_n11771__;
  assign new_new_n11773__ = ~new_new_n11705__ & ~new_new_n11772__;
  assign new_new_n11774__ = new_new_n11705__ & new_new_n11772__;
  assign new_new_n11775__ = ~new_new_n11773__ & ~new_new_n11774__;
  assign new_new_n11776__ = pi30 & pi39;
  assign new_new_n11777__ = pi28 & pi41;
  assign new_new_n11778__ = pi29 & pi40;
  assign new_new_n11779__ = ~new_new_n11777__ & ~new_new_n11778__;
  assign new_new_n11780__ = new_new_n11777__ & new_new_n11778__;
  assign new_new_n11781__ = ~new_new_n11779__ & ~new_new_n11780__;
  assign new_new_n11782__ = new_new_n11776__ & ~new_new_n11781__;
  assign new_new_n11783__ = ~new_new_n11776__ & new_new_n11781__;
  assign new_new_n11784__ = ~new_new_n11782__ & ~new_new_n11783__;
  assign new_new_n11785__ = pi19 & pi50;
  assign new_new_n11786__ = pi18 & pi51;
  assign new_new_n11787__ = pi17 & pi52;
  assign new_new_n11788__ = ~new_new_n11786__ & ~new_new_n11787__;
  assign new_new_n11789__ = new_new_n11786__ & new_new_n11787__;
  assign new_new_n11790__ = ~new_new_n11788__ & ~new_new_n11789__;
  assign new_new_n11791__ = new_new_n11785__ & ~new_new_n11790__;
  assign new_new_n11792__ = ~new_new_n11785__ & new_new_n11790__;
  assign new_new_n11793__ = ~new_new_n11791__ & ~new_new_n11792__;
  assign new_new_n11794__ = new_new_n11784__ & new_new_n11793__;
  assign new_new_n11795__ = ~new_new_n11784__ & ~new_new_n11793__;
  assign new_new_n11796__ = ~new_new_n11794__ & ~new_new_n11795__;
  assign new_new_n11797__ = ~new_new_n11570__ & ~new_new_n11573__;
  assign new_new_n11798__ = ~new_new_n11569__ & ~new_new_n11797__;
  assign new_new_n11799__ = new_new_n11796__ & ~new_new_n11798__;
  assign new_new_n11800__ = ~new_new_n11796__ & new_new_n11798__;
  assign new_new_n11801__ = ~new_new_n11799__ & ~new_new_n11800__;
  assign new_new_n11802__ = new_new_n11526__ & new_new_n11543__;
  assign new_new_n11803__ = ~new_new_n11528__ & ~new_new_n11802__;
  assign new_new_n11804__ = ~new_new_n11526__ & ~new_new_n11543__;
  assign new_new_n11805__ = ~new_new_n11803__ & ~new_new_n11804__;
  assign new_new_n11806__ = ~new_new_n11801__ & ~new_new_n11805__;
  assign new_new_n11807__ = new_new_n11801__ & new_new_n11805__;
  assign new_new_n11808__ = ~new_new_n11806__ & ~new_new_n11807__;
  assign new_new_n11809__ = pi07 & pi62;
  assign new_new_n11810__ = ~pi34 & pi35;
  assign new_new_n11811__ = ~new_new_n11809__ & new_new_n11810__;
  assign new_new_n11812__ = new_new_n11809__ & ~new_new_n11810__;
  assign new_new_n11813__ = ~new_new_n11811__ & ~new_new_n11812__;
  assign new_new_n11814__ = pi33 & pi36;
  assign new_new_n11815__ = pi31 & pi38;
  assign new_new_n11816__ = pi32 & pi37;
  assign new_new_n11817__ = ~new_new_n11815__ & ~new_new_n11816__;
  assign new_new_n11818__ = new_new_n11815__ & new_new_n11816__;
  assign new_new_n11819__ = ~new_new_n11817__ & ~new_new_n11818__;
  assign new_new_n11820__ = new_new_n11814__ & ~new_new_n11819__;
  assign new_new_n11821__ = ~new_new_n11814__ & new_new_n11819__;
  assign new_new_n11822__ = ~new_new_n11820__ & ~new_new_n11821__;
  assign new_new_n11823__ = pi20 & pi49;
  assign new_new_n11824__ = pi15 & pi54;
  assign new_new_n11825__ = pi16 & pi53;
  assign new_new_n11826__ = ~new_new_n11824__ & ~new_new_n11825__;
  assign new_new_n11827__ = new_new_n11824__ & new_new_n11825__;
  assign new_new_n11828__ = ~new_new_n11826__ & ~new_new_n11827__;
  assign new_new_n11829__ = new_new_n11823__ & ~new_new_n11828__;
  assign new_new_n11830__ = ~new_new_n11823__ & new_new_n11828__;
  assign new_new_n11831__ = ~new_new_n11829__ & ~new_new_n11830__;
  assign new_new_n11832__ = new_new_n11822__ & new_new_n11831__;
  assign new_new_n11833__ = ~new_new_n11822__ & ~new_new_n11831__;
  assign new_new_n11834__ = ~new_new_n11832__ & ~new_new_n11833__;
  assign new_new_n11835__ = new_new_n11813__ & new_new_n11834__;
  assign new_new_n11836__ = ~new_new_n11813__ & ~new_new_n11834__;
  assign new_new_n11837__ = ~new_new_n11835__ & ~new_new_n11836__;
  assign new_new_n11838__ = new_new_n11808__ & ~new_new_n11837__;
  assign new_new_n11839__ = ~new_new_n11808__ & new_new_n11837__;
  assign new_new_n11840__ = ~new_new_n11838__ & ~new_new_n11839__;
  assign new_new_n11841__ = new_new_n11775__ & ~new_new_n11840__;
  assign new_new_n11842__ = ~new_new_n11775__ & new_new_n11840__;
  assign new_new_n11843__ = ~new_new_n11841__ & ~new_new_n11842__;
  assign new_new_n11844__ = ~new_new_n11522__ & ~new_new_n11585__;
  assign new_new_n11845__ = ~new_new_n11523__ & ~new_new_n11844__;
  assign new_new_n11846__ = new_new_n11843__ & ~new_new_n11845__;
  assign new_new_n11847__ = ~new_new_n11843__ & new_new_n11845__;
  assign new_new_n11848__ = ~new_new_n11846__ & ~new_new_n11847__;
  assign new_new_n11849__ = ~new_new_n11449__ & ~new_new_n11453__;
  assign new_new_n11850__ = ~new_new_n11450__ & ~new_new_n11849__;
  assign new_new_n11851__ = new_new_n11848__ & ~new_new_n11850__;
  assign new_new_n11852__ = ~new_new_n11848__ & new_new_n11850__;
  assign new_new_n11853__ = ~new_new_n11851__ & ~new_new_n11852__;
  assign new_new_n11854__ = new_new_n11703__ & ~new_new_n11853__;
  assign new_new_n11855__ = ~new_new_n11703__ & new_new_n11853__;
  assign new_new_n11856__ = ~new_new_n11854__ & ~new_new_n11855__;
  assign new_new_n11857__ = new_new_n11468__ & ~new_new_n11596__;
  assign new_new_n11858__ = ~new_new_n11597__ & ~new_new_n11856__;
  assign new_new_n11859__ = ~new_new_n11857__ & new_new_n11858__;
  assign new_new_n11860__ = ~new_new_n11601__ & new_new_n11859__;
  assign new_new_n11861__ = new_new_n11328__ & new_new_n11467__;
  assign new_new_n11862__ = new_new_n11327__ & new_new_n11467__;
  assign new_new_n11863__ = ~new_new_n11327__ & ~new_new_n11467__;
  assign new_new_n11864__ = ~new_new_n11325__ & ~new_new_n11468__;
  assign new_new_n11865__ = ~new_new_n11863__ & new_new_n11864__;
  assign new_new_n11866__ = ~new_new_n11862__ & ~new_new_n11865__;
  assign new_new_n11867__ = new_new_n11588__ & ~new_new_n11866__;
  assign new_new_n11868__ = ~new_new_n11328__ & new_new_n11468__;
  assign new_new_n11869__ = new_new_n11329__ & ~new_new_n11467__;
  assign new_new_n11870__ = ~new_new_n11868__ & ~new_new_n11869__;
  assign new_new_n11871__ = ~new_new_n11588__ & ~new_new_n11870__;
  assign new_new_n11872__ = new_new_n11329__ & new_new_n11468__;
  assign new_new_n11873__ = new_new_n11856__ & ~new_new_n11861__;
  assign new_new_n11874__ = ~new_new_n11872__ & new_new_n11873__;
  assign new_new_n11875__ = ~new_new_n11871__ & new_new_n11874__;
  assign new_new_n11876__ = ~new_new_n11867__ & new_new_n11875__;
  assign po070 = ~new_new_n11860__ & ~new_new_n11876__;
  assign new_new_n11878__ = ~new_new_n11774__ & new_new_n11840__;
  assign new_new_n11879__ = ~new_new_n11773__ & ~new_new_n11878__;
  assign new_new_n11880__ = ~new_new_n11650__ & new_new_n11652__;
  assign new_new_n11881__ = ~new_new_n11649__ & ~new_new_n11880__;
  assign new_new_n11882__ = ~new_new_n11879__ & new_new_n11881__;
  assign new_new_n11883__ = new_new_n11879__ & ~new_new_n11881__;
  assign new_new_n11884__ = ~new_new_n11882__ & ~new_new_n11883__;
  assign new_new_n11885__ = ~new_new_n11608__ & ~new_new_n11612__;
  assign new_new_n11886__ = ~new_new_n11609__ & ~new_new_n11885__;
  assign new_new_n11887__ = ~new_new_n11741__ & ~new_new_n11769__;
  assign new_new_n11888__ = ~new_new_n11742__ & ~new_new_n11887__;
  assign new_new_n11889__ = ~new_new_n11886__ & new_new_n11888__;
  assign new_new_n11890__ = new_new_n11886__ & ~new_new_n11888__;
  assign new_new_n11891__ = ~new_new_n11889__ & ~new_new_n11890__;
  assign new_new_n11892__ = ~new_new_n11671__ & ~new_new_n11677__;
  assign new_new_n11893__ = ~new_new_n11676__ & ~new_new_n11892__;
  assign new_new_n11894__ = ~new_new_n11623__ & ~new_new_n11629__;
  assign new_new_n11895__ = ~new_new_n11622__ & ~new_new_n11894__;
  assign new_new_n11896__ = ~new_new_n11893__ & ~new_new_n11895__;
  assign new_new_n11897__ = new_new_n11893__ & new_new_n11895__;
  assign new_new_n11898__ = ~new_new_n11896__ & ~new_new_n11897__;
  assign new_new_n11899__ = ~new_new_n11708__ & ~new_new_n11712__;
  assign new_new_n11900__ = ~new_new_n11711__ & ~new_new_n11899__;
  assign new_new_n11901__ = ~new_new_n11746__ & ~new_new_n11750__;
  assign new_new_n11902__ = ~new_new_n11749__ & ~new_new_n11901__;
  assign new_new_n11903__ = ~new_new_n11758__ & ~new_new_n11762__;
  assign new_new_n11904__ = ~new_new_n11761__ & ~new_new_n11903__;
  assign new_new_n11905__ = ~new_new_n11902__ & ~new_new_n11904__;
  assign new_new_n11906__ = new_new_n11902__ & new_new_n11904__;
  assign new_new_n11907__ = ~new_new_n11905__ & ~new_new_n11906__;
  assign new_new_n11908__ = new_new_n11900__ & ~new_new_n11907__;
  assign new_new_n11909__ = ~new_new_n11900__ & new_new_n11907__;
  assign new_new_n11910__ = ~new_new_n11908__ & ~new_new_n11909__;
  assign new_new_n11911__ = new_new_n11898__ & new_new_n11910__;
  assign new_new_n11912__ = ~new_new_n11898__ & ~new_new_n11910__;
  assign new_new_n11913__ = ~new_new_n11911__ & ~new_new_n11912__;
  assign new_new_n11914__ = new_new_n11891__ & ~new_new_n11913__;
  assign new_new_n11915__ = ~new_new_n11891__ & new_new_n11913__;
  assign new_new_n11916__ = ~new_new_n11914__ & ~new_new_n11915__;
  assign new_new_n11917__ = new_new_n11884__ & ~new_new_n11916__;
  assign new_new_n11918__ = ~new_new_n11884__ & new_new_n11916__;
  assign new_new_n11919__ = ~new_new_n11917__ & ~new_new_n11918__;
  assign new_new_n11920__ = ~new_new_n11660__ & ~new_new_n11697__;
  assign new_new_n11921__ = ~new_new_n11661__ & ~new_new_n11920__;
  assign new_new_n11922__ = ~new_new_n11667__ & new_new_n11681__;
  assign new_new_n11923__ = ~new_new_n11668__ & ~new_new_n11922__;
  assign new_new_n11924__ = ~new_new_n11785__ & ~new_new_n11789__;
  assign new_new_n11925__ = ~new_new_n11788__ & ~new_new_n11924__;
  assign new_new_n11926__ = ~new_new_n11823__ & ~new_new_n11827__;
  assign new_new_n11927__ = ~new_new_n11826__ & ~new_new_n11926__;
  assign new_new_n11928__ = pi34 & pi36;
  assign new_new_n11929__ = pi32 & pi38;
  assign new_new_n11930__ = pi33 & pi37;
  assign new_new_n11931__ = ~new_new_n11929__ & ~new_new_n11930__;
  assign new_new_n11932__ = new_new_n11929__ & new_new_n11930__;
  assign new_new_n11933__ = ~new_new_n11931__ & ~new_new_n11932__;
  assign new_new_n11934__ = new_new_n11928__ & ~new_new_n11933__;
  assign new_new_n11935__ = ~new_new_n11928__ & new_new_n11933__;
  assign new_new_n11936__ = ~new_new_n11934__ & ~new_new_n11935__;
  assign new_new_n11937__ = ~new_new_n11927__ & new_new_n11936__;
  assign new_new_n11938__ = new_new_n11927__ & ~new_new_n11936__;
  assign new_new_n11939__ = ~new_new_n11937__ & ~new_new_n11938__;
  assign new_new_n11940__ = new_new_n11925__ & ~new_new_n11939__;
  assign new_new_n11941__ = ~new_new_n11925__ & new_new_n11939__;
  assign new_new_n11942__ = ~new_new_n11940__ & ~new_new_n11941__;
  assign new_new_n11943__ = new_new_n11923__ & ~new_new_n11942__;
  assign new_new_n11944__ = ~new_new_n11923__ & new_new_n11942__;
  assign new_new_n11945__ = ~new_new_n11943__ & ~new_new_n11944__;
  assign new_new_n11946__ = pi12 & pi58;
  assign new_new_n11947__ = pi13 & pi57;
  assign new_new_n11948__ = ~new_new_n11946__ & ~new_new_n11947__;
  assign new_new_n11949__ = new_new_n11946__ & new_new_n11947__;
  assign new_new_n11950__ = ~new_new_n11948__ & ~new_new_n11949__;
  assign new_new_n11951__ = new_new_n5783__ & ~new_new_n11950__;
  assign new_new_n11952__ = ~new_new_n5783__ & new_new_n11950__;
  assign new_new_n11953__ = ~new_new_n11951__ & ~new_new_n11952__;
  assign new_new_n11954__ = pi18 & pi52;
  assign new_new_n11955__ = pi17 & pi53;
  assign new_new_n11956__ = pi16 & pi54;
  assign new_new_n11957__ = ~new_new_n11955__ & ~new_new_n11956__;
  assign new_new_n11958__ = new_new_n11955__ & new_new_n11956__;
  assign new_new_n11959__ = ~new_new_n11957__ & ~new_new_n11958__;
  assign new_new_n11960__ = new_new_n11954__ & ~new_new_n11959__;
  assign new_new_n11961__ = ~new_new_n11954__ & new_new_n11959__;
  assign new_new_n11962__ = ~new_new_n11960__ & ~new_new_n11961__;
  assign new_new_n11963__ = new_new_n11953__ & new_new_n11962__;
  assign new_new_n11964__ = ~new_new_n11953__ & ~new_new_n11962__;
  assign new_new_n11965__ = ~new_new_n11963__ & ~new_new_n11964__;
  assign new_new_n11966__ = pi11 & pi59;
  assign new_new_n11967__ = pi09 & pi61;
  assign new_new_n11968__ = pi10 & pi60;
  assign new_new_n11969__ = ~new_new_n11967__ & ~new_new_n11968__;
  assign new_new_n11970__ = new_new_n11967__ & new_new_n11968__;
  assign new_new_n11971__ = ~new_new_n11969__ & ~new_new_n11970__;
  assign new_new_n11972__ = new_new_n11966__ & ~new_new_n11971__;
  assign new_new_n11973__ = ~new_new_n11966__ & new_new_n11971__;
  assign new_new_n11974__ = ~new_new_n11972__ & ~new_new_n11973__;
  assign new_new_n11975__ = new_new_n11965__ & ~new_new_n11974__;
  assign new_new_n11976__ = ~new_new_n11965__ & new_new_n11974__;
  assign new_new_n11977__ = ~new_new_n11975__ & ~new_new_n11976__;
  assign new_new_n11978__ = new_new_n11945__ & ~new_new_n11977__;
  assign new_new_n11979__ = ~new_new_n11945__ & new_new_n11977__;
  assign new_new_n11980__ = ~new_new_n11978__ & ~new_new_n11979__;
  assign new_new_n11981__ = new_new_n11617__ & new_new_n11642__;
  assign new_new_n11982__ = ~new_new_n11617__ & ~new_new_n11642__;
  assign new_new_n11983__ = ~new_new_n11624__ & ~new_new_n11629__;
  assign new_new_n11984__ = new_new_n11624__ & new_new_n11629__;
  assign new_new_n11985__ = ~new_new_n11983__ & ~new_new_n11984__;
  assign new_new_n11986__ = ~new_new_n11982__ & ~new_new_n11985__;
  assign new_new_n11987__ = ~new_new_n11981__ & ~new_new_n11986__;
  assign new_new_n11988__ = pi31 & pi39;
  assign new_new_n11989__ = pi29 & pi41;
  assign new_new_n11990__ = pi30 & pi40;
  assign new_new_n11991__ = ~new_new_n11989__ & ~new_new_n11990__;
  assign new_new_n11992__ = new_new_n11989__ & new_new_n11990__;
  assign new_new_n11993__ = ~new_new_n11991__ & ~new_new_n11992__;
  assign new_new_n11994__ = new_new_n11988__ & ~new_new_n11993__;
  assign new_new_n11995__ = ~new_new_n11988__ & new_new_n11993__;
  assign new_new_n11996__ = ~new_new_n11994__ & ~new_new_n11995__;
  assign new_new_n11997__ = pi28 & pi42;
  assign new_new_n11998__ = pi07 & pi63;
  assign new_new_n11999__ = ~new_new_n6164__ & ~new_new_n11998__;
  assign new_new_n12000__ = new_new_n6164__ & new_new_n11998__;
  assign new_new_n12001__ = ~new_new_n11999__ & ~new_new_n12000__;
  assign new_new_n12002__ = new_new_n11997__ & ~new_new_n12001__;
  assign new_new_n12003__ = ~new_new_n11997__ & new_new_n12001__;
  assign new_new_n12004__ = ~new_new_n12002__ & ~new_new_n12003__;
  assign new_new_n12005__ = new_new_n11996__ & new_new_n12004__;
  assign new_new_n12006__ = ~new_new_n11996__ & ~new_new_n12004__;
  assign new_new_n12007__ = ~new_new_n12005__ & ~new_new_n12006__;
  assign new_new_n12008__ = ~new_new_n11634__ & ~new_new_n11640__;
  assign new_new_n12009__ = new_new_n12007__ & ~new_new_n12008__;
  assign new_new_n12010__ = ~new_new_n12007__ & new_new_n12008__;
  assign new_new_n12011__ = ~new_new_n12009__ & ~new_new_n12010__;
  assign new_new_n12012__ = new_new_n11987__ & ~new_new_n12011__;
  assign new_new_n12013__ = ~new_new_n11987__ & new_new_n12011__;
  assign new_new_n12014__ = ~new_new_n12012__ & ~new_new_n12013__;
  assign new_new_n12015__ = pi27 & pi43;
  assign new_new_n12016__ = pi26 & pi44;
  assign new_new_n12017__ = pi25 & pi45;
  assign new_new_n12018__ = ~new_new_n12016__ & ~new_new_n12017__;
  assign new_new_n12019__ = new_new_n12016__ & new_new_n12017__;
  assign new_new_n12020__ = ~new_new_n12018__ & ~new_new_n12019__;
  assign new_new_n12021__ = new_new_n12015__ & ~new_new_n12020__;
  assign new_new_n12022__ = ~new_new_n12015__ & new_new_n12020__;
  assign new_new_n12023__ = ~new_new_n12021__ & ~new_new_n12022__;
  assign new_new_n12024__ = pi21 & pi49;
  assign new_new_n12025__ = pi20 & pi50;
  assign new_new_n12026__ = pi19 & pi51;
  assign new_new_n12027__ = ~new_new_n12025__ & ~new_new_n12026__;
  assign new_new_n12028__ = new_new_n12025__ & new_new_n12026__;
  assign new_new_n12029__ = ~new_new_n12027__ & ~new_new_n12028__;
  assign new_new_n12030__ = new_new_n12024__ & ~new_new_n12029__;
  assign new_new_n12031__ = ~new_new_n12024__ & new_new_n12029__;
  assign new_new_n12032__ = ~new_new_n12030__ & ~new_new_n12031__;
  assign new_new_n12033__ = pi22 & pi48;
  assign new_new_n12034__ = pi15 & pi55;
  assign new_new_n12035__ = pi14 & pi56;
  assign new_new_n12036__ = ~new_new_n12034__ & ~new_new_n12035__;
  assign new_new_n12037__ = new_new_n12034__ & new_new_n12035__;
  assign new_new_n12038__ = ~new_new_n12036__ & ~new_new_n12037__;
  assign new_new_n12039__ = new_new_n12033__ & ~new_new_n12038__;
  assign new_new_n12040__ = ~new_new_n12033__ & new_new_n12038__;
  assign new_new_n12041__ = ~new_new_n12039__ & ~new_new_n12040__;
  assign new_new_n12042__ = new_new_n12032__ & new_new_n12041__;
  assign new_new_n12043__ = ~new_new_n12032__ & ~new_new_n12041__;
  assign new_new_n12044__ = ~new_new_n12042__ & ~new_new_n12043__;
  assign new_new_n12045__ = new_new_n12023__ & ~new_new_n12044__;
  assign new_new_n12046__ = ~new_new_n12023__ & new_new_n12044__;
  assign new_new_n12047__ = ~new_new_n12045__ & ~new_new_n12046__;
  assign new_new_n12048__ = new_new_n12014__ & new_new_n12047__;
  assign new_new_n12049__ = ~new_new_n12014__ & ~new_new_n12047__;
  assign new_new_n12050__ = ~new_new_n12048__ & ~new_new_n12049__;
  assign new_new_n12051__ = ~new_new_n11980__ & new_new_n12050__;
  assign new_new_n12052__ = new_new_n11980__ & ~new_new_n12050__;
  assign new_new_n12053__ = ~new_new_n12051__ & ~new_new_n12052__;
  assign new_new_n12054__ = ~new_new_n11690__ & new_new_n11694__;
  assign new_new_n12055__ = ~new_new_n11691__ & ~new_new_n12054__;
  assign new_new_n12056__ = new_new_n12053__ & new_new_n12055__;
  assign new_new_n12057__ = ~new_new_n12053__ & ~new_new_n12055__;
  assign new_new_n12058__ = ~new_new_n12056__ & ~new_new_n12057__;
  assign new_new_n12059__ = ~new_new_n11921__ & ~new_new_n12058__;
  assign new_new_n12060__ = new_new_n11921__ & new_new_n12058__;
  assign new_new_n12061__ = ~new_new_n12059__ & ~new_new_n12060__;
  assign new_new_n12062__ = ~new_new_n11726__ & ~new_new_n11737__;
  assign new_new_n12063__ = ~new_new_n11727__ & ~new_new_n12062__;
  assign new_new_n12064__ = ~new_new_n11813__ & ~new_new_n11832__;
  assign new_new_n12065__ = ~new_new_n11833__ & ~new_new_n12064__;
  assign new_new_n12066__ = ~new_new_n11756__ & new_new_n11766__;
  assign new_new_n12067__ = ~new_new_n11755__ & ~new_new_n12066__;
  assign new_new_n12068__ = new_new_n12065__ & ~new_new_n12067__;
  assign new_new_n12069__ = ~new_new_n12065__ & new_new_n12067__;
  assign new_new_n12070__ = ~new_new_n12068__ & ~new_new_n12069__;
  assign new_new_n12071__ = ~new_new_n12063__ & ~new_new_n12070__;
  assign new_new_n12072__ = new_new_n12063__ & new_new_n12070__;
  assign new_new_n12073__ = ~new_new_n12071__ & ~new_new_n12072__;
  assign new_new_n12074__ = ~pi07 & ~pi34;
  assign new_new_n12075__ = ~new_new_n11814__ & ~new_new_n11818__;
  assign new_new_n12076__ = ~new_new_n11817__ & ~new_new_n12075__;
  assign new_new_n12077__ = pi34 & new_new_n12076__;
  assign new_new_n12078__ = ~pi62 & ~new_new_n12077__;
  assign new_new_n12079__ = ~pi08 & ~new_new_n12076__;
  assign new_new_n12080__ = pi08 & pi62;
  assign new_new_n12081__ = new_new_n12076__ & new_new_n12080__;
  assign new_new_n12082__ = pi35 & ~new_new_n12074__;
  assign new_new_n12083__ = ~new_new_n12079__ & new_new_n12082__;
  assign new_new_n12084__ = ~new_new_n12081__ & new_new_n12083__;
  assign new_new_n12085__ = ~new_new_n12078__ & new_new_n12084__;
  assign new_new_n12086__ = pi34 & pi35;
  assign new_new_n12087__ = new_new_n12076__ & ~new_new_n12080__;
  assign new_new_n12088__ = ~pi08 & ~new_new_n4603__;
  assign new_new_n12089__ = ~new_new_n4603__ & new_new_n12076__;
  assign new_new_n12090__ = pi62 & ~new_new_n12088__;
  assign new_new_n12091__ = ~new_new_n12089__ & new_new_n12090__;
  assign new_new_n12092__ = ~new_new_n12086__ & ~new_new_n12087__;
  assign new_new_n12093__ = ~new_new_n12091__ & new_new_n12092__;
  assign new_new_n12094__ = ~new_new_n12085__ & ~new_new_n12093__;
  assign new_new_n12095__ = ~new_new_n11794__ & new_new_n11798__;
  assign new_new_n12096__ = ~new_new_n11795__ & ~new_new_n12095__;
  assign new_new_n12097__ = new_new_n12094__ & ~new_new_n12096__;
  assign new_new_n12098__ = ~new_new_n12094__ & new_new_n12096__;
  assign new_new_n12099__ = ~new_new_n12097__ & ~new_new_n12098__;
  assign new_new_n12100__ = ~new_new_n11729__ & ~new_new_n11733__;
  assign new_new_n12101__ = ~new_new_n11732__ & ~new_new_n12100__;
  assign new_new_n12102__ = ~new_new_n11776__ & ~new_new_n11780__;
  assign new_new_n12103__ = ~new_new_n11779__ & ~new_new_n12102__;
  assign new_new_n12104__ = new_new_n12101__ & new_new_n12103__;
  assign new_new_n12105__ = ~new_new_n12101__ & ~new_new_n12103__;
  assign new_new_n12106__ = ~new_new_n11717__ & ~new_new_n11721__;
  assign new_new_n12107__ = ~new_new_n11720__ & ~new_new_n12106__;
  assign new_new_n12108__ = ~new_new_n12104__ & ~new_new_n12107__;
  assign new_new_n12109__ = ~new_new_n12105__ & ~new_new_n12108__;
  assign new_new_n12110__ = ~new_new_n12104__ & new_new_n12109__;
  assign new_new_n12111__ = ~new_new_n12105__ & new_new_n12108__;
  assign new_new_n12112__ = ~new_new_n12107__ & ~new_new_n12111__;
  assign new_new_n12113__ = ~new_new_n12110__ & ~new_new_n12112__;
  assign new_new_n12114__ = new_new_n12099__ & ~new_new_n12113__;
  assign new_new_n12115__ = ~new_new_n12099__ & new_new_n12113__;
  assign new_new_n12116__ = ~new_new_n12114__ & ~new_new_n12115__;
  assign new_new_n12117__ = ~new_new_n11806__ & new_new_n11837__;
  assign new_new_n12118__ = ~new_new_n11807__ & ~new_new_n12117__;
  assign new_new_n12119__ = ~new_new_n12116__ & new_new_n12118__;
  assign new_new_n12120__ = new_new_n12116__ & ~new_new_n12118__;
  assign new_new_n12121__ = ~new_new_n12119__ & ~new_new_n12120__;
  assign new_new_n12122__ = new_new_n12073__ & new_new_n12121__;
  assign new_new_n12123__ = ~new_new_n12073__ & ~new_new_n12121__;
  assign new_new_n12124__ = ~new_new_n12122__ & ~new_new_n12123__;
  assign new_new_n12125__ = new_new_n12061__ & ~new_new_n12124__;
  assign new_new_n12126__ = ~new_new_n12061__ & new_new_n12124__;
  assign new_new_n12127__ = ~new_new_n12125__ & ~new_new_n12126__;
  assign new_new_n12128__ = ~new_new_n11919__ & new_new_n12127__;
  assign new_new_n12129__ = new_new_n11919__ & ~new_new_n12127__;
  assign new_new_n12130__ = ~new_new_n12128__ & ~new_new_n12129__;
  assign new_new_n12131__ = ~new_new_n11701__ & ~new_new_n11853__;
  assign new_new_n12132__ = ~new_new_n11702__ & ~new_new_n12131__;
  assign new_new_n12133__ = new_new_n12130__ & ~new_new_n12132__;
  assign new_new_n12134__ = ~new_new_n12130__ & new_new_n12132__;
  assign new_new_n12135__ = ~new_new_n12133__ & ~new_new_n12134__;
  assign new_new_n12136__ = ~new_new_n11847__ & ~new_new_n11850__;
  assign new_new_n12137__ = ~new_new_n11846__ & ~new_new_n12136__;
  assign new_new_n12138__ = ~new_new_n11596__ & ~new_new_n11856__;
  assign new_new_n12139__ = new_new_n11596__ & new_new_n11856__;
  assign new_new_n12140__ = ~new_new_n11468__ & ~new_new_n12139__;
  assign new_new_n12141__ = ~new_new_n12138__ & ~new_new_n12140__;
  assign new_new_n12142__ = ~new_new_n11598__ & ~new_new_n11856__;
  assign new_new_n12143__ = ~new_new_n11599__ & ~new_new_n12142__;
  assign new_new_n12144__ = ~new_new_n11467__ & new_new_n12143__;
  assign new_new_n12145__ = ~new_new_n12141__ & ~new_new_n12144__;
  assign new_new_n12146__ = new_new_n12137__ & ~new_new_n12145__;
  assign new_new_n12147__ = ~new_new_n12137__ & new_new_n12145__;
  assign new_new_n12148__ = ~new_new_n12146__ & ~new_new_n12147__;
  assign new_new_n12149__ = new_new_n12135__ & new_new_n12148__;
  assign new_new_n12150__ = ~new_new_n12135__ & ~new_new_n12148__;
  assign po071 = ~new_new_n12149__ & ~new_new_n12150__;
  assign new_new_n12152__ = new_new_n12130__ & new_new_n12137__;
  assign new_new_n12153__ = ~new_new_n12128__ & ~new_new_n12152__;
  assign new_new_n12154__ = ~new_new_n12130__ & ~new_new_n12137__;
  assign new_new_n12155__ = ~new_new_n12152__ & ~new_new_n12154__;
  assign new_new_n12156__ = ~new_new_n12132__ & new_new_n12155__;
  assign new_new_n12157__ = new_new_n12145__ & ~new_new_n12156__;
  assign new_new_n12158__ = new_new_n12132__ & ~new_new_n12155__;
  assign new_new_n12159__ = ~new_new_n12157__ & ~new_new_n12158__;
  assign new_new_n12160__ = ~new_new_n12153__ & new_new_n12159__;
  assign new_new_n12161__ = new_new_n12153__ & ~new_new_n12159__;
  assign new_new_n12162__ = ~new_new_n12160__ & ~new_new_n12161__;
  assign new_new_n12163__ = ~new_new_n12060__ & ~new_new_n12124__;
  assign new_new_n12164__ = ~new_new_n12059__ & ~new_new_n12163__;
  assign new_new_n12165__ = ~new_new_n11882__ & ~new_new_n11916__;
  assign new_new_n12166__ = ~new_new_n11883__ & ~new_new_n12165__;
  assign new_new_n12167__ = ~new_new_n11896__ & ~new_new_n11910__;
  assign new_new_n12168__ = ~new_new_n11897__ & ~new_new_n12167__;
  assign new_new_n12169__ = pi09 & pi62;
  assign new_new_n12170__ = pi22 & pi49;
  assign new_new_n12171__ = new_new_n12169__ & ~new_new_n12170__;
  assign new_new_n12172__ = ~new_new_n12169__ & new_new_n12170__;
  assign new_new_n12173__ = ~new_new_n12171__ & ~new_new_n12172__;
  assign new_new_n12174__ = pi21 & pi50;
  assign new_new_n12175__ = pi19 & pi52;
  assign new_new_n12176__ = pi20 & pi51;
  assign new_new_n12177__ = ~new_new_n12175__ & ~new_new_n12176__;
  assign new_new_n12178__ = new_new_n12175__ & new_new_n12176__;
  assign new_new_n12179__ = ~new_new_n12177__ & ~new_new_n12178__;
  assign new_new_n12180__ = new_new_n12174__ & ~new_new_n12179__;
  assign new_new_n12181__ = ~new_new_n12174__ & new_new_n12179__;
  assign new_new_n12182__ = ~new_new_n12180__ & ~new_new_n12181__;
  assign new_new_n12183__ = pi33 & pi38;
  assign new_new_n12184__ = pi34 & pi37;
  assign new_new_n12185__ = ~new_new_n12183__ & ~new_new_n12184__;
  assign new_new_n12186__ = new_new_n12183__ & new_new_n12184__;
  assign new_new_n12187__ = ~new_new_n12185__ & ~new_new_n12186__;
  assign new_new_n12188__ = pi35 & pi36;
  assign new_new_n12189__ = ~new_new_n12187__ & new_new_n12188__;
  assign new_new_n12190__ = new_new_n12187__ & ~new_new_n12188__;
  assign new_new_n12191__ = ~new_new_n12189__ & ~new_new_n12190__;
  assign new_new_n12192__ = pi36 & ~new_new_n12191__;
  assign new_new_n12193__ = ~pi36 & ~new_new_n12187__;
  assign new_new_n12194__ = ~new_new_n12192__ & ~new_new_n12193__;
  assign new_new_n12195__ = new_new_n12182__ & ~new_new_n12194__;
  assign new_new_n12196__ = ~new_new_n12182__ & new_new_n12194__;
  assign new_new_n12197__ = ~new_new_n12195__ & ~new_new_n12196__;
  assign new_new_n12198__ = new_new_n12173__ & new_new_n12197__;
  assign new_new_n12199__ = ~new_new_n12173__ & ~new_new_n12197__;
  assign new_new_n12200__ = ~new_new_n12198__ & ~new_new_n12199__;
  assign new_new_n12201__ = ~new_new_n12168__ & ~new_new_n12200__;
  assign new_new_n12202__ = new_new_n12168__ & new_new_n12200__;
  assign new_new_n12203__ = ~new_new_n12201__ & ~new_new_n12202__;
  assign new_new_n12204__ = ~new_new_n11928__ & ~new_new_n11932__;
  assign new_new_n12205__ = ~new_new_n11931__ & ~new_new_n12204__;
  assign new_new_n12206__ = ~new_new_n11954__ & ~new_new_n11958__;
  assign new_new_n12207__ = ~new_new_n11957__ & ~new_new_n12206__;
  assign new_new_n12208__ = new_new_n12205__ & new_new_n12207__;
  assign new_new_n12209__ = ~new_new_n12205__ & ~new_new_n12207__;
  assign new_new_n12210__ = ~new_new_n12208__ & ~new_new_n12209__;
  assign new_new_n12211__ = pi11 & pi60;
  assign new_new_n12212__ = pi10 & pi61;
  assign new_new_n12213__ = pi08 & pi63;
  assign new_new_n12214__ = ~new_new_n12212__ & ~new_new_n12213__;
  assign new_new_n12215__ = new_new_n12212__ & new_new_n12213__;
  assign new_new_n12216__ = ~new_new_n12214__ & ~new_new_n12215__;
  assign new_new_n12217__ = new_new_n12211__ & ~new_new_n12216__;
  assign new_new_n12218__ = ~new_new_n12211__ & new_new_n12216__;
  assign new_new_n12219__ = ~new_new_n12217__ & ~new_new_n12218__;
  assign new_new_n12220__ = new_new_n12210__ & ~new_new_n12219__;
  assign new_new_n12221__ = ~new_new_n12210__ & new_new_n12219__;
  assign new_new_n12222__ = ~new_new_n12220__ & ~new_new_n12221__;
  assign new_new_n12223__ = new_new_n12203__ & ~new_new_n12222__;
  assign new_new_n12224__ = ~new_new_n12203__ & new_new_n12222__;
  assign new_new_n12225__ = ~new_new_n12223__ & ~new_new_n12224__;
  assign new_new_n12226__ = ~new_new_n12068__ & ~new_new_n12072__;
  assign new_new_n12227__ = pi26 & pi45;
  assign new_new_n12228__ = pi25 & pi46;
  assign new_new_n12229__ = pi24 & pi47;
  assign new_new_n12230__ = ~new_new_n12228__ & ~new_new_n12229__;
  assign new_new_n12231__ = new_new_n12228__ & new_new_n12229__;
  assign new_new_n12232__ = ~new_new_n12230__ & ~new_new_n12231__;
  assign new_new_n12233__ = new_new_n12227__ & ~new_new_n12232__;
  assign new_new_n12234__ = ~new_new_n12227__ & new_new_n12232__;
  assign new_new_n12235__ = ~new_new_n12233__ & ~new_new_n12234__;
  assign new_new_n12236__ = pi16 & pi55;
  assign new_new_n12237__ = pi15 & pi56;
  assign new_new_n12238__ = pi14 & pi57;
  assign new_new_n12239__ = ~new_new_n12237__ & ~new_new_n12238__;
  assign new_new_n12240__ = new_new_n12237__ & new_new_n12238__;
  assign new_new_n12241__ = ~new_new_n12239__ & ~new_new_n12240__;
  assign new_new_n12242__ = new_new_n12236__ & ~new_new_n12241__;
  assign new_new_n12243__ = ~new_new_n12236__ & new_new_n12241__;
  assign new_new_n12244__ = ~new_new_n12242__ & ~new_new_n12243__;
  assign new_new_n12245__ = ~new_new_n12235__ & ~new_new_n12244__;
  assign new_new_n12246__ = new_new_n12235__ & new_new_n12244__;
  assign new_new_n12247__ = ~new_new_n12245__ & ~new_new_n12246__;
  assign new_new_n12248__ = ~new_new_n12024__ & ~new_new_n12028__;
  assign new_new_n12249__ = ~new_new_n12027__ & ~new_new_n12248__;
  assign new_new_n12250__ = pi13 & pi58;
  assign new_new_n12251__ = pi12 & pi59;
  assign new_new_n12252__ = new_new_n12250__ & ~new_new_n12251__;
  assign new_new_n12253__ = ~new_new_n12250__ & new_new_n12251__;
  assign new_new_n12254__ = ~new_new_n12252__ & ~new_new_n12253__;
  assign new_new_n12255__ = new_new_n12249__ & new_new_n12254__;
  assign new_new_n12256__ = ~new_new_n12249__ & ~new_new_n12254__;
  assign new_new_n12257__ = ~new_new_n12255__ & ~new_new_n12256__;
  assign new_new_n12258__ = new_new_n12247__ & ~new_new_n12257__;
  assign new_new_n12259__ = ~new_new_n12247__ & new_new_n12257__;
  assign new_new_n12260__ = ~new_new_n12258__ & ~new_new_n12259__;
  assign new_new_n12261__ = new_new_n12226__ & new_new_n12260__;
  assign new_new_n12262__ = ~new_new_n12226__ & ~new_new_n12260__;
  assign new_new_n12263__ = ~new_new_n12261__ & ~new_new_n12262__;
  assign new_new_n12264__ = pi29 & pi42;
  assign new_new_n12265__ = pi28 & pi43;
  assign new_new_n12266__ = pi27 & pi44;
  assign new_new_n12267__ = ~new_new_n12265__ & ~new_new_n12266__;
  assign new_new_n12268__ = new_new_n12265__ & new_new_n12266__;
  assign new_new_n12269__ = ~new_new_n12267__ & ~new_new_n12268__;
  assign new_new_n12270__ = new_new_n12264__ & ~new_new_n12269__;
  assign new_new_n12271__ = ~new_new_n12264__ & new_new_n12269__;
  assign new_new_n12272__ = ~new_new_n12270__ & ~new_new_n12271__;
  assign new_new_n12273__ = pi23 & pi48;
  assign new_new_n12274__ = pi17 & pi54;
  assign new_new_n12275__ = pi18 & pi53;
  assign new_new_n12276__ = ~new_new_n12274__ & ~new_new_n12275__;
  assign new_new_n12277__ = new_new_n12274__ & new_new_n12275__;
  assign new_new_n12278__ = ~new_new_n12276__ & ~new_new_n12277__;
  assign new_new_n12279__ = new_new_n12273__ & ~new_new_n12278__;
  assign new_new_n12280__ = ~new_new_n12273__ & new_new_n12278__;
  assign new_new_n12281__ = ~new_new_n12279__ & ~new_new_n12280__;
  assign new_new_n12282__ = new_new_n12272__ & new_new_n12281__;
  assign new_new_n12283__ = ~new_new_n12272__ & ~new_new_n12281__;
  assign new_new_n12284__ = ~new_new_n12282__ & ~new_new_n12283__;
  assign new_new_n12285__ = pi32 & pi39;
  assign new_new_n12286__ = pi30 & pi41;
  assign new_new_n12287__ = pi31 & pi40;
  assign new_new_n12288__ = ~new_new_n12286__ & ~new_new_n12287__;
  assign new_new_n12289__ = new_new_n12286__ & new_new_n12287__;
  assign new_new_n12290__ = ~new_new_n12288__ & ~new_new_n12289__;
  assign new_new_n12291__ = new_new_n12285__ & ~new_new_n12290__;
  assign new_new_n12292__ = ~new_new_n12285__ & new_new_n12290__;
  assign new_new_n12293__ = ~new_new_n12291__ & ~new_new_n12292__;
  assign new_new_n12294__ = new_new_n12284__ & ~new_new_n12293__;
  assign new_new_n12295__ = ~new_new_n12284__ & new_new_n12293__;
  assign new_new_n12296__ = ~new_new_n12294__ & ~new_new_n12295__;
  assign new_new_n12297__ = new_new_n12263__ & ~new_new_n12296__;
  assign new_new_n12298__ = ~new_new_n12263__ & new_new_n12296__;
  assign new_new_n12299__ = ~new_new_n12297__ & ~new_new_n12298__;
  assign new_new_n12300__ = new_new_n12225__ & new_new_n12299__;
  assign new_new_n12301__ = ~new_new_n12225__ & ~new_new_n12299__;
  assign new_new_n12302__ = ~new_new_n12300__ & ~new_new_n12301__;
  assign new_new_n12303__ = ~new_new_n11890__ & ~new_new_n11913__;
  assign new_new_n12304__ = ~new_new_n11889__ & ~new_new_n12303__;
  assign new_new_n12305__ = new_new_n12302__ & new_new_n12304__;
  assign new_new_n12306__ = ~new_new_n12302__ & ~new_new_n12304__;
  assign new_new_n12307__ = ~new_new_n12305__ & ~new_new_n12306__;
  assign new_new_n12308__ = new_new_n12166__ & ~new_new_n12307__;
  assign new_new_n12309__ = ~new_new_n12166__ & new_new_n12307__;
  assign new_new_n12310__ = ~new_new_n12308__ & ~new_new_n12309__;
  assign new_new_n12311__ = ~new_new_n12012__ & ~new_new_n12047__;
  assign new_new_n12312__ = ~new_new_n12013__ & ~new_new_n12311__;
  assign new_new_n12313__ = ~new_new_n11963__ & ~new_new_n11974__;
  assign new_new_n12314__ = ~new_new_n11964__ & ~new_new_n12313__;
  assign new_new_n12315__ = ~new_new_n11900__ & ~new_new_n11906__;
  assign new_new_n12316__ = ~new_new_n11905__ & ~new_new_n12315__;
  assign new_new_n12317__ = ~new_new_n12023__ & ~new_new_n12042__;
  assign new_new_n12318__ = ~new_new_n12043__ & ~new_new_n12317__;
  assign new_new_n12319__ = ~new_new_n12316__ & new_new_n12318__;
  assign new_new_n12320__ = new_new_n12316__ & ~new_new_n12318__;
  assign new_new_n12321__ = ~new_new_n12319__ & ~new_new_n12320__;
  assign new_new_n12322__ = new_new_n12314__ & ~new_new_n12321__;
  assign new_new_n12323__ = ~new_new_n12314__ & new_new_n12321__;
  assign new_new_n12324__ = ~new_new_n12322__ & ~new_new_n12323__;
  assign new_new_n12325__ = new_new_n12312__ & new_new_n12324__;
  assign new_new_n12326__ = ~new_new_n12312__ & ~new_new_n12324__;
  assign new_new_n12327__ = ~new_new_n12325__ & ~new_new_n12326__;
  assign new_new_n12328__ = ~new_new_n11988__ & ~new_new_n11992__;
  assign new_new_n12329__ = ~new_new_n11991__ & ~new_new_n12328__;
  assign new_new_n12330__ = ~new_new_n11997__ & ~new_new_n12000__;
  assign new_new_n12331__ = ~new_new_n11999__ & ~new_new_n12330__;
  assign new_new_n12332__ = ~new_new_n12329__ & ~new_new_n12331__;
  assign new_new_n12333__ = new_new_n12329__ & new_new_n12331__;
  assign new_new_n12334__ = ~new_new_n12332__ & ~new_new_n12333__;
  assign new_new_n12335__ = ~new_new_n12033__ & ~new_new_n12037__;
  assign new_new_n12336__ = ~new_new_n12036__ & ~new_new_n12335__;
  assign new_new_n12337__ = ~new_new_n12334__ & new_new_n12336__;
  assign new_new_n12338__ = new_new_n12334__ & ~new_new_n12336__;
  assign new_new_n12339__ = ~new_new_n12337__ & ~new_new_n12338__;
  assign new_new_n12340__ = ~new_new_n12005__ & new_new_n12008__;
  assign new_new_n12341__ = ~new_new_n12006__ & ~new_new_n12340__;
  assign new_new_n12342__ = ~new_new_n12339__ & ~new_new_n12341__;
  assign new_new_n12343__ = new_new_n12339__ & new_new_n12341__;
  assign new_new_n12344__ = ~new_new_n12342__ & ~new_new_n12343__;
  assign new_new_n12345__ = ~new_new_n12015__ & ~new_new_n12019__;
  assign new_new_n12346__ = ~new_new_n12018__ & ~new_new_n12345__;
  assign new_new_n12347__ = ~new_new_n11966__ & ~new_new_n11970__;
  assign new_new_n12348__ = ~new_new_n11969__ & ~new_new_n12347__;
  assign new_new_n12349__ = ~new_new_n5783__ & ~new_new_n11949__;
  assign new_new_n12350__ = ~new_new_n11948__ & ~new_new_n12349__;
  assign new_new_n12351__ = new_new_n12348__ & new_new_n12350__;
  assign new_new_n12352__ = ~new_new_n12348__ & ~new_new_n12350__;
  assign new_new_n12353__ = ~new_new_n12351__ & ~new_new_n12352__;
  assign new_new_n12354__ = new_new_n12346__ & ~new_new_n12353__;
  assign new_new_n12355__ = ~new_new_n12346__ & new_new_n12353__;
  assign new_new_n12356__ = ~new_new_n12354__ & ~new_new_n12355__;
  assign new_new_n12357__ = new_new_n12344__ & ~new_new_n12356__;
  assign new_new_n12358__ = ~new_new_n12344__ & new_new_n12356__;
  assign new_new_n12359__ = ~new_new_n12357__ & ~new_new_n12358__;
  assign new_new_n12360__ = new_new_n12327__ & ~new_new_n12359__;
  assign new_new_n12361__ = ~new_new_n12327__ & new_new_n12359__;
  assign new_new_n12362__ = ~new_new_n12360__ & ~new_new_n12361__;
  assign new_new_n12363__ = new_new_n12310__ & ~new_new_n12362__;
  assign new_new_n12364__ = ~new_new_n12310__ & new_new_n12362__;
  assign new_new_n12365__ = ~new_new_n12363__ & ~new_new_n12364__;
  assign new_new_n12366__ = ~new_new_n12164__ & new_new_n12365__;
  assign new_new_n12367__ = new_new_n12164__ & ~new_new_n12365__;
  assign new_new_n12368__ = ~new_new_n12366__ & ~new_new_n12367__;
  assign new_new_n12369__ = ~new_new_n12052__ & ~new_new_n12055__;
  assign new_new_n12370__ = ~new_new_n12051__ & ~new_new_n12369__;
  assign new_new_n12371__ = new_new_n12073__ & ~new_new_n12119__;
  assign new_new_n12372__ = ~new_new_n12120__ & ~new_new_n12371__;
  assign new_new_n12373__ = ~new_new_n12370__ & new_new_n12372__;
  assign new_new_n12374__ = new_new_n12370__ & ~new_new_n12372__;
  assign new_new_n12375__ = ~new_new_n12373__ & ~new_new_n12374__;
  assign new_new_n12376__ = ~new_new_n12098__ & new_new_n12113__;
  assign new_new_n12377__ = ~new_new_n12097__ & ~new_new_n12376__;
  assign new_new_n12378__ = ~new_new_n11943__ & ~new_new_n11977__;
  assign new_new_n12379__ = ~new_new_n11944__ & ~new_new_n12378__;
  assign new_new_n12380__ = new_new_n12076__ & ~new_new_n12088__;
  assign new_new_n12381__ = new_new_n4803__ & ~new_new_n12074__;
  assign new_new_n12382__ = ~new_new_n12380__ & ~new_new_n12381__;
  assign new_new_n12383__ = pi62 & ~new_new_n12382__;
  assign new_new_n12384__ = new_new_n12076__ & new_new_n12086__;
  assign new_new_n12385__ = ~new_new_n12383__ & ~new_new_n12384__;
  assign new_new_n12386__ = ~new_new_n12109__ & new_new_n12385__;
  assign new_new_n12387__ = new_new_n12109__ & ~new_new_n12385__;
  assign new_new_n12388__ = ~new_new_n12386__ & ~new_new_n12387__;
  assign new_new_n12389__ = new_new_n11925__ & ~new_new_n11937__;
  assign new_new_n12390__ = ~new_new_n11938__ & ~new_new_n12389__;
  assign new_new_n12391__ = new_new_n12388__ & new_new_n12390__;
  assign new_new_n12392__ = ~new_new_n12388__ & ~new_new_n12390__;
  assign new_new_n12393__ = ~new_new_n12391__ & ~new_new_n12392__;
  assign new_new_n12394__ = new_new_n12379__ & ~new_new_n12393__;
  assign new_new_n12395__ = ~new_new_n12379__ & new_new_n12393__;
  assign new_new_n12396__ = ~new_new_n12394__ & ~new_new_n12395__;
  assign new_new_n12397__ = new_new_n12377__ & new_new_n12396__;
  assign new_new_n12398__ = ~new_new_n12377__ & ~new_new_n12396__;
  assign new_new_n12399__ = ~new_new_n12397__ & ~new_new_n12398__;
  assign new_new_n12400__ = new_new_n12375__ & ~new_new_n12399__;
  assign new_new_n12401__ = ~new_new_n12375__ & new_new_n12399__;
  assign new_new_n12402__ = ~new_new_n12400__ & ~new_new_n12401__;
  assign new_new_n12403__ = new_new_n12368__ & ~new_new_n12402__;
  assign new_new_n12404__ = ~new_new_n12368__ & new_new_n12402__;
  assign new_new_n12405__ = ~new_new_n12403__ & ~new_new_n12404__;
  assign new_new_n12406__ = new_new_n12162__ & new_new_n12405__;
  assign new_new_n12407__ = ~new_new_n12162__ & ~new_new_n12405__;
  assign po072 = new_new_n12406__ | new_new_n12407__;
  assign new_new_n12409__ = ~new_new_n12367__ & new_new_n12402__;
  assign new_new_n12410__ = ~new_new_n12366__ & ~new_new_n12409__;
  assign new_new_n12411__ = new_new_n12160__ & new_new_n12410__;
  assign new_new_n12412__ = new_new_n12366__ & new_new_n12402__;
  assign new_new_n12413__ = new_new_n12367__ & ~new_new_n12402__;
  assign new_new_n12414__ = ~new_new_n12412__ & ~new_new_n12413__;
  assign new_new_n12415__ = new_new_n12162__ & new_new_n12414__;
  assign new_new_n12416__ = new_new_n12161__ & ~new_new_n12410__;
  assign new_new_n12417__ = ~new_new_n12411__ & ~new_new_n12416__;
  assign new_new_n12418__ = ~new_new_n12415__ & new_new_n12417__;
  assign new_new_n12419__ = ~new_new_n12261__ & ~new_new_n12296__;
  assign new_new_n12420__ = ~new_new_n12262__ & ~new_new_n12419__;
  assign new_new_n12421__ = ~new_new_n12346__ & ~new_new_n12351__;
  assign new_new_n12422__ = ~new_new_n12352__ & ~new_new_n12421__;
  assign new_new_n12423__ = ~new_new_n12282__ & ~new_new_n12293__;
  assign new_new_n12424__ = ~new_new_n12283__ & ~new_new_n12423__;
  assign new_new_n12425__ = new_new_n12182__ & new_new_n12191__;
  assign new_new_n12426__ = ~new_new_n12182__ & ~new_new_n12191__;
  assign new_new_n12427__ = pi36 & new_new_n12173__;
  assign new_new_n12428__ = ~pi36 & ~new_new_n12173__;
  assign new_new_n12429__ = ~new_new_n12427__ & ~new_new_n12428__;
  assign new_new_n12430__ = ~new_new_n12426__ & new_new_n12429__;
  assign new_new_n12431__ = ~new_new_n12425__ & ~new_new_n12430__;
  assign new_new_n12432__ = new_new_n12424__ & ~new_new_n12431__;
  assign new_new_n12433__ = ~new_new_n12424__ & new_new_n12431__;
  assign new_new_n12434__ = ~new_new_n12432__ & ~new_new_n12433__;
  assign new_new_n12435__ = new_new_n12422__ & ~new_new_n12434__;
  assign new_new_n12436__ = ~new_new_n12422__ & new_new_n12434__;
  assign new_new_n12437__ = ~new_new_n12435__ & ~new_new_n12436__;
  assign new_new_n12438__ = new_new_n12420__ & ~new_new_n12437__;
  assign new_new_n12439__ = ~new_new_n12420__ & new_new_n12437__;
  assign new_new_n12440__ = ~new_new_n12438__ & ~new_new_n12439__;
  assign new_new_n12441__ = ~new_new_n12245__ & new_new_n12257__;
  assign new_new_n12442__ = ~new_new_n12246__ & ~new_new_n12441__;
  assign new_new_n12443__ = ~new_new_n12174__ & ~new_new_n12178__;
  assign new_new_n12444__ = ~new_new_n12177__ & ~new_new_n12443__;
  assign new_new_n12445__ = ~new_new_n12186__ & ~new_new_n12188__;
  assign new_new_n12446__ = ~new_new_n12185__ & ~new_new_n12445__;
  assign new_new_n12447__ = ~new_new_n12444__ & ~new_new_n12446__;
  assign new_new_n12448__ = new_new_n12444__ & new_new_n12446__;
  assign new_new_n12449__ = ~new_new_n12447__ & ~new_new_n12448__;
  assign new_new_n12450__ = ~pi36 & ~new_new_n12169__;
  assign new_new_n12451__ = new_new_n12170__ & ~new_new_n12450__;
  assign new_new_n12452__ = pi62 & new_new_n5347__;
  assign new_new_n12453__ = ~new_new_n12451__ & ~new_new_n12452__;
  assign new_new_n12454__ = new_new_n12449__ & ~new_new_n12453__;
  assign new_new_n12455__ = ~new_new_n12449__ & new_new_n12453__;
  assign new_new_n12456__ = ~new_new_n12454__ & ~new_new_n12455__;
  assign new_new_n12457__ = new_new_n12442__ & new_new_n12456__;
  assign new_new_n12458__ = ~new_new_n12442__ & ~new_new_n12456__;
  assign new_new_n12459__ = ~new_new_n12457__ & ~new_new_n12458__;
  assign new_new_n12460__ = ~new_new_n12285__ & ~new_new_n12289__;
  assign new_new_n12461__ = ~new_new_n12288__ & ~new_new_n12460__;
  assign new_new_n12462__ = ~new_new_n12264__ & ~new_new_n12268__;
  assign new_new_n12463__ = ~new_new_n12267__ & ~new_new_n12462__;
  assign new_new_n12464__ = ~new_new_n12273__ & ~new_new_n12277__;
  assign new_new_n12465__ = ~new_new_n12276__ & ~new_new_n12464__;
  assign new_new_n12466__ = ~new_new_n12463__ & ~new_new_n12465__;
  assign new_new_n12467__ = new_new_n12463__ & new_new_n12465__;
  assign new_new_n12468__ = ~new_new_n12466__ & ~new_new_n12467__;
  assign new_new_n12469__ = new_new_n12461__ & ~new_new_n12468__;
  assign new_new_n12470__ = ~new_new_n12461__ & new_new_n12468__;
  assign new_new_n12471__ = ~new_new_n12469__ & ~new_new_n12470__;
  assign new_new_n12472__ = ~new_new_n12459__ & new_new_n12471__;
  assign new_new_n12473__ = new_new_n12459__ & ~new_new_n12471__;
  assign new_new_n12474__ = ~new_new_n12472__ & ~new_new_n12473__;
  assign new_new_n12475__ = ~new_new_n12440__ & new_new_n12474__;
  assign new_new_n12476__ = new_new_n12440__ & ~new_new_n12474__;
  assign new_new_n12477__ = ~new_new_n12475__ & ~new_new_n12476__;
  assign new_new_n12478__ = ~new_new_n12373__ & new_new_n12399__;
  assign new_new_n12479__ = ~new_new_n12374__ & ~new_new_n12478__;
  assign new_new_n12480__ = new_new_n12477__ & ~new_new_n12479__;
  assign new_new_n12481__ = ~new_new_n12477__ & new_new_n12479__;
  assign new_new_n12482__ = ~new_new_n12480__ & ~new_new_n12481__;
  assign new_new_n12483__ = new_new_n12377__ & ~new_new_n12394__;
  assign new_new_n12484__ = ~new_new_n12395__ & ~new_new_n12483__;
  assign new_new_n12485__ = ~new_new_n12227__ & ~new_new_n12231__;
  assign new_new_n12486__ = ~new_new_n12230__ & ~new_new_n12485__;
  assign new_new_n12487__ = ~new_new_n12236__ & ~new_new_n12240__;
  assign new_new_n12488__ = ~new_new_n12239__ & ~new_new_n12487__;
  assign new_new_n12489__ = ~new_new_n12486__ & ~new_new_n12488__;
  assign new_new_n12490__ = new_new_n12486__ & new_new_n12488__;
  assign new_new_n12491__ = ~new_new_n12489__ & ~new_new_n12490__;
  assign new_new_n12492__ = ~new_new_n12211__ & ~new_new_n12215__;
  assign new_new_n12493__ = ~new_new_n12214__ & ~new_new_n12492__;
  assign new_new_n12494__ = ~new_new_n12491__ & new_new_n12493__;
  assign new_new_n12495__ = ~new_new_n12490__ & ~new_new_n12493__;
  assign new_new_n12496__ = ~new_new_n12489__ & new_new_n12495__;
  assign new_new_n12497__ = ~new_new_n12494__ & ~new_new_n12496__;
  assign new_new_n12498__ = ~new_new_n12386__ & ~new_new_n12390__;
  assign new_new_n12499__ = ~new_new_n12387__ & ~new_new_n12498__;
  assign new_new_n12500__ = new_new_n12497__ & new_new_n12499__;
  assign new_new_n12501__ = ~new_new_n12497__ & ~new_new_n12499__;
  assign new_new_n12502__ = ~new_new_n12500__ & ~new_new_n12501__;
  assign new_new_n12503__ = pi28 & pi44;
  assign new_new_n12504__ = pi27 & pi45;
  assign new_new_n12505__ = pi26 & pi46;
  assign new_new_n12506__ = ~new_new_n12504__ & ~new_new_n12505__;
  assign new_new_n12507__ = new_new_n12504__ & new_new_n12505__;
  assign new_new_n12508__ = ~new_new_n12506__ & ~new_new_n12507__;
  assign new_new_n12509__ = new_new_n12503__ & ~new_new_n12508__;
  assign new_new_n12510__ = ~new_new_n12503__ & new_new_n12508__;
  assign new_new_n12511__ = ~new_new_n12509__ & ~new_new_n12510__;
  assign new_new_n12512__ = pi34 & pi38;
  assign new_new_n12513__ = pi33 & pi39;
  assign new_new_n12514__ = pi19 & pi53;
  assign new_new_n12515__ = ~new_new_n12513__ & ~new_new_n12514__;
  assign new_new_n12516__ = new_new_n12513__ & new_new_n12514__;
  assign new_new_n12517__ = ~new_new_n12515__ & ~new_new_n12516__;
  assign new_new_n12518__ = new_new_n12512__ & ~new_new_n12517__;
  assign new_new_n12519__ = ~new_new_n12512__ & new_new_n12517__;
  assign new_new_n12520__ = ~new_new_n12518__ & ~new_new_n12519__;
  assign new_new_n12521__ = new_new_n12511__ & new_new_n12520__;
  assign new_new_n12522__ = ~new_new_n12511__ & ~new_new_n12520__;
  assign new_new_n12523__ = ~new_new_n12521__ & ~new_new_n12522__;
  assign new_new_n12524__ = pi15 & pi57;
  assign new_new_n12525__ = pi14 & pi58;
  assign new_new_n12526__ = pi13 & pi59;
  assign new_new_n12527__ = ~new_new_n12525__ & ~new_new_n12526__;
  assign new_new_n12528__ = new_new_n12525__ & new_new_n12526__;
  assign new_new_n12529__ = ~new_new_n12527__ & ~new_new_n12528__;
  assign new_new_n12530__ = new_new_n12524__ & ~new_new_n12529__;
  assign new_new_n12531__ = ~new_new_n12524__ & new_new_n12529__;
  assign new_new_n12532__ = ~new_new_n12530__ & ~new_new_n12531__;
  assign new_new_n12533__ = ~new_new_n12523__ & new_new_n12532__;
  assign new_new_n12534__ = new_new_n12523__ & ~new_new_n12532__;
  assign new_new_n12535__ = ~new_new_n12533__ & ~new_new_n12534__;
  assign new_new_n12536__ = new_new_n12502__ & new_new_n12535__;
  assign new_new_n12537__ = ~new_new_n12502__ & ~new_new_n12535__;
  assign new_new_n12538__ = ~new_new_n12536__ & ~new_new_n12537__;
  assign new_new_n12539__ = new_new_n12484__ & new_new_n12538__;
  assign new_new_n12540__ = ~new_new_n12484__ & ~new_new_n12538__;
  assign new_new_n12541__ = ~new_new_n12539__ & ~new_new_n12540__;
  assign new_new_n12542__ = pi35 & pi37;
  assign new_new_n12543__ = pi22 & pi50;
  assign new_new_n12544__ = pi21 & pi51;
  assign new_new_n12545__ = ~new_new_n12543__ & ~new_new_n12544__;
  assign new_new_n12546__ = new_new_n12543__ & new_new_n12544__;
  assign new_new_n12547__ = ~new_new_n12545__ & ~new_new_n12546__;
  assign new_new_n12548__ = new_new_n12542__ & ~new_new_n12547__;
  assign new_new_n12549__ = ~new_new_n12542__ & new_new_n12547__;
  assign new_new_n12550__ = ~new_new_n12548__ & ~new_new_n12549__;
  assign new_new_n12551__ = pi20 & pi52;
  assign new_new_n12552__ = pi18 & pi54;
  assign new_new_n12553__ = pi17 & pi55;
  assign new_new_n12554__ = ~new_new_n12552__ & ~new_new_n12553__;
  assign new_new_n12555__ = new_new_n12552__ & new_new_n12553__;
  assign new_new_n12556__ = ~new_new_n12554__ & ~new_new_n12555__;
  assign new_new_n12557__ = new_new_n12551__ & ~new_new_n12556__;
  assign new_new_n12558__ = ~new_new_n12551__ & new_new_n12556__;
  assign new_new_n12559__ = ~new_new_n12557__ & ~new_new_n12558__;
  assign new_new_n12560__ = new_new_n12550__ & new_new_n12559__;
  assign new_new_n12561__ = ~new_new_n12550__ & ~new_new_n12559__;
  assign new_new_n12562__ = ~new_new_n12560__ & ~new_new_n12561__;
  assign new_new_n12563__ = ~new_new_n12314__ & ~new_new_n12319__;
  assign new_new_n12564__ = ~new_new_n12320__ & ~new_new_n12563__;
  assign new_new_n12565__ = pi11 & pi61;
  assign new_new_n12566__ = pi10 & pi62;
  assign new_new_n12567__ = pi09 & pi63;
  assign new_new_n12568__ = ~new_new_n12566__ & ~new_new_n12567__;
  assign new_new_n12569__ = new_new_n12566__ & new_new_n12567__;
  assign new_new_n12570__ = ~new_new_n12568__ & ~new_new_n12569__;
  assign new_new_n12571__ = new_new_n12565__ & ~new_new_n12570__;
  assign new_new_n12572__ = ~new_new_n12565__ & new_new_n12570__;
  assign new_new_n12573__ = ~new_new_n12571__ & ~new_new_n12572__;
  assign new_new_n12574__ = pi25 & pi47;
  assign new_new_n12575__ = pi24 & pi48;
  assign new_new_n12576__ = pi12 & pi60;
  assign new_new_n12577__ = ~new_new_n12575__ & ~new_new_n12576__;
  assign new_new_n12578__ = new_new_n12575__ & new_new_n12576__;
  assign new_new_n12579__ = ~new_new_n12577__ & ~new_new_n12578__;
  assign new_new_n12580__ = new_new_n12574__ & ~new_new_n12579__;
  assign new_new_n12581__ = ~new_new_n12574__ & new_new_n12579__;
  assign new_new_n12582__ = ~new_new_n12580__ & ~new_new_n12581__;
  assign new_new_n12583__ = new_new_n12573__ & new_new_n12582__;
  assign new_new_n12584__ = ~new_new_n12573__ & ~new_new_n12582__;
  assign new_new_n12585__ = ~new_new_n12583__ & ~new_new_n12584__;
  assign new_new_n12586__ = ~new_new_n12250__ & ~new_new_n12251__;
  assign new_new_n12587__ = new_new_n12250__ & new_new_n12251__;
  assign new_new_n12588__ = ~new_new_n12249__ & ~new_new_n12587__;
  assign new_new_n12589__ = ~new_new_n12586__ & ~new_new_n12588__;
  assign new_new_n12590__ = new_new_n12585__ & ~new_new_n12589__;
  assign new_new_n12591__ = ~new_new_n12585__ & new_new_n12589__;
  assign new_new_n12592__ = ~new_new_n12590__ & ~new_new_n12591__;
  assign new_new_n12593__ = new_new_n12564__ & new_new_n12592__;
  assign new_new_n12594__ = ~new_new_n12564__ & ~new_new_n12592__;
  assign new_new_n12595__ = ~new_new_n12593__ & ~new_new_n12594__;
  assign new_new_n12596__ = pi32 & pi40;
  assign new_new_n12597__ = pi16 & pi56;
  assign new_new_n12598__ = pi23 & pi49;
  assign new_new_n12599__ = ~new_new_n12597__ & ~new_new_n12598__;
  assign new_new_n12600__ = new_new_n12597__ & new_new_n12598__;
  assign new_new_n12601__ = ~new_new_n12599__ & ~new_new_n12600__;
  assign new_new_n12602__ = new_new_n12596__ & ~new_new_n12601__;
  assign new_new_n12603__ = ~new_new_n12596__ & new_new_n12601__;
  assign new_new_n12604__ = ~new_new_n12602__ & ~new_new_n12603__;
  assign new_new_n12605__ = new_new_n12595__ & ~new_new_n12604__;
  assign new_new_n12606__ = ~new_new_n12595__ & new_new_n12604__;
  assign new_new_n12607__ = ~new_new_n12605__ & ~new_new_n12606__;
  assign new_new_n12608__ = new_new_n12562__ & new_new_n12607__;
  assign new_new_n12609__ = ~new_new_n12562__ & ~new_new_n12607__;
  assign new_new_n12610__ = ~new_new_n12608__ & ~new_new_n12609__;
  assign new_new_n12611__ = ~new_new_n12541__ & new_new_n12610__;
  assign new_new_n12612__ = new_new_n12541__ & ~new_new_n12610__;
  assign new_new_n12613__ = ~new_new_n12611__ & ~new_new_n12612__;
  assign new_new_n12614__ = ~new_new_n12482__ & new_new_n12613__;
  assign new_new_n12615__ = new_new_n12482__ & ~new_new_n12613__;
  assign new_new_n12616__ = ~new_new_n12614__ & ~new_new_n12615__;
  assign new_new_n12617__ = ~new_new_n12308__ & new_new_n12362__;
  assign new_new_n12618__ = ~new_new_n12309__ & ~new_new_n12617__;
  assign new_new_n12619__ = ~new_new_n12616__ & ~new_new_n12618__;
  assign new_new_n12620__ = new_new_n12616__ & new_new_n12618__;
  assign new_new_n12621__ = ~new_new_n12619__ & ~new_new_n12620__;
  assign new_new_n12622__ = ~new_new_n12326__ & new_new_n12359__;
  assign new_new_n12623__ = ~new_new_n12325__ & ~new_new_n12622__;
  assign new_new_n12624__ = ~new_new_n12202__ & new_new_n12222__;
  assign new_new_n12625__ = ~new_new_n12201__ & ~new_new_n12624__;
  assign new_new_n12626__ = ~new_new_n12333__ & ~new_new_n12336__;
  assign new_new_n12627__ = ~new_new_n12332__ & ~new_new_n12626__;
  assign new_new_n12628__ = pi31 & pi41;
  assign new_new_n12629__ = pi29 & pi43;
  assign new_new_n12630__ = pi30 & pi42;
  assign new_new_n12631__ = ~new_new_n12629__ & ~new_new_n12630__;
  assign new_new_n12632__ = new_new_n12629__ & new_new_n12630__;
  assign new_new_n12633__ = ~new_new_n12631__ & ~new_new_n12632__;
  assign new_new_n12634__ = new_new_n12628__ & ~new_new_n12633__;
  assign new_new_n12635__ = ~new_new_n12628__ & new_new_n12633__;
  assign new_new_n12636__ = ~new_new_n12634__ & ~new_new_n12635__;
  assign new_new_n12637__ = ~new_new_n12627__ & new_new_n12636__;
  assign new_new_n12638__ = new_new_n12627__ & ~new_new_n12636__;
  assign new_new_n12639__ = ~new_new_n12637__ & ~new_new_n12638__;
  assign new_new_n12640__ = ~new_new_n12209__ & ~new_new_n12219__;
  assign new_new_n12641__ = ~new_new_n12208__ & ~new_new_n12640__;
  assign new_new_n12642__ = new_new_n12639__ & ~new_new_n12641__;
  assign new_new_n12643__ = ~new_new_n12639__ & new_new_n12641__;
  assign new_new_n12644__ = ~new_new_n12642__ & ~new_new_n12643__;
  assign new_new_n12645__ = new_new_n12625__ & ~new_new_n12644__;
  assign new_new_n12646__ = ~new_new_n12625__ & new_new_n12644__;
  assign new_new_n12647__ = ~new_new_n12645__ & ~new_new_n12646__;
  assign new_new_n12648__ = ~new_new_n12343__ & ~new_new_n12356__;
  assign new_new_n12649__ = ~new_new_n12342__ & ~new_new_n12648__;
  assign new_new_n12650__ = new_new_n12647__ & new_new_n12649__;
  assign new_new_n12651__ = ~new_new_n12647__ & ~new_new_n12649__;
  assign new_new_n12652__ = ~new_new_n12650__ & ~new_new_n12651__;
  assign new_new_n12653__ = ~new_new_n12623__ & ~new_new_n12652__;
  assign new_new_n12654__ = new_new_n12623__ & new_new_n12652__;
  assign new_new_n12655__ = ~new_new_n12653__ & ~new_new_n12654__;
  assign new_new_n12656__ = ~new_new_n12300__ & ~new_new_n12304__;
  assign new_new_n12657__ = ~new_new_n12301__ & ~new_new_n12656__;
  assign new_new_n12658__ = new_new_n12655__ & new_new_n12657__;
  assign new_new_n12659__ = ~new_new_n12655__ & ~new_new_n12657__;
  assign new_new_n12660__ = ~new_new_n12658__ & ~new_new_n12659__;
  assign new_new_n12661__ = new_new_n12621__ & ~new_new_n12660__;
  assign new_new_n12662__ = ~new_new_n12621__ & new_new_n12660__;
  assign new_new_n12663__ = ~new_new_n12661__ & ~new_new_n12662__;
  assign new_new_n12664__ = ~new_new_n12418__ & ~new_new_n12663__;
  assign new_new_n12665__ = new_new_n12160__ & new_new_n12366__;
  assign new_new_n12666__ = new_new_n12160__ & new_new_n12365__;
  assign new_new_n12667__ = ~new_new_n12160__ & ~new_new_n12365__;
  assign new_new_n12668__ = ~new_new_n12161__ & ~new_new_n12164__;
  assign new_new_n12669__ = ~new_new_n12667__ & new_new_n12668__;
  assign new_new_n12670__ = ~new_new_n12666__ & ~new_new_n12669__;
  assign new_new_n12671__ = new_new_n12402__ & ~new_new_n12670__;
  assign new_new_n12672__ = new_new_n12161__ & ~new_new_n12366__;
  assign new_new_n12673__ = new_new_n12164__ & new_new_n12667__;
  assign new_new_n12674__ = ~new_new_n12672__ & ~new_new_n12673__;
  assign new_new_n12675__ = ~new_new_n12402__ & ~new_new_n12674__;
  assign new_new_n12676__ = new_new_n12161__ & new_new_n12367__;
  assign new_new_n12677__ = ~new_new_n12665__ & ~new_new_n12676__;
  assign new_new_n12678__ = ~new_new_n12671__ & new_new_n12677__;
  assign new_new_n12679__ = ~new_new_n12675__ & new_new_n12678__;
  assign new_new_n12680__ = new_new_n12663__ & ~new_new_n12679__;
  assign po073 = new_new_n12664__ | new_new_n12680__;
  assign new_new_n12682__ = ~new_new_n12501__ & ~new_new_n12535__;
  assign new_new_n12683__ = ~new_new_n12500__ & ~new_new_n12682__;
  assign new_new_n12684__ = ~new_new_n12489__ & ~new_new_n12495__;
  assign new_new_n12685__ = pi33 & pi40;
  assign new_new_n12686__ = pi32 & pi41;
  assign new_new_n12687__ = pi31 & pi42;
  assign new_new_n12688__ = ~new_new_n12686__ & ~new_new_n12687__;
  assign new_new_n12689__ = new_new_n12686__ & new_new_n12687__;
  assign new_new_n12690__ = ~new_new_n12688__ & ~new_new_n12689__;
  assign new_new_n12691__ = new_new_n12685__ & ~new_new_n12690__;
  assign new_new_n12692__ = ~new_new_n12685__ & new_new_n12690__;
  assign new_new_n12693__ = ~new_new_n12691__ & ~new_new_n12692__;
  assign new_new_n12694__ = ~new_new_n12684__ & new_new_n12693__;
  assign new_new_n12695__ = new_new_n12684__ & ~new_new_n12693__;
  assign new_new_n12696__ = ~new_new_n12694__ & ~new_new_n12695__;
  assign new_new_n12697__ = ~new_new_n12461__ & ~new_new_n12467__;
  assign new_new_n12698__ = ~new_new_n12466__ & ~new_new_n12697__;
  assign new_new_n12699__ = new_new_n12696__ & new_new_n12698__;
  assign new_new_n12700__ = ~new_new_n12696__ & ~new_new_n12698__;
  assign new_new_n12701__ = ~new_new_n12699__ & ~new_new_n12700__;
  assign new_new_n12702__ = ~new_new_n12683__ & ~new_new_n12701__;
  assign new_new_n12703__ = new_new_n12683__ & new_new_n12701__;
  assign new_new_n12704__ = ~new_new_n12702__ & ~new_new_n12703__;
  assign new_new_n12705__ = ~new_new_n12457__ & new_new_n12471__;
  assign new_new_n12706__ = ~new_new_n12458__ & ~new_new_n12705__;
  assign new_new_n12707__ = new_new_n12704__ & ~new_new_n12706__;
  assign new_new_n12708__ = ~new_new_n12704__ & new_new_n12706__;
  assign new_new_n12709__ = ~new_new_n12707__ & ~new_new_n12708__;
  assign new_new_n12710__ = ~new_new_n12439__ & new_new_n12474__;
  assign new_new_n12711__ = ~new_new_n12438__ & ~new_new_n12710__;
  assign new_new_n12712__ = ~new_new_n12709__ & ~new_new_n12711__;
  assign new_new_n12713__ = new_new_n12709__ & new_new_n12711__;
  assign new_new_n12714__ = ~new_new_n12712__ & ~new_new_n12713__;
  assign new_new_n12715__ = ~new_new_n12540__ & new_new_n12610__;
  assign new_new_n12716__ = ~new_new_n12539__ & ~new_new_n12715__;
  assign new_new_n12717__ = new_new_n12714__ & new_new_n12716__;
  assign new_new_n12718__ = ~new_new_n12714__ & ~new_new_n12716__;
  assign new_new_n12719__ = ~new_new_n12717__ & ~new_new_n12718__;
  assign new_new_n12720__ = ~new_new_n12481__ & new_new_n12613__;
  assign new_new_n12721__ = ~new_new_n12480__ & ~new_new_n12720__;
  assign new_new_n12722__ = new_new_n12719__ & ~new_new_n12721__;
  assign new_new_n12723__ = ~new_new_n12719__ & new_new_n12721__;
  assign new_new_n12724__ = ~new_new_n12722__ & ~new_new_n12723__;
  assign new_new_n12725__ = ~new_new_n12654__ & ~new_new_n12658__;
  assign new_new_n12726__ = ~new_new_n12521__ & ~new_new_n12532__;
  assign new_new_n12727__ = ~new_new_n12522__ & ~new_new_n12726__;
  assign new_new_n12728__ = ~new_new_n12584__ & ~new_new_n12589__;
  assign new_new_n12729__ = ~new_new_n12583__ & ~new_new_n12728__;
  assign new_new_n12730__ = ~new_new_n12447__ & ~new_new_n12453__;
  assign new_new_n12731__ = ~new_new_n12448__ & ~new_new_n12730__;
  assign new_new_n12732__ = ~new_new_n12729__ & new_new_n12731__;
  assign new_new_n12733__ = new_new_n12729__ & ~new_new_n12731__;
  assign new_new_n12734__ = ~new_new_n12732__ & ~new_new_n12733__;
  assign new_new_n12735__ = new_new_n12727__ & ~new_new_n12734__;
  assign new_new_n12736__ = ~new_new_n12727__ & new_new_n12734__;
  assign new_new_n12737__ = ~new_new_n12735__ & ~new_new_n12736__;
  assign new_new_n12738__ = new_new_n12595__ & new_new_n12604__;
  assign new_new_n12739__ = new_new_n12559__ & ~new_new_n12738__;
  assign new_new_n12740__ = ~new_new_n12559__ & ~new_new_n12605__;
  assign new_new_n12741__ = new_new_n12550__ & ~new_new_n12739__;
  assign new_new_n12742__ = ~new_new_n12740__ & new_new_n12741__;
  assign new_new_n12743__ = new_new_n12559__ & ~new_new_n12605__;
  assign new_new_n12744__ = ~new_new_n12559__ & ~new_new_n12738__;
  assign new_new_n12745__ = ~new_new_n12550__ & ~new_new_n12743__;
  assign new_new_n12746__ = ~new_new_n12744__ & new_new_n12745__;
  assign new_new_n12747__ = ~new_new_n12593__ & ~new_new_n12742__;
  assign new_new_n12748__ = ~new_new_n12746__ & new_new_n12747__;
  assign new_new_n12749__ = new_new_n12737__ & new_new_n12748__;
  assign new_new_n12750__ = ~new_new_n12737__ & ~new_new_n12748__;
  assign new_new_n12751__ = ~new_new_n12749__ & ~new_new_n12750__;
  assign new_new_n12752__ = ~new_new_n12565__ & ~new_new_n12569__;
  assign new_new_n12753__ = ~new_new_n12568__ & ~new_new_n12752__;
  assign new_new_n12754__ = ~new_new_n12551__ & ~new_new_n12555__;
  assign new_new_n12755__ = ~new_new_n12554__ & ~new_new_n12754__;
  assign new_new_n12756__ = ~new_new_n12574__ & ~new_new_n12578__;
  assign new_new_n12757__ = ~new_new_n12577__ & ~new_new_n12756__;
  assign new_new_n12758__ = pi13 & pi60;
  assign new_new_n12759__ = ~new_new_n12512__ & ~new_new_n12516__;
  assign new_new_n12760__ = ~new_new_n12515__ & ~new_new_n12759__;
  assign new_new_n12761__ = ~new_new_n12542__ & ~new_new_n12546__;
  assign new_new_n12762__ = ~new_new_n12545__ & ~new_new_n12761__;
  assign new_new_n12763__ = new_new_n12760__ & new_new_n12762__;
  assign new_new_n12764__ = ~new_new_n12760__ & ~new_new_n12762__;
  assign new_new_n12765__ = ~new_new_n12763__ & ~new_new_n12764__;
  assign new_new_n12766__ = new_new_n12758__ & ~new_new_n12765__;
  assign new_new_n12767__ = ~new_new_n12758__ & new_new_n12765__;
  assign new_new_n12768__ = ~new_new_n12766__ & ~new_new_n12767__;
  assign new_new_n12769__ = ~new_new_n12560__ & ~new_new_n12604__;
  assign new_new_n12770__ = ~new_new_n12561__ & ~new_new_n12769__;
  assign new_new_n12771__ = ~new_new_n12768__ & ~new_new_n12770__;
  assign new_new_n12772__ = new_new_n12768__ & new_new_n12770__;
  assign new_new_n12773__ = ~new_new_n12771__ & ~new_new_n12772__;
  assign new_new_n12774__ = new_new_n12757__ & new_new_n12773__;
  assign new_new_n12775__ = ~new_new_n12757__ & ~new_new_n12773__;
  assign new_new_n12776__ = ~new_new_n12774__ & ~new_new_n12775__;
  assign new_new_n12777__ = new_new_n12755__ & ~new_new_n12776__;
  assign new_new_n12778__ = ~new_new_n12755__ & new_new_n12776__;
  assign new_new_n12779__ = ~new_new_n12777__ & ~new_new_n12778__;
  assign new_new_n12780__ = new_new_n12753__ & new_new_n12779__;
  assign new_new_n12781__ = ~new_new_n12753__ & ~new_new_n12779__;
  assign new_new_n12782__ = ~new_new_n12780__ & ~new_new_n12781__;
  assign new_new_n12783__ = new_new_n12751__ & new_new_n12782__;
  assign new_new_n12784__ = ~new_new_n12751__ & ~new_new_n12782__;
  assign new_new_n12785__ = ~new_new_n12783__ & ~new_new_n12784__;
  assign new_new_n12786__ = ~new_new_n12725__ & new_new_n12785__;
  assign new_new_n12787__ = new_new_n12725__ & ~new_new_n12785__;
  assign new_new_n12788__ = ~new_new_n12786__ & ~new_new_n12787__;
  assign new_new_n12789__ = new_new_n12422__ & ~new_new_n12432__;
  assign new_new_n12790__ = ~new_new_n12433__ & ~new_new_n12789__;
  assign new_new_n12791__ = pi23 & pi50;
  assign new_new_n12792__ = pi11 & pi62;
  assign new_new_n12793__ = ~new_new_n12791__ & ~new_new_n12792__;
  assign new_new_n12794__ = new_new_n12791__ & new_new_n12792__;
  assign new_new_n12795__ = ~new_new_n12793__ & ~new_new_n12794__;
  assign new_new_n12796__ = pi37 & ~new_new_n12795__;
  assign new_new_n12797__ = ~pi37 & ~new_new_n12794__;
  assign new_new_n12798__ = ~new_new_n12793__ & new_new_n12797__;
  assign new_new_n12799__ = ~new_new_n12796__ & ~new_new_n12798__;
  assign new_new_n12800__ = pi22 & pi51;
  assign new_new_n12801__ = pi20 & pi53;
  assign new_new_n12802__ = pi21 & pi52;
  assign new_new_n12803__ = ~new_new_n12801__ & ~new_new_n12802__;
  assign new_new_n12804__ = new_new_n12801__ & new_new_n12802__;
  assign new_new_n12805__ = ~new_new_n12803__ & ~new_new_n12804__;
  assign new_new_n12806__ = new_new_n12800__ & ~new_new_n12805__;
  assign new_new_n12807__ = ~new_new_n12800__ & new_new_n12805__;
  assign new_new_n12808__ = ~new_new_n12806__ & ~new_new_n12807__;
  assign new_new_n12809__ = new_new_n12799__ & new_new_n12808__;
  assign new_new_n12810__ = ~new_new_n12799__ & ~new_new_n12808__;
  assign new_new_n12811__ = ~new_new_n12809__ & ~new_new_n12810__;
  assign new_new_n12812__ = pi19 & pi54;
  assign new_new_n12813__ = pi18 & pi55;
  assign new_new_n12814__ = ~new_new_n12812__ & ~new_new_n12813__;
  assign new_new_n12815__ = new_new_n12812__ & new_new_n12813__;
  assign new_new_n12816__ = ~new_new_n12814__ & ~new_new_n12815__;
  assign new_new_n12817__ = new_new_n6794__ & ~new_new_n12816__;
  assign new_new_n12818__ = ~new_new_n6794__ & new_new_n12816__;
  assign new_new_n12819__ = ~new_new_n12817__ & ~new_new_n12818__;
  assign new_new_n12820__ = new_new_n12811__ & ~new_new_n12819__;
  assign new_new_n12821__ = ~new_new_n12811__ & new_new_n12819__;
  assign new_new_n12822__ = ~new_new_n12820__ & ~new_new_n12821__;
  assign new_new_n12823__ = new_new_n12790__ & ~new_new_n12822__;
  assign new_new_n12824__ = ~new_new_n12790__ & new_new_n12822__;
  assign new_new_n12825__ = ~new_new_n12823__ & ~new_new_n12824__;
  assign new_new_n12826__ = ~new_new_n12596__ & ~new_new_n12600__;
  assign new_new_n12827__ = ~new_new_n12599__ & ~new_new_n12826__;
  assign new_new_n12828__ = pi27 & pi46;
  assign new_new_n12829__ = pi26 & pi47;
  assign new_new_n12830__ = pi17 & pi56;
  assign new_new_n12831__ = ~new_new_n12829__ & ~new_new_n12830__;
  assign new_new_n12832__ = new_new_n12829__ & new_new_n12830__;
  assign new_new_n12833__ = ~new_new_n12831__ & ~new_new_n12832__;
  assign new_new_n12834__ = new_new_n12828__ & ~new_new_n12833__;
  assign new_new_n12835__ = ~new_new_n12828__ & new_new_n12833__;
  assign new_new_n12836__ = ~new_new_n12834__ & ~new_new_n12835__;
  assign new_new_n12837__ = pi16 & pi57;
  assign new_new_n12838__ = pi14 & pi59;
  assign new_new_n12839__ = pi15 & pi58;
  assign new_new_n12840__ = ~new_new_n12838__ & ~new_new_n12839__;
  assign new_new_n12841__ = new_new_n12838__ & new_new_n12839__;
  assign new_new_n12842__ = ~new_new_n12840__ & ~new_new_n12841__;
  assign new_new_n12843__ = new_new_n12837__ & ~new_new_n12842__;
  assign new_new_n12844__ = ~new_new_n12837__ & new_new_n12842__;
  assign new_new_n12845__ = ~new_new_n12843__ & ~new_new_n12844__;
  assign new_new_n12846__ = new_new_n12836__ & new_new_n12845__;
  assign new_new_n12847__ = ~new_new_n12836__ & ~new_new_n12845__;
  assign new_new_n12848__ = new_new_n12827__ & ~new_new_n12846__;
  assign new_new_n12849__ = ~new_new_n12847__ & ~new_new_n12848__;
  assign new_new_n12850__ = ~new_new_n12846__ & new_new_n12849__;
  assign new_new_n12851__ = ~new_new_n12827__ & ~new_new_n12850__;
  assign new_new_n12852__ = ~new_new_n12847__ & new_new_n12848__;
  assign new_new_n12853__ = ~new_new_n12851__ & ~new_new_n12852__;
  assign new_new_n12854__ = new_new_n12825__ & ~new_new_n12853__;
  assign new_new_n12855__ = ~new_new_n12825__ & new_new_n12853__;
  assign new_new_n12856__ = ~new_new_n12854__ & ~new_new_n12855__;
  assign new_new_n12857__ = ~new_new_n12637__ & ~new_new_n12641__;
  assign new_new_n12858__ = ~new_new_n12638__ & ~new_new_n12857__;
  assign new_new_n12859__ = ~new_new_n12628__ & ~new_new_n12632__;
  assign new_new_n12860__ = ~new_new_n12631__ & ~new_new_n12859__;
  assign new_new_n12861__ = ~new_new_n12524__ & ~new_new_n12528__;
  assign new_new_n12862__ = ~new_new_n12527__ & ~new_new_n12861__;
  assign new_new_n12863__ = ~new_new_n12503__ & ~new_new_n12507__;
  assign new_new_n12864__ = ~new_new_n12506__ & ~new_new_n12863__;
  assign new_new_n12865__ = ~new_new_n12862__ & ~new_new_n12864__;
  assign new_new_n12866__ = new_new_n12862__ & new_new_n12864__;
  assign new_new_n12867__ = ~new_new_n12865__ & ~new_new_n12866__;
  assign new_new_n12868__ = new_new_n12860__ & ~new_new_n12867__;
  assign new_new_n12869__ = ~new_new_n12860__ & new_new_n12867__;
  assign new_new_n12870__ = ~new_new_n12868__ & ~new_new_n12869__;
  assign new_new_n12871__ = new_new_n12858__ & new_new_n12870__;
  assign new_new_n12872__ = ~new_new_n12858__ & ~new_new_n12870__;
  assign new_new_n12873__ = ~new_new_n12871__ & ~new_new_n12872__;
  assign new_new_n12874__ = pi36 & pi37;
  assign new_new_n12875__ = pi34 & pi39;
  assign new_new_n12876__ = pi35 & pi38;
  assign new_new_n12877__ = ~new_new_n12875__ & ~new_new_n12876__;
  assign new_new_n12878__ = new_new_n12875__ & new_new_n12876__;
  assign new_new_n12879__ = ~new_new_n12877__ & ~new_new_n12878__;
  assign new_new_n12880__ = new_new_n12874__ & ~new_new_n12879__;
  assign new_new_n12881__ = ~new_new_n12874__ & new_new_n12879__;
  assign new_new_n12882__ = ~new_new_n12880__ & ~new_new_n12881__;
  assign new_new_n12883__ = pi10 & pi63;
  assign new_new_n12884__ = pi12 & pi61;
  assign new_new_n12885__ = ~new_new_n12883__ & ~new_new_n12884__;
  assign new_new_n12886__ = new_new_n12883__ & new_new_n12884__;
  assign new_new_n12887__ = ~new_new_n12885__ & ~new_new_n12886__;
  assign new_new_n12888__ = new_new_n6170__ & ~new_new_n12887__;
  assign new_new_n12889__ = ~new_new_n6170__ & new_new_n12887__;
  assign new_new_n12890__ = ~new_new_n12888__ & ~new_new_n12889__;
  assign new_new_n12891__ = ~new_new_n12882__ & ~new_new_n12890__;
  assign new_new_n12892__ = new_new_n12882__ & new_new_n12890__;
  assign new_new_n12893__ = ~new_new_n12891__ & ~new_new_n12892__;
  assign new_new_n12894__ = pi30 & pi43;
  assign new_new_n12895__ = pi29 & pi44;
  assign new_new_n12896__ = pi28 & pi45;
  assign new_new_n12897__ = ~new_new_n12895__ & ~new_new_n12896__;
  assign new_new_n12898__ = new_new_n12895__ & new_new_n12896__;
  assign new_new_n12899__ = ~new_new_n12897__ & ~new_new_n12898__;
  assign new_new_n12900__ = new_new_n12894__ & ~new_new_n12899__;
  assign new_new_n12901__ = ~new_new_n12894__ & new_new_n12899__;
  assign new_new_n12902__ = ~new_new_n12900__ & ~new_new_n12901__;
  assign new_new_n12903__ = new_new_n12893__ & new_new_n12902__;
  assign new_new_n12904__ = ~new_new_n12893__ & ~new_new_n12902__;
  assign new_new_n12905__ = ~new_new_n12903__ & ~new_new_n12904__;
  assign new_new_n12906__ = new_new_n12873__ & ~new_new_n12905__;
  assign new_new_n12907__ = ~new_new_n12873__ & new_new_n12905__;
  assign new_new_n12908__ = ~new_new_n12906__ & ~new_new_n12907__;
  assign new_new_n12909__ = new_new_n12856__ & ~new_new_n12908__;
  assign new_new_n12910__ = ~new_new_n12856__ & new_new_n12908__;
  assign new_new_n12911__ = ~new_new_n12909__ & ~new_new_n12910__;
  assign new_new_n12912__ = ~new_new_n12646__ & new_new_n12649__;
  assign new_new_n12913__ = ~new_new_n12645__ & ~new_new_n12912__;
  assign new_new_n12914__ = new_new_n12911__ & new_new_n12913__;
  assign new_new_n12915__ = ~new_new_n12911__ & ~new_new_n12913__;
  assign new_new_n12916__ = ~new_new_n12914__ & ~new_new_n12915__;
  assign new_new_n12917__ = new_new_n12788__ & ~new_new_n12916__;
  assign new_new_n12918__ = ~new_new_n12788__ & new_new_n12916__;
  assign new_new_n12919__ = ~new_new_n12917__ & ~new_new_n12918__;
  assign new_new_n12920__ = ~new_new_n12160__ & new_new_n12410__;
  assign new_new_n12921__ = new_new_n12663__ & ~new_new_n12920__;
  assign new_new_n12922__ = ~new_new_n12413__ & new_new_n12663__;
  assign new_new_n12923__ = ~new_new_n12412__ & ~new_new_n12922__;
  assign new_new_n12924__ = ~new_new_n12161__ & ~new_new_n12923__;
  assign new_new_n12925__ = new_new_n12160__ & ~new_new_n12410__;
  assign new_new_n12926__ = ~new_new_n12924__ & ~new_new_n12925__;
  assign new_new_n12927__ = ~new_new_n12921__ & new_new_n12926__;
  assign new_new_n12928__ = ~new_new_n12919__ & ~new_new_n12927__;
  assign new_new_n12929__ = new_new_n12919__ & new_new_n12927__;
  assign new_new_n12930__ = ~new_new_n12928__ & ~new_new_n12929__;
  assign new_new_n12931__ = ~new_new_n12620__ & new_new_n12660__;
  assign new_new_n12932__ = ~new_new_n12619__ & ~new_new_n12931__;
  assign new_new_n12933__ = new_new_n12930__ & ~new_new_n12932__;
  assign new_new_n12934__ = ~new_new_n12930__ & new_new_n12932__;
  assign new_new_n12935__ = ~new_new_n12933__ & ~new_new_n12934__;
  assign new_new_n12936__ = new_new_n12724__ & new_new_n12935__;
  assign new_new_n12937__ = ~new_new_n12724__ & ~new_new_n12935__;
  assign po074 = new_new_n12936__ | new_new_n12937__;
  assign new_new_n12939__ = ~new_new_n12749__ & new_new_n12782__;
  assign new_new_n12940__ = ~new_new_n12750__ & ~new_new_n12939__;
  assign new_new_n12941__ = ~new_new_n12910__ & ~new_new_n12913__;
  assign new_new_n12942__ = ~new_new_n12909__ & ~new_new_n12941__;
  assign new_new_n12943__ = ~new_new_n12940__ & ~new_new_n12942__;
  assign new_new_n12944__ = new_new_n12940__ & new_new_n12942__;
  assign new_new_n12945__ = ~new_new_n12943__ & ~new_new_n12944__;
  assign new_new_n12946__ = new_new_n12755__ & ~new_new_n12757__;
  assign new_new_n12947__ = ~new_new_n12755__ & new_new_n12757__;
  assign new_new_n12948__ = ~new_new_n12946__ & ~new_new_n12947__;
  assign new_new_n12949__ = ~new_new_n12753__ & new_new_n12948__;
  assign new_new_n12950__ = new_new_n12753__ & ~new_new_n12948__;
  assign new_new_n12951__ = ~new_new_n12949__ & ~new_new_n12950__;
  assign new_new_n12952__ = new_new_n12773__ & new_new_n12951__;
  assign new_new_n12953__ = ~new_new_n12771__ & ~new_new_n12952__;
  assign new_new_n12954__ = ~new_new_n12758__ & ~new_new_n12763__;
  assign new_new_n12955__ = ~new_new_n12764__ & ~new_new_n12954__;
  assign new_new_n12956__ = ~new_new_n12755__ & ~new_new_n12757__;
  assign new_new_n12957__ = new_new_n12755__ & new_new_n12757__;
  assign new_new_n12958__ = ~new_new_n12753__ & ~new_new_n12957__;
  assign new_new_n12959__ = ~new_new_n12956__ & ~new_new_n12958__;
  assign new_new_n12960__ = new_new_n12955__ & new_new_n12959__;
  assign new_new_n12961__ = ~new_new_n12955__ & ~new_new_n12959__;
  assign new_new_n12962__ = ~new_new_n12960__ & ~new_new_n12961__;
  assign new_new_n12963__ = ~new_new_n12849__ & new_new_n12962__;
  assign new_new_n12964__ = new_new_n12849__ & ~new_new_n12962__;
  assign new_new_n12965__ = ~new_new_n12963__ & ~new_new_n12964__;
  assign new_new_n12966__ = new_new_n12727__ & ~new_new_n12733__;
  assign new_new_n12967__ = ~new_new_n12732__ & ~new_new_n12966__;
  assign new_new_n12968__ = new_new_n12965__ & new_new_n12967__;
  assign new_new_n12969__ = ~new_new_n12965__ & ~new_new_n12967__;
  assign new_new_n12970__ = ~new_new_n12968__ & ~new_new_n12969__;
  assign new_new_n12971__ = new_new_n12953__ & new_new_n12970__;
  assign new_new_n12972__ = ~new_new_n12953__ & ~new_new_n12970__;
  assign new_new_n12973__ = ~new_new_n12971__ & ~new_new_n12972__;
  assign new_new_n12974__ = new_new_n12945__ & ~new_new_n12973__;
  assign new_new_n12975__ = ~new_new_n12945__ & new_new_n12973__;
  assign new_new_n12976__ = ~new_new_n12974__ & ~new_new_n12975__;
  assign new_new_n12977__ = ~new_new_n12713__ & ~new_new_n12716__;
  assign new_new_n12978__ = ~new_new_n12712__ & ~new_new_n12977__;
  assign new_new_n12979__ = ~new_new_n12695__ & ~new_new_n12698__;
  assign new_new_n12980__ = ~new_new_n12694__ & ~new_new_n12979__;
  assign new_new_n12981__ = ~new_new_n12685__ & ~new_new_n12689__;
  assign new_new_n12982__ = ~new_new_n12688__ & ~new_new_n12981__;
  assign new_new_n12983__ = ~new_new_n12874__ & ~new_new_n12878__;
  assign new_new_n12984__ = ~new_new_n12877__ & ~new_new_n12983__;
  assign new_new_n12985__ = pi16 & pi58;
  assign new_new_n12986__ = pi15 & pi59;
  assign new_new_n12987__ = pi14 & pi60;
  assign new_new_n12988__ = ~new_new_n12986__ & ~new_new_n12987__;
  assign new_new_n12989__ = new_new_n12986__ & new_new_n12987__;
  assign new_new_n12990__ = ~new_new_n12988__ & ~new_new_n12989__;
  assign new_new_n12991__ = new_new_n12985__ & ~new_new_n12990__;
  assign new_new_n12992__ = ~new_new_n12985__ & new_new_n12990__;
  assign new_new_n12993__ = ~new_new_n12991__ & ~new_new_n12992__;
  assign new_new_n12994__ = ~new_new_n12984__ & new_new_n12993__;
  assign new_new_n12995__ = new_new_n12984__ & ~new_new_n12993__;
  assign new_new_n12996__ = ~new_new_n12994__ & ~new_new_n12995__;
  assign new_new_n12997__ = new_new_n12982__ & new_new_n12996__;
  assign new_new_n12998__ = ~new_new_n12982__ & ~new_new_n12996__;
  assign new_new_n12999__ = ~new_new_n12997__ & ~new_new_n12998__;
  assign new_new_n13000__ = new_new_n12980__ & new_new_n12999__;
  assign new_new_n13001__ = ~new_new_n12810__ & new_new_n12819__;
  assign new_new_n13002__ = ~new_new_n12980__ & ~new_new_n12999__;
  assign new_new_n13003__ = ~new_new_n12809__ & ~new_new_n13001__;
  assign new_new_n13004__ = ~new_new_n13002__ & new_new_n13003__;
  assign new_new_n13005__ = ~new_new_n13000__ & new_new_n13004__;
  assign new_new_n13006__ = new_new_n12808__ & new_new_n13000__;
  assign new_new_n13007__ = new_new_n12819__ & new_new_n13002__;
  assign new_new_n13008__ = ~new_new_n13006__ & ~new_new_n13007__;
  assign new_new_n13009__ = new_new_n12799__ & ~new_new_n13008__;
  assign new_new_n13010__ = new_new_n12808__ & new_new_n13002__;
  assign new_new_n13011__ = new_new_n12811__ & new_new_n13000__;
  assign new_new_n13012__ = ~new_new_n13010__ & ~new_new_n13011__;
  assign new_new_n13013__ = new_new_n12822__ & ~new_new_n13012__;
  assign new_new_n13014__ = ~new_new_n13005__ & ~new_new_n13009__;
  assign new_new_n13015__ = ~new_new_n13013__ & new_new_n13014__;
  assign new_new_n13016__ = ~new_new_n12871__ & ~new_new_n12905__;
  assign new_new_n13017__ = ~new_new_n12872__ & ~new_new_n13016__;
  assign new_new_n13018__ = ~new_new_n13015__ & new_new_n13017__;
  assign new_new_n13019__ = new_new_n13015__ & ~new_new_n13017__;
  assign new_new_n13020__ = ~new_new_n13018__ & ~new_new_n13019__;
  assign new_new_n13021__ = ~new_new_n12824__ & ~new_new_n12853__;
  assign new_new_n13022__ = ~new_new_n12823__ & ~new_new_n13021__;
  assign new_new_n13023__ = new_new_n13020__ & new_new_n13022__;
  assign new_new_n13024__ = ~new_new_n13020__ & ~new_new_n13022__;
  assign new_new_n13025__ = ~new_new_n13023__ & ~new_new_n13024__;
  assign new_new_n13026__ = new_new_n12978__ & ~new_new_n13025__;
  assign new_new_n13027__ = ~new_new_n12978__ & new_new_n13025__;
  assign new_new_n13028__ = ~new_new_n13026__ & ~new_new_n13027__;
  assign new_new_n13029__ = ~new_new_n12892__ & ~new_new_n12902__;
  assign new_new_n13030__ = ~new_new_n12891__ & ~new_new_n13029__;
  assign new_new_n13031__ = ~new_new_n12837__ & ~new_new_n12841__;
  assign new_new_n13032__ = ~new_new_n12840__ & ~new_new_n13031__;
  assign new_new_n13033__ = ~new_new_n12894__ & ~new_new_n12898__;
  assign new_new_n13034__ = ~new_new_n12897__ & ~new_new_n13033__;
  assign new_new_n13035__ = ~new_new_n12828__ & ~new_new_n12832__;
  assign new_new_n13036__ = ~new_new_n12831__ & ~new_new_n13035__;
  assign new_new_n13037__ = ~new_new_n13034__ & ~new_new_n13036__;
  assign new_new_n13038__ = new_new_n13034__ & new_new_n13036__;
  assign new_new_n13039__ = ~new_new_n13037__ & ~new_new_n13038__;
  assign new_new_n13040__ = new_new_n13032__ & ~new_new_n13039__;
  assign new_new_n13041__ = ~new_new_n13032__ & new_new_n13039__;
  assign new_new_n13042__ = ~new_new_n13040__ & ~new_new_n13041__;
  assign new_new_n13043__ = new_new_n13030__ & new_new_n13042__;
  assign new_new_n13044__ = ~new_new_n13030__ & ~new_new_n13042__;
  assign new_new_n13045__ = ~new_new_n13043__ & ~new_new_n13044__;
  assign new_new_n13046__ = ~new_new_n6170__ & ~new_new_n12886__;
  assign new_new_n13047__ = ~new_new_n12885__ & ~new_new_n13046__;
  assign new_new_n13048__ = ~new_new_n6794__ & ~new_new_n12815__;
  assign new_new_n13049__ = ~new_new_n12814__ & ~new_new_n13048__;
  assign new_new_n13050__ = ~new_new_n12800__ & ~new_new_n12804__;
  assign new_new_n13051__ = ~new_new_n12803__ & ~new_new_n13050__;
  assign new_new_n13052__ = new_new_n13049__ & new_new_n13051__;
  assign new_new_n13053__ = ~new_new_n13049__ & ~new_new_n13051__;
  assign new_new_n13054__ = ~new_new_n13047__ & ~new_new_n13052__;
  assign new_new_n13055__ = ~new_new_n13053__ & ~new_new_n13054__;
  assign new_new_n13056__ = ~new_new_n13052__ & new_new_n13055__;
  assign new_new_n13057__ = new_new_n13047__ & ~new_new_n13056__;
  assign new_new_n13058__ = ~new_new_n13053__ & new_new_n13054__;
  assign new_new_n13059__ = ~new_new_n13057__ & ~new_new_n13058__;
  assign new_new_n13060__ = new_new_n13045__ & ~new_new_n13059__;
  assign new_new_n13061__ = ~new_new_n13045__ & new_new_n13059__;
  assign new_new_n13062__ = ~new_new_n13060__ & ~new_new_n13061__;
  assign new_new_n13063__ = ~new_new_n12703__ & ~new_new_n12706__;
  assign new_new_n13064__ = ~new_new_n12702__ & ~new_new_n13063__;
  assign new_new_n13065__ = pi28 & pi46;
  assign new_new_n13066__ = pi27 & pi47;
  assign new_new_n13067__ = pi26 & pi48;
  assign new_new_n13068__ = ~new_new_n13066__ & ~new_new_n13067__;
  assign new_new_n13069__ = new_new_n13066__ & new_new_n13067__;
  assign new_new_n13070__ = ~new_new_n13068__ & ~new_new_n13069__;
  assign new_new_n13071__ = new_new_n13065__ & ~new_new_n13070__;
  assign new_new_n13072__ = ~new_new_n13065__ & new_new_n13070__;
  assign new_new_n13073__ = ~new_new_n13071__ & ~new_new_n13072__;
  assign new_new_n13074__ = pi33 & pi41;
  assign new_new_n13075__ = pi25 & pi49;
  assign new_new_n13076__ = pi18 & pi56;
  assign new_new_n13077__ = ~new_new_n13075__ & ~new_new_n13076__;
  assign new_new_n13078__ = new_new_n13075__ & new_new_n13076__;
  assign new_new_n13079__ = ~new_new_n13077__ & ~new_new_n13078__;
  assign new_new_n13080__ = new_new_n13074__ & ~new_new_n13079__;
  assign new_new_n13081__ = ~new_new_n13074__ & new_new_n13079__;
  assign new_new_n13082__ = ~new_new_n13080__ & ~new_new_n13081__;
  assign new_new_n13083__ = new_new_n13073__ & new_new_n13082__;
  assign new_new_n13084__ = ~new_new_n13073__ & ~new_new_n13082__;
  assign new_new_n13085__ = ~new_new_n13083__ & ~new_new_n13084__;
  assign new_new_n13086__ = pi32 & pi42;
  assign new_new_n13087__ = pi31 & pi43;
  assign new_new_n13088__ = pi11 & pi63;
  assign new_new_n13089__ = ~new_new_n13087__ & ~new_new_n13088__;
  assign new_new_n13090__ = new_new_n13087__ & new_new_n13088__;
  assign new_new_n13091__ = ~new_new_n13089__ & ~new_new_n13090__;
  assign new_new_n13092__ = new_new_n13086__ & ~new_new_n13091__;
  assign new_new_n13093__ = ~new_new_n13086__ & new_new_n13091__;
  assign new_new_n13094__ = ~new_new_n13092__ & ~new_new_n13093__;
  assign new_new_n13095__ = new_new_n13085__ & ~new_new_n13094__;
  assign new_new_n13096__ = ~new_new_n13085__ & new_new_n13094__;
  assign new_new_n13097__ = ~new_new_n13095__ & ~new_new_n13096__;
  assign new_new_n13098__ = pi22 & pi52;
  assign new_new_n13099__ = pi21 & pi53;
  assign new_new_n13100__ = pi19 & pi55;
  assign new_new_n13101__ = ~new_new_n13099__ & ~new_new_n13100__;
  assign new_new_n13102__ = new_new_n13099__ & new_new_n13100__;
  assign new_new_n13103__ = ~new_new_n13101__ & ~new_new_n13102__;
  assign new_new_n13104__ = new_new_n13098__ & ~new_new_n13103__;
  assign new_new_n13105__ = ~new_new_n13098__ & new_new_n13103__;
  assign new_new_n13106__ = ~new_new_n13104__ & ~new_new_n13105__;
  assign new_new_n13107__ = pi35 & pi39;
  assign new_new_n13108__ = pi34 & pi40;
  assign new_new_n13109__ = pi20 & pi54;
  assign new_new_n13110__ = ~new_new_n13108__ & ~new_new_n13109__;
  assign new_new_n13111__ = new_new_n13108__ & new_new_n13109__;
  assign new_new_n13112__ = ~new_new_n13110__ & ~new_new_n13111__;
  assign new_new_n13113__ = new_new_n13107__ & ~new_new_n13112__;
  assign new_new_n13114__ = ~new_new_n13107__ & new_new_n13112__;
  assign new_new_n13115__ = ~new_new_n13113__ & ~new_new_n13114__;
  assign new_new_n13116__ = ~new_new_n13106__ & ~new_new_n13115__;
  assign new_new_n13117__ = new_new_n13106__ & new_new_n13115__;
  assign new_new_n13118__ = ~new_new_n13116__ & ~new_new_n13117__;
  assign new_new_n13119__ = pi36 & pi38;
  assign new_new_n13120__ = pi24 & pi50;
  assign new_new_n13121__ = pi23 & pi51;
  assign new_new_n13122__ = ~new_new_n13120__ & ~new_new_n13121__;
  assign new_new_n13123__ = new_new_n13120__ & new_new_n13121__;
  assign new_new_n13124__ = ~new_new_n13122__ & ~new_new_n13123__;
  assign new_new_n13125__ = new_new_n13119__ & ~new_new_n13124__;
  assign new_new_n13126__ = ~new_new_n13119__ & new_new_n13124__;
  assign new_new_n13127__ = ~new_new_n13125__ & ~new_new_n13126__;
  assign new_new_n13128__ = ~new_new_n13118__ & new_new_n13127__;
  assign new_new_n13129__ = new_new_n13118__ & ~new_new_n13127__;
  assign new_new_n13130__ = ~new_new_n13128__ & ~new_new_n13129__;
  assign new_new_n13131__ = ~new_new_n12860__ & ~new_new_n12866__;
  assign new_new_n13132__ = ~new_new_n12865__ & ~new_new_n13131__;
  assign new_new_n13133__ = pi13 & pi61;
  assign new_new_n13134__ = pi12 & pi62;
  assign new_new_n13135__ = ~new_new_n13133__ & ~new_new_n13134__;
  assign new_new_n13136__ = new_new_n13133__ & new_new_n13134__;
  assign new_new_n13137__ = ~new_new_n13135__ & ~new_new_n13136__;
  assign new_new_n13138__ = ~new_new_n12793__ & ~new_new_n12797__;
  assign new_new_n13139__ = ~new_new_n13137__ & new_new_n13138__;
  assign new_new_n13140__ = new_new_n13137__ & ~new_new_n13138__;
  assign new_new_n13141__ = ~new_new_n13139__ & ~new_new_n13140__;
  assign new_new_n13142__ = pi30 & pi44;
  assign new_new_n13143__ = pi29 & pi45;
  assign new_new_n13144__ = pi17 & pi57;
  assign new_new_n13145__ = ~new_new_n13143__ & ~new_new_n13144__;
  assign new_new_n13146__ = new_new_n13143__ & new_new_n13144__;
  assign new_new_n13147__ = ~new_new_n13145__ & ~new_new_n13146__;
  assign new_new_n13148__ = new_new_n13142__ & ~new_new_n13147__;
  assign new_new_n13149__ = ~new_new_n13142__ & new_new_n13147__;
  assign new_new_n13150__ = ~new_new_n13148__ & ~new_new_n13149__;
  assign new_new_n13151__ = new_new_n13141__ & new_new_n13150__;
  assign new_new_n13152__ = ~new_new_n13141__ & ~new_new_n13150__;
  assign new_new_n13153__ = ~new_new_n13151__ & ~new_new_n13152__;
  assign new_new_n13154__ = new_new_n13132__ & new_new_n13153__;
  assign new_new_n13155__ = ~new_new_n13132__ & ~new_new_n13153__;
  assign new_new_n13156__ = ~new_new_n13154__ & ~new_new_n13155__;
  assign new_new_n13157__ = ~new_new_n13130__ & ~new_new_n13156__;
  assign new_new_n13158__ = new_new_n13130__ & new_new_n13156__;
  assign new_new_n13159__ = ~new_new_n13157__ & ~new_new_n13158__;
  assign new_new_n13160__ = new_new_n13097__ & new_new_n13159__;
  assign new_new_n13161__ = ~new_new_n13097__ & ~new_new_n13159__;
  assign new_new_n13162__ = ~new_new_n13160__ & ~new_new_n13161__;
  assign new_new_n13163__ = ~new_new_n13064__ & ~new_new_n13162__;
  assign new_new_n13164__ = new_new_n13064__ & new_new_n13162__;
  assign new_new_n13165__ = new_new_n13062__ & ~new_new_n13163__;
  assign new_new_n13166__ = ~new_new_n13164__ & ~new_new_n13165__;
  assign new_new_n13167__ = ~new_new_n13163__ & new_new_n13166__;
  assign new_new_n13168__ = ~new_new_n13062__ & ~new_new_n13167__;
  assign new_new_n13169__ = ~new_new_n13164__ & new_new_n13165__;
  assign new_new_n13170__ = ~new_new_n13168__ & ~new_new_n13169__;
  assign new_new_n13171__ = new_new_n13028__ & ~new_new_n13170__;
  assign new_new_n13172__ = ~new_new_n13028__ & new_new_n13170__;
  assign new_new_n13173__ = ~new_new_n13171__ & ~new_new_n13172__;
  assign new_new_n13174__ = new_new_n12976__ & ~new_new_n13173__;
  assign new_new_n13175__ = ~new_new_n12976__ & new_new_n13173__;
  assign new_new_n13176__ = ~new_new_n13174__ & ~new_new_n13175__;
  assign new_new_n13177__ = ~new_new_n12786__ & new_new_n12916__;
  assign new_new_n13178__ = ~new_new_n12787__ & ~new_new_n13177__;
  assign new_new_n13179__ = new_new_n13176__ & ~new_new_n13178__;
  assign new_new_n13180__ = ~new_new_n13176__ & new_new_n13178__;
  assign new_new_n13181__ = ~new_new_n13179__ & ~new_new_n13180__;
  assign new_new_n13182__ = ~new_new_n12721__ & ~new_new_n12932__;
  assign new_new_n13183__ = new_new_n12721__ & new_new_n12932__;
  assign new_new_n13184__ = ~new_new_n13182__ & ~new_new_n13183__;
  assign new_new_n13185__ = ~new_new_n12724__ & ~new_new_n13184__;
  assign new_new_n13186__ = new_new_n12930__ & ~new_new_n13185__;
  assign new_new_n13187__ = ~new_new_n12723__ & ~new_new_n12932__;
  assign new_new_n13188__ = ~new_new_n12722__ & ~new_new_n13187__;
  assign new_new_n13189__ = ~new_new_n12929__ & new_new_n13188__;
  assign new_new_n13190__ = ~new_new_n12928__ & ~new_new_n13188__;
  assign new_new_n13191__ = ~new_new_n13189__ & ~new_new_n13190__;
  assign new_new_n13192__ = ~new_new_n13181__ & ~new_new_n13186__;
  assign new_new_n13193__ = ~new_new_n13191__ & new_new_n13192__;
  assign new_new_n13194__ = new_new_n12929__ & ~new_new_n12932__;
  assign new_new_n13195__ = ~new_new_n12721__ & new_new_n13194__;
  assign new_new_n13196__ = ~new_new_n12929__ & new_new_n12932__;
  assign new_new_n13197__ = ~new_new_n12721__ & ~new_new_n12928__;
  assign new_new_n13198__ = ~new_new_n13196__ & new_new_n13197__;
  assign new_new_n13199__ = ~new_new_n13194__ & ~new_new_n13198__;
  assign new_new_n13200__ = new_new_n12719__ & ~new_new_n13199__;
  assign new_new_n13201__ = new_new_n12928__ & new_new_n13183__;
  assign new_new_n13202__ = new_new_n12928__ & ~new_new_n13182__;
  assign new_new_n13203__ = new_new_n12721__ & new_new_n13196__;
  assign new_new_n13204__ = ~new_new_n13202__ & ~new_new_n13203__;
  assign new_new_n13205__ = ~new_new_n12719__ & ~new_new_n13204__;
  assign new_new_n13206__ = new_new_n13181__ & ~new_new_n13201__;
  assign new_new_n13207__ = ~new_new_n13195__ & new_new_n13206__;
  assign new_new_n13208__ = ~new_new_n13200__ & new_new_n13207__;
  assign new_new_n13209__ = ~new_new_n13205__ & new_new_n13208__;
  assign po075 = ~new_new_n13193__ & ~new_new_n13209__;
  assign new_new_n13211__ = ~new_new_n12953__ & ~new_new_n12969__;
  assign new_new_n13212__ = ~new_new_n12968__ & ~new_new_n13211__;
  assign new_new_n13213__ = ~new_new_n13117__ & ~new_new_n13127__;
  assign new_new_n13214__ = ~new_new_n13116__ & ~new_new_n13213__;
  assign new_new_n13215__ = ~new_new_n13083__ & ~new_new_n13094__;
  assign new_new_n13216__ = ~new_new_n13084__ & ~new_new_n13215__;
  assign new_new_n13217__ = ~new_new_n13142__ & ~new_new_n13146__;
  assign new_new_n13218__ = ~new_new_n13145__ & ~new_new_n13217__;
  assign new_new_n13219__ = ~new_new_n12985__ & ~new_new_n12989__;
  assign new_new_n13220__ = ~new_new_n12988__ & ~new_new_n13219__;
  assign new_new_n13221__ = ~new_new_n13065__ & ~new_new_n13069__;
  assign new_new_n13222__ = ~new_new_n13068__ & ~new_new_n13221__;
  assign new_new_n13223__ = new_new_n13220__ & new_new_n13222__;
  assign new_new_n13224__ = ~new_new_n13220__ & ~new_new_n13222__;
  assign new_new_n13225__ = ~new_new_n13223__ & ~new_new_n13224__;
  assign new_new_n13226__ = new_new_n13218__ & ~new_new_n13225__;
  assign new_new_n13227__ = ~new_new_n13218__ & new_new_n13225__;
  assign new_new_n13228__ = ~new_new_n13226__ & ~new_new_n13227__;
  assign new_new_n13229__ = new_new_n13216__ & new_new_n13228__;
  assign new_new_n13230__ = ~new_new_n13216__ & ~new_new_n13228__;
  assign new_new_n13231__ = ~new_new_n13229__ & ~new_new_n13230__;
  assign new_new_n13232__ = new_new_n13214__ & new_new_n13231__;
  assign new_new_n13233__ = ~new_new_n13214__ & ~new_new_n13231__;
  assign new_new_n13234__ = ~new_new_n13232__ & ~new_new_n13233__;
  assign new_new_n13235__ = new_new_n13212__ & new_new_n13234__;
  assign new_new_n13236__ = ~new_new_n13212__ & ~new_new_n13234__;
  assign new_new_n13237__ = ~new_new_n13235__ & ~new_new_n13236__;
  assign new_new_n13238__ = ~new_new_n12960__ & ~new_new_n12963__;
  assign new_new_n13239__ = pi13 & pi62;
  assign new_new_n13240__ = ~pi37 & pi38;
  assign new_new_n13241__ = ~new_new_n13239__ & new_new_n13240__;
  assign new_new_n13242__ = new_new_n13239__ & ~new_new_n13240__;
  assign new_new_n13243__ = ~new_new_n13241__ & ~new_new_n13242__;
  assign new_new_n13244__ = pi36 & pi39;
  assign new_new_n13245__ = pi35 & pi40;
  assign new_new_n13246__ = pi23 & pi52;
  assign new_new_n13247__ = ~new_new_n13245__ & ~new_new_n13246__;
  assign new_new_n13248__ = new_new_n13245__ & new_new_n13246__;
  assign new_new_n13249__ = ~new_new_n13247__ & ~new_new_n13248__;
  assign new_new_n13250__ = new_new_n13244__ & ~new_new_n13249__;
  assign new_new_n13251__ = ~new_new_n13244__ & new_new_n13249__;
  assign new_new_n13252__ = ~new_new_n13250__ & ~new_new_n13251__;
  assign new_new_n13253__ = pi30 & pi45;
  assign new_new_n13254__ = pi12 & pi63;
  assign new_new_n13255__ = pi19 & pi56;
  assign new_new_n13256__ = ~new_new_n13254__ & ~new_new_n13255__;
  assign new_new_n13257__ = new_new_n13254__ & new_new_n13255__;
  assign new_new_n13258__ = ~new_new_n13256__ & ~new_new_n13257__;
  assign new_new_n13259__ = new_new_n13253__ & ~new_new_n13258__;
  assign new_new_n13260__ = ~new_new_n13253__ & new_new_n13258__;
  assign new_new_n13261__ = ~new_new_n13259__ & ~new_new_n13260__;
  assign new_new_n13262__ = new_new_n13252__ & new_new_n13261__;
  assign new_new_n13263__ = ~new_new_n13252__ & ~new_new_n13261__;
  assign new_new_n13264__ = ~new_new_n13262__ & ~new_new_n13263__;
  assign new_new_n13265__ = new_new_n13243__ & new_new_n13264__;
  assign new_new_n13266__ = ~new_new_n13243__ & ~new_new_n13264__;
  assign new_new_n13267__ = ~new_new_n13265__ & ~new_new_n13266__;
  assign new_new_n13268__ = ~new_new_n13238__ & ~new_new_n13267__;
  assign new_new_n13269__ = new_new_n13238__ & new_new_n13267__;
  assign new_new_n13270__ = ~new_new_n13268__ & ~new_new_n13269__;
  assign new_new_n13271__ = pi16 & pi59;
  assign new_new_n13272__ = pi15 & pi60;
  assign new_new_n13273__ = pi14 & pi61;
  assign new_new_n13274__ = ~new_new_n13272__ & ~new_new_n13273__;
  assign new_new_n13275__ = new_new_n13272__ & new_new_n13273__;
  assign new_new_n13276__ = ~new_new_n13274__ & ~new_new_n13275__;
  assign new_new_n13277__ = new_new_n13271__ & ~new_new_n13276__;
  assign new_new_n13278__ = ~new_new_n13271__ & new_new_n13276__;
  assign new_new_n13279__ = ~new_new_n13277__ & ~new_new_n13278__;
  assign new_new_n13280__ = pi29 & pi46;
  assign new_new_n13281__ = pi27 & pi48;
  assign new_new_n13282__ = pi28 & pi47;
  assign new_new_n13283__ = ~new_new_n13281__ & ~new_new_n13282__;
  assign new_new_n13284__ = new_new_n13281__ & new_new_n13282__;
  assign new_new_n13285__ = ~new_new_n13283__ & ~new_new_n13284__;
  assign new_new_n13286__ = new_new_n13280__ & ~new_new_n13285__;
  assign new_new_n13287__ = ~new_new_n13280__ & new_new_n13285__;
  assign new_new_n13288__ = ~new_new_n13286__ & ~new_new_n13287__;
  assign new_new_n13289__ = new_new_n13279__ & new_new_n13288__;
  assign new_new_n13290__ = ~new_new_n13279__ & ~new_new_n13288__;
  assign new_new_n13291__ = ~new_new_n13289__ & ~new_new_n13290__;
  assign new_new_n13292__ = pi26 & pi49;
  assign new_new_n13293__ = pi18 & pi57;
  assign new_new_n13294__ = pi17 & pi58;
  assign new_new_n13295__ = ~new_new_n13293__ & ~new_new_n13294__;
  assign new_new_n13296__ = new_new_n13293__ & new_new_n13294__;
  assign new_new_n13297__ = ~new_new_n13295__ & ~new_new_n13296__;
  assign new_new_n13298__ = new_new_n13292__ & ~new_new_n13297__;
  assign new_new_n13299__ = ~new_new_n13292__ & new_new_n13297__;
  assign new_new_n13300__ = ~new_new_n13298__ & ~new_new_n13299__;
  assign new_new_n13301__ = ~new_new_n13291__ & new_new_n13300__;
  assign new_new_n13302__ = new_new_n13291__ & ~new_new_n13300__;
  assign new_new_n13303__ = ~new_new_n13301__ & ~new_new_n13302__;
  assign new_new_n13304__ = new_new_n13270__ & ~new_new_n13303__;
  assign new_new_n13305__ = ~new_new_n13270__ & new_new_n13303__;
  assign new_new_n13306__ = ~new_new_n13304__ & ~new_new_n13305__;
  assign new_new_n13307__ = new_new_n13237__ & ~new_new_n13306__;
  assign new_new_n13308__ = ~new_new_n13237__ & new_new_n13306__;
  assign new_new_n13309__ = ~new_new_n13307__ & ~new_new_n13308__;
  assign new_new_n13310__ = ~new_new_n12943__ & ~new_new_n12973__;
  assign new_new_n13311__ = ~new_new_n12944__ & ~new_new_n13310__;
  assign new_new_n13312__ = ~new_new_n13309__ & new_new_n13311__;
  assign new_new_n13313__ = new_new_n13309__ & ~new_new_n13311__;
  assign new_new_n13314__ = ~new_new_n13312__ & ~new_new_n13313__;
  assign new_new_n13315__ = new_new_n13132__ & ~new_new_n13151__;
  assign new_new_n13316__ = ~new_new_n13152__ & ~new_new_n13315__;
  assign new_new_n13317__ = ~new_new_n13098__ & ~new_new_n13102__;
  assign new_new_n13318__ = ~new_new_n13101__ & ~new_new_n13317__;
  assign new_new_n13319__ = ~new_new_n13136__ & ~new_new_n13138__;
  assign new_new_n13320__ = ~new_new_n13135__ & ~new_new_n13319__;
  assign new_new_n13321__ = ~new_new_n13318__ & new_new_n13320__;
  assign new_new_n13322__ = new_new_n13318__ & ~new_new_n13320__;
  assign new_new_n13323__ = ~new_new_n13321__ & ~new_new_n13322__;
  assign new_new_n13324__ = new_new_n13316__ & ~new_new_n13323__;
  assign new_new_n13325__ = ~new_new_n13316__ & new_new_n13323__;
  assign new_new_n13326__ = ~new_new_n13324__ & ~new_new_n13325__;
  assign new_new_n13327__ = ~new_new_n13119__ & ~new_new_n13123__;
  assign new_new_n13328__ = ~new_new_n13122__ & ~new_new_n13327__;
  assign new_new_n13329__ = ~new_new_n13107__ & ~new_new_n13111__;
  assign new_new_n13330__ = ~new_new_n13110__ & ~new_new_n13329__;
  assign new_new_n13331__ = new_new_n13328__ & new_new_n13330__;
  assign new_new_n13332__ = ~new_new_n13328__ & ~new_new_n13330__;
  assign new_new_n13333__ = ~new_new_n13331__ & ~new_new_n13332__;
  assign new_new_n13334__ = ~new_new_n13086__ & ~new_new_n13090__;
  assign new_new_n13335__ = ~new_new_n13089__ & ~new_new_n13334__;
  assign new_new_n13336__ = ~new_new_n13074__ & ~new_new_n13078__;
  assign new_new_n13337__ = ~new_new_n13077__ & ~new_new_n13336__;
  assign new_new_n13338__ = new_new_n13335__ & ~new_new_n13337__;
  assign new_new_n13339__ = ~new_new_n13335__ & new_new_n13337__;
  assign new_new_n13340__ = ~new_new_n13338__ & ~new_new_n13339__;
  assign new_new_n13341__ = new_new_n13333__ & ~new_new_n13340__;
  assign new_new_n13342__ = ~new_new_n13333__ & new_new_n13340__;
  assign new_new_n13343__ = ~new_new_n13341__ & ~new_new_n13342__;
  assign new_new_n13344__ = new_new_n13326__ & new_new_n13343__;
  assign new_new_n13345__ = ~new_new_n13326__ & ~new_new_n13343__;
  assign new_new_n13346__ = ~new_new_n13344__ & ~new_new_n13345__;
  assign new_new_n13347__ = ~new_new_n13097__ & ~new_new_n13158__;
  assign new_new_n13348__ = ~new_new_n13157__ & ~new_new_n13347__;
  assign new_new_n13349__ = ~new_new_n13346__ & new_new_n13348__;
  assign new_new_n13350__ = new_new_n13346__ & ~new_new_n13348__;
  assign new_new_n13351__ = ~new_new_n13349__ & ~new_new_n13350__;
  assign new_new_n13352__ = ~new_new_n13032__ & ~new_new_n13038__;
  assign new_new_n13353__ = ~new_new_n13037__ & ~new_new_n13352__;
  assign new_new_n13354__ = new_new_n13055__ & new_new_n13353__;
  assign new_new_n13355__ = ~new_new_n13055__ & ~new_new_n13353__;
  assign new_new_n13356__ = ~new_new_n13354__ & ~new_new_n13355__;
  assign new_new_n13357__ = ~new_new_n12982__ & ~new_new_n12995__;
  assign new_new_n13358__ = ~new_new_n12994__ & ~new_new_n13357__;
  assign new_new_n13359__ = new_new_n13356__ & ~new_new_n13358__;
  assign new_new_n13360__ = ~new_new_n13356__ & new_new_n13358__;
  assign new_new_n13361__ = ~new_new_n13359__ & ~new_new_n13360__;
  assign new_new_n13362__ = ~new_new_n13351__ & new_new_n13361__;
  assign new_new_n13363__ = new_new_n13351__ & ~new_new_n13361__;
  assign new_new_n13364__ = ~new_new_n13362__ & ~new_new_n13363__;
  assign new_new_n13365__ = new_new_n13314__ & new_new_n13364__;
  assign new_new_n13366__ = ~new_new_n13314__ & ~new_new_n13364__;
  assign new_new_n13367__ = ~new_new_n13365__ & ~new_new_n13366__;
  assign new_new_n13368__ = new_new_n12929__ & ~new_new_n13188__;
  assign new_new_n13369__ = ~new_new_n13181__ & ~new_new_n13189__;
  assign new_new_n13370__ = ~new_new_n12719__ & new_new_n13183__;
  assign new_new_n13371__ = ~new_new_n13181__ & ~new_new_n13370__;
  assign new_new_n13372__ = new_new_n12719__ & new_new_n13182__;
  assign new_new_n13373__ = ~new_new_n13371__ & ~new_new_n13372__;
  assign new_new_n13374__ = ~new_new_n12928__ & ~new_new_n13373__;
  assign new_new_n13375__ = ~new_new_n13368__ & ~new_new_n13374__;
  assign new_new_n13376__ = ~new_new_n13369__ & new_new_n13375__;
  assign new_new_n13377__ = new_new_n13367__ & new_new_n13376__;
  assign new_new_n13378__ = ~new_new_n13367__ & ~new_new_n13376__;
  assign new_new_n13379__ = ~new_new_n13377__ & ~new_new_n13378__;
  assign new_new_n13380__ = ~new_new_n13175__ & ~new_new_n13178__;
  assign new_new_n13381__ = ~new_new_n13174__ & ~new_new_n13380__;
  assign new_new_n13382__ = ~new_new_n13027__ & ~new_new_n13170__;
  assign new_new_n13383__ = ~new_new_n13026__ & ~new_new_n13382__;
  assign new_new_n13384__ = ~new_new_n13381__ & new_new_n13383__;
  assign new_new_n13385__ = new_new_n13381__ & ~new_new_n13383__;
  assign new_new_n13386__ = ~new_new_n13384__ & ~new_new_n13385__;
  assign new_new_n13387__ = ~new_new_n13043__ & ~new_new_n13059__;
  assign new_new_n13388__ = ~new_new_n13044__ & ~new_new_n13387__;
  assign new_new_n13389__ = ~new_new_n13000__ & ~new_new_n13004__;
  assign new_new_n13390__ = ~new_new_n13388__ & ~new_new_n13389__;
  assign new_new_n13391__ = new_new_n13388__ & new_new_n13389__;
  assign new_new_n13392__ = ~new_new_n13390__ & ~new_new_n13391__;
  assign new_new_n13393__ = pi34 & pi41;
  assign new_new_n13394__ = pi20 & pi55;
  assign new_new_n13395__ = pi25 & pi50;
  assign new_new_n13396__ = ~new_new_n13394__ & ~new_new_n13395__;
  assign new_new_n13397__ = new_new_n13394__ & new_new_n13395__;
  assign new_new_n13398__ = ~new_new_n13396__ & ~new_new_n13397__;
  assign new_new_n13399__ = new_new_n13393__ & ~new_new_n13398__;
  assign new_new_n13400__ = ~new_new_n13393__ & new_new_n13398__;
  assign new_new_n13401__ = ~new_new_n13399__ & ~new_new_n13400__;
  assign new_new_n13402__ = pi24 & pi51;
  assign new_new_n13403__ = pi22 & pi53;
  assign new_new_n13404__ = pi21 & pi54;
  assign new_new_n13405__ = ~new_new_n13403__ & ~new_new_n13404__;
  assign new_new_n13406__ = new_new_n13403__ & new_new_n13404__;
  assign new_new_n13407__ = ~new_new_n13405__ & ~new_new_n13406__;
  assign new_new_n13408__ = new_new_n13402__ & ~new_new_n13407__;
  assign new_new_n13409__ = ~new_new_n13402__ & new_new_n13407__;
  assign new_new_n13410__ = ~new_new_n13408__ & ~new_new_n13409__;
  assign new_new_n13411__ = new_new_n13401__ & new_new_n13410__;
  assign new_new_n13412__ = ~new_new_n13401__ & ~new_new_n13410__;
  assign new_new_n13413__ = ~new_new_n13411__ & ~new_new_n13412__;
  assign new_new_n13414__ = pi33 & pi42;
  assign new_new_n13415__ = pi32 & pi43;
  assign new_new_n13416__ = pi31 & pi44;
  assign new_new_n13417__ = ~new_new_n13415__ & ~new_new_n13416__;
  assign new_new_n13418__ = new_new_n13415__ & new_new_n13416__;
  assign new_new_n13419__ = ~new_new_n13417__ & ~new_new_n13418__;
  assign new_new_n13420__ = new_new_n13414__ & ~new_new_n13419__;
  assign new_new_n13421__ = ~new_new_n13414__ & new_new_n13419__;
  assign new_new_n13422__ = ~new_new_n13420__ & ~new_new_n13421__;
  assign new_new_n13423__ = new_new_n13413__ & ~new_new_n13422__;
  assign new_new_n13424__ = ~new_new_n13413__ & new_new_n13422__;
  assign new_new_n13425__ = ~new_new_n13423__ & ~new_new_n13424__;
  assign new_new_n13426__ = new_new_n13392__ & ~new_new_n13425__;
  assign new_new_n13427__ = ~new_new_n13392__ & new_new_n13425__;
  assign new_new_n13428__ = ~new_new_n13426__ & ~new_new_n13427__;
  assign new_new_n13429__ = new_new_n13166__ & new_new_n13428__;
  assign new_new_n13430__ = ~new_new_n13166__ & ~new_new_n13428__;
  assign new_new_n13431__ = ~new_new_n13429__ & ~new_new_n13430__;
  assign new_new_n13432__ = ~new_new_n13019__ & ~new_new_n13022__;
  assign new_new_n13433__ = ~new_new_n13018__ & ~new_new_n13432__;
  assign new_new_n13434__ = new_new_n13431__ & ~new_new_n13433__;
  assign new_new_n13435__ = ~new_new_n13431__ & new_new_n13433__;
  assign new_new_n13436__ = ~new_new_n13434__ & ~new_new_n13435__;
  assign new_new_n13437__ = new_new_n13386__ & ~new_new_n13436__;
  assign new_new_n13438__ = ~new_new_n13386__ & new_new_n13436__;
  assign new_new_n13439__ = ~new_new_n13437__ & ~new_new_n13438__;
  assign new_new_n13440__ = new_new_n13379__ & new_new_n13439__;
  assign new_new_n13441__ = ~new_new_n13379__ & ~new_new_n13439__;
  assign po076 = ~new_new_n13440__ & ~new_new_n13441__;
  assign new_new_n13443__ = new_new_n13384__ & ~new_new_n13436__;
  assign new_new_n13444__ = new_new_n13385__ & new_new_n13436__;
  assign new_new_n13445__ = ~new_new_n13443__ & ~new_new_n13444__;
  assign new_new_n13446__ = new_new_n13379__ & new_new_n13445__;
  assign new_new_n13447__ = ~new_new_n13385__ & ~new_new_n13436__;
  assign new_new_n13448__ = ~new_new_n13384__ & ~new_new_n13447__;
  assign new_new_n13449__ = new_new_n13378__ & ~new_new_n13448__;
  assign new_new_n13450__ = new_new_n13377__ & new_new_n13448__;
  assign new_new_n13451__ = ~new_new_n13449__ & ~new_new_n13450__;
  assign new_new_n13452__ = ~new_new_n13446__ & new_new_n13451__;
  assign new_new_n13453__ = ~new_new_n13312__ & new_new_n13364__;
  assign new_new_n13454__ = ~new_new_n13313__ & ~new_new_n13453__;
  assign new_new_n13455__ = ~new_new_n13235__ & ~new_new_n13306__;
  assign new_new_n13456__ = ~new_new_n13236__ & ~new_new_n13455__;
  assign new_new_n13457__ = ~new_new_n13214__ & ~new_new_n13229__;
  assign new_new_n13458__ = ~new_new_n13230__ & ~new_new_n13457__;
  assign new_new_n13459__ = new_new_n13320__ & new_new_n13340__;
  assign new_new_n13460__ = ~new_new_n13320__ & ~new_new_n13340__;
  assign new_new_n13461__ = ~new_new_n13459__ & ~new_new_n13460__;
  assign new_new_n13462__ = new_new_n13316__ & new_new_n13461__;
  assign new_new_n13463__ = ~new_new_n13316__ & ~new_new_n13461__;
  assign new_new_n13464__ = ~new_new_n13318__ & new_new_n13333__;
  assign new_new_n13465__ = new_new_n13318__ & ~new_new_n13333__;
  assign new_new_n13466__ = ~new_new_n13464__ & ~new_new_n13465__;
  assign new_new_n13467__ = ~new_new_n13463__ & new_new_n13466__;
  assign new_new_n13468__ = ~new_new_n13462__ & ~new_new_n13467__;
  assign new_new_n13469__ = new_new_n13458__ & ~new_new_n13468__;
  assign new_new_n13470__ = ~new_new_n13458__ & new_new_n13468__;
  assign new_new_n13471__ = ~new_new_n13469__ & ~new_new_n13470__;
  assign new_new_n13472__ = pi32 & pi44;
  assign new_new_n13473__ = pi31 & pi45;
  assign new_new_n13474__ = pi13 & pi63;
  assign new_new_n13475__ = ~new_new_n13473__ & ~new_new_n13474__;
  assign new_new_n13476__ = new_new_n13473__ & new_new_n13474__;
  assign new_new_n13477__ = ~new_new_n13475__ & ~new_new_n13476__;
  assign new_new_n13478__ = new_new_n13472__ & ~new_new_n13477__;
  assign new_new_n13479__ = ~new_new_n13472__ & new_new_n13477__;
  assign new_new_n13480__ = ~new_new_n13478__ & ~new_new_n13479__;
  assign new_new_n13481__ = pi33 & pi43;
  assign new_new_n13482__ = pi23 & pi53;
  assign new_new_n13483__ = pi19 & pi57;
  assign new_new_n13484__ = ~new_new_n13482__ & ~new_new_n13483__;
  assign new_new_n13485__ = new_new_n13482__ & new_new_n13483__;
  assign new_new_n13486__ = ~new_new_n13484__ & ~new_new_n13485__;
  assign new_new_n13487__ = new_new_n13481__ & ~new_new_n13486__;
  assign new_new_n13488__ = ~new_new_n13481__ & new_new_n13486__;
  assign new_new_n13489__ = ~new_new_n13487__ & ~new_new_n13488__;
  assign new_new_n13490__ = pi22 & pi54;
  assign new_new_n13491__ = pi21 & pi55;
  assign new_new_n13492__ = pi20 & pi56;
  assign new_new_n13493__ = ~new_new_n13491__ & ~new_new_n13492__;
  assign new_new_n13494__ = new_new_n13491__ & new_new_n13492__;
  assign new_new_n13495__ = ~new_new_n13493__ & ~new_new_n13494__;
  assign new_new_n13496__ = new_new_n13490__ & ~new_new_n13495__;
  assign new_new_n13497__ = ~new_new_n13490__ & new_new_n13495__;
  assign new_new_n13498__ = ~new_new_n13496__ & ~new_new_n13497__;
  assign new_new_n13499__ = new_new_n13489__ & new_new_n13498__;
  assign new_new_n13500__ = ~new_new_n13489__ & ~new_new_n13498__;
  assign new_new_n13501__ = ~new_new_n13499__ & ~new_new_n13500__;
  assign new_new_n13502__ = new_new_n13480__ & ~new_new_n13501__;
  assign new_new_n13503__ = ~new_new_n13480__ & new_new_n13501__;
  assign new_new_n13504__ = ~new_new_n13502__ & ~new_new_n13503__;
  assign new_new_n13505__ = new_new_n13471__ & new_new_n13504__;
  assign new_new_n13506__ = ~new_new_n13471__ & ~new_new_n13504__;
  assign new_new_n13507__ = ~new_new_n13505__ & ~new_new_n13506__;
  assign new_new_n13508__ = ~new_new_n13456__ & new_new_n13507__;
  assign new_new_n13509__ = new_new_n13456__ & ~new_new_n13507__;
  assign new_new_n13510__ = ~new_new_n13508__ & ~new_new_n13509__;
  assign new_new_n13511__ = ~new_new_n13349__ & new_new_n13361__;
  assign new_new_n13512__ = ~new_new_n13350__ & ~new_new_n13511__;
  assign new_new_n13513__ = new_new_n13510__ & new_new_n13512__;
  assign new_new_n13514__ = ~new_new_n13510__ & ~new_new_n13512__;
  assign new_new_n13515__ = ~new_new_n13513__ & ~new_new_n13514__;
  assign new_new_n13516__ = ~new_new_n13454__ & new_new_n13515__;
  assign new_new_n13517__ = new_new_n13454__ & ~new_new_n13515__;
  assign new_new_n13518__ = ~new_new_n13516__ & ~new_new_n13517__;
  assign new_new_n13519__ = ~new_new_n13430__ & ~new_new_n13433__;
  assign new_new_n13520__ = ~new_new_n13429__ & ~new_new_n13519__;
  assign new_new_n13521__ = ~new_new_n13318__ & ~new_new_n13331__;
  assign new_new_n13522__ = ~new_new_n13332__ & ~new_new_n13521__;
  assign new_new_n13523__ = ~new_new_n13218__ & ~new_new_n13223__;
  assign new_new_n13524__ = ~new_new_n13224__ & ~new_new_n13523__;
  assign new_new_n13525__ = ~new_new_n13320__ & ~new_new_n13337__;
  assign new_new_n13526__ = new_new_n13320__ & new_new_n13337__;
  assign new_new_n13527__ = ~new_new_n13335__ & ~new_new_n13526__;
  assign new_new_n13528__ = ~new_new_n13525__ & ~new_new_n13527__;
  assign new_new_n13529__ = ~new_new_n13524__ & ~new_new_n13528__;
  assign new_new_n13530__ = new_new_n13524__ & new_new_n13528__;
  assign new_new_n13531__ = ~new_new_n13529__ & ~new_new_n13530__;
  assign new_new_n13532__ = new_new_n13522__ & ~new_new_n13531__;
  assign new_new_n13533__ = ~new_new_n13522__ & new_new_n13531__;
  assign new_new_n13534__ = ~new_new_n13532__ & ~new_new_n13533__;
  assign new_new_n13535__ = ~new_new_n13411__ & ~new_new_n13422__;
  assign new_new_n13536__ = ~new_new_n13412__ & ~new_new_n13535__;
  assign new_new_n13537__ = ~new_new_n13280__ & ~new_new_n13284__;
  assign new_new_n13538__ = ~new_new_n13283__ & ~new_new_n13537__;
  assign new_new_n13539__ = ~new_new_n13253__ & ~new_new_n13257__;
  assign new_new_n13540__ = ~new_new_n13256__ & ~new_new_n13539__;
  assign new_new_n13541__ = ~new_new_n13538__ & ~new_new_n13540__;
  assign new_new_n13542__ = new_new_n13538__ & new_new_n13540__;
  assign new_new_n13543__ = ~new_new_n13541__ & ~new_new_n13542__;
  assign new_new_n13544__ = new_new_n13536__ & ~new_new_n13543__;
  assign new_new_n13545__ = ~new_new_n13536__ & new_new_n13543__;
  assign new_new_n13546__ = ~new_new_n13544__ & ~new_new_n13545__;
  assign new_new_n13547__ = ~new_new_n13393__ & ~new_new_n13397__;
  assign new_new_n13548__ = ~new_new_n13396__ & ~new_new_n13547__;
  assign new_new_n13549__ = ~new_new_n13244__ & ~new_new_n13248__;
  assign new_new_n13550__ = ~new_new_n13247__ & ~new_new_n13549__;
  assign new_new_n13551__ = ~pi14 & ~new_new_n13550__;
  assign new_new_n13552__ = ~pi62 & ~new_new_n13550__;
  assign new_new_n13553__ = ~new_new_n13551__ & ~new_new_n13552__;
  assign new_new_n13554__ = pi37 & ~new_new_n13553__;
  assign new_new_n13555__ = pi14 & new_new_n13550__;
  assign new_new_n13556__ = ~new_new_n13551__ & ~new_new_n13555__;
  assign new_new_n13557__ = pi13 & ~new_new_n13556__;
  assign new_new_n13558__ = pi37 & new_new_n13555__;
  assign new_new_n13559__ = ~new_new_n13557__ & ~new_new_n13558__;
  assign new_new_n13560__ = pi62 & ~new_new_n13559__;
  assign new_new_n13561__ = ~new_new_n13554__ & ~new_new_n13560__;
  assign new_new_n13562__ = pi38 & ~new_new_n13561__;
  assign new_new_n13563__ = ~new_new_n6746__ & ~new_new_n13555__;
  assign new_new_n13564__ = pi62 & ~new_new_n13563__;
  assign new_new_n13565__ = pi37 & pi38;
  assign new_new_n13566__ = new_new_n13553__ & ~new_new_n13565__;
  assign new_new_n13567__ = ~new_new_n13564__ & new_new_n13566__;
  assign new_new_n13568__ = ~new_new_n13562__ & ~new_new_n13567__;
  assign new_new_n13569__ = new_new_n13548__ & ~new_new_n13568__;
  assign new_new_n13570__ = ~new_new_n13548__ & new_new_n13568__;
  assign new_new_n13571__ = ~new_new_n13569__ & ~new_new_n13570__;
  assign new_new_n13572__ = new_new_n13546__ & new_new_n13571__;
  assign new_new_n13573__ = ~new_new_n13546__ & ~new_new_n13571__;
  assign new_new_n13574__ = ~new_new_n13572__ & ~new_new_n13573__;
  assign new_new_n13575__ = ~new_new_n13534__ & new_new_n13574__;
  assign new_new_n13576__ = new_new_n13534__ & ~new_new_n13574__;
  assign new_new_n13577__ = ~new_new_n13575__ & ~new_new_n13576__;
  assign new_new_n13578__ = ~new_new_n13269__ & new_new_n13303__;
  assign new_new_n13579__ = ~new_new_n13268__ & ~new_new_n13578__;
  assign new_new_n13580__ = new_new_n13577__ & new_new_n13579__;
  assign new_new_n13581__ = ~new_new_n13577__ & ~new_new_n13579__;
  assign new_new_n13582__ = ~new_new_n13580__ & ~new_new_n13581__;
  assign new_new_n13583__ = new_new_n13520__ & ~new_new_n13582__;
  assign new_new_n13584__ = ~new_new_n13520__ & new_new_n13582__;
  assign new_new_n13585__ = ~new_new_n13583__ & ~new_new_n13584__;
  assign new_new_n13586__ = ~new_new_n13271__ & ~new_new_n13275__;
  assign new_new_n13587__ = ~new_new_n13274__ & ~new_new_n13586__;
  assign new_new_n13588__ = ~new_new_n13414__ & ~new_new_n13418__;
  assign new_new_n13589__ = ~new_new_n13417__ & ~new_new_n13588__;
  assign new_new_n13590__ = ~new_new_n13587__ & ~new_new_n13589__;
  assign new_new_n13591__ = new_new_n13587__ & new_new_n13589__;
  assign new_new_n13592__ = ~new_new_n13590__ & ~new_new_n13591__;
  assign new_new_n13593__ = ~new_new_n13292__ & ~new_new_n13296__;
  assign new_new_n13594__ = ~new_new_n13295__ & ~new_new_n13593__;
  assign new_new_n13595__ = ~new_new_n13592__ & new_new_n13594__;
  assign new_new_n13596__ = ~new_new_n13591__ & ~new_new_n13594__;
  assign new_new_n13597__ = ~new_new_n13590__ & new_new_n13596__;
  assign new_new_n13598__ = ~new_new_n13595__ & ~new_new_n13597__;
  assign new_new_n13599__ = ~new_new_n13243__ & ~new_new_n13262__;
  assign new_new_n13600__ = ~new_new_n13263__ & ~new_new_n13599__;
  assign new_new_n13601__ = ~new_new_n13289__ & ~new_new_n13300__;
  assign new_new_n13602__ = ~new_new_n13290__ & ~new_new_n13601__;
  assign new_new_n13603__ = new_new_n13600__ & new_new_n13602__;
  assign new_new_n13604__ = ~new_new_n13600__ & ~new_new_n13602__;
  assign new_new_n13605__ = ~new_new_n13603__ & ~new_new_n13604__;
  assign new_new_n13606__ = ~new_new_n13598__ & new_new_n13605__;
  assign new_new_n13607__ = new_new_n13598__ & ~new_new_n13605__;
  assign new_new_n13608__ = ~new_new_n13606__ & ~new_new_n13607__;
  assign new_new_n13609__ = ~new_new_n13390__ & ~new_new_n13425__;
  assign new_new_n13610__ = ~new_new_n13391__ & ~new_new_n13609__;
  assign new_new_n13611__ = ~new_new_n13608__ & ~new_new_n13610__;
  assign new_new_n13612__ = new_new_n13608__ & new_new_n13610__;
  assign new_new_n13613__ = ~new_new_n13611__ & ~new_new_n13612__;
  assign new_new_n13614__ = ~new_new_n13354__ & ~new_new_n13358__;
  assign new_new_n13615__ = ~new_new_n13355__ & ~new_new_n13614__;
  assign new_new_n13616__ = pi37 & pi39;
  assign new_new_n13617__ = pi25 & pi51;
  assign new_new_n13618__ = pi24 & pi52;
  assign new_new_n13619__ = ~new_new_n13617__ & ~new_new_n13618__;
  assign new_new_n13620__ = new_new_n13617__ & new_new_n13618__;
  assign new_new_n13621__ = ~new_new_n13619__ & ~new_new_n13620__;
  assign new_new_n13622__ = new_new_n13616__ & ~new_new_n13621__;
  assign new_new_n13623__ = ~new_new_n13616__ & new_new_n13621__;
  assign new_new_n13624__ = ~new_new_n13622__ & ~new_new_n13623__;
  assign new_new_n13625__ = pi30 & pi46;
  assign new_new_n13626__ = pi28 & pi48;
  assign new_new_n13627__ = pi29 & pi47;
  assign new_new_n13628__ = ~new_new_n13626__ & ~new_new_n13627__;
  assign new_new_n13629__ = new_new_n13626__ & new_new_n13627__;
  assign new_new_n13630__ = ~new_new_n13628__ & ~new_new_n13629__;
  assign new_new_n13631__ = new_new_n13625__ & ~new_new_n13630__;
  assign new_new_n13632__ = ~new_new_n13625__ & new_new_n13630__;
  assign new_new_n13633__ = ~new_new_n13631__ & ~new_new_n13632__;
  assign new_new_n13634__ = new_new_n13624__ & new_new_n13633__;
  assign new_new_n13635__ = ~new_new_n13624__ & ~new_new_n13633__;
  assign new_new_n13636__ = ~new_new_n13634__ & ~new_new_n13635__;
  assign new_new_n13637__ = pi36 & pi40;
  assign new_new_n13638__ = pi35 & pi41;
  assign new_new_n13639__ = pi34 & pi42;
  assign new_new_n13640__ = ~new_new_n13638__ & ~new_new_n13639__;
  assign new_new_n13641__ = new_new_n13638__ & new_new_n13639__;
  assign new_new_n13642__ = ~new_new_n13640__ & ~new_new_n13641__;
  assign new_new_n13643__ = new_new_n13637__ & ~new_new_n13642__;
  assign new_new_n13644__ = ~new_new_n13637__ & new_new_n13642__;
  assign new_new_n13645__ = ~new_new_n13643__ & ~new_new_n13644__;
  assign new_new_n13646__ = ~new_new_n13636__ & new_new_n13645__;
  assign new_new_n13647__ = new_new_n13636__ & ~new_new_n13645__;
  assign new_new_n13648__ = ~new_new_n13646__ & ~new_new_n13647__;
  assign new_new_n13649__ = new_new_n13615__ & new_new_n13648__;
  assign new_new_n13650__ = ~new_new_n13615__ & ~new_new_n13648__;
  assign new_new_n13651__ = ~new_new_n13649__ & ~new_new_n13650__;
  assign new_new_n13652__ = pi27 & pi49;
  assign new_new_n13653__ = pi18 & pi58;
  assign new_new_n13654__ = ~new_new_n6799__ & ~new_new_n13653__;
  assign new_new_n13655__ = new_new_n6799__ & new_new_n13653__;
  assign new_new_n13656__ = ~new_new_n13654__ & ~new_new_n13655__;
  assign new_new_n13657__ = new_new_n13652__ & ~new_new_n13656__;
  assign new_new_n13658__ = ~new_new_n13652__ & new_new_n13656__;
  assign new_new_n13659__ = ~new_new_n13657__ & ~new_new_n13658__;
  assign new_new_n13660__ = pi17 & pi59;
  assign new_new_n13661__ = pi15 & pi61;
  assign new_new_n13662__ = pi16 & pi60;
  assign new_new_n13663__ = ~new_new_n13661__ & ~new_new_n13662__;
  assign new_new_n13664__ = new_new_n13661__ & new_new_n13662__;
  assign new_new_n13665__ = ~new_new_n13663__ & ~new_new_n13664__;
  assign new_new_n13666__ = new_new_n13660__ & ~new_new_n13665__;
  assign new_new_n13667__ = ~new_new_n13660__ & new_new_n13665__;
  assign new_new_n13668__ = ~new_new_n13666__ & ~new_new_n13667__;
  assign new_new_n13669__ = new_new_n13659__ & new_new_n13668__;
  assign new_new_n13670__ = ~new_new_n13659__ & ~new_new_n13668__;
  assign new_new_n13671__ = ~new_new_n13669__ & ~new_new_n13670__;
  assign new_new_n13672__ = ~new_new_n13402__ & ~new_new_n13406__;
  assign new_new_n13673__ = ~new_new_n13405__ & ~new_new_n13672__;
  assign new_new_n13674__ = new_new_n13671__ & ~new_new_n13673__;
  assign new_new_n13675__ = ~new_new_n13671__ & new_new_n13673__;
  assign new_new_n13676__ = ~new_new_n13674__ & ~new_new_n13675__;
  assign new_new_n13677__ = new_new_n13651__ & new_new_n13676__;
  assign new_new_n13678__ = ~new_new_n13651__ & ~new_new_n13676__;
  assign new_new_n13679__ = ~new_new_n13677__ & ~new_new_n13678__;
  assign new_new_n13680__ = new_new_n13613__ & ~new_new_n13679__;
  assign new_new_n13681__ = ~new_new_n13613__ & new_new_n13679__;
  assign new_new_n13682__ = ~new_new_n13680__ & ~new_new_n13681__;
  assign new_new_n13683__ = new_new_n13585__ & ~new_new_n13682__;
  assign new_new_n13684__ = ~new_new_n13585__ & new_new_n13682__;
  assign new_new_n13685__ = ~new_new_n13683__ & ~new_new_n13684__;
  assign new_new_n13686__ = new_new_n13518__ & new_new_n13685__;
  assign new_new_n13687__ = ~new_new_n13518__ & ~new_new_n13685__;
  assign new_new_n13688__ = ~new_new_n13686__ & ~new_new_n13687__;
  assign new_new_n13689__ = ~new_new_n13452__ & new_new_n13688__;
  assign new_new_n13690__ = ~new_new_n13367__ & new_new_n13436__;
  assign new_new_n13691__ = ~new_new_n13376__ & new_new_n13690__;
  assign new_new_n13692__ = new_new_n13381__ & new_new_n13691__;
  assign new_new_n13693__ = new_new_n13367__ & ~new_new_n13436__;
  assign new_new_n13694__ = ~new_new_n13376__ & ~new_new_n13693__;
  assign new_new_n13695__ = ~new_new_n13690__ & ~new_new_n13694__;
  assign new_new_n13696__ = ~new_new_n13381__ & new_new_n13695__;
  assign new_new_n13697__ = new_new_n13376__ & new_new_n13693__;
  assign new_new_n13698__ = ~new_new_n13696__ & ~new_new_n13697__;
  assign new_new_n13699__ = new_new_n13383__ & ~new_new_n13698__;
  assign new_new_n13700__ = ~new_new_n13381__ & ~new_new_n13691__;
  assign new_new_n13701__ = ~new_new_n13383__ & ~new_new_n13695__;
  assign new_new_n13702__ = ~new_new_n13700__ & new_new_n13701__;
  assign new_new_n13703__ = new_new_n13376__ & ~new_new_n13381__;
  assign new_new_n13704__ = new_new_n13693__ & new_new_n13703__;
  assign new_new_n13705__ = ~new_new_n13692__ & ~new_new_n13704__;
  assign new_new_n13706__ = ~new_new_n13702__ & new_new_n13705__;
  assign new_new_n13707__ = ~new_new_n13699__ & new_new_n13706__;
  assign new_new_n13708__ = ~new_new_n13688__ & ~new_new_n13707__;
  assign po077 = new_new_n13689__ | new_new_n13708__;
  assign new_new_n13710__ = ~new_new_n13376__ & new_new_n13381__;
  assign new_new_n13711__ = ~new_new_n13688__ & ~new_new_n13710__;
  assign new_new_n13712__ = ~new_new_n13383__ & ~new_new_n13711__;
  assign new_new_n13713__ = new_new_n13688__ & ~new_new_n13703__;
  assign new_new_n13714__ = ~new_new_n13690__ & ~new_new_n13713__;
  assign new_new_n13715__ = ~new_new_n13712__ & new_new_n13714__;
  assign new_new_n13716__ = new_new_n13688__ & ~new_new_n13693__;
  assign new_new_n13717__ = ~new_new_n13688__ & new_new_n13693__;
  assign new_new_n13718__ = ~new_new_n13376__ & ~new_new_n13384__;
  assign new_new_n13719__ = ~new_new_n13385__ & ~new_new_n13718__;
  assign new_new_n13720__ = ~new_new_n13717__ & ~new_new_n13719__;
  assign new_new_n13721__ = ~new_new_n13716__ & ~new_new_n13720__;
  assign new_new_n13722__ = ~new_new_n13715__ & ~new_new_n13721__;
  assign new_new_n13723__ = ~new_new_n13517__ & ~new_new_n13685__;
  assign new_new_n13724__ = ~new_new_n13516__ & ~new_new_n13723__;
  assign new_new_n13725__ = ~new_new_n13722__ & ~new_new_n13724__;
  assign new_new_n13726__ = new_new_n13722__ & new_new_n13724__;
  assign new_new_n13727__ = ~new_new_n13725__ & ~new_new_n13726__;
  assign new_new_n13728__ = ~new_new_n13583__ & ~new_new_n13682__;
  assign new_new_n13729__ = ~new_new_n13584__ & ~new_new_n13728__;
  assign new_new_n13730__ = ~new_new_n13611__ & ~new_new_n13679__;
  assign new_new_n13731__ = ~new_new_n13612__ & ~new_new_n13730__;
  assign new_new_n13732__ = ~new_new_n13576__ & ~new_new_n13579__;
  assign new_new_n13733__ = ~new_new_n13575__ & ~new_new_n13732__;
  assign new_new_n13734__ = ~new_new_n13731__ & ~new_new_n13733__;
  assign new_new_n13735__ = new_new_n13731__ & new_new_n13733__;
  assign new_new_n13736__ = ~new_new_n13734__ & ~new_new_n13735__;
  assign new_new_n13737__ = ~new_new_n13598__ & ~new_new_n13603__;
  assign new_new_n13738__ = ~new_new_n13604__ & ~new_new_n13737__;
  assign new_new_n13739__ = new_new_n13536__ & new_new_n13568__;
  assign new_new_n13740__ = ~new_new_n13536__ & ~new_new_n13568__;
  assign new_new_n13741__ = ~new_new_n13543__ & new_new_n13548__;
  assign new_new_n13742__ = new_new_n13543__ & ~new_new_n13548__;
  assign new_new_n13743__ = ~new_new_n13741__ & ~new_new_n13742__;
  assign new_new_n13744__ = ~new_new_n13740__ & new_new_n13743__;
  assign new_new_n13745__ = ~new_new_n13739__ & ~new_new_n13744__;
  assign new_new_n13746__ = new_new_n13738__ & ~new_new_n13745__;
  assign new_new_n13747__ = ~new_new_n13738__ & new_new_n13745__;
  assign new_new_n13748__ = ~new_new_n13746__ & ~new_new_n13747__;
  assign new_new_n13749__ = pi34 & pi43;
  assign new_new_n13750__ = pi22 & pi55;
  assign new_new_n13751__ = ~new_new_n6942__ & ~new_new_n13750__;
  assign new_new_n13752__ = new_new_n6942__ & new_new_n13750__;
  assign new_new_n13753__ = ~new_new_n13751__ & ~new_new_n13752__;
  assign new_new_n13754__ = new_new_n13749__ & ~new_new_n13753__;
  assign new_new_n13755__ = ~new_new_n13749__ & new_new_n13753__;
  assign new_new_n13756__ = ~new_new_n13754__ & ~new_new_n13755__;
  assign new_new_n13757__ = pi25 & pi52;
  assign new_new_n13758__ = pi24 & pi53;
  assign new_new_n13759__ = pi23 & pi54;
  assign new_new_n13760__ = ~new_new_n13758__ & ~new_new_n13759__;
  assign new_new_n13761__ = new_new_n13758__ & new_new_n13759__;
  assign new_new_n13762__ = ~new_new_n13760__ & ~new_new_n13761__;
  assign new_new_n13763__ = new_new_n13757__ & ~new_new_n13762__;
  assign new_new_n13764__ = ~new_new_n13757__ & new_new_n13762__;
  assign new_new_n13765__ = ~new_new_n13763__ & ~new_new_n13764__;
  assign new_new_n13766__ = new_new_n13756__ & new_new_n13765__;
  assign new_new_n13767__ = ~new_new_n13756__ & ~new_new_n13765__;
  assign new_new_n13768__ = ~new_new_n13766__ & ~new_new_n13767__;
  assign new_new_n13769__ = pi33 & pi44;
  assign new_new_n13770__ = pi16 & pi61;
  assign new_new_n13771__ = pi32 & pi45;
  assign new_new_n13772__ = ~new_new_n13770__ & ~new_new_n13771__;
  assign new_new_n13773__ = new_new_n13770__ & new_new_n13771__;
  assign new_new_n13774__ = ~new_new_n13772__ & ~new_new_n13773__;
  assign new_new_n13775__ = new_new_n13769__ & ~new_new_n13774__;
  assign new_new_n13776__ = ~new_new_n13769__ & new_new_n13774__;
  assign new_new_n13777__ = ~new_new_n13775__ & ~new_new_n13776__;
  assign new_new_n13778__ = new_new_n13768__ & ~new_new_n13777__;
  assign new_new_n13779__ = ~new_new_n13768__ & new_new_n13777__;
  assign new_new_n13780__ = ~new_new_n13778__ & ~new_new_n13779__;
  assign new_new_n13781__ = new_new_n13748__ & ~new_new_n13780__;
  assign new_new_n13782__ = ~new_new_n13748__ & new_new_n13780__;
  assign new_new_n13783__ = ~new_new_n13781__ & ~new_new_n13782__;
  assign new_new_n13784__ = new_new_n13736__ & ~new_new_n13783__;
  assign new_new_n13785__ = ~new_new_n13736__ & new_new_n13783__;
  assign new_new_n13786__ = ~new_new_n13784__ & ~new_new_n13785__;
  assign new_new_n13787__ = new_new_n13729__ & new_new_n13786__;
  assign new_new_n13788__ = ~new_new_n13729__ & ~new_new_n13786__;
  assign new_new_n13789__ = ~new_new_n13787__ & ~new_new_n13788__;
  assign new_new_n13790__ = ~new_new_n13508__ & ~new_new_n13512__;
  assign new_new_n13791__ = ~new_new_n13509__ & ~new_new_n13790__;
  assign new_new_n13792__ = ~new_new_n13590__ & ~new_new_n13596__;
  assign new_new_n13793__ = ~new_new_n13542__ & ~new_new_n13548__;
  assign new_new_n13794__ = ~new_new_n13541__ & ~new_new_n13793__;
  assign new_new_n13795__ = ~new_new_n13616__ & ~new_new_n13620__;
  assign new_new_n13796__ = ~new_new_n13619__ & ~new_new_n13795__;
  assign new_new_n13797__ = pi18 & pi59;
  assign new_new_n13798__ = pi17 & pi60;
  assign new_new_n13799__ = ~new_new_n13797__ & ~new_new_n13798__;
  assign new_new_n13800__ = new_new_n13797__ & new_new_n13798__;
  assign new_new_n13801__ = ~new_new_n13799__ & ~new_new_n13800__;
  assign new_new_n13802__ = new_new_n13796__ & ~new_new_n13801__;
  assign new_new_n13803__ = ~new_new_n13796__ & new_new_n13801__;
  assign new_new_n13804__ = ~new_new_n13802__ & ~new_new_n13803__;
  assign new_new_n13805__ = new_new_n13794__ & ~new_new_n13804__;
  assign new_new_n13806__ = ~new_new_n13794__ & new_new_n13804__;
  assign new_new_n13807__ = ~new_new_n13805__ & ~new_new_n13806__;
  assign new_new_n13808__ = new_new_n13792__ & ~new_new_n13807__;
  assign new_new_n13809__ = ~new_new_n13792__ & new_new_n13807__;
  assign new_new_n13810__ = ~new_new_n13808__ & ~new_new_n13809__;
  assign new_new_n13811__ = ~new_new_n13480__ & ~new_new_n13499__;
  assign new_new_n13812__ = ~new_new_n13500__ & ~new_new_n13811__;
  assign new_new_n13813__ = ~new_new_n13481__ & ~new_new_n13485__;
  assign new_new_n13814__ = ~new_new_n13484__ & ~new_new_n13813__;
  assign new_new_n13815__ = new_new_n13812__ & ~new_new_n13814__;
  assign new_new_n13816__ = ~new_new_n13812__ & new_new_n13814__;
  assign new_new_n13817__ = ~new_new_n13815__ & ~new_new_n13816__;
  assign new_new_n13818__ = ~new_new_n13625__ & ~new_new_n13629__;
  assign new_new_n13819__ = ~new_new_n13628__ & ~new_new_n13818__;
  assign new_new_n13820__ = ~new_new_n13472__ & ~new_new_n13476__;
  assign new_new_n13821__ = ~new_new_n13475__ & ~new_new_n13820__;
  assign new_new_n13822__ = ~new_new_n13819__ & ~new_new_n13821__;
  assign new_new_n13823__ = new_new_n13819__ & new_new_n13821__;
  assign new_new_n13824__ = ~new_new_n13822__ & ~new_new_n13823__;
  assign new_new_n13825__ = ~new_new_n13490__ & ~new_new_n13494__;
  assign new_new_n13826__ = ~new_new_n13493__ & ~new_new_n13825__;
  assign new_new_n13827__ = ~new_new_n13660__ & ~new_new_n13664__;
  assign new_new_n13828__ = ~new_new_n13663__ & ~new_new_n13827__;
  assign new_new_n13829__ = ~new_new_n13652__ & ~new_new_n13655__;
  assign new_new_n13830__ = ~new_new_n13654__ & ~new_new_n13829__;
  assign new_new_n13831__ = new_new_n13828__ & ~new_new_n13830__;
  assign new_new_n13832__ = ~new_new_n13828__ & new_new_n13830__;
  assign new_new_n13833__ = ~new_new_n13831__ & ~new_new_n13832__;
  assign new_new_n13834__ = new_new_n13826__ & new_new_n13833__;
  assign new_new_n13835__ = ~new_new_n13826__ & ~new_new_n13833__;
  assign new_new_n13836__ = ~new_new_n13834__ & ~new_new_n13835__;
  assign new_new_n13837__ = new_new_n13824__ & ~new_new_n13836__;
  assign new_new_n13838__ = ~new_new_n13824__ & new_new_n13836__;
  assign new_new_n13839__ = ~new_new_n13837__ & ~new_new_n13838__;
  assign new_new_n13840__ = new_new_n13817__ & new_new_n13839__;
  assign new_new_n13841__ = ~new_new_n13817__ & ~new_new_n13839__;
  assign new_new_n13842__ = ~new_new_n13840__ & ~new_new_n13841__;
  assign new_new_n13843__ = new_new_n13810__ & ~new_new_n13842__;
  assign new_new_n13844__ = ~new_new_n13810__ & new_new_n13842__;
  assign new_new_n13845__ = ~new_new_n13843__ & ~new_new_n13844__;
  assign new_new_n13846__ = ~new_new_n13650__ & ~new_new_n13676__;
  assign new_new_n13847__ = ~new_new_n13649__ & ~new_new_n13846__;
  assign new_new_n13848__ = new_new_n13845__ & ~new_new_n13847__;
  assign new_new_n13849__ = ~new_new_n13845__ & new_new_n13847__;
  assign new_new_n13850__ = ~new_new_n13848__ & ~new_new_n13849__;
  assign new_new_n13851__ = ~new_new_n13791__ & ~new_new_n13850__;
  assign new_new_n13852__ = new_new_n13791__ & new_new_n13850__;
  assign new_new_n13853__ = ~new_new_n13851__ & ~new_new_n13852__;
  assign new_new_n13854__ = ~new_new_n13634__ & ~new_new_n13645__;
  assign new_new_n13855__ = ~new_new_n13635__ & ~new_new_n13854__;
  assign new_new_n13856__ = pi13 & ~new_new_n13551__;
  assign new_new_n13857__ = ~new_new_n6759__ & ~new_new_n13856__;
  assign new_new_n13858__ = pi38 & ~new_new_n13857__;
  assign new_new_n13859__ = ~new_new_n13555__ & ~new_new_n13858__;
  assign new_new_n13860__ = pi62 & ~new_new_n13859__;
  assign new_new_n13861__ = new_new_n13550__ & new_new_n13565__;
  assign new_new_n13862__ = ~new_new_n13860__ & ~new_new_n13861__;
  assign new_new_n13863__ = ~new_new_n13669__ & new_new_n13673__;
  assign new_new_n13864__ = ~new_new_n13670__ & ~new_new_n13863__;
  assign new_new_n13865__ = ~new_new_n13862__ & ~new_new_n13864__;
  assign new_new_n13866__ = new_new_n13862__ & new_new_n13864__;
  assign new_new_n13867__ = ~new_new_n13865__ & ~new_new_n13866__;
  assign new_new_n13868__ = ~new_new_n13855__ & new_new_n13867__;
  assign new_new_n13869__ = new_new_n13855__ & ~new_new_n13867__;
  assign new_new_n13870__ = ~new_new_n13868__ & ~new_new_n13869__;
  assign new_new_n13871__ = ~new_new_n13522__ & ~new_new_n13530__;
  assign new_new_n13872__ = ~new_new_n13529__ & ~new_new_n13871__;
  assign new_new_n13873__ = pi31 & pi46;
  assign new_new_n13874__ = pi30 & pi47;
  assign new_new_n13875__ = pi14 & pi63;
  assign new_new_n13876__ = ~new_new_n13874__ & ~new_new_n13875__;
  assign new_new_n13877__ = new_new_n13874__ & new_new_n13875__;
  assign new_new_n13878__ = ~new_new_n13876__ & ~new_new_n13877__;
  assign new_new_n13879__ = new_new_n13873__ & ~new_new_n13878__;
  assign new_new_n13880__ = ~new_new_n13873__ & new_new_n13878__;
  assign new_new_n13881__ = ~new_new_n13879__ & ~new_new_n13880__;
  assign new_new_n13882__ = pi37 & pi40;
  assign new_new_n13883__ = pi35 & pi42;
  assign new_new_n13884__ = pi36 & pi41;
  assign new_new_n13885__ = ~new_new_n13883__ & ~new_new_n13884__;
  assign new_new_n13886__ = new_new_n13883__ & new_new_n13884__;
  assign new_new_n13887__ = ~new_new_n13885__ & ~new_new_n13886__;
  assign new_new_n13888__ = new_new_n13882__ & ~new_new_n13887__;
  assign new_new_n13889__ = ~new_new_n13882__ & new_new_n13887__;
  assign new_new_n13890__ = ~new_new_n13888__ & ~new_new_n13889__;
  assign new_new_n13891__ = new_new_n13881__ & new_new_n13890__;
  assign new_new_n13892__ = ~new_new_n13881__ & ~new_new_n13890__;
  assign new_new_n13893__ = ~new_new_n13891__ & ~new_new_n13892__;
  assign new_new_n13894__ = pi15 & pi62;
  assign new_new_n13895__ = ~pi38 & pi39;
  assign new_new_n13896__ = new_new_n13894__ & ~new_new_n13895__;
  assign new_new_n13897__ = ~new_new_n13894__ & new_new_n13895__;
  assign new_new_n13898__ = ~new_new_n13896__ & ~new_new_n13897__;
  assign new_new_n13899__ = new_new_n13893__ & ~new_new_n13898__;
  assign new_new_n13900__ = ~new_new_n13893__ & new_new_n13898__;
  assign new_new_n13901__ = ~new_new_n13899__ & ~new_new_n13900__;
  assign new_new_n13902__ = ~new_new_n13872__ & ~new_new_n13901__;
  assign new_new_n13903__ = new_new_n13872__ & new_new_n13901__;
  assign new_new_n13904__ = ~new_new_n13902__ & ~new_new_n13903__;
  assign new_new_n13905__ = ~new_new_n13637__ & ~new_new_n13641__;
  assign new_new_n13906__ = ~new_new_n13640__ & ~new_new_n13905__;
  assign new_new_n13907__ = pi21 & pi56;
  assign new_new_n13908__ = pi20 & pi57;
  assign new_new_n13909__ = pi19 & pi58;
  assign new_new_n13910__ = ~new_new_n13908__ & ~new_new_n13909__;
  assign new_new_n13911__ = new_new_n13908__ & new_new_n13909__;
  assign new_new_n13912__ = ~new_new_n13910__ & ~new_new_n13911__;
  assign new_new_n13913__ = new_new_n13907__ & ~new_new_n13912__;
  assign new_new_n13914__ = ~new_new_n13907__ & new_new_n13912__;
  assign new_new_n13915__ = ~new_new_n13913__ & ~new_new_n13914__;
  assign new_new_n13916__ = ~new_new_n13906__ & new_new_n13915__;
  assign new_new_n13917__ = new_new_n13906__ & ~new_new_n13915__;
  assign new_new_n13918__ = ~new_new_n13916__ & ~new_new_n13917__;
  assign new_new_n13919__ = pi29 & pi48;
  assign new_new_n13920__ = pi28 & pi49;
  assign new_new_n13921__ = pi27 & pi50;
  assign new_new_n13922__ = ~new_new_n13920__ & ~new_new_n13921__;
  assign new_new_n13923__ = new_new_n13920__ & new_new_n13921__;
  assign new_new_n13924__ = ~new_new_n13922__ & ~new_new_n13923__;
  assign new_new_n13925__ = new_new_n13919__ & ~new_new_n13924__;
  assign new_new_n13926__ = ~new_new_n13919__ & new_new_n13924__;
  assign new_new_n13927__ = ~new_new_n13925__ & ~new_new_n13926__;
  assign new_new_n13928__ = new_new_n13918__ & new_new_n13927__;
  assign new_new_n13929__ = ~new_new_n13918__ & ~new_new_n13927__;
  assign new_new_n13930__ = ~new_new_n13928__ & ~new_new_n13929__;
  assign new_new_n13931__ = new_new_n13904__ & ~new_new_n13930__;
  assign new_new_n13932__ = ~new_new_n13904__ & new_new_n13930__;
  assign new_new_n13933__ = ~new_new_n13931__ & ~new_new_n13932__;
  assign new_new_n13934__ = ~new_new_n13470__ & ~new_new_n13504__;
  assign new_new_n13935__ = ~new_new_n13469__ & ~new_new_n13934__;
  assign new_new_n13936__ = ~new_new_n13933__ & ~new_new_n13935__;
  assign new_new_n13937__ = new_new_n13933__ & new_new_n13935__;
  assign new_new_n13938__ = ~new_new_n13936__ & ~new_new_n13937__;
  assign new_new_n13939__ = new_new_n13870__ & new_new_n13938__;
  assign new_new_n13940__ = ~new_new_n13870__ & ~new_new_n13938__;
  assign new_new_n13941__ = ~new_new_n13939__ & ~new_new_n13940__;
  assign new_new_n13942__ = new_new_n13853__ & new_new_n13941__;
  assign new_new_n13943__ = ~new_new_n13853__ & ~new_new_n13941__;
  assign new_new_n13944__ = ~new_new_n13942__ & ~new_new_n13943__;
  assign new_new_n13945__ = new_new_n13789__ & ~new_new_n13944__;
  assign new_new_n13946__ = ~new_new_n13789__ & new_new_n13944__;
  assign new_new_n13947__ = ~new_new_n13945__ & ~new_new_n13946__;
  assign new_new_n13948__ = new_new_n13727__ & new_new_n13947__;
  assign new_new_n13949__ = ~new_new_n13727__ & ~new_new_n13947__;
  assign po078 = new_new_n13948__ | new_new_n13949__;
  assign new_new_n13951__ = ~new_new_n13843__ & ~new_new_n13847__;
  assign new_new_n13952__ = ~new_new_n13844__ & ~new_new_n13951__;
  assign new_new_n13953__ = ~new_new_n13865__ & ~new_new_n13868__;
  assign new_new_n13954__ = pi21 & pi57;
  assign new_new_n13955__ = pi18 & pi60;
  assign new_new_n13956__ = pi19 & pi59;
  assign new_new_n13957__ = ~new_new_n13955__ & ~new_new_n13956__;
  assign new_new_n13958__ = new_new_n13955__ & new_new_n13956__;
  assign new_new_n13959__ = ~new_new_n13957__ & ~new_new_n13958__;
  assign new_new_n13960__ = new_new_n13954__ & ~new_new_n13959__;
  assign new_new_n13961__ = ~new_new_n13954__ & new_new_n13959__;
  assign new_new_n13962__ = ~new_new_n13960__ & ~new_new_n13961__;
  assign new_new_n13963__ = pi29 & pi49;
  assign new_new_n13964__ = pi28 & pi50;
  assign new_new_n13965__ = pi27 & pi51;
  assign new_new_n13966__ = ~new_new_n13964__ & ~new_new_n13965__;
  assign new_new_n13967__ = new_new_n13964__ & new_new_n13965__;
  assign new_new_n13968__ = ~new_new_n13966__ & ~new_new_n13967__;
  assign new_new_n13969__ = new_new_n13963__ & ~new_new_n13968__;
  assign new_new_n13970__ = ~new_new_n13963__ & new_new_n13968__;
  assign new_new_n13971__ = ~new_new_n13969__ & ~new_new_n13970__;
  assign new_new_n13972__ = new_new_n13962__ & new_new_n13971__;
  assign new_new_n13973__ = ~new_new_n13962__ & ~new_new_n13971__;
  assign new_new_n13974__ = ~new_new_n13972__ & ~new_new_n13973__;
  assign new_new_n13975__ = pi17 & pi61;
  assign new_new_n13976__ = pi16 & pi62;
  assign new_new_n13977__ = pi15 & pi63;
  assign new_new_n13978__ = ~new_new_n13976__ & ~new_new_n13977__;
  assign new_new_n13979__ = new_new_n13976__ & new_new_n13977__;
  assign new_new_n13980__ = ~new_new_n13978__ & ~new_new_n13979__;
  assign new_new_n13981__ = new_new_n13975__ & ~new_new_n13980__;
  assign new_new_n13982__ = ~new_new_n13975__ & new_new_n13980__;
  assign new_new_n13983__ = ~new_new_n13981__ & ~new_new_n13982__;
  assign new_new_n13984__ = ~new_new_n13974__ & new_new_n13983__;
  assign new_new_n13985__ = new_new_n13974__ & ~new_new_n13983__;
  assign new_new_n13986__ = ~new_new_n13984__ & ~new_new_n13985__;
  assign new_new_n13987__ = ~new_new_n13953__ & new_new_n13986__;
  assign new_new_n13988__ = new_new_n13953__ & ~new_new_n13986__;
  assign new_new_n13989__ = ~new_new_n13987__ & ~new_new_n13988__;
  assign new_new_n13990__ = pi34 & pi44;
  assign new_new_n13991__ = pi33 & pi45;
  assign new_new_n13992__ = pi32 & pi46;
  assign new_new_n13993__ = ~new_new_n13991__ & ~new_new_n13992__;
  assign new_new_n13994__ = new_new_n13991__ & new_new_n13992__;
  assign new_new_n13995__ = ~new_new_n13993__ & ~new_new_n13994__;
  assign new_new_n13996__ = new_new_n13990__ & ~new_new_n13995__;
  assign new_new_n13997__ = ~new_new_n13990__ & new_new_n13995__;
  assign new_new_n13998__ = ~new_new_n13996__ & ~new_new_n13997__;
  assign new_new_n13999__ = pi25 & pi53;
  assign new_new_n14000__ = pi24 & pi54;
  assign new_new_n14001__ = pi22 & pi56;
  assign new_new_n14002__ = ~new_new_n14000__ & ~new_new_n14001__;
  assign new_new_n14003__ = new_new_n14000__ & new_new_n14001__;
  assign new_new_n14004__ = ~new_new_n14002__ & ~new_new_n14003__;
  assign new_new_n14005__ = new_new_n13999__ & ~new_new_n14004__;
  assign new_new_n14006__ = ~new_new_n13999__ & new_new_n14004__;
  assign new_new_n14007__ = ~new_new_n14005__ & ~new_new_n14006__;
  assign new_new_n14008__ = new_new_n13998__ & new_new_n14007__;
  assign new_new_n14009__ = ~new_new_n13998__ & ~new_new_n14007__;
  assign new_new_n14010__ = pi31 & pi47;
  assign new_new_n14011__ = pi20 & pi58;
  assign new_new_n14012__ = pi30 & pi48;
  assign new_new_n14013__ = ~new_new_n14011__ & ~new_new_n14012__;
  assign new_new_n14014__ = new_new_n14011__ & new_new_n14012__;
  assign new_new_n14015__ = ~new_new_n14013__ & ~new_new_n14014__;
  assign new_new_n14016__ = new_new_n14010__ & ~new_new_n14015__;
  assign new_new_n14017__ = ~new_new_n14010__ & new_new_n14015__;
  assign new_new_n14018__ = ~new_new_n14016__ & ~new_new_n14017__;
  assign new_new_n14019__ = ~new_new_n14008__ & ~new_new_n14018__;
  assign new_new_n14020__ = ~new_new_n14009__ & ~new_new_n14019__;
  assign new_new_n14021__ = ~new_new_n14008__ & new_new_n14020__;
  assign new_new_n14022__ = ~new_new_n14009__ & new_new_n14019__;
  assign new_new_n14023__ = ~new_new_n14018__ & ~new_new_n14022__;
  assign new_new_n14024__ = ~new_new_n14021__ & ~new_new_n14023__;
  assign new_new_n14025__ = new_new_n13989__ & ~new_new_n14024__;
  assign new_new_n14026__ = ~new_new_n13989__ & new_new_n14024__;
  assign new_new_n14027__ = ~new_new_n14025__ & ~new_new_n14026__;
  assign new_new_n14028__ = ~new_new_n13952__ & new_new_n14027__;
  assign new_new_n14029__ = new_new_n13952__ & ~new_new_n14027__;
  assign new_new_n14030__ = ~new_new_n14028__ & ~new_new_n14029__;
  assign new_new_n14031__ = ~new_new_n13870__ & ~new_new_n13937__;
  assign new_new_n14032__ = ~new_new_n13936__ & ~new_new_n14031__;
  assign new_new_n14033__ = new_new_n14030__ & new_new_n14032__;
  assign new_new_n14034__ = ~new_new_n14030__ & ~new_new_n14032__;
  assign new_new_n14035__ = ~new_new_n14033__ & ~new_new_n14034__;
  assign new_new_n14036__ = ~new_new_n13852__ & ~new_new_n13941__;
  assign new_new_n14037__ = ~new_new_n13851__ & ~new_new_n14036__;
  assign new_new_n14038__ = ~new_new_n14035__ & ~new_new_n14037__;
  assign new_new_n14039__ = new_new_n14035__ & new_new_n14037__;
  assign new_new_n14040__ = ~new_new_n14038__ & ~new_new_n14039__;
  assign new_new_n14041__ = ~new_new_n13891__ & ~new_new_n13898__;
  assign new_new_n14042__ = ~new_new_n13892__ & ~new_new_n14041__;
  assign new_new_n14043__ = ~new_new_n13766__ & ~new_new_n13777__;
  assign new_new_n14044__ = ~new_new_n13767__ & ~new_new_n14043__;
  assign new_new_n14045__ = new_new_n14042__ & new_new_n14044__;
  assign new_new_n14046__ = ~new_new_n14042__ & ~new_new_n14044__;
  assign new_new_n14047__ = ~new_new_n14045__ & ~new_new_n14046__;
  assign new_new_n14048__ = ~new_new_n13916__ & ~new_new_n13927__;
  assign new_new_n14049__ = ~new_new_n13917__ & ~new_new_n14048__;
  assign new_new_n14050__ = new_new_n14047__ & ~new_new_n14049__;
  assign new_new_n14051__ = ~new_new_n14047__ & new_new_n14049__;
  assign new_new_n14052__ = ~new_new_n14050__ & ~new_new_n14051__;
  assign new_new_n14053__ = ~new_new_n13769__ & ~new_new_n13773__;
  assign new_new_n14054__ = ~new_new_n13772__ & ~new_new_n14053__;
  assign new_new_n14055__ = ~new_new_n13873__ & ~new_new_n13877__;
  assign new_new_n14056__ = ~new_new_n13876__ & ~new_new_n14055__;
  assign new_new_n14057__ = ~new_new_n14054__ & ~new_new_n14056__;
  assign new_new_n14058__ = new_new_n14054__ & new_new_n14056__;
  assign new_new_n14059__ = ~new_new_n14057__ & ~new_new_n14058__;
  assign new_new_n14060__ = ~new_new_n13919__ & ~new_new_n13923__;
  assign new_new_n14061__ = ~new_new_n13922__ & ~new_new_n14060__;
  assign new_new_n14062__ = ~new_new_n14059__ & new_new_n14061__;
  assign new_new_n14063__ = new_new_n14059__ & ~new_new_n14061__;
  assign new_new_n14064__ = ~new_new_n14062__ & ~new_new_n14063__;
  assign new_new_n14065__ = ~pi38 & ~new_new_n13894__;
  assign new_new_n14066__ = pi39 & ~new_new_n14065__;
  assign new_new_n14067__ = ~new_new_n13757__ & ~new_new_n13761__;
  assign new_new_n14068__ = ~new_new_n13760__ & ~new_new_n14067__;
  assign new_new_n14069__ = ~new_new_n13882__ & ~new_new_n13886__;
  assign new_new_n14070__ = ~new_new_n13885__ & ~new_new_n14069__;
  assign new_new_n14071__ = new_new_n14068__ & new_new_n14070__;
  assign new_new_n14072__ = ~new_new_n14068__ & ~new_new_n14070__;
  assign new_new_n14073__ = ~new_new_n14071__ & ~new_new_n14072__;
  assign new_new_n14074__ = new_new_n14066__ & ~new_new_n14073__;
  assign new_new_n14075__ = ~new_new_n14066__ & new_new_n14073__;
  assign new_new_n14076__ = ~new_new_n14074__ & ~new_new_n14075__;
  assign new_new_n14077__ = ~new_new_n13814__ & ~new_new_n13830__;
  assign new_new_n14078__ = new_new_n13814__ & new_new_n13830__;
  assign new_new_n14079__ = ~new_new_n13828__ & ~new_new_n14078__;
  assign new_new_n14080__ = ~new_new_n14077__ & ~new_new_n14079__;
  assign new_new_n14081__ = new_new_n14076__ & ~new_new_n14080__;
  assign new_new_n14082__ = ~new_new_n14076__ & new_new_n14080__;
  assign new_new_n14083__ = ~new_new_n14081__ & ~new_new_n14082__;
  assign new_new_n14084__ = new_new_n14064__ & new_new_n14083__;
  assign new_new_n14085__ = ~new_new_n14064__ & ~new_new_n14083__;
  assign new_new_n14086__ = ~new_new_n14084__ & ~new_new_n14085__;
  assign new_new_n14087__ = new_new_n14052__ & ~new_new_n14086__;
  assign new_new_n14088__ = ~new_new_n14052__ & new_new_n14086__;
  assign new_new_n14089__ = ~new_new_n14087__ & ~new_new_n14088__;
  assign new_new_n14090__ = new_new_n13824__ & ~new_new_n13826__;
  assign new_new_n14091__ = ~new_new_n13824__ & new_new_n13826__;
  assign new_new_n14092__ = ~new_new_n14090__ & ~new_new_n14091__;
  assign new_new_n14093__ = new_new_n13812__ & new_new_n14092__;
  assign new_new_n14094__ = ~new_new_n13812__ & ~new_new_n14092__;
  assign new_new_n14095__ = new_new_n13814__ & new_new_n13833__;
  assign new_new_n14096__ = ~new_new_n13814__ & ~new_new_n13833__;
  assign new_new_n14097__ = ~new_new_n14095__ & ~new_new_n14096__;
  assign new_new_n14098__ = ~new_new_n14094__ & new_new_n14097__;
  assign new_new_n14099__ = ~new_new_n14093__ & ~new_new_n14098__;
  assign new_new_n14100__ = new_new_n14089__ & ~new_new_n14099__;
  assign new_new_n14101__ = ~new_new_n14089__ & new_new_n14099__;
  assign new_new_n14102__ = ~new_new_n14100__ & ~new_new_n14101__;
  assign new_new_n14103__ = ~new_new_n13735__ & ~new_new_n13783__;
  assign new_new_n14104__ = ~new_new_n13734__ & ~new_new_n14103__;
  assign new_new_n14105__ = ~new_new_n13903__ & new_new_n13930__;
  assign new_new_n14106__ = ~new_new_n13902__ & ~new_new_n14105__;
  assign new_new_n14107__ = new_new_n13792__ & ~new_new_n13806__;
  assign new_new_n14108__ = ~new_new_n13805__ & ~new_new_n14107__;
  assign new_new_n14109__ = ~new_new_n13823__ & ~new_new_n13826__;
  assign new_new_n14110__ = ~new_new_n13822__ & ~new_new_n14109__;
  assign new_new_n14111__ = pi36 & pi42;
  assign new_new_n14112__ = pi35 & pi43;
  assign new_new_n14113__ = pi23 & pi55;
  assign new_new_n14114__ = ~new_new_n14112__ & ~new_new_n14113__;
  assign new_new_n14115__ = new_new_n14112__ & new_new_n14113__;
  assign new_new_n14116__ = ~new_new_n14114__ & ~new_new_n14115__;
  assign new_new_n14117__ = new_new_n14111__ & ~new_new_n14116__;
  assign new_new_n14118__ = ~new_new_n14111__ & new_new_n14116__;
  assign new_new_n14119__ = ~new_new_n14117__ & ~new_new_n14118__;
  assign new_new_n14120__ = pi38 & pi40;
  assign new_new_n14121__ = pi37 & pi41;
  assign new_new_n14122__ = pi26 & pi52;
  assign new_new_n14123__ = ~new_new_n14121__ & ~new_new_n14122__;
  assign new_new_n14124__ = new_new_n14121__ & new_new_n14122__;
  assign new_new_n14125__ = ~new_new_n14123__ & ~new_new_n14124__;
  assign new_new_n14126__ = new_new_n14120__ & ~new_new_n14125__;
  assign new_new_n14127__ = ~new_new_n14120__ & new_new_n14125__;
  assign new_new_n14128__ = ~new_new_n14126__ & ~new_new_n14127__;
  assign new_new_n14129__ = ~new_new_n14119__ & ~new_new_n14128__;
  assign new_new_n14130__ = new_new_n14119__ & new_new_n14128__;
  assign new_new_n14131__ = ~new_new_n14129__ & ~new_new_n14130__;
  assign new_new_n14132__ = new_new_n14110__ & new_new_n14131__;
  assign new_new_n14133__ = ~new_new_n14110__ & ~new_new_n14131__;
  assign new_new_n14134__ = ~new_new_n14132__ & ~new_new_n14133__;
  assign new_new_n14135__ = new_new_n14108__ & ~new_new_n14134__;
  assign new_new_n14136__ = ~new_new_n14108__ & new_new_n14134__;
  assign new_new_n14137__ = ~new_new_n14135__ & ~new_new_n14136__;
  assign new_new_n14138__ = ~new_new_n13749__ & ~new_new_n13752__;
  assign new_new_n14139__ = ~new_new_n13751__ & ~new_new_n14138__;
  assign new_new_n14140__ = ~new_new_n13796__ & ~new_new_n13800__;
  assign new_new_n14141__ = ~new_new_n13799__ & ~new_new_n14140__;
  assign new_new_n14142__ = ~new_new_n14139__ & ~new_new_n14141__;
  assign new_new_n14143__ = new_new_n14139__ & new_new_n14141__;
  assign new_new_n14144__ = ~new_new_n14142__ & ~new_new_n14143__;
  assign new_new_n14145__ = ~new_new_n13907__ & ~new_new_n13911__;
  assign new_new_n14146__ = ~new_new_n13910__ & ~new_new_n14145__;
  assign new_new_n14147__ = new_new_n14144__ & ~new_new_n14146__;
  assign new_new_n14148__ = ~new_new_n14144__ & new_new_n14146__;
  assign new_new_n14149__ = ~new_new_n14147__ & ~new_new_n14148__;
  assign new_new_n14150__ = new_new_n14137__ & ~new_new_n14149__;
  assign new_new_n14151__ = ~new_new_n14137__ & new_new_n14149__;
  assign new_new_n14152__ = ~new_new_n14150__ & ~new_new_n14151__;
  assign new_new_n14153__ = new_new_n14106__ & new_new_n14152__;
  assign new_new_n14154__ = ~new_new_n14106__ & ~new_new_n14152__;
  assign new_new_n14155__ = ~new_new_n14153__ & ~new_new_n14154__;
  assign new_new_n14156__ = ~new_new_n13747__ & ~new_new_n13780__;
  assign new_new_n14157__ = ~new_new_n13746__ & ~new_new_n14156__;
  assign new_new_n14158__ = new_new_n14155__ & ~new_new_n14157__;
  assign new_new_n14159__ = ~new_new_n14155__ & new_new_n14157__;
  assign new_new_n14160__ = ~new_new_n14158__ & ~new_new_n14159__;
  assign new_new_n14161__ = ~new_new_n14104__ & ~new_new_n14160__;
  assign new_new_n14162__ = new_new_n14104__ & new_new_n14160__;
  assign new_new_n14163__ = ~new_new_n14161__ & ~new_new_n14162__;
  assign new_new_n14164__ = ~new_new_n14102__ & new_new_n14163__;
  assign new_new_n14165__ = new_new_n14102__ & ~new_new_n14163__;
  assign new_new_n14166__ = ~new_new_n14164__ & ~new_new_n14165__;
  assign new_new_n14167__ = new_new_n14040__ & new_new_n14166__;
  assign new_new_n14168__ = ~new_new_n14040__ & ~new_new_n14166__;
  assign new_new_n14169__ = ~new_new_n14167__ & ~new_new_n14168__;
  assign new_new_n14170__ = new_new_n13787__ & new_new_n13944__;
  assign new_new_n14171__ = new_new_n13788__ & ~new_new_n13944__;
  assign new_new_n14172__ = ~new_new_n14170__ & ~new_new_n14171__;
  assign new_new_n14173__ = new_new_n13727__ & new_new_n14172__;
  assign new_new_n14174__ = ~new_new_n13788__ & new_new_n13944__;
  assign new_new_n14175__ = ~new_new_n13787__ & ~new_new_n14174__;
  assign new_new_n14176__ = new_new_n13726__ & ~new_new_n14175__;
  assign new_new_n14177__ = new_new_n13725__ & new_new_n14175__;
  assign new_new_n14178__ = ~new_new_n14176__ & ~new_new_n14177__;
  assign new_new_n14179__ = ~new_new_n14173__ & new_new_n14178__;
  assign new_new_n14180__ = ~new_new_n14169__ & ~new_new_n14179__;
  assign new_new_n14181__ = new_new_n13725__ & new_new_n13787__;
  assign new_new_n14182__ = new_new_n13725__ & new_new_n13729__;
  assign new_new_n14183__ = ~new_new_n13725__ & ~new_new_n13729__;
  assign new_new_n14184__ = ~new_new_n13726__ & new_new_n13786__;
  assign new_new_n14185__ = ~new_new_n14183__ & new_new_n14184__;
  assign new_new_n14186__ = ~new_new_n14182__ & ~new_new_n14185__;
  assign new_new_n14187__ = new_new_n13944__ & ~new_new_n14186__;
  assign new_new_n14188__ = new_new_n13726__ & ~new_new_n13787__;
  assign new_new_n14189__ = ~new_new_n13786__ & new_new_n14183__;
  assign new_new_n14190__ = ~new_new_n14188__ & ~new_new_n14189__;
  assign new_new_n14191__ = ~new_new_n13944__ & ~new_new_n14190__;
  assign new_new_n14192__ = new_new_n13726__ & new_new_n13788__;
  assign new_new_n14193__ = ~new_new_n14181__ & ~new_new_n14192__;
  assign new_new_n14194__ = ~new_new_n14187__ & new_new_n14193__;
  assign new_new_n14195__ = ~new_new_n14191__ & new_new_n14194__;
  assign new_new_n14196__ = new_new_n14169__ & ~new_new_n14195__;
  assign po079 = new_new_n14180__ | new_new_n14196__;
  assign new_new_n14198__ = new_new_n13788__ & ~new_new_n14169__;
  assign new_new_n14199__ = ~new_new_n13788__ & new_new_n14169__;
  assign new_new_n14200__ = ~new_new_n13725__ & ~new_new_n13944__;
  assign new_new_n14201__ = ~new_new_n13726__ & ~new_new_n14200__;
  assign new_new_n14202__ = ~new_new_n14199__ & ~new_new_n14201__;
  assign new_new_n14203__ = ~new_new_n13726__ & new_new_n14169__;
  assign new_new_n14204__ = ~new_new_n13725__ & ~new_new_n14169__;
  assign new_new_n14205__ = new_new_n13944__ & ~new_new_n14204__;
  assign new_new_n14206__ = ~new_new_n13787__ & ~new_new_n14203__;
  assign new_new_n14207__ = ~new_new_n14205__ & new_new_n14206__;
  assign new_new_n14208__ = ~new_new_n14198__ & ~new_new_n14202__;
  assign new_new_n14209__ = ~new_new_n14207__ & new_new_n14208__;
  assign new_new_n14210__ = ~new_new_n14039__ & ~new_new_n14166__;
  assign new_new_n14211__ = ~new_new_n14038__ & ~new_new_n14210__;
  assign new_new_n14212__ = ~new_new_n14209__ & ~new_new_n14211__;
  assign new_new_n14213__ = new_new_n14209__ & new_new_n14211__;
  assign new_new_n14214__ = ~new_new_n14212__ & ~new_new_n14213__;
  assign new_new_n14215__ = ~new_new_n14064__ & ~new_new_n14081__;
  assign new_new_n14216__ = ~new_new_n14082__ & ~new_new_n14215__;
  assign new_new_n14217__ = pi33 & pi46;
  assign new_new_n14218__ = pi32 & pi47;
  assign new_new_n14219__ = pi31 & pi48;
  assign new_new_n14220__ = ~new_new_n14218__ & ~new_new_n14219__;
  assign new_new_n14221__ = new_new_n14218__ & new_new_n14219__;
  assign new_new_n14222__ = ~new_new_n14220__ & ~new_new_n14221__;
  assign new_new_n14223__ = new_new_n14217__ & ~new_new_n14222__;
  assign new_new_n14224__ = ~new_new_n14217__ & new_new_n14222__;
  assign new_new_n14225__ = ~new_new_n14223__ & ~new_new_n14224__;
  assign new_new_n14226__ = pi21 & pi58;
  assign new_new_n14227__ = pi19 & pi60;
  assign new_new_n14228__ = pi20 & pi59;
  assign new_new_n14229__ = ~new_new_n14227__ & ~new_new_n14228__;
  assign new_new_n14230__ = new_new_n14227__ & new_new_n14228__;
  assign new_new_n14231__ = ~new_new_n14229__ & ~new_new_n14230__;
  assign new_new_n14232__ = new_new_n14226__ & ~new_new_n14231__;
  assign new_new_n14233__ = ~new_new_n14226__ & new_new_n14231__;
  assign new_new_n14234__ = ~new_new_n14232__ & ~new_new_n14233__;
  assign new_new_n14235__ = new_new_n14225__ & new_new_n14234__;
  assign new_new_n14236__ = ~new_new_n14225__ & ~new_new_n14234__;
  assign new_new_n14237__ = ~new_new_n14235__ & ~new_new_n14236__;
  assign new_new_n14238__ = pi30 & pi49;
  assign new_new_n14239__ = pi29 & pi50;
  assign new_new_n14240__ = pi22 & pi57;
  assign new_new_n14241__ = ~new_new_n14239__ & ~new_new_n14240__;
  assign new_new_n14242__ = new_new_n14239__ & new_new_n14240__;
  assign new_new_n14243__ = ~new_new_n14241__ & ~new_new_n14242__;
  assign new_new_n14244__ = new_new_n14238__ & ~new_new_n14243__;
  assign new_new_n14245__ = ~new_new_n14238__ & new_new_n14243__;
  assign new_new_n14246__ = ~new_new_n14244__ & ~new_new_n14245__;
  assign new_new_n14247__ = ~new_new_n14237__ & new_new_n14246__;
  assign new_new_n14248__ = new_new_n14237__ & ~new_new_n14246__;
  assign new_new_n14249__ = ~new_new_n14247__ & ~new_new_n14248__;
  assign new_new_n14250__ = ~new_new_n14216__ & new_new_n14249__;
  assign new_new_n14251__ = new_new_n14216__ & ~new_new_n14249__;
  assign new_new_n14252__ = ~new_new_n14250__ & ~new_new_n14251__;
  assign new_new_n14253__ = pi39 & pi40;
  assign new_new_n14254__ = pi38 & pi41;
  assign new_new_n14255__ = pi37 & pi42;
  assign new_new_n14256__ = ~new_new_n14254__ & ~new_new_n14255__;
  assign new_new_n14257__ = new_new_n14254__ & new_new_n14255__;
  assign new_new_n14258__ = ~new_new_n14256__ & ~new_new_n14257__;
  assign new_new_n14259__ = new_new_n14253__ & ~new_new_n14258__;
  assign new_new_n14260__ = ~new_new_n14253__ & new_new_n14258__;
  assign new_new_n14261__ = ~new_new_n14259__ & ~new_new_n14260__;
  assign new_new_n14262__ = pi28 & pi51;
  assign new_new_n14263__ = pi17 & pi62;
  assign new_new_n14264__ = ~new_new_n14262__ & ~new_new_n14263__;
  assign new_new_n14265__ = new_new_n14262__ & new_new_n14263__;
  assign new_new_n14266__ = ~new_new_n14264__ & ~new_new_n14265__;
  assign new_new_n14267__ = pi40 & ~new_new_n14266__;
  assign new_new_n14268__ = ~pi40 & ~new_new_n14265__;
  assign new_new_n14269__ = ~new_new_n14264__ & new_new_n14268__;
  assign new_new_n14270__ = ~new_new_n14267__ & ~new_new_n14269__;
  assign new_new_n14271__ = pi25 & pi54;
  assign new_new_n14272__ = pi24 & pi55;
  assign new_new_n14273__ = ~new_new_n14271__ & ~new_new_n14272__;
  assign new_new_n14274__ = new_new_n14271__ & new_new_n14272__;
  assign new_new_n14275__ = ~new_new_n14273__ & ~new_new_n14274__;
  assign new_new_n14276__ = new_new_n7755__ & ~new_new_n14275__;
  assign new_new_n14277__ = ~new_new_n7755__ & new_new_n14275__;
  assign new_new_n14278__ = ~new_new_n14276__ & ~new_new_n14277__;
  assign new_new_n14279__ = new_new_n14270__ & new_new_n14278__;
  assign new_new_n14280__ = ~new_new_n14270__ & ~new_new_n14278__;
  assign new_new_n14281__ = ~new_new_n14279__ & ~new_new_n14280__;
  assign new_new_n14282__ = ~new_new_n14261__ & new_new_n14281__;
  assign new_new_n14283__ = new_new_n14261__ & ~new_new_n14281__;
  assign new_new_n14284__ = ~new_new_n14282__ & ~new_new_n14283__;
  assign new_new_n14285__ = new_new_n14252__ & ~new_new_n14284__;
  assign new_new_n14286__ = ~new_new_n14252__ & new_new_n14284__;
  assign new_new_n14287__ = ~new_new_n14285__ & ~new_new_n14286__;
  assign new_new_n14288__ = ~new_new_n14087__ & ~new_new_n14099__;
  assign new_new_n14289__ = ~new_new_n14088__ & ~new_new_n14288__;
  assign new_new_n14290__ = new_new_n14287__ & ~new_new_n14289__;
  assign new_new_n14291__ = ~new_new_n14287__ & new_new_n14289__;
  assign new_new_n14292__ = ~new_new_n14290__ & ~new_new_n14291__;
  assign new_new_n14293__ = ~new_new_n14135__ & ~new_new_n14149__;
  assign new_new_n14294__ = ~new_new_n14136__ & ~new_new_n14293__;
  assign new_new_n14295__ = ~new_new_n14058__ & ~new_new_n14061__;
  assign new_new_n14296__ = ~new_new_n14057__ & ~new_new_n14295__;
  assign new_new_n14297__ = ~new_new_n13972__ & ~new_new_n13983__;
  assign new_new_n14298__ = ~new_new_n13973__ & ~new_new_n14297__;
  assign new_new_n14299__ = ~new_new_n14066__ & ~new_new_n14071__;
  assign new_new_n14300__ = ~new_new_n14072__ & ~new_new_n14299__;
  assign new_new_n14301__ = ~new_new_n14298__ & new_new_n14300__;
  assign new_new_n14302__ = new_new_n14298__ & ~new_new_n14300__;
  assign new_new_n14303__ = ~new_new_n14301__ & ~new_new_n14302__;
  assign new_new_n14304__ = ~new_new_n14296__ & ~new_new_n14303__;
  assign new_new_n14305__ = new_new_n14296__ & new_new_n14303__;
  assign new_new_n14306__ = ~new_new_n14304__ & ~new_new_n14305__;
  assign new_new_n14307__ = new_new_n14294__ & ~new_new_n14306__;
  assign new_new_n14308__ = ~new_new_n14294__ & new_new_n14306__;
  assign new_new_n14309__ = ~new_new_n14307__ & ~new_new_n14308__;
  assign new_new_n14310__ = ~new_new_n14045__ & ~new_new_n14049__;
  assign new_new_n14311__ = ~new_new_n14046__ & ~new_new_n14310__;
  assign new_new_n14312__ = new_new_n14309__ & ~new_new_n14311__;
  assign new_new_n14313__ = ~new_new_n14309__ & new_new_n14311__;
  assign new_new_n14314__ = ~new_new_n14312__ & ~new_new_n14313__;
  assign new_new_n14315__ = new_new_n14292__ & ~new_new_n14314__;
  assign new_new_n14316__ = ~new_new_n14292__ & new_new_n14314__;
  assign new_new_n14317__ = ~new_new_n14315__ & ~new_new_n14316__;
  assign new_new_n14318__ = new_new_n14102__ & ~new_new_n14161__;
  assign new_new_n14319__ = ~new_new_n14162__ & ~new_new_n14318__;
  assign new_new_n14320__ = ~new_new_n14153__ & ~new_new_n14157__;
  assign new_new_n14321__ = ~new_new_n14154__ & ~new_new_n14320__;
  assign new_new_n14322__ = ~new_new_n14028__ & ~new_new_n14032__;
  assign new_new_n14323__ = ~new_new_n14029__ & ~new_new_n14322__;
  assign new_new_n14324__ = ~new_new_n14321__ & ~new_new_n14323__;
  assign new_new_n14325__ = new_new_n14321__ & new_new_n14323__;
  assign new_new_n14326__ = ~new_new_n14324__ & ~new_new_n14325__;
  assign new_new_n14327__ = ~new_new_n13987__ & new_new_n14024__;
  assign new_new_n14328__ = ~new_new_n13988__ & ~new_new_n14327__;
  assign new_new_n14329__ = ~new_new_n13954__ & ~new_new_n13958__;
  assign new_new_n14330__ = ~new_new_n13957__ & ~new_new_n14329__;
  assign new_new_n14331__ = ~new_new_n13963__ & ~new_new_n13967__;
  assign new_new_n14332__ = ~new_new_n13966__ & ~new_new_n14331__;
  assign new_new_n14333__ = ~new_new_n13999__ & ~new_new_n14003__;
  assign new_new_n14334__ = ~new_new_n14002__ & ~new_new_n14333__;
  assign new_new_n14335__ = ~new_new_n14332__ & ~new_new_n14334__;
  assign new_new_n14336__ = new_new_n14332__ & new_new_n14334__;
  assign new_new_n14337__ = ~new_new_n14335__ & ~new_new_n14336__;
  assign new_new_n14338__ = new_new_n14330__ & ~new_new_n14337__;
  assign new_new_n14339__ = ~new_new_n14330__ & new_new_n14337__;
  assign new_new_n14340__ = ~new_new_n14338__ & ~new_new_n14339__;
  assign new_new_n14341__ = ~new_new_n14143__ & ~new_new_n14146__;
  assign new_new_n14342__ = ~new_new_n14142__ & ~new_new_n14341__;
  assign new_new_n14343__ = pi36 & pi43;
  assign new_new_n14344__ = pi23 & pi56;
  assign new_new_n14345__ = pi27 & pi52;
  assign new_new_n14346__ = ~new_new_n14344__ & ~new_new_n14345__;
  assign new_new_n14347__ = new_new_n14344__ & new_new_n14345__;
  assign new_new_n14348__ = ~new_new_n14346__ & ~new_new_n14347__;
  assign new_new_n14349__ = new_new_n14343__ & ~new_new_n14348__;
  assign new_new_n14350__ = ~new_new_n14343__ & new_new_n14348__;
  assign new_new_n14351__ = ~new_new_n14349__ & ~new_new_n14350__;
  assign new_new_n14352__ = pi35 & pi44;
  assign new_new_n14353__ = pi16 & pi63;
  assign new_new_n14354__ = pi34 & pi45;
  assign new_new_n14355__ = ~new_new_n14353__ & ~new_new_n14354__;
  assign new_new_n14356__ = new_new_n14353__ & new_new_n14354__;
  assign new_new_n14357__ = ~new_new_n14355__ & ~new_new_n14356__;
  assign new_new_n14358__ = new_new_n14352__ & ~new_new_n14357__;
  assign new_new_n14359__ = ~new_new_n14352__ & new_new_n14357__;
  assign new_new_n14360__ = ~new_new_n14358__ & ~new_new_n14359__;
  assign new_new_n14361__ = new_new_n14351__ & new_new_n14360__;
  assign new_new_n14362__ = ~new_new_n14351__ & ~new_new_n14360__;
  assign new_new_n14363__ = ~new_new_n14361__ & ~new_new_n14362__;
  assign new_new_n14364__ = new_new_n14342__ & new_new_n14363__;
  assign new_new_n14365__ = ~new_new_n14342__ & ~new_new_n14363__;
  assign new_new_n14366__ = ~new_new_n14364__ & ~new_new_n14365__;
  assign new_new_n14367__ = ~new_new_n14340__ & new_new_n14366__;
  assign new_new_n14368__ = new_new_n14340__ & ~new_new_n14366__;
  assign new_new_n14369__ = ~new_new_n14367__ & ~new_new_n14368__;
  assign new_new_n14370__ = new_new_n14110__ & ~new_new_n14130__;
  assign new_new_n14371__ = ~new_new_n14129__ & ~new_new_n14370__;
  assign new_new_n14372__ = new_new_n14369__ & ~new_new_n14371__;
  assign new_new_n14373__ = ~new_new_n14369__ & new_new_n14371__;
  assign new_new_n14374__ = ~new_new_n14372__ & ~new_new_n14373__;
  assign new_new_n14375__ = ~new_new_n14328__ & ~new_new_n14374__;
  assign new_new_n14376__ = new_new_n14328__ & new_new_n14374__;
  assign new_new_n14377__ = ~new_new_n14375__ & ~new_new_n14376__;
  assign new_new_n14378__ = pi18 & pi61;
  assign new_new_n14379__ = ~new_new_n14111__ & ~new_new_n14115__;
  assign new_new_n14380__ = ~new_new_n14114__ & ~new_new_n14379__;
  assign new_new_n14381__ = ~new_new_n14120__ & ~new_new_n14124__;
  assign new_new_n14382__ = ~new_new_n14123__ & ~new_new_n14381__;
  assign new_new_n14383__ = new_new_n14380__ & new_new_n14382__;
  assign new_new_n14384__ = ~new_new_n14380__ & ~new_new_n14382__;
  assign new_new_n14385__ = ~new_new_n14383__ & ~new_new_n14384__;
  assign new_new_n14386__ = new_new_n14378__ & ~new_new_n14385__;
  assign new_new_n14387__ = ~new_new_n14378__ & new_new_n14385__;
  assign new_new_n14388__ = ~new_new_n14386__ & ~new_new_n14387__;
  assign new_new_n14389__ = ~new_new_n14020__ & ~new_new_n14388__;
  assign new_new_n14390__ = new_new_n14020__ & new_new_n14388__;
  assign new_new_n14391__ = ~new_new_n14389__ & ~new_new_n14390__;
  assign new_new_n14392__ = ~new_new_n13990__ & ~new_new_n13994__;
  assign new_new_n14393__ = ~new_new_n13993__ & ~new_new_n14392__;
  assign new_new_n14394__ = ~new_new_n13975__ & ~new_new_n13979__;
  assign new_new_n14395__ = ~new_new_n13978__ & ~new_new_n14394__;
  assign new_new_n14396__ = ~new_new_n14010__ & ~new_new_n14014__;
  assign new_new_n14397__ = ~new_new_n14013__ & ~new_new_n14396__;
  assign new_new_n14398__ = ~new_new_n14395__ & ~new_new_n14397__;
  assign new_new_n14399__ = new_new_n14395__ & new_new_n14397__;
  assign new_new_n14400__ = ~new_new_n14398__ & ~new_new_n14399__;
  assign new_new_n14401__ = new_new_n14393__ & ~new_new_n14400__;
  assign new_new_n14402__ = ~new_new_n14393__ & new_new_n14400__;
  assign new_new_n14403__ = ~new_new_n14401__ & ~new_new_n14402__;
  assign new_new_n14404__ = new_new_n14391__ & new_new_n14403__;
  assign new_new_n14405__ = ~new_new_n14391__ & ~new_new_n14403__;
  assign new_new_n14406__ = ~new_new_n14404__ & ~new_new_n14405__;
  assign new_new_n14407__ = new_new_n14377__ & ~new_new_n14406__;
  assign new_new_n14408__ = ~new_new_n14377__ & new_new_n14406__;
  assign new_new_n14409__ = ~new_new_n14407__ & ~new_new_n14408__;
  assign new_new_n14410__ = new_new_n14326__ & new_new_n14409__;
  assign new_new_n14411__ = ~new_new_n14326__ & ~new_new_n14409__;
  assign new_new_n14412__ = ~new_new_n14410__ & ~new_new_n14411__;
  assign new_new_n14413__ = new_new_n14319__ & new_new_n14412__;
  assign new_new_n14414__ = ~new_new_n14319__ & ~new_new_n14412__;
  assign new_new_n14415__ = ~new_new_n14413__ & ~new_new_n14414__;
  assign new_new_n14416__ = ~new_new_n14317__ & new_new_n14415__;
  assign new_new_n14417__ = new_new_n14317__ & ~new_new_n14415__;
  assign new_new_n14418__ = ~new_new_n14416__ & ~new_new_n14417__;
  assign new_new_n14419__ = new_new_n14214__ & new_new_n14418__;
  assign new_new_n14420__ = ~new_new_n14214__ & ~new_new_n14418__;
  assign po080 = ~new_new_n14419__ & ~new_new_n14420__;
  assign new_new_n14422__ = ~new_new_n14325__ & ~new_new_n14409__;
  assign new_new_n14423__ = ~new_new_n14324__ & ~new_new_n14422__;
  assign new_new_n14424__ = ~new_new_n14376__ & new_new_n14406__;
  assign new_new_n14425__ = ~new_new_n14375__ & ~new_new_n14424__;
  assign new_new_n14426__ = pi38 & pi42;
  assign new_new_n14427__ = pi25 & pi55;
  assign new_new_n14428__ = pi37 & pi43;
  assign new_new_n14429__ = ~new_new_n14427__ & ~new_new_n14428__;
  assign new_new_n14430__ = new_new_n14427__ & new_new_n14428__;
  assign new_new_n14431__ = ~new_new_n14429__ & ~new_new_n14430__;
  assign new_new_n14432__ = new_new_n14426__ & ~new_new_n14431__;
  assign new_new_n14433__ = ~new_new_n14426__ & new_new_n14431__;
  assign new_new_n14434__ = ~new_new_n14432__ & ~new_new_n14433__;
  assign new_new_n14435__ = pi26 & pi54;
  assign new_new_n14436__ = pi23 & pi57;
  assign new_new_n14437__ = pi24 & pi56;
  assign new_new_n14438__ = ~new_new_n14436__ & ~new_new_n14437__;
  assign new_new_n14439__ = new_new_n14436__ & new_new_n14437__;
  assign new_new_n14440__ = ~new_new_n14438__ & ~new_new_n14439__;
  assign new_new_n14441__ = new_new_n14435__ & ~new_new_n14440__;
  assign new_new_n14442__ = ~new_new_n14435__ & new_new_n14440__;
  assign new_new_n14443__ = ~new_new_n14441__ & ~new_new_n14442__;
  assign new_new_n14444__ = new_new_n14434__ & new_new_n14443__;
  assign new_new_n14445__ = ~new_new_n14434__ & ~new_new_n14443__;
  assign new_new_n14446__ = ~new_new_n14444__ & ~new_new_n14445__;
  assign new_new_n14447__ = pi39 & pi41;
  assign new_new_n14448__ = pi28 & pi52;
  assign new_new_n14449__ = pi27 & pi53;
  assign new_new_n14450__ = ~new_new_n14448__ & ~new_new_n14449__;
  assign new_new_n14451__ = new_new_n14448__ & new_new_n14449__;
  assign new_new_n14452__ = ~new_new_n14450__ & ~new_new_n14451__;
  assign new_new_n14453__ = new_new_n14447__ & ~new_new_n14452__;
  assign new_new_n14454__ = ~new_new_n14447__ & new_new_n14452__;
  assign new_new_n14455__ = ~new_new_n14453__ & ~new_new_n14454__;
  assign new_new_n14456__ = ~new_new_n14446__ & new_new_n14455__;
  assign new_new_n14457__ = new_new_n14446__ & ~new_new_n14455__;
  assign new_new_n14458__ = ~new_new_n14456__ & ~new_new_n14457__;
  assign new_new_n14459__ = pi36 & pi44;
  assign new_new_n14460__ = pi35 & pi45;
  assign new_new_n14461__ = pi34 & pi46;
  assign new_new_n14462__ = ~new_new_n14460__ & ~new_new_n14461__;
  assign new_new_n14463__ = new_new_n14460__ & new_new_n14461__;
  assign new_new_n14464__ = ~new_new_n14462__ & ~new_new_n14463__;
  assign new_new_n14465__ = new_new_n14459__ & ~new_new_n14464__;
  assign new_new_n14466__ = ~new_new_n14459__ & new_new_n14464__;
  assign new_new_n14467__ = ~new_new_n14465__ & ~new_new_n14466__;
  assign new_new_n14468__ = pi33 & pi47;
  assign new_new_n14469__ = pi29 & pi51;
  assign new_new_n14470__ = pi17 & pi63;
  assign new_new_n14471__ = ~new_new_n14469__ & ~new_new_n14470__;
  assign new_new_n14472__ = new_new_n14469__ & new_new_n14470__;
  assign new_new_n14473__ = ~new_new_n14471__ & ~new_new_n14472__;
  assign new_new_n14474__ = new_new_n14468__ & ~new_new_n14473__;
  assign new_new_n14475__ = ~new_new_n14468__ & new_new_n14473__;
  assign new_new_n14476__ = ~new_new_n14474__ & ~new_new_n14475__;
  assign new_new_n14477__ = new_new_n14467__ & new_new_n14476__;
  assign new_new_n14478__ = ~new_new_n14467__ & ~new_new_n14476__;
  assign new_new_n14479__ = ~new_new_n14477__ & ~new_new_n14478__;
  assign new_new_n14480__ = pi18 & pi62;
  assign new_new_n14481__ = pi19 & pi61;
  assign new_new_n14482__ = ~new_new_n14264__ & ~new_new_n14268__;
  assign new_new_n14483__ = new_new_n14481__ & new_new_n14482__;
  assign new_new_n14484__ = ~new_new_n14481__ & ~new_new_n14482__;
  assign new_new_n14485__ = ~new_new_n14483__ & ~new_new_n14484__;
  assign new_new_n14486__ = new_new_n14480__ & ~new_new_n14485__;
  assign new_new_n14487__ = ~new_new_n14480__ & new_new_n14485__;
  assign new_new_n14488__ = ~new_new_n14486__ & ~new_new_n14487__;
  assign new_new_n14489__ = new_new_n14479__ & ~new_new_n14488__;
  assign new_new_n14490__ = ~new_new_n14479__ & new_new_n14488__;
  assign new_new_n14491__ = ~new_new_n14489__ & ~new_new_n14490__;
  assign new_new_n14492__ = ~new_new_n14458__ & ~new_new_n14491__;
  assign new_new_n14493__ = new_new_n14458__ & new_new_n14491__;
  assign new_new_n14494__ = ~new_new_n14492__ & ~new_new_n14493__;
  assign new_new_n14495__ = pi32 & pi48;
  assign new_new_n14496__ = pi30 & pi50;
  assign new_new_n14497__ = pi31 & pi49;
  assign new_new_n14498__ = ~new_new_n14496__ & ~new_new_n14497__;
  assign new_new_n14499__ = new_new_n14496__ & new_new_n14497__;
  assign new_new_n14500__ = ~new_new_n14498__ & ~new_new_n14499__;
  assign new_new_n14501__ = new_new_n14495__ & ~new_new_n14500__;
  assign new_new_n14502__ = ~new_new_n14495__ & new_new_n14500__;
  assign new_new_n14503__ = ~new_new_n14501__ & ~new_new_n14502__;
  assign new_new_n14504__ = ~new_new_n14253__ & ~new_new_n14257__;
  assign new_new_n14505__ = ~new_new_n14256__ & ~new_new_n14504__;
  assign new_new_n14506__ = pi22 & pi58;
  assign new_new_n14507__ = pi20 & pi60;
  assign new_new_n14508__ = pi21 & pi59;
  assign new_new_n14509__ = ~new_new_n14507__ & ~new_new_n14508__;
  assign new_new_n14510__ = new_new_n14507__ & new_new_n14508__;
  assign new_new_n14511__ = ~new_new_n14509__ & ~new_new_n14510__;
  assign new_new_n14512__ = new_new_n14506__ & ~new_new_n14511__;
  assign new_new_n14513__ = ~new_new_n14506__ & new_new_n14511__;
  assign new_new_n14514__ = ~new_new_n14512__ & ~new_new_n14513__;
  assign new_new_n14515__ = new_new_n14505__ & ~new_new_n14514__;
  assign new_new_n14516__ = ~new_new_n14505__ & new_new_n14514__;
  assign new_new_n14517__ = ~new_new_n14515__ & ~new_new_n14516__;
  assign new_new_n14518__ = new_new_n14503__ & new_new_n14517__;
  assign new_new_n14519__ = ~new_new_n14503__ & ~new_new_n14517__;
  assign new_new_n14520__ = ~new_new_n14518__ & ~new_new_n14519__;
  assign new_new_n14521__ = new_new_n14494__ & ~new_new_n14520__;
  assign new_new_n14522__ = ~new_new_n14494__ & new_new_n14520__;
  assign new_new_n14523__ = ~new_new_n14521__ & ~new_new_n14522__;
  assign new_new_n14524__ = ~new_new_n14425__ & ~new_new_n14523__;
  assign new_new_n14525__ = new_new_n14425__ & new_new_n14523__;
  assign new_new_n14526__ = ~new_new_n14524__ & ~new_new_n14525__;
  assign new_new_n14527__ = ~new_new_n14307__ & ~new_new_n14311__;
  assign new_new_n14528__ = ~new_new_n14308__ & ~new_new_n14527__;
  assign new_new_n14529__ = new_new_n14526__ & ~new_new_n14528__;
  assign new_new_n14530__ = ~new_new_n14526__ & new_new_n14528__;
  assign new_new_n14531__ = ~new_new_n14529__ & ~new_new_n14530__;
  assign new_new_n14532__ = new_new_n14423__ & new_new_n14531__;
  assign new_new_n14533__ = ~new_new_n14423__ & ~new_new_n14531__;
  assign new_new_n14534__ = ~new_new_n14532__ & ~new_new_n14533__;
  assign new_new_n14535__ = new_new_n14317__ & ~new_new_n14413__;
  assign new_new_n14536__ = ~new_new_n14414__ & ~new_new_n14535__;
  assign new_new_n14537__ = ~new_new_n14213__ & ~new_new_n14418__;
  assign new_new_n14538__ = ~new_new_n14212__ & ~new_new_n14537__;
  assign new_new_n14539__ = ~new_new_n14536__ & ~new_new_n14538__;
  assign new_new_n14540__ = new_new_n14536__ & new_new_n14538__;
  assign new_new_n14541__ = ~new_new_n14539__ & ~new_new_n14540__;
  assign new_new_n14542__ = ~new_new_n14290__ & new_new_n14314__;
  assign new_new_n14543__ = ~new_new_n14291__ & ~new_new_n14542__;
  assign new_new_n14544__ = ~new_new_n14390__ & ~new_new_n14403__;
  assign new_new_n14545__ = ~new_new_n14389__ & ~new_new_n14544__;
  assign new_new_n14546__ = ~new_new_n14393__ & ~new_new_n14399__;
  assign new_new_n14547__ = ~new_new_n14398__ & ~new_new_n14546__;
  assign new_new_n14548__ = ~new_new_n14330__ & ~new_new_n14336__;
  assign new_new_n14549__ = ~new_new_n14335__ & ~new_new_n14548__;
  assign new_new_n14550__ = ~new_new_n14378__ & ~new_new_n14383__;
  assign new_new_n14551__ = ~new_new_n14384__ & ~new_new_n14550__;
  assign new_new_n14552__ = ~new_new_n14549__ & ~new_new_n14551__;
  assign new_new_n14553__ = new_new_n14549__ & new_new_n14551__;
  assign new_new_n14554__ = ~new_new_n14552__ & ~new_new_n14553__;
  assign new_new_n14555__ = new_new_n14547__ & ~new_new_n14554__;
  assign new_new_n14556__ = ~new_new_n14547__ & new_new_n14554__;
  assign new_new_n14557__ = ~new_new_n14555__ & ~new_new_n14556__;
  assign new_new_n14558__ = ~new_new_n14545__ & ~new_new_n14557__;
  assign new_new_n14559__ = new_new_n14545__ & new_new_n14557__;
  assign new_new_n14560__ = ~new_new_n14558__ & ~new_new_n14559__;
  assign new_new_n14561__ = ~new_new_n14367__ & new_new_n14371__;
  assign new_new_n14562__ = ~new_new_n14368__ & ~new_new_n14561__;
  assign new_new_n14563__ = new_new_n14560__ & new_new_n14562__;
  assign new_new_n14564__ = ~new_new_n14560__ & ~new_new_n14562__;
  assign new_new_n14565__ = ~new_new_n14563__ & ~new_new_n14564__;
  assign new_new_n14566__ = ~new_new_n14543__ & new_new_n14565__;
  assign new_new_n14567__ = new_new_n14543__ & ~new_new_n14565__;
  assign new_new_n14568__ = ~new_new_n14566__ & ~new_new_n14567__;
  assign new_new_n14569__ = ~new_new_n14251__ & new_new_n14284__;
  assign new_new_n14570__ = ~new_new_n14250__ & ~new_new_n14569__;
  assign new_new_n14571__ = ~new_new_n14261__ & ~new_new_n14279__;
  assign new_new_n14572__ = ~new_new_n14280__ & ~new_new_n14571__;
  assign new_new_n14573__ = ~new_new_n14235__ & ~new_new_n14246__;
  assign new_new_n14574__ = ~new_new_n14236__ & ~new_new_n14573__;
  assign new_new_n14575__ = new_new_n14572__ & ~new_new_n14574__;
  assign new_new_n14576__ = ~new_new_n14572__ & new_new_n14574__;
  assign new_new_n14577__ = ~new_new_n14575__ & ~new_new_n14576__;
  assign new_new_n14578__ = ~new_new_n14226__ & ~new_new_n14230__;
  assign new_new_n14579__ = ~new_new_n14229__ & ~new_new_n14578__;
  assign new_new_n14580__ = ~new_new_n14217__ & ~new_new_n14221__;
  assign new_new_n14581__ = ~new_new_n14220__ & ~new_new_n14580__;
  assign new_new_n14582__ = ~new_new_n14238__ & ~new_new_n14242__;
  assign new_new_n14583__ = ~new_new_n14241__ & ~new_new_n14582__;
  assign new_new_n14584__ = ~new_new_n14581__ & ~new_new_n14583__;
  assign new_new_n14585__ = new_new_n14581__ & new_new_n14583__;
  assign new_new_n14586__ = ~new_new_n14584__ & ~new_new_n14585__;
  assign new_new_n14587__ = new_new_n14579__ & ~new_new_n14586__;
  assign new_new_n14588__ = ~new_new_n14579__ & new_new_n14586__;
  assign new_new_n14589__ = ~new_new_n14587__ & ~new_new_n14588__;
  assign new_new_n14590__ = new_new_n14577__ & new_new_n14589__;
  assign new_new_n14591__ = ~new_new_n14577__ & ~new_new_n14589__;
  assign new_new_n14592__ = ~new_new_n14590__ & ~new_new_n14591__;
  assign new_new_n14593__ = new_new_n14342__ & ~new_new_n14361__;
  assign new_new_n14594__ = ~new_new_n14362__ & ~new_new_n14593__;
  assign new_new_n14595__ = ~new_new_n14296__ & ~new_new_n14301__;
  assign new_new_n14596__ = ~new_new_n14302__ & ~new_new_n14595__;
  assign new_new_n14597__ = new_new_n14594__ & ~new_new_n14596__;
  assign new_new_n14598__ = ~new_new_n14594__ & new_new_n14596__;
  assign new_new_n14599__ = ~new_new_n14597__ & ~new_new_n14598__;
  assign new_new_n14600__ = ~new_new_n14352__ & ~new_new_n14356__;
  assign new_new_n14601__ = ~new_new_n14355__ & ~new_new_n14600__;
  assign new_new_n14602__ = ~new_new_n14343__ & ~new_new_n14347__;
  assign new_new_n14603__ = ~new_new_n14346__ & ~new_new_n14602__;
  assign new_new_n14604__ = ~new_new_n7755__ & ~new_new_n14274__;
  assign new_new_n14605__ = ~new_new_n14273__ & ~new_new_n14604__;
  assign new_new_n14606__ = new_new_n14603__ & new_new_n14605__;
  assign new_new_n14607__ = ~new_new_n14603__ & ~new_new_n14605__;
  assign new_new_n14608__ = ~new_new_n14606__ & ~new_new_n14607__;
  assign new_new_n14609__ = new_new_n14601__ & ~new_new_n14608__;
  assign new_new_n14610__ = ~new_new_n14601__ & new_new_n14608__;
  assign new_new_n14611__ = ~new_new_n14609__ & ~new_new_n14610__;
  assign new_new_n14612__ = new_new_n14599__ & ~new_new_n14611__;
  assign new_new_n14613__ = ~new_new_n14599__ & new_new_n14611__;
  assign new_new_n14614__ = ~new_new_n14612__ & ~new_new_n14613__;
  assign new_new_n14615__ = new_new_n14592__ & new_new_n14614__;
  assign new_new_n14616__ = ~new_new_n14592__ & ~new_new_n14614__;
  assign new_new_n14617__ = ~new_new_n14615__ & ~new_new_n14616__;
  assign new_new_n14618__ = ~new_new_n14570__ & new_new_n14617__;
  assign new_new_n14619__ = new_new_n14570__ & ~new_new_n14617__;
  assign new_new_n14620__ = ~new_new_n14618__ & ~new_new_n14619__;
  assign new_new_n14621__ = new_new_n14568__ & new_new_n14620__;
  assign new_new_n14622__ = ~new_new_n14568__ & ~new_new_n14620__;
  assign new_new_n14623__ = ~new_new_n14621__ & ~new_new_n14622__;
  assign new_new_n14624__ = new_new_n14541__ & ~new_new_n14623__;
  assign new_new_n14625__ = ~new_new_n14541__ & new_new_n14623__;
  assign new_new_n14626__ = ~new_new_n14624__ & ~new_new_n14625__;
  assign new_new_n14627__ = new_new_n14534__ & new_new_n14626__;
  assign new_new_n14628__ = ~new_new_n14534__ & ~new_new_n14626__;
  assign po081 = new_new_n14627__ | new_new_n14628__;
  assign new_new_n14630__ = ~new_new_n14566__ & ~new_new_n14620__;
  assign new_new_n14631__ = ~new_new_n14567__ & ~new_new_n14630__;
  assign new_new_n14632__ = new_new_n14572__ & new_new_n14589__;
  assign new_new_n14633__ = ~new_new_n14574__ & ~new_new_n14632__;
  assign new_new_n14634__ = ~new_new_n14572__ & ~new_new_n14589__;
  assign new_new_n14635__ = ~new_new_n14633__ & ~new_new_n14634__;
  assign new_new_n14636__ = ~new_new_n14601__ & ~new_new_n14606__;
  assign new_new_n14637__ = ~new_new_n14607__ & ~new_new_n14636__;
  assign new_new_n14638__ = ~new_new_n14579__ & ~new_new_n14585__;
  assign new_new_n14639__ = ~new_new_n14584__ & ~new_new_n14638__;
  assign new_new_n14640__ = pi39 & pi42;
  assign new_new_n14641__ = pi38 & pi43;
  assign new_new_n14642__ = pi27 & pi54;
  assign new_new_n14643__ = ~new_new_n14641__ & ~new_new_n14642__;
  assign new_new_n14644__ = new_new_n14641__ & new_new_n14642__;
  assign new_new_n14645__ = ~new_new_n14643__ & ~new_new_n14644__;
  assign new_new_n14646__ = new_new_n14640__ & ~new_new_n14645__;
  assign new_new_n14647__ = ~new_new_n14640__ & new_new_n14645__;
  assign new_new_n14648__ = ~new_new_n14646__ & ~new_new_n14647__;
  assign new_new_n14649__ = ~new_new_n14639__ & new_new_n14648__;
  assign new_new_n14650__ = new_new_n14639__ & ~new_new_n14648__;
  assign new_new_n14651__ = ~new_new_n14649__ & ~new_new_n14650__;
  assign new_new_n14652__ = new_new_n14637__ & ~new_new_n14651__;
  assign new_new_n14653__ = ~new_new_n14637__ & new_new_n14651__;
  assign new_new_n14654__ = ~new_new_n14652__ & ~new_new_n14653__;
  assign new_new_n14655__ = ~new_new_n14635__ & ~new_new_n14654__;
  assign new_new_n14656__ = new_new_n14635__ & new_new_n14654__;
  assign new_new_n14657__ = ~new_new_n14655__ & ~new_new_n14656__;
  assign new_new_n14658__ = ~new_new_n14525__ & new_new_n14528__;
  assign new_new_n14659__ = ~new_new_n14524__ & ~new_new_n14658__;
  assign new_new_n14660__ = ~new_new_n14444__ & ~new_new_n14455__;
  assign new_new_n14661__ = ~new_new_n14445__ & ~new_new_n14660__;
  assign new_new_n14662__ = new_new_n14503__ & ~new_new_n14515__;
  assign new_new_n14663__ = ~new_new_n14516__ & ~new_new_n14662__;
  assign new_new_n14664__ = ~new_new_n14426__ & ~new_new_n14430__;
  assign new_new_n14665__ = ~new_new_n14429__ & ~new_new_n14664__;
  assign new_new_n14666__ = ~new_new_n14447__ & ~new_new_n14451__;
  assign new_new_n14667__ = ~new_new_n14450__ & ~new_new_n14666__;
  assign new_new_n14668__ = ~new_new_n14435__ & ~new_new_n14439__;
  assign new_new_n14669__ = ~new_new_n14438__ & ~new_new_n14668__;
  assign new_new_n14670__ = ~new_new_n14667__ & ~new_new_n14669__;
  assign new_new_n14671__ = new_new_n14667__ & new_new_n14669__;
  assign new_new_n14672__ = ~new_new_n14670__ & ~new_new_n14671__;
  assign new_new_n14673__ = new_new_n14665__ & ~new_new_n14672__;
  assign new_new_n14674__ = ~new_new_n14665__ & new_new_n14672__;
  assign new_new_n14675__ = ~new_new_n14673__ & ~new_new_n14674__;
  assign new_new_n14676__ = new_new_n14663__ & ~new_new_n14675__;
  assign new_new_n14677__ = ~new_new_n14663__ & new_new_n14675__;
  assign new_new_n14678__ = ~new_new_n14676__ & ~new_new_n14677__;
  assign new_new_n14679__ = new_new_n14661__ & ~new_new_n14678__;
  assign new_new_n14680__ = ~new_new_n14661__ & new_new_n14678__;
  assign new_new_n14681__ = ~new_new_n14679__ & ~new_new_n14680__;
  assign new_new_n14682__ = ~new_new_n14459__ & ~new_new_n14463__;
  assign new_new_n14683__ = ~new_new_n14462__ & ~new_new_n14682__;
  assign new_new_n14684__ = ~new_new_n14480__ & ~new_new_n14483__;
  assign new_new_n14685__ = ~new_new_n14484__ & ~new_new_n14684__;
  assign new_new_n14686__ = ~new_new_n14683__ & ~new_new_n14685__;
  assign new_new_n14687__ = new_new_n14683__ & new_new_n14685__;
  assign new_new_n14688__ = ~new_new_n14686__ & ~new_new_n14687__;
  assign new_new_n14689__ = pi32 & pi49;
  assign new_new_n14690__ = pi31 & pi50;
  assign new_new_n14691__ = pi30 & pi51;
  assign new_new_n14692__ = ~new_new_n14690__ & ~new_new_n14691__;
  assign new_new_n14693__ = new_new_n14690__ & new_new_n14691__;
  assign new_new_n14694__ = ~new_new_n14692__ & ~new_new_n14693__;
  assign new_new_n14695__ = new_new_n14689__ & ~new_new_n14694__;
  assign new_new_n14696__ = ~new_new_n14689__ & new_new_n14694__;
  assign new_new_n14697__ = ~new_new_n14695__ & ~new_new_n14696__;
  assign new_new_n14698__ = new_new_n14688__ & new_new_n14697__;
  assign new_new_n14699__ = ~new_new_n14688__ & ~new_new_n14697__;
  assign new_new_n14700__ = ~new_new_n14698__ & ~new_new_n14699__;
  assign new_new_n14701__ = new_new_n14681__ & ~new_new_n14700__;
  assign new_new_n14702__ = ~new_new_n14681__ & new_new_n14700__;
  assign new_new_n14703__ = ~new_new_n14701__ & ~new_new_n14702__;
  assign new_new_n14704__ = ~new_new_n14495__ & ~new_new_n14499__;
  assign new_new_n14705__ = ~new_new_n14498__ & ~new_new_n14704__;
  assign new_new_n14706__ = ~new_new_n14506__ & ~new_new_n14510__;
  assign new_new_n14707__ = ~new_new_n14509__ & ~new_new_n14706__;
  assign new_new_n14708__ = ~new_new_n14705__ & ~new_new_n14707__;
  assign new_new_n14709__ = new_new_n14705__ & new_new_n14707__;
  assign new_new_n14710__ = ~new_new_n14708__ & ~new_new_n14709__;
  assign new_new_n14711__ = ~new_new_n14468__ & ~new_new_n14472__;
  assign new_new_n14712__ = ~new_new_n14471__ & ~new_new_n14711__;
  assign new_new_n14713__ = ~new_new_n14710__ & new_new_n14712__;
  assign new_new_n14714__ = new_new_n14710__ & ~new_new_n14712__;
  assign new_new_n14715__ = ~new_new_n14713__ & ~new_new_n14714__;
  assign new_new_n14716__ = ~new_new_n14477__ & ~new_new_n14488__;
  assign new_new_n14717__ = ~new_new_n14478__ & ~new_new_n14716__;
  assign new_new_n14718__ = ~new_new_n14715__ & ~new_new_n14717__;
  assign new_new_n14719__ = new_new_n14715__ & new_new_n14717__;
  assign new_new_n14720__ = ~new_new_n14718__ & ~new_new_n14719__;
  assign new_new_n14721__ = ~new_new_n14493__ & new_new_n14520__;
  assign new_new_n14722__ = ~new_new_n14492__ & ~new_new_n14721__;
  assign new_new_n14723__ = new_new_n14720__ & ~new_new_n14722__;
  assign new_new_n14724__ = ~new_new_n14720__ & new_new_n14722__;
  assign new_new_n14725__ = ~new_new_n14723__ & ~new_new_n14724__;
  assign new_new_n14726__ = new_new_n14703__ & new_new_n14725__;
  assign new_new_n14727__ = ~new_new_n14703__ & ~new_new_n14725__;
  assign new_new_n14728__ = ~new_new_n14726__ & ~new_new_n14727__;
  assign new_new_n14729__ = ~new_new_n14659__ & new_new_n14728__;
  assign new_new_n14730__ = new_new_n14659__ & ~new_new_n14728__;
  assign new_new_n14731__ = ~new_new_n14729__ & ~new_new_n14730__;
  assign new_new_n14732__ = ~new_new_n14598__ & new_new_n14611__;
  assign new_new_n14733__ = ~new_new_n14597__ & ~new_new_n14732__;
  assign new_new_n14734__ = new_new_n14731__ & ~new_new_n14733__;
  assign new_new_n14735__ = ~new_new_n14731__ & new_new_n14733__;
  assign new_new_n14736__ = ~new_new_n14734__ & ~new_new_n14735__;
  assign new_new_n14737__ = new_new_n14657__ & new_new_n14736__;
  assign new_new_n14738__ = ~new_new_n14657__ & ~new_new_n14736__;
  assign new_new_n14739__ = ~new_new_n14737__ & ~new_new_n14738__;
  assign new_new_n14740__ = ~new_new_n14631__ & new_new_n14739__;
  assign new_new_n14741__ = new_new_n14631__ & ~new_new_n14739__;
  assign new_new_n14742__ = ~new_new_n14740__ & ~new_new_n14741__;
  assign new_new_n14743__ = ~new_new_n14570__ & ~new_new_n14616__;
  assign new_new_n14744__ = ~new_new_n14615__ & ~new_new_n14743__;
  assign new_new_n14745__ = ~new_new_n14547__ & ~new_new_n14553__;
  assign new_new_n14746__ = ~new_new_n14552__ & ~new_new_n14745__;
  assign new_new_n14747__ = pi34 & pi47;
  assign new_new_n14748__ = pi24 & pi57;
  assign new_new_n14749__ = pi33 & pi48;
  assign new_new_n14750__ = ~new_new_n14748__ & ~new_new_n14749__;
  assign new_new_n14751__ = new_new_n14748__ & new_new_n14749__;
  assign new_new_n14752__ = ~new_new_n14750__ & ~new_new_n14751__;
  assign new_new_n14753__ = new_new_n14747__ & ~new_new_n14752__;
  assign new_new_n14754__ = ~new_new_n14747__ & new_new_n14752__;
  assign new_new_n14755__ = ~new_new_n14753__ & ~new_new_n14754__;
  assign new_new_n14756__ = pi25 & pi56;
  assign new_new_n14757__ = pi23 & pi58;
  assign new_new_n14758__ = pi22 & pi59;
  assign new_new_n14759__ = ~new_new_n14757__ & ~new_new_n14758__;
  assign new_new_n14760__ = new_new_n14757__ & new_new_n14758__;
  assign new_new_n14761__ = ~new_new_n14759__ & ~new_new_n14760__;
  assign new_new_n14762__ = new_new_n14756__ & ~new_new_n14761__;
  assign new_new_n14763__ = ~new_new_n14756__ & new_new_n14761__;
  assign new_new_n14764__ = ~new_new_n14762__ & ~new_new_n14763__;
  assign new_new_n14765__ = new_new_n14755__ & new_new_n14764__;
  assign new_new_n14766__ = ~new_new_n14755__ & ~new_new_n14764__;
  assign new_new_n14767__ = ~new_new_n14765__ & ~new_new_n14766__;
  assign new_new_n14768__ = pi19 & pi62;
  assign new_new_n14769__ = ~pi40 & pi41;
  assign new_new_n14770__ = new_new_n14768__ & ~new_new_n14769__;
  assign new_new_n14771__ = ~new_new_n14768__ & new_new_n14769__;
  assign new_new_n14772__ = ~new_new_n14770__ & ~new_new_n14771__;
  assign new_new_n14773__ = ~new_new_n14767__ & new_new_n14772__;
  assign new_new_n14774__ = new_new_n14767__ & ~new_new_n14772__;
  assign new_new_n14775__ = ~new_new_n14773__ & ~new_new_n14774__;
  assign new_new_n14776__ = new_new_n14746__ & new_new_n14775__;
  assign new_new_n14777__ = ~new_new_n14746__ & ~new_new_n14775__;
  assign new_new_n14778__ = ~new_new_n14776__ & ~new_new_n14777__;
  assign new_new_n14779__ = pi37 & pi44;
  assign new_new_n14780__ = pi35 & pi46;
  assign new_new_n14781__ = pi36 & pi45;
  assign new_new_n14782__ = ~new_new_n14780__ & ~new_new_n14781__;
  assign new_new_n14783__ = new_new_n14780__ & new_new_n14781__;
  assign new_new_n14784__ = ~new_new_n14782__ & ~new_new_n14783__;
  assign new_new_n14785__ = new_new_n14779__ & ~new_new_n14784__;
  assign new_new_n14786__ = ~new_new_n14779__ & new_new_n14784__;
  assign new_new_n14787__ = ~new_new_n14785__ & ~new_new_n14786__;
  assign new_new_n14788__ = pi29 & pi52;
  assign new_new_n14789__ = pi28 & pi53;
  assign new_new_n14790__ = pi26 & pi55;
  assign new_new_n14791__ = ~new_new_n14789__ & ~new_new_n14790__;
  assign new_new_n14792__ = new_new_n14789__ & new_new_n14790__;
  assign new_new_n14793__ = ~new_new_n14791__ & ~new_new_n14792__;
  assign new_new_n14794__ = new_new_n14788__ & ~new_new_n14793__;
  assign new_new_n14795__ = ~new_new_n14788__ & new_new_n14793__;
  assign new_new_n14796__ = ~new_new_n14794__ & ~new_new_n14795__;
  assign new_new_n14797__ = ~new_new_n14787__ & ~new_new_n14796__;
  assign new_new_n14798__ = new_new_n14787__ & new_new_n14796__;
  assign new_new_n14799__ = ~new_new_n14797__ & ~new_new_n14798__;
  assign new_new_n14800__ = pi21 & pi60;
  assign new_new_n14801__ = pi20 & pi61;
  assign new_new_n14802__ = pi18 & pi63;
  assign new_new_n14803__ = ~new_new_n14801__ & ~new_new_n14802__;
  assign new_new_n14804__ = new_new_n14801__ & new_new_n14802__;
  assign new_new_n14805__ = ~new_new_n14803__ & ~new_new_n14804__;
  assign new_new_n14806__ = new_new_n14800__ & ~new_new_n14805__;
  assign new_new_n14807__ = ~new_new_n14800__ & new_new_n14805__;
  assign new_new_n14808__ = ~new_new_n14806__ & ~new_new_n14807__;
  assign new_new_n14809__ = new_new_n14799__ & ~new_new_n14808__;
  assign new_new_n14810__ = ~new_new_n14799__ & new_new_n14808__;
  assign new_new_n14811__ = ~new_new_n14809__ & ~new_new_n14810__;
  assign new_new_n14812__ = new_new_n14778__ & ~new_new_n14811__;
  assign new_new_n14813__ = ~new_new_n14778__ & new_new_n14811__;
  assign new_new_n14814__ = ~new_new_n14812__ & ~new_new_n14813__;
  assign new_new_n14815__ = new_new_n14744__ & new_new_n14814__;
  assign new_new_n14816__ = ~new_new_n14744__ & ~new_new_n14814__;
  assign new_new_n14817__ = ~new_new_n14815__ & ~new_new_n14816__;
  assign new_new_n14818__ = ~new_new_n14558__ & ~new_new_n14562__;
  assign new_new_n14819__ = ~new_new_n14559__ & ~new_new_n14818__;
  assign new_new_n14820__ = new_new_n14817__ & ~new_new_n14819__;
  assign new_new_n14821__ = ~new_new_n14817__ & new_new_n14819__;
  assign new_new_n14822__ = ~new_new_n14820__ & ~new_new_n14821__;
  assign new_new_n14823__ = new_new_n14742__ & ~new_new_n14822__;
  assign new_new_n14824__ = ~new_new_n14742__ & new_new_n14822__;
  assign new_new_n14825__ = ~new_new_n14823__ & ~new_new_n14824__;
  assign new_new_n14826__ = new_new_n14532__ & new_new_n14623__;
  assign new_new_n14827__ = new_new_n14533__ & ~new_new_n14623__;
  assign new_new_n14828__ = ~new_new_n14826__ & ~new_new_n14827__;
  assign new_new_n14829__ = new_new_n14541__ & new_new_n14828__;
  assign new_new_n14830__ = ~new_new_n14532__ & ~new_new_n14623__;
  assign new_new_n14831__ = ~new_new_n14533__ & ~new_new_n14830__;
  assign new_new_n14832__ = new_new_n14540__ & ~new_new_n14831__;
  assign new_new_n14833__ = new_new_n14539__ & new_new_n14831__;
  assign new_new_n14834__ = ~new_new_n14832__ & ~new_new_n14833__;
  assign new_new_n14835__ = ~new_new_n14829__ & new_new_n14834__;
  assign new_new_n14836__ = ~new_new_n14825__ & ~new_new_n14835__;
  assign new_new_n14837__ = ~new_new_n14531__ & ~new_new_n14538__;
  assign new_new_n14838__ = ~new_new_n14536__ & new_new_n14837__;
  assign new_new_n14839__ = ~new_new_n14423__ & new_new_n14838__;
  assign new_new_n14840__ = ~new_new_n14531__ & ~new_new_n14540__;
  assign new_new_n14841__ = ~new_new_n14539__ & ~new_new_n14840__;
  assign new_new_n14842__ = new_new_n14423__ & new_new_n14841__;
  assign new_new_n14843__ = new_new_n14531__ & new_new_n14538__;
  assign new_new_n14844__ = new_new_n14536__ & new_new_n14843__;
  assign new_new_n14845__ = ~new_new_n14842__ & ~new_new_n14844__;
  assign new_new_n14846__ = new_new_n14623__ & ~new_new_n14845__;
  assign new_new_n14847__ = ~new_new_n14423__ & ~new_new_n14841__;
  assign new_new_n14848__ = ~new_new_n14838__ & ~new_new_n14847__;
  assign new_new_n14849__ = ~new_new_n14623__ & ~new_new_n14848__;
  assign new_new_n14850__ = new_new_n14423__ & new_new_n14536__;
  assign new_new_n14851__ = new_new_n14843__ & new_new_n14850__;
  assign new_new_n14852__ = ~new_new_n14839__ & ~new_new_n14851__;
  assign new_new_n14853__ = ~new_new_n14846__ & new_new_n14852__;
  assign new_new_n14854__ = ~new_new_n14849__ & new_new_n14853__;
  assign new_new_n14855__ = new_new_n14825__ & ~new_new_n14854__;
  assign po082 = new_new_n14836__ | new_new_n14855__;
  assign new_new_n14857__ = ~new_new_n14741__ & new_new_n14822__;
  assign new_new_n14858__ = ~new_new_n14740__ & ~new_new_n14857__;
  assign new_new_n14859__ = ~new_new_n14423__ & ~new_new_n14536__;
  assign new_new_n14860__ = new_new_n14623__ & ~new_new_n14859__;
  assign new_new_n14861__ = new_new_n14825__ & ~new_new_n14837__;
  assign new_new_n14862__ = ~new_new_n14850__ & ~new_new_n14860__;
  assign new_new_n14863__ = ~new_new_n14861__ & new_new_n14862__;
  assign new_new_n14864__ = ~new_new_n14623__ & new_new_n14859__;
  assign new_new_n14865__ = new_new_n14825__ & ~new_new_n14864__;
  assign new_new_n14866__ = new_new_n14623__ & new_new_n14850__;
  assign new_new_n14867__ = ~new_new_n14865__ & ~new_new_n14866__;
  assign new_new_n14868__ = ~new_new_n14843__ & new_new_n14867__;
  assign new_new_n14869__ = ~new_new_n14825__ & new_new_n14837__;
  assign new_new_n14870__ = ~new_new_n14868__ & ~new_new_n14869__;
  assign new_new_n14871__ = ~new_new_n14863__ & new_new_n14870__;
  assign new_new_n14872__ = new_new_n14858__ & new_new_n14871__;
  assign new_new_n14873__ = ~new_new_n14858__ & ~new_new_n14871__;
  assign new_new_n14874__ = ~new_new_n14872__ & ~new_new_n14873__;
  assign new_new_n14875__ = new_new_n14657__ & ~new_new_n14733__;
  assign new_new_n14876__ = ~new_new_n14657__ & new_new_n14733__;
  assign new_new_n14877__ = ~new_new_n14875__ & ~new_new_n14876__;
  assign new_new_n14878__ = ~new_new_n14730__ & new_new_n14877__;
  assign new_new_n14879__ = ~new_new_n14729__ & ~new_new_n14878__;
  assign new_new_n14880__ = ~new_new_n14661__ & ~new_new_n14677__;
  assign new_new_n14881__ = ~new_new_n14676__ & ~new_new_n14880__;
  assign new_new_n14882__ = ~new_new_n14700__ & ~new_new_n14719__;
  assign new_new_n14883__ = ~new_new_n14718__ & ~new_new_n14882__;
  assign new_new_n14884__ = new_new_n14881__ & new_new_n14883__;
  assign new_new_n14885__ = ~new_new_n14881__ & ~new_new_n14883__;
  assign new_new_n14886__ = ~new_new_n14884__ & ~new_new_n14885__;
  assign new_new_n14887__ = ~new_new_n14709__ & ~new_new_n14712__;
  assign new_new_n14888__ = ~new_new_n14708__ & ~new_new_n14887__;
  assign new_new_n14889__ = ~new_new_n14665__ & ~new_new_n14671__;
  assign new_new_n14890__ = ~new_new_n14670__ & ~new_new_n14889__;
  assign new_new_n14891__ = ~new_new_n14888__ & ~new_new_n14890__;
  assign new_new_n14892__ = new_new_n14888__ & new_new_n14890__;
  assign new_new_n14893__ = ~new_new_n14891__ & ~new_new_n14892__;
  assign new_new_n14894__ = pi25 & pi57;
  assign new_new_n14895__ = ~new_new_n8363__ & ~new_new_n14894__;
  assign new_new_n14896__ = new_new_n8363__ & new_new_n14894__;
  assign new_new_n14897__ = ~new_new_n14895__ & ~new_new_n14896__;
  assign new_new_n14898__ = new_new_n7761__ & ~new_new_n14897__;
  assign new_new_n14899__ = ~new_new_n7761__ & new_new_n14897__;
  assign new_new_n14900__ = ~new_new_n14898__ & ~new_new_n14899__;
  assign new_new_n14901__ = new_new_n14893__ & new_new_n14900__;
  assign new_new_n14902__ = ~new_new_n14893__ & ~new_new_n14900__;
  assign new_new_n14903__ = ~new_new_n14901__ & ~new_new_n14902__;
  assign new_new_n14904__ = new_new_n14886__ & ~new_new_n14903__;
  assign new_new_n14905__ = ~new_new_n14886__ & new_new_n14903__;
  assign new_new_n14906__ = ~new_new_n14904__ & ~new_new_n14905__;
  assign new_new_n14907__ = ~new_new_n14776__ & ~new_new_n14811__;
  assign new_new_n14908__ = ~new_new_n14777__ & ~new_new_n14907__;
  assign new_new_n14909__ = ~new_new_n14765__ & ~new_new_n14772__;
  assign new_new_n14910__ = ~new_new_n14766__ & ~new_new_n14909__;
  assign new_new_n14911__ = ~new_new_n14640__ & ~new_new_n14644__;
  assign new_new_n14912__ = ~new_new_n14643__ & ~new_new_n14911__;
  assign new_new_n14913__ = pi63 & new_new_n14912__;
  assign new_new_n14914__ = pi19 & new_new_n14913__;
  assign new_new_n14915__ = ~pi63 & ~new_new_n14912__;
  assign new_new_n14916__ = ~pi19 & ~new_new_n14912__;
  assign new_new_n14917__ = ~new_new_n14915__ & ~new_new_n14916__;
  assign new_new_n14918__ = ~new_new_n14914__ & new_new_n14917__;
  assign new_new_n14919__ = pi40 & ~new_new_n14918__;
  assign new_new_n14920__ = ~pi40 & new_new_n14913__;
  assign new_new_n14921__ = pi19 & new_new_n14915__;
  assign new_new_n14922__ = ~new_new_n14920__ & ~new_new_n14921__;
  assign new_new_n14923__ = pi62 & ~new_new_n14922__;
  assign new_new_n14924__ = ~new_new_n14919__ & ~new_new_n14923__;
  assign new_new_n14925__ = pi41 & ~new_new_n14924__;
  assign new_new_n14926__ = pi40 & pi41;
  assign new_new_n14927__ = pi41 & pi62;
  assign new_new_n14928__ = ~new_new_n14913__ & ~new_new_n14927__;
  assign new_new_n14929__ = pi19 & ~new_new_n14928__;
  assign new_new_n14930__ = new_new_n14917__ & ~new_new_n14926__;
  assign new_new_n14931__ = ~new_new_n14929__ & new_new_n14930__;
  assign new_new_n14932__ = ~new_new_n14925__ & ~new_new_n14931__;
  assign new_new_n14933__ = new_new_n14910__ & new_new_n14932__;
  assign new_new_n14934__ = ~new_new_n14686__ & ~new_new_n14697__;
  assign new_new_n14935__ = ~new_new_n14910__ & ~new_new_n14932__;
  assign new_new_n14936__ = ~new_new_n14687__ & ~new_new_n14934__;
  assign new_new_n14937__ = ~new_new_n14935__ & new_new_n14936__;
  assign new_new_n14938__ = ~new_new_n14933__ & new_new_n14937__;
  assign new_new_n14939__ = new_new_n14683__ & new_new_n14933__;
  assign new_new_n14940__ = ~new_new_n14697__ & new_new_n14935__;
  assign new_new_n14941__ = ~new_new_n14939__ & ~new_new_n14940__;
  assign new_new_n14942__ = new_new_n14685__ & ~new_new_n14941__;
  assign new_new_n14943__ = new_new_n14683__ & new_new_n14935__;
  assign new_new_n14944__ = new_new_n14688__ & new_new_n14933__;
  assign new_new_n14945__ = ~new_new_n14943__ & ~new_new_n14944__;
  assign new_new_n14946__ = new_new_n14700__ & ~new_new_n14945__;
  assign new_new_n14947__ = ~new_new_n14938__ & ~new_new_n14942__;
  assign new_new_n14948__ = ~new_new_n14946__ & new_new_n14947__;
  assign new_new_n14949__ = new_new_n14908__ & ~new_new_n14948__;
  assign new_new_n14950__ = ~new_new_n14908__ & new_new_n14948__;
  assign new_new_n14951__ = ~new_new_n14949__ & ~new_new_n14950__;
  assign new_new_n14952__ = ~new_new_n14779__ & ~new_new_n14783__;
  assign new_new_n14953__ = ~new_new_n14782__ & ~new_new_n14952__;
  assign new_new_n14954__ = ~new_new_n14798__ & ~new_new_n14808__;
  assign new_new_n14955__ = ~new_new_n14797__ & ~new_new_n14954__;
  assign new_new_n14956__ = new_new_n14953__ & ~new_new_n14955__;
  assign new_new_n14957__ = ~new_new_n14953__ & new_new_n14955__;
  assign new_new_n14958__ = ~new_new_n14956__ & ~new_new_n14957__;
  assign new_new_n14959__ = ~new_new_n14756__ & ~new_new_n14760__;
  assign new_new_n14960__ = ~new_new_n14759__ & ~new_new_n14959__;
  assign new_new_n14961__ = ~new_new_n14689__ & ~new_new_n14693__;
  assign new_new_n14962__ = ~new_new_n14692__ & ~new_new_n14961__;
  assign new_new_n14963__ = ~new_new_n14747__ & ~new_new_n14751__;
  assign new_new_n14964__ = ~new_new_n14750__ & ~new_new_n14963__;
  assign new_new_n14965__ = ~new_new_n14788__ & ~new_new_n14792__;
  assign new_new_n14966__ = ~new_new_n14791__ & ~new_new_n14965__;
  assign new_new_n14967__ = new_new_n14964__ & new_new_n14966__;
  assign new_new_n14968__ = ~new_new_n14964__ & ~new_new_n14966__;
  assign new_new_n14969__ = ~new_new_n14962__ & ~new_new_n14967__;
  assign new_new_n14970__ = ~new_new_n14968__ & ~new_new_n14969__;
  assign new_new_n14971__ = ~new_new_n14967__ & new_new_n14970__;
  assign new_new_n14972__ = new_new_n14962__ & ~new_new_n14971__;
  assign new_new_n14973__ = ~new_new_n14968__ & new_new_n14969__;
  assign new_new_n14974__ = ~new_new_n14972__ & ~new_new_n14973__;
  assign new_new_n14975__ = ~new_new_n14800__ & ~new_new_n14804__;
  assign new_new_n14976__ = ~new_new_n14803__ & ~new_new_n14975__;
  assign new_new_n14977__ = new_new_n14974__ & ~new_new_n14976__;
  assign new_new_n14978__ = ~new_new_n14974__ & new_new_n14976__;
  assign new_new_n14979__ = ~new_new_n14977__ & ~new_new_n14978__;
  assign new_new_n14980__ = new_new_n14960__ & ~new_new_n14979__;
  assign new_new_n14981__ = ~new_new_n14960__ & new_new_n14979__;
  assign new_new_n14982__ = ~new_new_n14980__ & ~new_new_n14981__;
  assign new_new_n14983__ = new_new_n14958__ & new_new_n14982__;
  assign new_new_n14984__ = ~new_new_n14958__ & ~new_new_n14982__;
  assign new_new_n14985__ = ~new_new_n14983__ & ~new_new_n14984__;
  assign new_new_n14986__ = ~new_new_n14951__ & new_new_n14985__;
  assign new_new_n14987__ = new_new_n14951__ & ~new_new_n14985__;
  assign new_new_n14988__ = ~new_new_n14986__ & ~new_new_n14987__;
  assign new_new_n14989__ = new_new_n14906__ & new_new_n14988__;
  assign new_new_n14990__ = ~new_new_n14906__ & ~new_new_n14988__;
  assign new_new_n14991__ = ~new_new_n14989__ & ~new_new_n14990__;
  assign new_new_n14992__ = ~new_new_n14816__ & ~new_new_n14819__;
  assign new_new_n14993__ = ~new_new_n14815__ & ~new_new_n14992__;
  assign new_new_n14994__ = new_new_n14991__ & ~new_new_n14993__;
  assign new_new_n14995__ = ~new_new_n14991__ & new_new_n14993__;
  assign new_new_n14996__ = ~new_new_n14994__ & ~new_new_n14995__;
  assign new_new_n14997__ = new_new_n14879__ & ~new_new_n14996__;
  assign new_new_n14998__ = ~new_new_n14879__ & new_new_n14996__;
  assign new_new_n14999__ = ~new_new_n14997__ & ~new_new_n14998__;
  assign new_new_n15000__ = ~new_new_n14656__ & new_new_n14733__;
  assign new_new_n15001__ = ~new_new_n14655__ & ~new_new_n15000__;
  assign new_new_n15002__ = ~new_new_n14681__ & ~new_new_n14722__;
  assign new_new_n15003__ = new_new_n14681__ & new_new_n14722__;
  assign new_new_n15004__ = new_new_n14700__ & new_new_n14720__;
  assign new_new_n15005__ = ~new_new_n14700__ & ~new_new_n14720__;
  assign new_new_n15006__ = ~new_new_n15004__ & ~new_new_n15005__;
  assign new_new_n15007__ = ~new_new_n15003__ & new_new_n15006__;
  assign new_new_n15008__ = ~new_new_n15002__ & ~new_new_n15007__;
  assign new_new_n15009__ = ~new_new_n15001__ & new_new_n15008__;
  assign new_new_n15010__ = new_new_n15001__ & ~new_new_n15008__;
  assign new_new_n15011__ = ~new_new_n15009__ & ~new_new_n15010__;
  assign new_new_n15012__ = new_new_n14637__ & ~new_new_n14649__;
  assign new_new_n15013__ = ~new_new_n14650__ & ~new_new_n15012__;
  assign new_new_n15014__ = pi37 & pi45;
  assign new_new_n15015__ = pi36 & pi46;
  assign new_new_n15016__ = pi35 & pi47;
  assign new_new_n15017__ = ~new_new_n15015__ & ~new_new_n15016__;
  assign new_new_n15018__ = new_new_n15015__ & new_new_n15016__;
  assign new_new_n15019__ = ~new_new_n15017__ & ~new_new_n15018__;
  assign new_new_n15020__ = new_new_n15014__ & ~new_new_n15019__;
  assign new_new_n15021__ = ~new_new_n15014__ & new_new_n15019__;
  assign new_new_n15022__ = ~new_new_n15020__ & ~new_new_n15021__;
  assign new_new_n15023__ = pi39 & pi43;
  assign new_new_n15024__ = pi26 & pi56;
  assign new_new_n15025__ = pi38 & pi44;
  assign new_new_n15026__ = ~new_new_n15024__ & ~new_new_n15025__;
  assign new_new_n15027__ = new_new_n15024__ & new_new_n15025__;
  assign new_new_n15028__ = ~new_new_n15026__ & ~new_new_n15027__;
  assign new_new_n15029__ = new_new_n15023__ & ~new_new_n15028__;
  assign new_new_n15030__ = ~new_new_n15023__ & new_new_n15028__;
  assign new_new_n15031__ = ~new_new_n15029__ & ~new_new_n15030__;
  assign new_new_n15032__ = new_new_n15022__ & new_new_n15031__;
  assign new_new_n15033__ = ~new_new_n15022__ & ~new_new_n15031__;
  assign new_new_n15034__ = ~new_new_n15032__ & ~new_new_n15033__;
  assign new_new_n15035__ = pi40 & pi42;
  assign new_new_n15036__ = pi30 & pi52;
  assign new_new_n15037__ = pi29 & pi53;
  assign new_new_n15038__ = ~new_new_n15036__ & ~new_new_n15037__;
  assign new_new_n15039__ = new_new_n15036__ & new_new_n15037__;
  assign new_new_n15040__ = ~new_new_n15038__ & ~new_new_n15039__;
  assign new_new_n15041__ = new_new_n15035__ & ~new_new_n15040__;
  assign new_new_n15042__ = ~new_new_n15035__ & new_new_n15040__;
  assign new_new_n15043__ = ~new_new_n15041__ & ~new_new_n15042__;
  assign new_new_n15044__ = new_new_n15034__ & ~new_new_n15043__;
  assign new_new_n15045__ = ~new_new_n15034__ & new_new_n15043__;
  assign new_new_n15046__ = ~new_new_n15044__ & ~new_new_n15045__;
  assign new_new_n15047__ = ~new_new_n15013__ & new_new_n15046__;
  assign new_new_n15048__ = new_new_n15013__ & ~new_new_n15046__;
  assign new_new_n15049__ = ~new_new_n15047__ & ~new_new_n15048__;
  assign new_new_n15050__ = pi24 & pi58;
  assign new_new_n15051__ = pi23 & pi59;
  assign new_new_n15052__ = pi22 & pi60;
  assign new_new_n15053__ = ~new_new_n15051__ & ~new_new_n15052__;
  assign new_new_n15054__ = new_new_n15051__ & new_new_n15052__;
  assign new_new_n15055__ = ~new_new_n15053__ & ~new_new_n15054__;
  assign new_new_n15056__ = new_new_n15050__ & ~new_new_n15055__;
  assign new_new_n15057__ = ~new_new_n15050__ & new_new_n15055__;
  assign new_new_n15058__ = ~new_new_n15056__ & ~new_new_n15057__;
  assign new_new_n15059__ = pi34 & pi48;
  assign new_new_n15060__ = pi33 & pi49;
  assign new_new_n15061__ = pi32 & pi50;
  assign new_new_n15062__ = ~new_new_n15060__ & ~new_new_n15061__;
  assign new_new_n15063__ = new_new_n15060__ & new_new_n15061__;
  assign new_new_n15064__ = ~new_new_n15062__ & ~new_new_n15063__;
  assign new_new_n15065__ = new_new_n15059__ & ~new_new_n15064__;
  assign new_new_n15066__ = ~new_new_n15059__ & new_new_n15064__;
  assign new_new_n15067__ = ~new_new_n15065__ & ~new_new_n15066__;
  assign new_new_n15068__ = new_new_n15058__ & new_new_n15067__;
  assign new_new_n15069__ = ~new_new_n15058__ & ~new_new_n15067__;
  assign new_new_n15070__ = ~new_new_n15068__ & ~new_new_n15069__;
  assign new_new_n15071__ = pi31 & pi51;
  assign new_new_n15072__ = pi21 & pi61;
  assign new_new_n15073__ = pi20 & pi62;
  assign new_new_n15074__ = ~new_new_n15072__ & ~new_new_n15073__;
  assign new_new_n15075__ = new_new_n15072__ & new_new_n15073__;
  assign new_new_n15076__ = ~new_new_n15074__ & ~new_new_n15075__;
  assign new_new_n15077__ = new_new_n15071__ & ~new_new_n15076__;
  assign new_new_n15078__ = ~new_new_n15071__ & new_new_n15076__;
  assign new_new_n15079__ = ~new_new_n15077__ & ~new_new_n15078__;
  assign new_new_n15080__ = ~new_new_n15070__ & new_new_n15079__;
  assign new_new_n15081__ = new_new_n15070__ & ~new_new_n15079__;
  assign new_new_n15082__ = ~new_new_n15080__ & ~new_new_n15081__;
  assign new_new_n15083__ = new_new_n15049__ & new_new_n15082__;
  assign new_new_n15084__ = ~new_new_n15049__ & ~new_new_n15082__;
  assign new_new_n15085__ = ~new_new_n15083__ & ~new_new_n15084__;
  assign new_new_n15086__ = new_new_n15011__ & ~new_new_n15085__;
  assign new_new_n15087__ = ~new_new_n15011__ & new_new_n15085__;
  assign new_new_n15088__ = ~new_new_n15086__ & ~new_new_n15087__;
  assign new_new_n15089__ = new_new_n14999__ & ~new_new_n15088__;
  assign new_new_n15090__ = ~new_new_n14999__ & new_new_n15088__;
  assign new_new_n15091__ = ~new_new_n15089__ & ~new_new_n15090__;
  assign new_new_n15092__ = new_new_n14874__ & new_new_n15091__;
  assign new_new_n15093__ = ~new_new_n14874__ & ~new_new_n15091__;
  assign po083 = ~new_new_n15092__ & ~new_new_n15093__;
  assign new_new_n15095__ = ~new_new_n14998__ & ~new_new_n15088__;
  assign new_new_n15096__ = ~new_new_n14997__ & ~new_new_n15095__;
  assign new_new_n15097__ = new_new_n14872__ & new_new_n15096__;
  assign new_new_n15098__ = new_new_n14998__ & new_new_n15088__;
  assign new_new_n15099__ = new_new_n14997__ & ~new_new_n15088__;
  assign new_new_n15100__ = ~new_new_n15098__ & ~new_new_n15099__;
  assign new_new_n15101__ = new_new_n14874__ & new_new_n15100__;
  assign new_new_n15102__ = new_new_n14873__ & ~new_new_n15096__;
  assign new_new_n15103__ = ~new_new_n15097__ & ~new_new_n15102__;
  assign new_new_n15104__ = ~new_new_n15101__ & new_new_n15103__;
  assign new_new_n15105__ = ~new_new_n14989__ & ~new_new_n14993__;
  assign new_new_n15106__ = ~new_new_n14990__ & ~new_new_n15105__;
  assign new_new_n15107__ = ~new_new_n14949__ & new_new_n14985__;
  assign new_new_n15108__ = ~new_new_n14950__ & ~new_new_n15107__;
  assign new_new_n15109__ = ~new_new_n14885__ & new_new_n14903__;
  assign new_new_n15110__ = ~new_new_n14884__ & ~new_new_n15109__;
  assign new_new_n15111__ = ~new_new_n15108__ & ~new_new_n15110__;
  assign new_new_n15112__ = new_new_n15108__ & new_new_n15110__;
  assign new_new_n15113__ = ~new_new_n15111__ & ~new_new_n15112__;
  assign new_new_n15114__ = pi38 & pi45;
  assign new_new_n15115__ = pi36 & pi47;
  assign new_new_n15116__ = pi37 & pi46;
  assign new_new_n15117__ = ~new_new_n15115__ & ~new_new_n15116__;
  assign new_new_n15118__ = new_new_n15115__ & new_new_n15116__;
  assign new_new_n15119__ = ~new_new_n15117__ & ~new_new_n15118__;
  assign new_new_n15120__ = new_new_n15114__ & ~new_new_n15119__;
  assign new_new_n15121__ = ~new_new_n15114__ & new_new_n15119__;
  assign new_new_n15122__ = ~new_new_n15120__ & ~new_new_n15121__;
  assign new_new_n15123__ = pi27 & pi56;
  assign new_new_n15124__ = pi20 & pi63;
  assign new_new_n15125__ = pi22 & pi61;
  assign new_new_n15126__ = ~new_new_n15124__ & ~new_new_n15125__;
  assign new_new_n15127__ = new_new_n15124__ & new_new_n15125__;
  assign new_new_n15128__ = ~new_new_n15126__ & ~new_new_n15127__;
  assign new_new_n15129__ = new_new_n15123__ & ~new_new_n15128__;
  assign new_new_n15130__ = ~new_new_n15123__ & new_new_n15128__;
  assign new_new_n15131__ = ~new_new_n15129__ & ~new_new_n15130__;
  assign new_new_n15132__ = new_new_n15122__ & new_new_n15131__;
  assign new_new_n15133__ = ~new_new_n15122__ & ~new_new_n15131__;
  assign new_new_n15134__ = ~new_new_n15132__ & ~new_new_n15133__;
  assign new_new_n15135__ = pi32 & pi51;
  assign new_new_n15136__ = pi26 & pi57;
  assign new_new_n15137__ = pi25 & pi58;
  assign new_new_n15138__ = ~new_new_n15136__ & ~new_new_n15137__;
  assign new_new_n15139__ = new_new_n15136__ & new_new_n15137__;
  assign new_new_n15140__ = ~new_new_n15138__ & ~new_new_n15139__;
  assign new_new_n15141__ = new_new_n15135__ & ~new_new_n15140__;
  assign new_new_n15142__ = ~new_new_n15135__ & new_new_n15140__;
  assign new_new_n15143__ = ~new_new_n15141__ & ~new_new_n15142__;
  assign new_new_n15144__ = new_new_n15134__ & ~new_new_n15143__;
  assign new_new_n15145__ = ~new_new_n15134__ & new_new_n15143__;
  assign new_new_n15146__ = ~new_new_n15144__ & ~new_new_n15145__;
  assign new_new_n15147__ = ~new_new_n14892__ & new_new_n14900__;
  assign new_new_n15148__ = ~new_new_n14891__ & ~new_new_n15147__;
  assign new_new_n15149__ = new_new_n15146__ & new_new_n15148__;
  assign new_new_n15150__ = ~new_new_n15146__ & ~new_new_n15148__;
  assign new_new_n15151__ = ~new_new_n15149__ & ~new_new_n15150__;
  assign new_new_n15152__ = pi40 & pi43;
  assign new_new_n15153__ = pi39 & pi44;
  assign new_new_n15154__ = pi29 & pi54;
  assign new_new_n15155__ = ~new_new_n15153__ & ~new_new_n15154__;
  assign new_new_n15156__ = new_new_n15153__ & new_new_n15154__;
  assign new_new_n15157__ = ~new_new_n15155__ & ~new_new_n15156__;
  assign new_new_n15158__ = new_new_n15152__ & ~new_new_n15157__;
  assign new_new_n15159__ = ~new_new_n15152__ & new_new_n15157__;
  assign new_new_n15160__ = ~new_new_n15158__ & ~new_new_n15159__;
  assign new_new_n15161__ = pi35 & pi48;
  assign new_new_n15162__ = pi33 & pi50;
  assign new_new_n15163__ = pi34 & pi49;
  assign new_new_n15164__ = ~new_new_n15162__ & ~new_new_n15163__;
  assign new_new_n15165__ = new_new_n15162__ & new_new_n15163__;
  assign new_new_n15166__ = ~new_new_n15164__ & ~new_new_n15165__;
  assign new_new_n15167__ = new_new_n15161__ & ~new_new_n15166__;
  assign new_new_n15168__ = ~new_new_n15161__ & new_new_n15166__;
  assign new_new_n15169__ = ~new_new_n15167__ & ~new_new_n15168__;
  assign new_new_n15170__ = new_new_n15160__ & new_new_n15169__;
  assign new_new_n15171__ = ~new_new_n15160__ & ~new_new_n15169__;
  assign new_new_n15172__ = ~new_new_n15170__ & ~new_new_n15171__;
  assign new_new_n15173__ = pi21 & pi62;
  assign new_new_n15174__ = ~pi41 & pi42;
  assign new_new_n15175__ = new_new_n15173__ & ~new_new_n15174__;
  assign new_new_n15176__ = ~new_new_n15173__ & new_new_n15174__;
  assign new_new_n15177__ = ~new_new_n15175__ & ~new_new_n15176__;
  assign new_new_n15178__ = new_new_n15172__ & ~new_new_n15177__;
  assign new_new_n15179__ = ~new_new_n15172__ & new_new_n15177__;
  assign new_new_n15180__ = ~new_new_n15178__ & ~new_new_n15179__;
  assign new_new_n15181__ = new_new_n15151__ & ~new_new_n15180__;
  assign new_new_n15182__ = ~new_new_n15151__ & new_new_n15180__;
  assign new_new_n15183__ = ~new_new_n15181__ & ~new_new_n15182__;
  assign new_new_n15184__ = new_new_n15113__ & ~new_new_n15183__;
  assign new_new_n15185__ = ~new_new_n15113__ & new_new_n15183__;
  assign new_new_n15186__ = ~new_new_n15184__ & ~new_new_n15185__;
  assign new_new_n15187__ = new_new_n15106__ & new_new_n15186__;
  assign new_new_n15188__ = ~new_new_n15106__ & ~new_new_n15186__;
  assign new_new_n15189__ = ~new_new_n15187__ & ~new_new_n15188__;
  assign new_new_n15190__ = new_new_n14955__ & new_new_n14974__;
  assign new_new_n15191__ = ~new_new_n14955__ & ~new_new_n14974__;
  assign new_new_n15192__ = ~new_new_n14953__ & ~new_new_n14976__;
  assign new_new_n15193__ = new_new_n14953__ & new_new_n14976__;
  assign new_new_n15194__ = ~new_new_n15192__ & ~new_new_n15193__;
  assign new_new_n15195__ = ~new_new_n14960__ & ~new_new_n15194__;
  assign new_new_n15196__ = new_new_n14960__ & new_new_n15194__;
  assign new_new_n15197__ = ~new_new_n15195__ & ~new_new_n15196__;
  assign new_new_n15198__ = ~new_new_n15191__ & ~new_new_n15197__;
  assign new_new_n15199__ = ~new_new_n15190__ & ~new_new_n15198__;
  assign new_new_n15200__ = ~new_new_n15071__ & ~new_new_n15075__;
  assign new_new_n15201__ = ~new_new_n15074__ & ~new_new_n15200__;
  assign new_new_n15202__ = ~new_new_n15059__ & ~new_new_n15063__;
  assign new_new_n15203__ = ~new_new_n15062__ & ~new_new_n15202__;
  assign new_new_n15204__ = ~new_new_n15201__ & ~new_new_n15203__;
  assign new_new_n15205__ = new_new_n15201__ & new_new_n15203__;
  assign new_new_n15206__ = ~new_new_n15204__ & ~new_new_n15205__;
  assign new_new_n15207__ = ~new_new_n7761__ & ~new_new_n14896__;
  assign new_new_n15208__ = ~new_new_n14895__ & ~new_new_n15207__;
  assign new_new_n15209__ = ~new_new_n15206__ & new_new_n15208__;
  assign new_new_n15210__ = ~new_new_n15205__ & ~new_new_n15208__;
  assign new_new_n15211__ = ~new_new_n15204__ & new_new_n15210__;
  assign new_new_n15212__ = ~new_new_n15209__ & ~new_new_n15211__;
  assign new_new_n15213__ = ~new_new_n15032__ & ~new_new_n15043__;
  assign new_new_n15214__ = ~new_new_n15033__ & ~new_new_n15213__;
  assign new_new_n15215__ = ~new_new_n15014__ & ~new_new_n15018__;
  assign new_new_n15216__ = ~new_new_n15017__ & ~new_new_n15215__;
  assign new_new_n15217__ = ~new_new_n15023__ & ~new_new_n15027__;
  assign new_new_n15218__ = ~new_new_n15026__ & ~new_new_n15217__;
  assign new_new_n15219__ = ~new_new_n15050__ & ~new_new_n15054__;
  assign new_new_n15220__ = ~new_new_n15053__ & ~new_new_n15219__;
  assign new_new_n15221__ = new_new_n15218__ & new_new_n15220__;
  assign new_new_n15222__ = ~new_new_n15218__ & ~new_new_n15220__;
  assign new_new_n15223__ = ~new_new_n15221__ & ~new_new_n15222__;
  assign new_new_n15224__ = new_new_n15216__ & ~new_new_n15223__;
  assign new_new_n15225__ = ~new_new_n15216__ & new_new_n15223__;
  assign new_new_n15226__ = ~new_new_n15224__ & ~new_new_n15225__;
  assign new_new_n15227__ = new_new_n15214__ & new_new_n15226__;
  assign new_new_n15228__ = ~new_new_n15214__ & ~new_new_n15226__;
  assign new_new_n15229__ = ~new_new_n15227__ & ~new_new_n15228__;
  assign new_new_n15230__ = ~new_new_n15212__ & new_new_n15229__;
  assign new_new_n15231__ = new_new_n15212__ & ~new_new_n15229__;
  assign new_new_n15232__ = ~new_new_n15230__ & ~new_new_n15231__;
  assign new_new_n15233__ = new_new_n15199__ & new_new_n15232__;
  assign new_new_n15234__ = ~new_new_n15199__ & ~new_new_n15232__;
  assign new_new_n15235__ = ~new_new_n15233__ & ~new_new_n15234__;
  assign new_new_n15236__ = ~new_new_n15047__ & ~new_new_n15082__;
  assign new_new_n15237__ = ~new_new_n15048__ & ~new_new_n15236__;
  assign new_new_n15238__ = new_new_n15235__ & ~new_new_n15237__;
  assign new_new_n15239__ = ~new_new_n15235__ & new_new_n15237__;
  assign new_new_n15240__ = ~new_new_n15238__ & ~new_new_n15239__;
  assign new_new_n15241__ = ~new_new_n14933__ & ~new_new_n14937__;
  assign new_new_n15242__ = ~new_new_n15068__ & ~new_new_n15079__;
  assign new_new_n15243__ = ~new_new_n15069__ & ~new_new_n15242__;
  assign new_new_n15244__ = ~new_new_n14970__ & new_new_n15243__;
  assign new_new_n15245__ = new_new_n14970__ & ~new_new_n15243__;
  assign new_new_n15246__ = ~new_new_n15244__ & ~new_new_n15245__;
  assign new_new_n15247__ = ~new_new_n14960__ & ~new_new_n15193__;
  assign new_new_n15248__ = ~new_new_n15192__ & ~new_new_n15247__;
  assign new_new_n15249__ = new_new_n15246__ & ~new_new_n15248__;
  assign new_new_n15250__ = ~new_new_n15246__ & new_new_n15248__;
  assign new_new_n15251__ = ~new_new_n15249__ & ~new_new_n15250__;
  assign new_new_n15252__ = ~new_new_n15241__ & new_new_n15251__;
  assign new_new_n15253__ = new_new_n15241__ & ~new_new_n15251__;
  assign new_new_n15254__ = ~new_new_n15252__ & ~new_new_n15253__;
  assign new_new_n15255__ = ~new_new_n15035__ & ~new_new_n15039__;
  assign new_new_n15256__ = ~new_new_n15038__ & ~new_new_n15255__;
  assign new_new_n15257__ = pi23 & pi60;
  assign new_new_n15258__ = pi24 & pi59;
  assign new_new_n15259__ = ~new_new_n15257__ & ~new_new_n15258__;
  assign new_new_n15260__ = new_new_n15257__ & new_new_n15258__;
  assign new_new_n15261__ = ~new_new_n15259__ & ~new_new_n15260__;
  assign new_new_n15262__ = new_new_n15256__ & ~new_new_n15261__;
  assign new_new_n15263__ = ~new_new_n15256__ & new_new_n15261__;
  assign new_new_n15264__ = ~new_new_n15262__ & ~new_new_n15263__;
  assign new_new_n15265__ = ~pi40 & ~new_new_n14768__;
  assign new_new_n15266__ = pi41 & ~new_new_n15265__;
  assign new_new_n15267__ = new_new_n14917__ & new_new_n15266__;
  assign new_new_n15268__ = ~new_new_n14914__ & ~new_new_n15267__;
  assign new_new_n15269__ = ~new_new_n15264__ & ~new_new_n15268__;
  assign new_new_n15270__ = new_new_n15264__ & new_new_n15268__;
  assign new_new_n15271__ = ~new_new_n15269__ & ~new_new_n15270__;
  assign new_new_n15272__ = pi31 & pi52;
  assign new_new_n15273__ = pi28 & pi55;
  assign new_new_n15274__ = pi30 & pi53;
  assign new_new_n15275__ = ~new_new_n15273__ & ~new_new_n15274__;
  assign new_new_n15276__ = new_new_n15273__ & new_new_n15274__;
  assign new_new_n15277__ = ~new_new_n15275__ & ~new_new_n15276__;
  assign new_new_n15278__ = new_new_n15272__ & ~new_new_n15277__;
  assign new_new_n15279__ = ~new_new_n15272__ & new_new_n15277__;
  assign new_new_n15280__ = ~new_new_n15278__ & ~new_new_n15279__;
  assign new_new_n15281__ = ~new_new_n15271__ & new_new_n15280__;
  assign new_new_n15282__ = new_new_n15271__ & ~new_new_n15280__;
  assign new_new_n15283__ = ~new_new_n15281__ & ~new_new_n15282__;
  assign new_new_n15284__ = new_new_n15254__ & new_new_n15283__;
  assign new_new_n15285__ = ~new_new_n15254__ & ~new_new_n15283__;
  assign new_new_n15286__ = ~new_new_n15284__ & ~new_new_n15285__;
  assign new_new_n15287__ = ~new_new_n15240__ & new_new_n15286__;
  assign new_new_n15288__ = new_new_n15240__ & ~new_new_n15286__;
  assign new_new_n15289__ = ~new_new_n15287__ & ~new_new_n15288__;
  assign new_new_n15290__ = ~new_new_n15009__ & ~new_new_n15085__;
  assign new_new_n15291__ = ~new_new_n15010__ & ~new_new_n15290__;
  assign new_new_n15292__ = new_new_n15289__ & ~new_new_n15291__;
  assign new_new_n15293__ = ~new_new_n15289__ & new_new_n15291__;
  assign new_new_n15294__ = ~new_new_n15292__ & ~new_new_n15293__;
  assign new_new_n15295__ = new_new_n15189__ & new_new_n15294__;
  assign new_new_n15296__ = ~new_new_n15189__ & ~new_new_n15294__;
  assign new_new_n15297__ = ~new_new_n15295__ & ~new_new_n15296__;
  assign new_new_n15298__ = ~new_new_n15104__ & new_new_n15297__;
  assign new_new_n15299__ = new_new_n14872__ & ~new_new_n14996__;
  assign new_new_n15300__ = new_new_n14879__ & new_new_n15299__;
  assign new_new_n15301__ = ~new_new_n14872__ & new_new_n14996__;
  assign new_new_n15302__ = ~new_new_n14873__ & new_new_n14879__;
  assign new_new_n15303__ = ~new_new_n15301__ & new_new_n15302__;
  assign new_new_n15304__ = ~new_new_n15299__ & ~new_new_n15303__;
  assign new_new_n15305__ = ~new_new_n15088__ & ~new_new_n15304__;
  assign new_new_n15306__ = new_new_n14873__ & new_new_n14998__;
  assign new_new_n15307__ = new_new_n14873__ & ~new_new_n14997__;
  assign new_new_n15308__ = ~new_new_n14879__ & new_new_n15301__;
  assign new_new_n15309__ = ~new_new_n15307__ & ~new_new_n15308__;
  assign new_new_n15310__ = new_new_n15088__ & ~new_new_n15309__;
  assign new_new_n15311__ = ~new_new_n15300__ & ~new_new_n15306__;
  assign new_new_n15312__ = ~new_new_n15305__ & new_new_n15311__;
  assign new_new_n15313__ = ~new_new_n15310__ & new_new_n15312__;
  assign new_new_n15314__ = ~new_new_n15297__ & ~new_new_n15313__;
  assign po084 = new_new_n15298__ | new_new_n15314__;
  assign new_new_n15316__ = ~new_new_n14873__ & ~new_new_n15297__;
  assign new_new_n15317__ = new_new_n15096__ & ~new_new_n15316__;
  assign new_new_n15318__ = ~new_new_n15099__ & new_new_n15297__;
  assign new_new_n15319__ = ~new_new_n15098__ & ~new_new_n15318__;
  assign new_new_n15320__ = ~new_new_n14872__ & ~new_new_n15319__;
  assign new_new_n15321__ = new_new_n14873__ & new_new_n15297__;
  assign new_new_n15322__ = ~new_new_n15320__ & ~new_new_n15321__;
  assign new_new_n15323__ = ~new_new_n15317__ & new_new_n15322__;
  assign new_new_n15324__ = ~new_new_n15288__ & new_new_n15291__;
  assign new_new_n15325__ = ~new_new_n15287__ & ~new_new_n15324__;
  assign new_new_n15326__ = ~new_new_n15253__ & ~new_new_n15283__;
  assign new_new_n15327__ = ~new_new_n15252__ & ~new_new_n15326__;
  assign new_new_n15328__ = ~new_new_n15245__ & ~new_new_n15248__;
  assign new_new_n15329__ = ~new_new_n15244__ & ~new_new_n15328__;
  assign new_new_n15330__ = ~new_new_n15269__ & new_new_n15280__;
  assign new_new_n15331__ = ~new_new_n15270__ & ~new_new_n15330__;
  assign new_new_n15332__ = new_new_n15329__ & new_new_n15331__;
  assign new_new_n15333__ = ~new_new_n15329__ & ~new_new_n15331__;
  assign new_new_n15334__ = ~new_new_n15332__ & ~new_new_n15333__;
  assign new_new_n15335__ = ~new_new_n15256__ & ~new_new_n15260__;
  assign new_new_n15336__ = ~new_new_n15259__ & ~new_new_n15335__;
  assign new_new_n15337__ = pi32 & pi52;
  assign new_new_n15338__ = pi26 & pi58;
  assign new_new_n15339__ = pi31 & pi53;
  assign new_new_n15340__ = ~new_new_n15338__ & ~new_new_n15339__;
  assign new_new_n15341__ = new_new_n15338__ & new_new_n15339__;
  assign new_new_n15342__ = ~new_new_n15340__ & ~new_new_n15341__;
  assign new_new_n15343__ = new_new_n15337__ & ~new_new_n15342__;
  assign new_new_n15344__ = ~new_new_n15337__ & new_new_n15342__;
  assign new_new_n15345__ = ~new_new_n15343__ & ~new_new_n15344__;
  assign new_new_n15346__ = ~new_new_n15336__ & new_new_n15345__;
  assign new_new_n15347__ = new_new_n15336__ & ~new_new_n15345__;
  assign new_new_n15348__ = ~new_new_n15346__ & ~new_new_n15347__;
  assign new_new_n15349__ = ~new_new_n15123__ & ~new_new_n15127__;
  assign new_new_n15350__ = ~new_new_n15126__ & ~new_new_n15349__;
  assign new_new_n15351__ = new_new_n15348__ & new_new_n15350__;
  assign new_new_n15352__ = ~new_new_n15348__ & ~new_new_n15350__;
  assign new_new_n15353__ = ~new_new_n15351__ & ~new_new_n15352__;
  assign new_new_n15354__ = new_new_n15334__ & ~new_new_n15353__;
  assign new_new_n15355__ = ~new_new_n15334__ & new_new_n15353__;
  assign new_new_n15356__ = ~new_new_n15354__ & ~new_new_n15355__;
  assign new_new_n15357__ = new_new_n15327__ & ~new_new_n15356__;
  assign new_new_n15358__ = ~new_new_n15327__ & new_new_n15356__;
  assign new_new_n15359__ = ~new_new_n15357__ & ~new_new_n15358__;
  assign new_new_n15360__ = pi36 & pi48;
  assign new_new_n15361__ = pi34 & pi50;
  assign new_new_n15362__ = pi35 & pi49;
  assign new_new_n15363__ = ~new_new_n15361__ & ~new_new_n15362__;
  assign new_new_n15364__ = new_new_n15361__ & new_new_n15362__;
  assign new_new_n15365__ = ~new_new_n15363__ & ~new_new_n15364__;
  assign new_new_n15366__ = new_new_n15360__ & ~new_new_n15365__;
  assign new_new_n15367__ = ~new_new_n15360__ & new_new_n15365__;
  assign new_new_n15368__ = ~new_new_n15366__ & ~new_new_n15367__;
  assign new_new_n15369__ = pi33 & pi51;
  assign new_new_n15370__ = pi24 & pi60;
  assign new_new_n15371__ = pi25 & pi59;
  assign new_new_n15372__ = ~new_new_n15370__ & ~new_new_n15371__;
  assign new_new_n15373__ = new_new_n15370__ & new_new_n15371__;
  assign new_new_n15374__ = ~new_new_n15372__ & ~new_new_n15373__;
  assign new_new_n15375__ = new_new_n15369__ & ~new_new_n15374__;
  assign new_new_n15376__ = ~new_new_n15369__ & new_new_n15374__;
  assign new_new_n15377__ = ~new_new_n15375__ & ~new_new_n15376__;
  assign new_new_n15378__ = new_new_n15368__ & new_new_n15377__;
  assign new_new_n15379__ = ~new_new_n15368__ & ~new_new_n15377__;
  assign new_new_n15380__ = ~new_new_n15378__ & ~new_new_n15379__;
  assign new_new_n15381__ = pi23 & pi61;
  assign new_new_n15382__ = pi22 & pi62;
  assign new_new_n15383__ = pi21 & pi63;
  assign new_new_n15384__ = ~new_new_n15382__ & ~new_new_n15383__;
  assign new_new_n15385__ = new_new_n15382__ & new_new_n15383__;
  assign new_new_n15386__ = ~new_new_n15384__ & ~new_new_n15385__;
  assign new_new_n15387__ = new_new_n15381__ & ~new_new_n15386__;
  assign new_new_n15388__ = ~new_new_n15381__ & new_new_n15386__;
  assign new_new_n15389__ = ~new_new_n15387__ & ~new_new_n15388__;
  assign new_new_n15390__ = new_new_n15380__ & ~new_new_n15389__;
  assign new_new_n15391__ = ~new_new_n15380__ & new_new_n15389__;
  assign new_new_n15392__ = ~new_new_n15390__ & ~new_new_n15391__;
  assign new_new_n15393__ = ~new_new_n15161__ & ~new_new_n15165__;
  assign new_new_n15394__ = ~new_new_n15164__ & ~new_new_n15393__;
  assign new_new_n15395__ = ~new_new_n15114__ & ~new_new_n15118__;
  assign new_new_n15396__ = ~new_new_n15117__ & ~new_new_n15395__;
  assign new_new_n15397__ = ~new_new_n15394__ & ~new_new_n15396__;
  assign new_new_n15398__ = new_new_n15394__ & new_new_n15396__;
  assign new_new_n15399__ = ~new_new_n15397__ & ~new_new_n15398__;
  assign new_new_n15400__ = ~new_new_n15135__ & ~new_new_n15139__;
  assign new_new_n15401__ = ~new_new_n15138__ & ~new_new_n15400__;
  assign new_new_n15402__ = ~new_new_n15399__ & new_new_n15401__;
  assign new_new_n15403__ = ~new_new_n15398__ & ~new_new_n15401__;
  assign new_new_n15404__ = ~new_new_n15397__ & new_new_n15403__;
  assign new_new_n15405__ = ~new_new_n15402__ & ~new_new_n15404__;
  assign new_new_n15406__ = ~new_new_n15216__ & ~new_new_n15221__;
  assign new_new_n15407__ = ~new_new_n15222__ & ~new_new_n15406__;
  assign new_new_n15408__ = ~new_new_n15204__ & ~new_new_n15210__;
  assign new_new_n15409__ = new_new_n15407__ & ~new_new_n15408__;
  assign new_new_n15410__ = ~new_new_n15407__ & new_new_n15408__;
  assign new_new_n15411__ = ~new_new_n15409__ & ~new_new_n15410__;
  assign new_new_n15412__ = new_new_n15405__ & new_new_n15411__;
  assign new_new_n15413__ = ~new_new_n15405__ & ~new_new_n15411__;
  assign new_new_n15414__ = ~new_new_n15412__ & ~new_new_n15413__;
  assign new_new_n15415__ = new_new_n15392__ & new_new_n15414__;
  assign new_new_n15416__ = ~new_new_n15392__ & ~new_new_n15414__;
  assign new_new_n15417__ = ~new_new_n15415__ & ~new_new_n15416__;
  assign new_new_n15418__ = pi41 & pi43;
  assign new_new_n15419__ = pi40 & pi44;
  assign new_new_n15420__ = pi39 & pi45;
  assign new_new_n15421__ = ~new_new_n15419__ & ~new_new_n15420__;
  assign new_new_n15422__ = new_new_n15419__ & new_new_n15420__;
  assign new_new_n15423__ = ~new_new_n15421__ & ~new_new_n15422__;
  assign new_new_n15424__ = new_new_n15418__ & ~new_new_n15423__;
  assign new_new_n15425__ = ~new_new_n15418__ & new_new_n15423__;
  assign new_new_n15426__ = ~new_new_n15424__ & ~new_new_n15425__;
  assign new_new_n15427__ = pi38 & pi46;
  assign new_new_n15428__ = pi29 & pi55;
  assign new_new_n15429__ = pi28 & pi56;
  assign new_new_n15430__ = ~new_new_n15428__ & ~new_new_n15429__;
  assign new_new_n15431__ = new_new_n15428__ & new_new_n15429__;
  assign new_new_n15432__ = ~new_new_n15430__ & ~new_new_n15431__;
  assign new_new_n15433__ = new_new_n15427__ & ~new_new_n15432__;
  assign new_new_n15434__ = ~new_new_n15427__ & new_new_n15432__;
  assign new_new_n15435__ = ~new_new_n15433__ & ~new_new_n15434__;
  assign new_new_n15436__ = new_new_n15426__ & new_new_n15435__;
  assign new_new_n15437__ = ~new_new_n15426__ & ~new_new_n15435__;
  assign new_new_n15438__ = ~new_new_n15436__ & ~new_new_n15437__;
  assign new_new_n15439__ = pi37 & pi47;
  assign new_new_n15440__ = pi27 & pi57;
  assign new_new_n15441__ = pi30 & pi54;
  assign new_new_n15442__ = ~new_new_n15440__ & ~new_new_n15441__;
  assign new_new_n15443__ = new_new_n15440__ & new_new_n15441__;
  assign new_new_n15444__ = ~new_new_n15442__ & ~new_new_n15443__;
  assign new_new_n15445__ = new_new_n15439__ & ~new_new_n15444__;
  assign new_new_n15446__ = ~new_new_n15439__ & new_new_n15444__;
  assign new_new_n15447__ = ~new_new_n15445__ & ~new_new_n15446__;
  assign new_new_n15448__ = new_new_n15438__ & ~new_new_n15447__;
  assign new_new_n15449__ = ~new_new_n15438__ & new_new_n15447__;
  assign new_new_n15450__ = ~new_new_n15448__ & ~new_new_n15449__;
  assign new_new_n15451__ = new_new_n15417__ & ~new_new_n15450__;
  assign new_new_n15452__ = ~new_new_n15417__ & new_new_n15450__;
  assign new_new_n15453__ = ~new_new_n15451__ & ~new_new_n15452__;
  assign new_new_n15454__ = new_new_n15359__ & ~new_new_n15453__;
  assign new_new_n15455__ = ~new_new_n15359__ & new_new_n15453__;
  assign new_new_n15456__ = ~new_new_n15454__ & ~new_new_n15455__;
  assign new_new_n15457__ = ~new_new_n15325__ & new_new_n15456__;
  assign new_new_n15458__ = new_new_n15325__ & ~new_new_n15456__;
  assign new_new_n15459__ = ~new_new_n15457__ & ~new_new_n15458__;
  assign new_new_n15460__ = ~new_new_n15233__ & ~new_new_n15237__;
  assign new_new_n15461__ = ~new_new_n15234__ & ~new_new_n15460__;
  assign new_new_n15462__ = ~new_new_n15112__ & new_new_n15183__;
  assign new_new_n15463__ = ~new_new_n15111__ & ~new_new_n15462__;
  assign new_new_n15464__ = ~new_new_n15461__ & ~new_new_n15463__;
  assign new_new_n15465__ = new_new_n15461__ & new_new_n15463__;
  assign new_new_n15466__ = ~new_new_n15464__ & ~new_new_n15465__;
  assign new_new_n15467__ = ~new_new_n15132__ & ~new_new_n15143__;
  assign new_new_n15468__ = ~new_new_n15133__ & ~new_new_n15467__;
  assign new_new_n15469__ = ~pi41 & ~new_new_n15173__;
  assign new_new_n15470__ = pi42 & ~new_new_n15469__;
  assign new_new_n15471__ = ~new_new_n15152__ & ~new_new_n15156__;
  assign new_new_n15472__ = ~new_new_n15155__ & ~new_new_n15471__;
  assign new_new_n15473__ = ~new_new_n15272__ & ~new_new_n15276__;
  assign new_new_n15474__ = ~new_new_n15275__ & ~new_new_n15473__;
  assign new_new_n15475__ = new_new_n15472__ & new_new_n15474__;
  assign new_new_n15476__ = ~new_new_n15472__ & ~new_new_n15474__;
  assign new_new_n15477__ = ~new_new_n15475__ & ~new_new_n15476__;
  assign new_new_n15478__ = new_new_n15470__ & ~new_new_n15477__;
  assign new_new_n15479__ = ~new_new_n15470__ & new_new_n15477__;
  assign new_new_n15480__ = ~new_new_n15478__ & ~new_new_n15479__;
  assign new_new_n15481__ = new_new_n15468__ & new_new_n15480__;
  assign new_new_n15482__ = ~new_new_n15468__ & ~new_new_n15480__;
  assign new_new_n15483__ = ~new_new_n15481__ & ~new_new_n15482__;
  assign new_new_n15484__ = ~new_new_n15170__ & ~new_new_n15177__;
  assign new_new_n15485__ = ~new_new_n15171__ & ~new_new_n15484__;
  assign new_new_n15486__ = ~new_new_n15150__ & new_new_n15180__;
  assign new_new_n15487__ = ~new_new_n15149__ & ~new_new_n15486__;
  assign new_new_n15488__ = ~new_new_n15485__ & new_new_n15487__;
  assign new_new_n15489__ = new_new_n15485__ & ~new_new_n15487__;
  assign new_new_n15490__ = ~new_new_n15488__ & ~new_new_n15489__;
  assign new_new_n15491__ = ~new_new_n15212__ & ~new_new_n15227__;
  assign new_new_n15492__ = ~new_new_n15228__ & ~new_new_n15491__;
  assign new_new_n15493__ = new_new_n15490__ & ~new_new_n15492__;
  assign new_new_n15494__ = ~new_new_n15490__ & new_new_n15492__;
  assign new_new_n15495__ = ~new_new_n15493__ & ~new_new_n15494__;
  assign new_new_n15496__ = new_new_n15483__ & new_new_n15495__;
  assign new_new_n15497__ = ~new_new_n15483__ & ~new_new_n15495__;
  assign new_new_n15498__ = ~new_new_n15496__ & ~new_new_n15497__;
  assign new_new_n15499__ = new_new_n15466__ & ~new_new_n15498__;
  assign new_new_n15500__ = ~new_new_n15466__ & new_new_n15498__;
  assign new_new_n15501__ = ~new_new_n15499__ & ~new_new_n15500__;
  assign new_new_n15502__ = new_new_n15459__ & new_new_n15501__;
  assign new_new_n15503__ = ~new_new_n15459__ & ~new_new_n15501__;
  assign new_new_n15504__ = ~new_new_n15502__ & ~new_new_n15503__;
  assign new_new_n15505__ = ~new_new_n15323__ & ~new_new_n15504__;
  assign new_new_n15506__ = new_new_n15323__ & new_new_n15504__;
  assign new_new_n15507__ = ~new_new_n15505__ & ~new_new_n15506__;
  assign new_new_n15508__ = ~new_new_n15188__ & ~new_new_n15294__;
  assign new_new_n15509__ = ~new_new_n15187__ & ~new_new_n15508__;
  assign new_new_n15510__ = ~new_new_n15507__ & new_new_n15509__;
  assign new_new_n15511__ = ~new_new_n15505__ & ~new_new_n15509__;
  assign new_new_n15512__ = ~new_new_n15506__ & new_new_n15511__;
  assign po085 = ~new_new_n15510__ & ~new_new_n15512__;
  assign new_new_n15514__ = ~new_new_n15506__ & ~new_new_n15511__;
  assign new_new_n15515__ = ~new_new_n15457__ & ~new_new_n15501__;
  assign new_new_n15516__ = ~new_new_n15458__ & ~new_new_n15515__;
  assign new_new_n15517__ = ~new_new_n15514__ & new_new_n15516__;
  assign new_new_n15518__ = new_new_n15514__ & ~new_new_n15516__;
  assign new_new_n15519__ = ~new_new_n15517__ & ~new_new_n15518__;
  assign new_new_n15520__ = ~new_new_n15357__ & new_new_n15453__;
  assign new_new_n15521__ = ~new_new_n15358__ & ~new_new_n15520__;
  assign new_new_n15522__ = new_new_n15483__ & new_new_n15485__;
  assign new_new_n15523__ = ~new_new_n15483__ & ~new_new_n15485__;
  assign new_new_n15524__ = ~new_new_n15522__ & ~new_new_n15523__;
  assign new_new_n15525__ = new_new_n15492__ & new_new_n15524__;
  assign new_new_n15526__ = ~new_new_n15487__ & ~new_new_n15525__;
  assign new_new_n15527__ = ~new_new_n15492__ & ~new_new_n15524__;
  assign new_new_n15528__ = ~new_new_n15526__ & ~new_new_n15527__;
  assign new_new_n15529__ = new_new_n15521__ & ~new_new_n15528__;
  assign new_new_n15530__ = ~new_new_n15521__ & new_new_n15528__;
  assign new_new_n15531__ = ~new_new_n15529__ & ~new_new_n15530__;
  assign new_new_n15532__ = ~new_new_n15332__ & ~new_new_n15353__;
  assign new_new_n15533__ = ~new_new_n15333__ & ~new_new_n15532__;
  assign new_new_n15534__ = ~new_new_n15397__ & ~new_new_n15403__;
  assign new_new_n15535__ = ~new_new_n15470__ & ~new_new_n15475__;
  assign new_new_n15536__ = ~new_new_n15476__ & ~new_new_n15535__;
  assign new_new_n15537__ = ~new_new_n15534__ & ~new_new_n15536__;
  assign new_new_n15538__ = new_new_n15534__ & new_new_n15536__;
  assign new_new_n15539__ = ~new_new_n15537__ & ~new_new_n15538__;
  assign new_new_n15540__ = ~new_new_n15346__ & new_new_n15350__;
  assign new_new_n15541__ = ~new_new_n15347__ & ~new_new_n15540__;
  assign new_new_n15542__ = new_new_n15539__ & ~new_new_n15541__;
  assign new_new_n15543__ = ~new_new_n15539__ & new_new_n15541__;
  assign new_new_n15544__ = ~new_new_n15542__ & ~new_new_n15543__;
  assign new_new_n15545__ = new_new_n15533__ & new_new_n15544__;
  assign new_new_n15546__ = ~new_new_n15533__ & ~new_new_n15544__;
  assign new_new_n15547__ = ~new_new_n15545__ & ~new_new_n15546__;
  assign new_new_n15548__ = ~new_new_n15416__ & new_new_n15450__;
  assign new_new_n15549__ = ~new_new_n15415__ & ~new_new_n15548__;
  assign new_new_n15550__ = new_new_n15547__ & ~new_new_n15549__;
  assign new_new_n15551__ = ~new_new_n15547__ & new_new_n15549__;
  assign new_new_n15552__ = ~new_new_n15550__ & ~new_new_n15551__;
  assign new_new_n15553__ = new_new_n15531__ & ~new_new_n15552__;
  assign new_new_n15554__ = ~new_new_n15531__ & new_new_n15552__;
  assign new_new_n15555__ = ~new_new_n15553__ & ~new_new_n15554__;
  assign new_new_n15556__ = ~new_new_n15378__ & ~new_new_n15389__;
  assign new_new_n15557__ = ~new_new_n15379__ & ~new_new_n15556__;
  assign new_new_n15558__ = ~new_new_n15436__ & ~new_new_n15447__;
  assign new_new_n15559__ = ~new_new_n15437__ & ~new_new_n15558__;
  assign new_new_n15560__ = ~new_new_n15557__ & ~new_new_n15559__;
  assign new_new_n15561__ = new_new_n15557__ & new_new_n15559__;
  assign new_new_n15562__ = ~new_new_n15560__ & ~new_new_n15561__;
  assign new_new_n15563__ = ~new_new_n15381__ & ~new_new_n15385__;
  assign new_new_n15564__ = ~new_new_n15384__ & ~new_new_n15563__;
  assign new_new_n15565__ = ~new_new_n15369__ & ~new_new_n15373__;
  assign new_new_n15566__ = ~new_new_n15372__ & ~new_new_n15565__;
  assign new_new_n15567__ = ~new_new_n15360__ & ~new_new_n15364__;
  assign new_new_n15568__ = ~new_new_n15363__ & ~new_new_n15567__;
  assign new_new_n15569__ = ~new_new_n15566__ & ~new_new_n15568__;
  assign new_new_n15570__ = new_new_n15566__ & new_new_n15568__;
  assign new_new_n15571__ = ~new_new_n15569__ & ~new_new_n15570__;
  assign new_new_n15572__ = new_new_n15564__ & ~new_new_n15571__;
  assign new_new_n15573__ = ~new_new_n15564__ & new_new_n15571__;
  assign new_new_n15574__ = ~new_new_n15572__ & ~new_new_n15573__;
  assign new_new_n15575__ = new_new_n15562__ & new_new_n15574__;
  assign new_new_n15576__ = ~new_new_n15562__ & ~new_new_n15574__;
  assign new_new_n15577__ = ~new_new_n15575__ & ~new_new_n15576__;
  assign new_new_n15578__ = ~new_new_n15481__ & ~new_new_n15522__;
  assign new_new_n15579__ = pi23 & pi62;
  assign new_new_n15580__ = ~pi42 & pi43;
  assign new_new_n15581__ = ~new_new_n15579__ & new_new_n15580__;
  assign new_new_n15582__ = new_new_n15579__ & ~new_new_n15580__;
  assign new_new_n15583__ = ~new_new_n15581__ & ~new_new_n15582__;
  assign new_new_n15584__ = pi31 & pi54;
  assign new_new_n15585__ = pi30 & pi55;
  assign new_new_n15586__ = ~new_new_n8458__ & ~new_new_n15585__;
  assign new_new_n15587__ = new_new_n8458__ & new_new_n15585__;
  assign new_new_n15588__ = ~new_new_n15586__ & ~new_new_n15587__;
  assign new_new_n15589__ = new_new_n15584__ & ~new_new_n15588__;
  assign new_new_n15590__ = ~new_new_n15584__ & new_new_n15588__;
  assign new_new_n15591__ = ~new_new_n15589__ & ~new_new_n15590__;
  assign new_new_n15592__ = pi38 & pi47;
  assign new_new_n15593__ = pi36 & pi49;
  assign new_new_n15594__ = pi37 & pi48;
  assign new_new_n15595__ = ~new_new_n15593__ & ~new_new_n15594__;
  assign new_new_n15596__ = new_new_n15593__ & new_new_n15594__;
  assign new_new_n15597__ = ~new_new_n15595__ & ~new_new_n15596__;
  assign new_new_n15598__ = new_new_n15592__ & ~new_new_n15597__;
  assign new_new_n15599__ = ~new_new_n15592__ & new_new_n15597__;
  assign new_new_n15600__ = ~new_new_n15598__ & ~new_new_n15599__;
  assign new_new_n15601__ = new_new_n15591__ & new_new_n15600__;
  assign new_new_n15602__ = ~new_new_n15591__ & ~new_new_n15600__;
  assign new_new_n15603__ = ~new_new_n15601__ & ~new_new_n15602__;
  assign new_new_n15604__ = new_new_n15583__ & ~new_new_n15603__;
  assign new_new_n15605__ = ~new_new_n15583__ & new_new_n15603__;
  assign new_new_n15606__ = ~new_new_n15604__ & ~new_new_n15605__;
  assign new_new_n15607__ = ~new_new_n15578__ & ~new_new_n15606__;
  assign new_new_n15608__ = new_new_n15578__ & new_new_n15606__;
  assign new_new_n15609__ = ~new_new_n15607__ & ~new_new_n15608__;
  assign new_new_n15610__ = pi34 & pi51;
  assign new_new_n15611__ = pi33 & pi52;
  assign new_new_n15612__ = pi32 & pi53;
  assign new_new_n15613__ = ~new_new_n15611__ & ~new_new_n15612__;
  assign new_new_n15614__ = new_new_n15611__ & new_new_n15612__;
  assign new_new_n15615__ = ~new_new_n15613__ & ~new_new_n15614__;
  assign new_new_n15616__ = new_new_n15610__ & ~new_new_n15615__;
  assign new_new_n15617__ = ~new_new_n15610__ & new_new_n15615__;
  assign new_new_n15618__ = ~new_new_n15616__ & ~new_new_n15617__;
  assign new_new_n15619__ = pi41 & pi44;
  assign new_new_n15620__ = pi40 & pi45;
  assign new_new_n15621__ = pi39 & pi46;
  assign new_new_n15622__ = ~new_new_n15620__ & ~new_new_n15621__;
  assign new_new_n15623__ = new_new_n15620__ & new_new_n15621__;
  assign new_new_n15624__ = ~new_new_n15622__ & ~new_new_n15623__;
  assign new_new_n15625__ = new_new_n15619__ & ~new_new_n15624__;
  assign new_new_n15626__ = ~new_new_n15619__ & new_new_n15624__;
  assign new_new_n15627__ = ~new_new_n15625__ & ~new_new_n15626__;
  assign new_new_n15628__ = new_new_n15618__ & new_new_n15627__;
  assign new_new_n15629__ = ~new_new_n15618__ & ~new_new_n15627__;
  assign new_new_n15630__ = ~new_new_n15628__ & ~new_new_n15629__;
  assign new_new_n15631__ = pi35 & pi50;
  assign new_new_n15632__ = pi22 & pi63;
  assign new_new_n15633__ = pi28 & pi57;
  assign new_new_n15634__ = ~new_new_n15632__ & ~new_new_n15633__;
  assign new_new_n15635__ = new_new_n15632__ & new_new_n15633__;
  assign new_new_n15636__ = ~new_new_n15634__ & ~new_new_n15635__;
  assign new_new_n15637__ = new_new_n15631__ & ~new_new_n15636__;
  assign new_new_n15638__ = ~new_new_n15631__ & new_new_n15636__;
  assign new_new_n15639__ = ~new_new_n15637__ & ~new_new_n15638__;
  assign new_new_n15640__ = ~new_new_n15630__ & new_new_n15639__;
  assign new_new_n15641__ = new_new_n15630__ & ~new_new_n15639__;
  assign new_new_n15642__ = ~new_new_n15640__ & ~new_new_n15641__;
  assign new_new_n15643__ = new_new_n15609__ & new_new_n15642__;
  assign new_new_n15644__ = ~new_new_n15609__ & ~new_new_n15642__;
  assign new_new_n15645__ = ~new_new_n15643__ & ~new_new_n15644__;
  assign new_new_n15646__ = ~new_new_n15577__ & new_new_n15645__;
  assign new_new_n15647__ = new_new_n15577__ & ~new_new_n15645__;
  assign new_new_n15648__ = ~new_new_n15646__ & ~new_new_n15647__;
  assign new_new_n15649__ = ~new_new_n15337__ & ~new_new_n15341__;
  assign new_new_n15650__ = ~new_new_n15340__ & ~new_new_n15649__;
  assign new_new_n15651__ = pi27 & pi58;
  assign new_new_n15652__ = pi26 & pi59;
  assign new_new_n15653__ = pi25 & pi60;
  assign new_new_n15654__ = ~new_new_n15652__ & ~new_new_n15653__;
  assign new_new_n15655__ = new_new_n15652__ & new_new_n15653__;
  assign new_new_n15656__ = ~new_new_n15654__ & ~new_new_n15655__;
  assign new_new_n15657__ = new_new_n15651__ & ~new_new_n15656__;
  assign new_new_n15658__ = ~new_new_n15651__ & new_new_n15656__;
  assign new_new_n15659__ = ~new_new_n15657__ & ~new_new_n15658__;
  assign new_new_n15660__ = ~new_new_n15650__ & new_new_n15659__;
  assign new_new_n15661__ = new_new_n15650__ & ~new_new_n15659__;
  assign new_new_n15662__ = ~new_new_n15660__ & ~new_new_n15661__;
  assign new_new_n15663__ = ~new_new_n15439__ & ~new_new_n15443__;
  assign new_new_n15664__ = ~new_new_n15442__ & ~new_new_n15663__;
  assign new_new_n15665__ = new_new_n15662__ & ~new_new_n15664__;
  assign new_new_n15666__ = ~new_new_n15662__ & new_new_n15664__;
  assign new_new_n15667__ = ~new_new_n15665__ & ~new_new_n15666__;
  assign new_new_n15668__ = new_new_n15405__ & ~new_new_n15407__;
  assign new_new_n15669__ = new_new_n15408__ & ~new_new_n15668__;
  assign new_new_n15670__ = ~new_new_n15405__ & new_new_n15407__;
  assign new_new_n15671__ = ~new_new_n15669__ & ~new_new_n15670__;
  assign new_new_n15672__ = ~new_new_n15667__ & ~new_new_n15671__;
  assign new_new_n15673__ = new_new_n15667__ & new_new_n15671__;
  assign new_new_n15674__ = ~new_new_n15672__ & ~new_new_n15673__;
  assign new_new_n15675__ = ~new_new_n15427__ & ~new_new_n15431__;
  assign new_new_n15676__ = ~new_new_n15430__ & ~new_new_n15675__;
  assign new_new_n15677__ = ~new_new_n15418__ & ~new_new_n15422__;
  assign new_new_n15678__ = ~new_new_n15421__ & ~new_new_n15677__;
  assign new_new_n15679__ = pi24 & pi61;
  assign new_new_n15680__ = new_new_n15678__ & ~new_new_n15679__;
  assign new_new_n15681__ = ~new_new_n15678__ & new_new_n15679__;
  assign new_new_n15682__ = ~new_new_n15680__ & ~new_new_n15681__;
  assign new_new_n15683__ = new_new_n15676__ & new_new_n15682__;
  assign new_new_n15684__ = ~new_new_n15676__ & ~new_new_n15682__;
  assign new_new_n15685__ = ~new_new_n15683__ & ~new_new_n15684__;
  assign new_new_n15686__ = new_new_n15674__ & new_new_n15685__;
  assign new_new_n15687__ = ~new_new_n15674__ & ~new_new_n15685__;
  assign new_new_n15688__ = ~new_new_n15686__ & ~new_new_n15687__;
  assign new_new_n15689__ = new_new_n15648__ & ~new_new_n15688__;
  assign new_new_n15690__ = ~new_new_n15648__ & new_new_n15688__;
  assign new_new_n15691__ = ~new_new_n15689__ & ~new_new_n15690__;
  assign new_new_n15692__ = ~new_new_n15555__ & new_new_n15691__;
  assign new_new_n15693__ = new_new_n15555__ & ~new_new_n15691__;
  assign new_new_n15694__ = ~new_new_n15692__ & ~new_new_n15693__;
  assign new_new_n15695__ = ~new_new_n15465__ & new_new_n15498__;
  assign new_new_n15696__ = ~new_new_n15464__ & ~new_new_n15695__;
  assign new_new_n15697__ = new_new_n15694__ & ~new_new_n15696__;
  assign new_new_n15698__ = ~new_new_n15694__ & new_new_n15696__;
  assign new_new_n15699__ = ~new_new_n15697__ & ~new_new_n15698__;
  assign new_new_n15700__ = new_new_n15519__ & new_new_n15699__;
  assign new_new_n15701__ = ~new_new_n15519__ & ~new_new_n15699__;
  assign po086 = new_new_n15700__ | new_new_n15701__;
  assign new_new_n15703__ = ~new_new_n15628__ & ~new_new_n15639__;
  assign new_new_n15704__ = ~new_new_n15629__ & ~new_new_n15703__;
  assign new_new_n15705__ = ~new_new_n15583__ & ~new_new_n15601__;
  assign new_new_n15706__ = ~new_new_n15602__ & ~new_new_n15705__;
  assign new_new_n15707__ = ~new_new_n15660__ & new_new_n15664__;
  assign new_new_n15708__ = ~new_new_n15661__ & ~new_new_n15707__;
  assign new_new_n15709__ = new_new_n15706__ & new_new_n15708__;
  assign new_new_n15710__ = ~new_new_n15706__ & ~new_new_n15708__;
  assign new_new_n15711__ = ~new_new_n15709__ & ~new_new_n15710__;
  assign new_new_n15712__ = new_new_n15704__ & ~new_new_n15711__;
  assign new_new_n15713__ = ~new_new_n15704__ & new_new_n15711__;
  assign new_new_n15714__ = ~new_new_n15712__ & ~new_new_n15713__;
  assign new_new_n15715__ = new_new_n15518__ & new_new_n15693__;
  assign new_new_n15716__ = new_new_n15517__ & ~new_new_n15693__;
  assign new_new_n15717__ = ~new_new_n15518__ & ~new_new_n15555__;
  assign new_new_n15718__ = new_new_n15691__ & new_new_n15717__;
  assign new_new_n15719__ = ~new_new_n15716__ & ~new_new_n15718__;
  assign new_new_n15720__ = new_new_n15696__ & ~new_new_n15719__;
  assign new_new_n15721__ = new_new_n15517__ & new_new_n15692__;
  assign new_new_n15722__ = new_new_n15518__ & new_new_n15555__;
  assign new_new_n15723__ = ~new_new_n15517__ & ~new_new_n15691__;
  assign new_new_n15724__ = ~new_new_n15722__ & ~new_new_n15723__;
  assign new_new_n15725__ = ~new_new_n15696__ & ~new_new_n15717__;
  assign new_new_n15726__ = ~new_new_n15724__ & new_new_n15725__;
  assign new_new_n15727__ = ~new_new_n15715__ & ~new_new_n15721__;
  assign new_new_n15728__ = ~new_new_n15726__ & new_new_n15727__;
  assign new_new_n15729__ = ~new_new_n15720__ & new_new_n15728__;
  assign new_new_n15730__ = ~new_new_n15608__ & ~new_new_n15642__;
  assign new_new_n15731__ = ~new_new_n15607__ & ~new_new_n15730__;
  assign new_new_n15732__ = ~new_new_n15673__ & ~new_new_n15685__;
  assign new_new_n15733__ = ~new_new_n15672__ & ~new_new_n15732__;
  assign new_new_n15734__ = new_new_n15731__ & ~new_new_n15733__;
  assign new_new_n15735__ = ~new_new_n15731__ & new_new_n15733__;
  assign new_new_n15736__ = ~new_new_n15734__ & ~new_new_n15735__;
  assign new_new_n15737__ = ~new_new_n15564__ & ~new_new_n15570__;
  assign new_new_n15738__ = ~new_new_n15569__ & ~new_new_n15737__;
  assign new_new_n15739__ = pi25 & pi62;
  assign new_new_n15740__ = new_new_n15679__ & new_new_n15739__;
  assign new_new_n15741__ = pi25 & pi61;
  assign new_new_n15742__ = pi42 & new_new_n15741__;
  assign new_new_n15743__ = ~pi62 & ~new_new_n15742__;
  assign new_new_n15744__ = ~pi24 & ~new_new_n15741__;
  assign new_new_n15745__ = ~pi23 & ~pi42;
  assign new_new_n15746__ = pi43 & ~new_new_n15745__;
  assign new_new_n15747__ = ~new_new_n15740__ & new_new_n15746__;
  assign new_new_n15748__ = ~new_new_n15744__ & new_new_n15747__;
  assign new_new_n15749__ = ~new_new_n15743__ & new_new_n15748__;
  assign new_new_n15750__ = pi42 & pi43;
  assign new_new_n15751__ = pi24 & ~new_new_n15741__;
  assign new_new_n15752__ = ~new_new_n10893__ & ~new_new_n15751__;
  assign new_new_n15753__ = pi62 & ~new_new_n15752__;
  assign new_new_n15754__ = pi24 & pi62;
  assign new_new_n15755__ = new_new_n15741__ & ~new_new_n15754__;
  assign new_new_n15756__ = ~new_new_n15750__ & ~new_new_n15755__;
  assign new_new_n15757__ = ~new_new_n15753__ & new_new_n15756__;
  assign new_new_n15758__ = ~new_new_n15749__ & ~new_new_n15757__;
  assign new_new_n15759__ = ~new_new_n15678__ & ~new_new_n15679__;
  assign new_new_n15760__ = new_new_n15678__ & new_new_n15679__;
  assign new_new_n15761__ = ~new_new_n15676__ & ~new_new_n15760__;
  assign new_new_n15762__ = ~new_new_n15759__ & ~new_new_n15761__;
  assign new_new_n15763__ = new_new_n15758__ & new_new_n15762__;
  assign new_new_n15764__ = ~new_new_n15758__ & ~new_new_n15762__;
  assign new_new_n15765__ = ~new_new_n15738__ & ~new_new_n15763__;
  assign new_new_n15766__ = ~new_new_n15764__ & ~new_new_n15765__;
  assign new_new_n15767__ = ~new_new_n15763__ & new_new_n15766__;
  assign new_new_n15768__ = new_new_n15738__ & ~new_new_n15767__;
  assign new_new_n15769__ = ~new_new_n15764__ & new_new_n15765__;
  assign new_new_n15770__ = ~new_new_n15768__ & ~new_new_n15769__;
  assign new_new_n15771__ = new_new_n15736__ & ~new_new_n15770__;
  assign new_new_n15772__ = ~new_new_n15736__ & new_new_n15770__;
  assign new_new_n15773__ = ~new_new_n15771__ & ~new_new_n15772__;
  assign new_new_n15774__ = ~new_new_n15545__ & new_new_n15549__;
  assign new_new_n15775__ = ~new_new_n15546__ & ~new_new_n15774__;
  assign new_new_n15776__ = new_new_n15773__ & new_new_n15775__;
  assign new_new_n15777__ = ~new_new_n15773__ & ~new_new_n15775__;
  assign new_new_n15778__ = ~new_new_n15776__ & ~new_new_n15777__;
  assign new_new_n15779__ = ~new_new_n15646__ & new_new_n15688__;
  assign new_new_n15780__ = ~new_new_n15647__ & ~new_new_n15779__;
  assign new_new_n15781__ = new_new_n15778__ & ~new_new_n15780__;
  assign new_new_n15782__ = ~new_new_n15778__ & new_new_n15780__;
  assign new_new_n15783__ = ~new_new_n15781__ & ~new_new_n15782__;
  assign new_new_n15784__ = ~new_new_n15530__ & new_new_n15552__;
  assign new_new_n15785__ = ~new_new_n15529__ & ~new_new_n15784__;
  assign new_new_n15786__ = new_new_n15783__ & new_new_n15785__;
  assign new_new_n15787__ = ~new_new_n15783__ & ~new_new_n15785__;
  assign new_new_n15788__ = ~new_new_n15786__ & ~new_new_n15787__;
  assign new_new_n15789__ = ~new_new_n15610__ & ~new_new_n15614__;
  assign new_new_n15790__ = ~new_new_n15613__ & ~new_new_n15789__;
  assign new_new_n15791__ = ~new_new_n15584__ & ~new_new_n15587__;
  assign new_new_n15792__ = ~new_new_n15586__ & ~new_new_n15791__;
  assign new_new_n15793__ = ~new_new_n15619__ & ~new_new_n15623__;
  assign new_new_n15794__ = ~new_new_n15622__ & ~new_new_n15793__;
  assign new_new_n15795__ = new_new_n15792__ & new_new_n15794__;
  assign new_new_n15796__ = ~new_new_n15792__ & ~new_new_n15794__;
  assign new_new_n15797__ = ~new_new_n15795__ & ~new_new_n15796__;
  assign new_new_n15798__ = new_new_n15790__ & ~new_new_n15797__;
  assign new_new_n15799__ = ~new_new_n15790__ & new_new_n15797__;
  assign new_new_n15800__ = ~new_new_n15798__ & ~new_new_n15799__;
  assign new_new_n15801__ = ~new_new_n15592__ & ~new_new_n15596__;
  assign new_new_n15802__ = ~new_new_n15595__ & ~new_new_n15801__;
  assign new_new_n15803__ = ~new_new_n15631__ & ~new_new_n15635__;
  assign new_new_n15804__ = ~new_new_n15634__ & ~new_new_n15803__;
  assign new_new_n15805__ = ~new_new_n15651__ & ~new_new_n15655__;
  assign new_new_n15806__ = ~new_new_n15654__ & ~new_new_n15805__;
  assign new_new_n15807__ = new_new_n15804__ & ~new_new_n15806__;
  assign new_new_n15808__ = ~new_new_n15804__ & new_new_n15806__;
  assign new_new_n15809__ = ~new_new_n15807__ & ~new_new_n15808__;
  assign new_new_n15810__ = new_new_n15802__ & new_new_n15809__;
  assign new_new_n15811__ = ~new_new_n15802__ & ~new_new_n15809__;
  assign new_new_n15812__ = ~new_new_n15810__ & ~new_new_n15811__;
  assign new_new_n15813__ = ~new_new_n15537__ & ~new_new_n15541__;
  assign new_new_n15814__ = ~new_new_n15538__ & ~new_new_n15813__;
  assign new_new_n15815__ = new_new_n15812__ & ~new_new_n15814__;
  assign new_new_n15816__ = ~new_new_n15812__ & new_new_n15814__;
  assign new_new_n15817__ = ~new_new_n15815__ & ~new_new_n15816__;
  assign new_new_n15818__ = new_new_n15800__ & new_new_n15817__;
  assign new_new_n15819__ = ~new_new_n15800__ & ~new_new_n15817__;
  assign new_new_n15820__ = ~new_new_n15818__ & ~new_new_n15819__;
  assign new_new_n15821__ = new_new_n15788__ & ~new_new_n15820__;
  assign new_new_n15822__ = ~new_new_n15788__ & new_new_n15820__;
  assign new_new_n15823__ = ~new_new_n15821__ & ~new_new_n15822__;
  assign new_new_n15824__ = ~new_new_n15729__ & new_new_n15823__;
  assign new_new_n15825__ = ~new_new_n15693__ & new_new_n15696__;
  assign new_new_n15826__ = ~new_new_n15692__ & ~new_new_n15825__;
  assign new_new_n15827__ = ~new_new_n15518__ & ~new_new_n15826__;
  assign new_new_n15828__ = ~new_new_n15517__ & new_new_n15826__;
  assign new_new_n15829__ = ~new_new_n15827__ & ~new_new_n15828__;
  assign new_new_n15830__ = new_new_n15693__ & ~new_new_n15696__;
  assign new_new_n15831__ = new_new_n15692__ & new_new_n15696__;
  assign new_new_n15832__ = ~new_new_n15830__ & ~new_new_n15831__;
  assign new_new_n15833__ = new_new_n15519__ & new_new_n15832__;
  assign new_new_n15834__ = ~new_new_n15829__ & ~new_new_n15833__;
  assign new_new_n15835__ = ~new_new_n15823__ & ~new_new_n15834__;
  assign new_new_n15836__ = ~new_new_n15824__ & ~new_new_n15835__;
  assign new_new_n15837__ = new_new_n15714__ & ~new_new_n15836__;
  assign new_new_n15838__ = ~new_new_n15714__ & new_new_n15836__;
  assign new_new_n15839__ = ~new_new_n15837__ & ~new_new_n15838__;
  assign new_new_n15840__ = pi40 & pi46;
  assign new_new_n15841__ = pi30 & pi56;
  assign new_new_n15842__ = pi39 & pi47;
  assign new_new_n15843__ = ~new_new_n15841__ & ~new_new_n15842__;
  assign new_new_n15844__ = new_new_n15841__ & new_new_n15842__;
  assign new_new_n15845__ = ~new_new_n15843__ & ~new_new_n15844__;
  assign new_new_n15846__ = new_new_n15840__ & ~new_new_n15845__;
  assign new_new_n15847__ = ~new_new_n15840__ & new_new_n15845__;
  assign new_new_n15848__ = ~new_new_n15846__ & ~new_new_n15847__;
  assign new_new_n15849__ = pi42 & pi44;
  assign new_new_n15850__ = pi41 & pi45;
  assign new_new_n15851__ = pi32 & pi54;
  assign new_new_n15852__ = ~new_new_n15850__ & ~new_new_n15851__;
  assign new_new_n15853__ = new_new_n15850__ & new_new_n15851__;
  assign new_new_n15854__ = ~new_new_n15852__ & ~new_new_n15853__;
  assign new_new_n15855__ = new_new_n15849__ & ~new_new_n15854__;
  assign new_new_n15856__ = ~new_new_n15849__ & new_new_n15854__;
  assign new_new_n15857__ = ~new_new_n15855__ & ~new_new_n15856__;
  assign new_new_n15858__ = new_new_n15848__ & new_new_n15857__;
  assign new_new_n15859__ = ~new_new_n15848__ & ~new_new_n15857__;
  assign new_new_n15860__ = ~new_new_n15858__ & ~new_new_n15859__;
  assign new_new_n15861__ = ~new_new_n15561__ & ~new_new_n15574__;
  assign new_new_n15862__ = ~new_new_n15560__ & ~new_new_n15861__;
  assign new_new_n15863__ = pi38 & pi48;
  assign new_new_n15864__ = pi31 & pi55;
  assign new_new_n15865__ = ~new_new_n8460__ & ~new_new_n15864__;
  assign new_new_n15866__ = new_new_n8460__ & new_new_n15864__;
  assign new_new_n15867__ = ~new_new_n15865__ & ~new_new_n15866__;
  assign new_new_n15868__ = new_new_n15863__ & ~new_new_n15867__;
  assign new_new_n15869__ = ~new_new_n15863__ & new_new_n15867__;
  assign new_new_n15870__ = ~new_new_n15868__ & ~new_new_n15869__;
  assign new_new_n15871__ = pi37 & pi49;
  assign new_new_n15872__ = pi23 & pi63;
  assign new_new_n15873__ = pi36 & pi50;
  assign new_new_n15874__ = ~new_new_n15872__ & ~new_new_n15873__;
  assign new_new_n15875__ = new_new_n15872__ & new_new_n15873__;
  assign new_new_n15876__ = ~new_new_n15874__ & ~new_new_n15875__;
  assign new_new_n15877__ = new_new_n15871__ & ~new_new_n15876__;
  assign new_new_n15878__ = ~new_new_n15871__ & new_new_n15876__;
  assign new_new_n15879__ = ~new_new_n15877__ & ~new_new_n15878__;
  assign new_new_n15880__ = new_new_n15870__ & new_new_n15879__;
  assign new_new_n15881__ = ~new_new_n15870__ & ~new_new_n15879__;
  assign new_new_n15882__ = ~new_new_n15880__ & ~new_new_n15881__;
  assign new_new_n15883__ = pi35 & pi51;
  assign new_new_n15884__ = pi33 & pi53;
  assign new_new_n15885__ = pi34 & pi52;
  assign new_new_n15886__ = ~new_new_n15884__ & ~new_new_n15885__;
  assign new_new_n15887__ = new_new_n15884__ & new_new_n15885__;
  assign new_new_n15888__ = ~new_new_n15886__ & ~new_new_n15887__;
  assign new_new_n15889__ = new_new_n15883__ & ~new_new_n15888__;
  assign new_new_n15890__ = ~new_new_n15883__ & new_new_n15888__;
  assign new_new_n15891__ = ~new_new_n15889__ & ~new_new_n15890__;
  assign new_new_n15892__ = new_new_n15882__ & ~new_new_n15891__;
  assign new_new_n15893__ = ~new_new_n15882__ & new_new_n15891__;
  assign new_new_n15894__ = ~new_new_n15892__ & ~new_new_n15893__;
  assign new_new_n15895__ = ~new_new_n15862__ & new_new_n15894__;
  assign new_new_n15896__ = new_new_n15862__ & ~new_new_n15894__;
  assign new_new_n15897__ = ~new_new_n15895__ & ~new_new_n15896__;
  assign new_new_n15898__ = pi28 & pi58;
  assign new_new_n15899__ = pi26 & pi60;
  assign new_new_n15900__ = pi27 & pi59;
  assign new_new_n15901__ = ~new_new_n15899__ & ~new_new_n15900__;
  assign new_new_n15902__ = new_new_n15899__ & new_new_n15900__;
  assign new_new_n15903__ = ~new_new_n15901__ & ~new_new_n15902__;
  assign new_new_n15904__ = new_new_n15898__ & ~new_new_n15903__;
  assign new_new_n15905__ = ~new_new_n15898__ & new_new_n15903__;
  assign new_new_n15906__ = ~new_new_n15904__ & ~new_new_n15905__;
  assign new_new_n15907__ = new_new_n15897__ & ~new_new_n15906__;
  assign new_new_n15908__ = ~new_new_n15897__ & new_new_n15906__;
  assign new_new_n15909__ = ~new_new_n15907__ & ~new_new_n15908__;
  assign new_new_n15910__ = new_new_n15860__ & new_new_n15909__;
  assign new_new_n15911__ = ~new_new_n15860__ & ~new_new_n15909__;
  assign new_new_n15912__ = ~new_new_n15910__ & ~new_new_n15911__;
  assign new_new_n15913__ = new_new_n15839__ & new_new_n15912__;
  assign new_new_n15914__ = ~new_new_n15839__ & ~new_new_n15912__;
  assign po087 = new_new_n15913__ | new_new_n15914__;
  assign new_new_n15916__ = ~new_new_n15827__ & po087;
  assign new_new_n15917__ = new_new_n15518__ & new_new_n15826__;
  assign new_new_n15918__ = ~new_new_n15830__ & ~po087;
  assign new_new_n15919__ = ~new_new_n15517__ & ~new_new_n15831__;
  assign new_new_n15920__ = ~new_new_n15918__ & new_new_n15919__;
  assign new_new_n15921__ = ~new_new_n15916__ & ~new_new_n15917__;
  assign new_new_n15922__ = ~new_new_n15920__ & new_new_n15921__;
  assign new_new_n15923__ = new_new_n15714__ & new_new_n15820__;
  assign new_new_n15924__ = ~new_new_n15714__ & ~new_new_n15820__;
  assign new_new_n15925__ = ~new_new_n15923__ & ~new_new_n15924__;
  assign new_new_n15926__ = new_new_n15912__ & ~new_new_n15925__;
  assign new_new_n15927__ = ~new_new_n15912__ & new_new_n15925__;
  assign new_new_n15928__ = ~new_new_n15926__ & ~new_new_n15927__;
  assign new_new_n15929__ = new_new_n15788__ & new_new_n15928__;
  assign new_new_n15930__ = ~new_new_n15786__ & ~new_new_n15929__;
  assign new_new_n15931__ = ~new_new_n15922__ & ~new_new_n15930__;
  assign new_new_n15932__ = new_new_n15922__ & new_new_n15930__;
  assign new_new_n15933__ = ~new_new_n15931__ & ~new_new_n15932__;
  assign new_new_n15934__ = ~new_new_n15776__ & ~new_new_n15780__;
  assign new_new_n15935__ = ~new_new_n15777__ & ~new_new_n15934__;
  assign new_new_n15936__ = new_new_n15797__ & ~new_new_n15802__;
  assign new_new_n15937__ = ~new_new_n15797__ & new_new_n15802__;
  assign new_new_n15938__ = ~new_new_n15936__ & ~new_new_n15937__;
  assign new_new_n15939__ = new_new_n15814__ & new_new_n15938__;
  assign new_new_n15940__ = ~new_new_n15814__ & ~new_new_n15938__;
  assign new_new_n15941__ = new_new_n15790__ & new_new_n15809__;
  assign new_new_n15942__ = ~new_new_n15790__ & ~new_new_n15809__;
  assign new_new_n15943__ = ~new_new_n15941__ & ~new_new_n15942__;
  assign new_new_n15944__ = ~new_new_n15940__ & new_new_n15943__;
  assign new_new_n15945__ = ~new_new_n15939__ & ~new_new_n15944__;
  assign new_new_n15946__ = ~new_new_n15898__ & ~new_new_n15902__;
  assign new_new_n15947__ = ~new_new_n15901__ & ~new_new_n15946__;
  assign new_new_n15948__ = ~new_new_n15871__ & ~new_new_n15875__;
  assign new_new_n15949__ = ~new_new_n15874__ & ~new_new_n15948__;
  assign new_new_n15950__ = ~new_new_n15947__ & ~new_new_n15949__;
  assign new_new_n15951__ = new_new_n15947__ & new_new_n15949__;
  assign new_new_n15952__ = ~new_new_n15950__ & ~new_new_n15951__;
  assign new_new_n15953__ = ~new_new_n15883__ & ~new_new_n15887__;
  assign new_new_n15954__ = ~new_new_n15886__ & ~new_new_n15953__;
  assign new_new_n15955__ = ~new_new_n15952__ & new_new_n15954__;
  assign new_new_n15956__ = ~new_new_n15951__ & ~new_new_n15954__;
  assign new_new_n15957__ = ~new_new_n15950__ & new_new_n15956__;
  assign new_new_n15958__ = ~new_new_n15955__ & ~new_new_n15957__;
  assign new_new_n15959__ = ~new_new_n15766__ & new_new_n15958__;
  assign new_new_n15960__ = new_new_n15766__ & ~new_new_n15958__;
  assign new_new_n15961__ = ~new_new_n15959__ & ~new_new_n15960__;
  assign new_new_n15962__ = ~new_new_n15840__ & ~new_new_n15844__;
  assign new_new_n15963__ = ~new_new_n15843__ & ~new_new_n15962__;
  assign new_new_n15964__ = ~new_new_n15849__ & ~new_new_n15853__;
  assign new_new_n15965__ = ~new_new_n15852__ & ~new_new_n15964__;
  assign new_new_n15966__ = ~new_new_n15863__ & ~new_new_n15866__;
  assign new_new_n15967__ = ~new_new_n15865__ & ~new_new_n15966__;
  assign new_new_n15968__ = new_new_n15965__ & new_new_n15967__;
  assign new_new_n15969__ = ~new_new_n15965__ & ~new_new_n15967__;
  assign new_new_n15970__ = ~new_new_n15968__ & ~new_new_n15969__;
  assign new_new_n15971__ = new_new_n15963__ & ~new_new_n15970__;
  assign new_new_n15972__ = ~new_new_n15963__ & new_new_n15970__;
  assign new_new_n15973__ = ~new_new_n15971__ & ~new_new_n15972__;
  assign new_new_n15974__ = new_new_n15961__ & ~new_new_n15973__;
  assign new_new_n15975__ = ~new_new_n15961__ & new_new_n15973__;
  assign new_new_n15976__ = ~new_new_n15974__ & ~new_new_n15975__;
  assign new_new_n15977__ = new_new_n15945__ & new_new_n15976__;
  assign new_new_n15978__ = ~new_new_n15945__ & ~new_new_n15976__;
  assign new_new_n15979__ = ~new_new_n15977__ & ~new_new_n15978__;
  assign new_new_n15980__ = ~new_new_n15704__ & ~new_new_n15709__;
  assign new_new_n15981__ = ~new_new_n15710__ & ~new_new_n15980__;
  assign new_new_n15982__ = new_new_n15979__ & ~new_new_n15981__;
  assign new_new_n15983__ = ~new_new_n15979__ & new_new_n15981__;
  assign new_new_n15984__ = ~new_new_n15982__ & ~new_new_n15983__;
  assign new_new_n15985__ = ~pi43 & pi44;
  assign new_new_n15986__ = new_new_n15739__ & ~new_new_n15985__;
  assign new_new_n15987__ = ~new_new_n15739__ & new_new_n15985__;
  assign new_new_n15988__ = ~new_new_n15986__ & ~new_new_n15987__;
  assign new_new_n15989__ = pi40 & pi47;
  assign new_new_n15990__ = pi33 & pi54;
  assign new_new_n15991__ = pi31 & pi56;
  assign new_new_n15992__ = ~new_new_n15990__ & ~new_new_n15991__;
  assign new_new_n15993__ = new_new_n15990__ & new_new_n15991__;
  assign new_new_n15994__ = ~new_new_n15992__ & ~new_new_n15993__;
  assign new_new_n15995__ = new_new_n15989__ & ~new_new_n15994__;
  assign new_new_n15996__ = ~new_new_n15989__ & new_new_n15994__;
  assign new_new_n15997__ = ~new_new_n15995__ & ~new_new_n15996__;
  assign new_new_n15998__ = new_new_n15988__ & new_new_n15997__;
  assign new_new_n15999__ = ~new_new_n15988__ & ~new_new_n15997__;
  assign new_new_n16000__ = ~new_new_n15998__ & ~new_new_n15999__;
  assign new_new_n16001__ = ~new_new_n15790__ & ~new_new_n15806__;
  assign new_new_n16002__ = new_new_n15790__ & new_new_n15806__;
  assign new_new_n16003__ = ~new_new_n15804__ & ~new_new_n16002__;
  assign new_new_n16004__ = ~new_new_n16001__ & ~new_new_n16003__;
  assign new_new_n16005__ = new_new_n16000__ & new_new_n16004__;
  assign new_new_n16006__ = ~new_new_n16000__ & ~new_new_n16004__;
  assign new_new_n16007__ = ~new_new_n16005__ & ~new_new_n16006__;
  assign new_new_n16008__ = pi36 & pi51;
  assign new_new_n16009__ = pi35 & pi52;
  assign new_new_n16010__ = pi29 & pi58;
  assign new_new_n16011__ = ~new_new_n16009__ & ~new_new_n16010__;
  assign new_new_n16012__ = new_new_n16009__ & new_new_n16010__;
  assign new_new_n16013__ = ~new_new_n16011__ & ~new_new_n16012__;
  assign new_new_n16014__ = new_new_n16008__ & ~new_new_n16013__;
  assign new_new_n16015__ = ~new_new_n16008__ & new_new_n16013__;
  assign new_new_n16016__ = ~new_new_n16014__ & ~new_new_n16015__;
  assign new_new_n16017__ = pi34 & pi53;
  assign new_new_n16018__ = pi30 & pi57;
  assign new_new_n16019__ = pi28 & pi59;
  assign new_new_n16020__ = ~new_new_n16018__ & ~new_new_n16019__;
  assign new_new_n16021__ = new_new_n16018__ & new_new_n16019__;
  assign new_new_n16022__ = ~new_new_n16020__ & ~new_new_n16021__;
  assign new_new_n16023__ = new_new_n16017__ & ~new_new_n16022__;
  assign new_new_n16024__ = ~new_new_n16017__ & new_new_n16022__;
  assign new_new_n16025__ = ~new_new_n16023__ & ~new_new_n16024__;
  assign new_new_n16026__ = new_new_n16016__ & new_new_n16025__;
  assign new_new_n16027__ = ~new_new_n16016__ & ~new_new_n16025__;
  assign new_new_n16028__ = ~new_new_n16026__ & ~new_new_n16027__;
  assign new_new_n16029__ = pi23 & ~new_new_n15744__;
  assign new_new_n16030__ = ~new_new_n10892__ & ~new_new_n16029__;
  assign new_new_n16031__ = pi43 & ~new_new_n16030__;
  assign new_new_n16032__ = pi25 & new_new_n15679__;
  assign new_new_n16033__ = ~new_new_n16031__ & ~new_new_n16032__;
  assign new_new_n16034__ = pi62 & ~new_new_n16033__;
  assign new_new_n16035__ = pi43 & new_new_n15742__;
  assign new_new_n16036__ = ~new_new_n16034__ & ~new_new_n16035__;
  assign new_new_n16037__ = new_new_n16028__ & ~new_new_n16036__;
  assign new_new_n16038__ = ~new_new_n16028__ & new_new_n16036__;
  assign new_new_n16039__ = ~new_new_n16037__ & ~new_new_n16038__;
  assign new_new_n16040__ = pi39 & pi48;
  assign new_new_n16041__ = pi37 & pi50;
  assign new_new_n16042__ = pi38 & pi49;
  assign new_new_n16043__ = ~new_new_n16041__ & ~new_new_n16042__;
  assign new_new_n16044__ = new_new_n16041__ & new_new_n16042__;
  assign new_new_n16045__ = ~new_new_n16043__ & ~new_new_n16044__;
  assign new_new_n16046__ = new_new_n16040__ & ~new_new_n16045__;
  assign new_new_n16047__ = ~new_new_n16040__ & new_new_n16045__;
  assign new_new_n16048__ = ~new_new_n16046__ & ~new_new_n16047__;
  assign new_new_n16049__ = pi42 & pi45;
  assign new_new_n16050__ = pi41 & pi46;
  assign new_new_n16051__ = pi32 & pi55;
  assign new_new_n16052__ = ~new_new_n16050__ & ~new_new_n16051__;
  assign new_new_n16053__ = new_new_n16050__ & new_new_n16051__;
  assign new_new_n16054__ = ~new_new_n16052__ & ~new_new_n16053__;
  assign new_new_n16055__ = new_new_n16049__ & ~new_new_n16054__;
  assign new_new_n16056__ = ~new_new_n16049__ & new_new_n16054__;
  assign new_new_n16057__ = ~new_new_n16055__ & ~new_new_n16056__;
  assign new_new_n16058__ = new_new_n16048__ & new_new_n16057__;
  assign new_new_n16059__ = ~new_new_n16048__ & ~new_new_n16057__;
  assign new_new_n16060__ = ~new_new_n16058__ & ~new_new_n16059__;
  assign new_new_n16061__ = pi27 & pi60;
  assign new_new_n16062__ = pi26 & pi61;
  assign new_new_n16063__ = pi24 & pi63;
  assign new_new_n16064__ = ~new_new_n16062__ & ~new_new_n16063__;
  assign new_new_n16065__ = new_new_n16062__ & new_new_n16063__;
  assign new_new_n16066__ = ~new_new_n16064__ & ~new_new_n16065__;
  assign new_new_n16067__ = new_new_n16061__ & ~new_new_n16066__;
  assign new_new_n16068__ = ~new_new_n16061__ & new_new_n16066__;
  assign new_new_n16069__ = ~new_new_n16067__ & ~new_new_n16068__;
  assign new_new_n16070__ = new_new_n16060__ & ~new_new_n16069__;
  assign new_new_n16071__ = ~new_new_n16060__ & new_new_n16069__;
  assign new_new_n16072__ = ~new_new_n16070__ & ~new_new_n16071__;
  assign new_new_n16073__ = new_new_n16039__ & new_new_n16072__;
  assign new_new_n16074__ = ~new_new_n16039__ & ~new_new_n16072__;
  assign new_new_n16075__ = ~new_new_n16073__ & ~new_new_n16074__;
  assign new_new_n16076__ = new_new_n16007__ & new_new_n16075__;
  assign new_new_n16077__ = ~new_new_n16007__ & ~new_new_n16075__;
  assign new_new_n16078__ = ~new_new_n16076__ & ~new_new_n16077__;
  assign new_new_n16079__ = new_new_n15984__ & new_new_n16078__;
  assign new_new_n16080__ = ~new_new_n15984__ & ~new_new_n16078__;
  assign new_new_n16081__ = ~new_new_n16079__ & ~new_new_n16080__;
  assign new_new_n16082__ = new_new_n15912__ & ~new_new_n15924__;
  assign new_new_n16083__ = ~new_new_n15923__ & ~new_new_n16082__;
  assign new_new_n16084__ = new_new_n16081__ & ~new_new_n16083__;
  assign new_new_n16085__ = ~new_new_n16081__ & new_new_n16083__;
  assign new_new_n16086__ = ~new_new_n16084__ & ~new_new_n16085__;
  assign new_new_n16087__ = new_new_n15935__ & new_new_n16086__;
  assign new_new_n16088__ = ~new_new_n15935__ & ~new_new_n16086__;
  assign new_new_n16089__ = ~new_new_n16087__ & ~new_new_n16088__;
  assign new_new_n16090__ = ~new_new_n15734__ & new_new_n15770__;
  assign new_new_n16091__ = ~new_new_n15735__ & ~new_new_n16090__;
  assign new_new_n16092__ = ~new_new_n15858__ & ~new_new_n15906__;
  assign new_new_n16093__ = ~new_new_n15859__ & ~new_new_n16092__;
  assign new_new_n16094__ = new_new_n15895__ & new_new_n16093__;
  assign new_new_n16095__ = new_new_n15858__ & new_new_n15906__;
  assign new_new_n16096__ = new_new_n15859__ & ~new_new_n15906__;
  assign new_new_n16097__ = ~new_new_n16095__ & ~new_new_n16096__;
  assign new_new_n16098__ = new_new_n15897__ & new_new_n16097__;
  assign new_new_n16099__ = new_new_n15896__ & ~new_new_n16093__;
  assign new_new_n16100__ = ~new_new_n16094__ & ~new_new_n16099__;
  assign new_new_n16101__ = ~new_new_n16098__ & new_new_n16100__;
  assign new_new_n16102__ = new_new_n16091__ & ~new_new_n16101__;
  assign new_new_n16103__ = new_new_n15859__ & new_new_n15895__;
  assign new_new_n16104__ = ~new_new_n15857__ & new_new_n15895__;
  assign new_new_n16105__ = new_new_n15857__ & ~new_new_n15895__;
  assign new_new_n16106__ = ~new_new_n15848__ & ~new_new_n15896__;
  assign new_new_n16107__ = ~new_new_n16105__ & new_new_n16106__;
  assign new_new_n16108__ = ~new_new_n16104__ & ~new_new_n16107__;
  assign new_new_n16109__ = ~new_new_n15906__ & ~new_new_n16108__;
  assign new_new_n16110__ = new_new_n15858__ & new_new_n15896__;
  assign new_new_n16111__ = ~new_new_n15859__ & new_new_n15896__;
  assign new_new_n16112__ = new_new_n15858__ & ~new_new_n15895__;
  assign new_new_n16113__ = ~new_new_n16111__ & ~new_new_n16112__;
  assign new_new_n16114__ = new_new_n15906__ & ~new_new_n16113__;
  assign new_new_n16115__ = ~new_new_n16103__ & ~new_new_n16110__;
  assign new_new_n16116__ = ~new_new_n16114__ & new_new_n16115__;
  assign new_new_n16117__ = ~new_new_n16109__ & new_new_n16116__;
  assign new_new_n16118__ = ~new_new_n16091__ & ~new_new_n16117__;
  assign new_new_n16119__ = ~new_new_n16102__ & ~new_new_n16118__;
  assign new_new_n16120__ = ~new_new_n15795__ & ~new_new_n15802__;
  assign new_new_n16121__ = ~new_new_n15796__ & ~new_new_n16120__;
  assign new_new_n16122__ = ~new_new_n15880__ & ~new_new_n15891__;
  assign new_new_n16123__ = ~new_new_n15881__ & ~new_new_n16122__;
  assign new_new_n16124__ = ~new_new_n16121__ & new_new_n16123__;
  assign new_new_n16125__ = new_new_n16121__ & ~new_new_n16123__;
  assign new_new_n16126__ = ~new_new_n16124__ & ~new_new_n16125__;
  assign new_new_n16127__ = new_new_n16119__ & new_new_n16126__;
  assign new_new_n16128__ = ~new_new_n16119__ & ~new_new_n16126__;
  assign new_new_n16129__ = ~new_new_n16127__ & ~new_new_n16128__;
  assign new_new_n16130__ = new_new_n16089__ & ~new_new_n16129__;
  assign new_new_n16131__ = ~new_new_n16089__ & new_new_n16129__;
  assign new_new_n16132__ = ~new_new_n16130__ & ~new_new_n16131__;
  assign new_new_n16133__ = new_new_n15933__ & new_new_n16132__;
  assign new_new_n16134__ = ~new_new_n15933__ & ~new_new_n16132__;
  assign po088 = new_new_n16133__ | new_new_n16134__;
  assign new_new_n16136__ = ~new_new_n16087__ & ~new_new_n16129__;
  assign new_new_n16137__ = ~new_new_n16088__ & ~new_new_n16136__;
  assign new_new_n16138__ = ~new_new_n15977__ & new_new_n15981__;
  assign new_new_n16139__ = ~new_new_n15978__ & ~new_new_n16138__;
  assign new_new_n16140__ = ~new_new_n16093__ & ~new_new_n16119__;
  assign new_new_n16141__ = ~new_new_n16123__ & ~new_new_n16140__;
  assign new_new_n16142__ = new_new_n16093__ & new_new_n16119__;
  assign new_new_n16143__ = new_new_n16123__ & ~new_new_n16142__;
  assign new_new_n16144__ = new_new_n16121__ & ~new_new_n16141__;
  assign new_new_n16145__ = ~new_new_n16143__ & new_new_n16144__;
  assign new_new_n16146__ = ~new_new_n16123__ & ~new_new_n16142__;
  assign new_new_n16147__ = new_new_n16123__ & ~new_new_n16140__;
  assign new_new_n16148__ = ~new_new_n16121__ & ~new_new_n16146__;
  assign new_new_n16149__ = ~new_new_n16147__ & new_new_n16148__;
  assign new_new_n16150__ = new_new_n16091__ & ~new_new_n16140__;
  assign new_new_n16151__ = ~new_new_n16142__ & new_new_n16150__;
  assign new_new_n16152__ = ~new_new_n16145__ & ~new_new_n16151__;
  assign new_new_n16153__ = ~new_new_n16149__ & new_new_n16152__;
  assign new_new_n16154__ = new_new_n16139__ & ~new_new_n16153__;
  assign new_new_n16155__ = ~new_new_n16139__ & new_new_n16153__;
  assign new_new_n16156__ = ~new_new_n16154__ & ~new_new_n16155__;
  assign new_new_n16157__ = ~new_new_n16026__ & ~new_new_n16036__;
  assign new_new_n16158__ = ~new_new_n16027__ & ~new_new_n16157__;
  assign new_new_n16159__ = ~new_new_n15950__ & ~new_new_n15956__;
  assign new_new_n16160__ = ~new_new_n16158__ & new_new_n16159__;
  assign new_new_n16161__ = new_new_n16158__ & ~new_new_n16159__;
  assign new_new_n16162__ = ~new_new_n16160__ & ~new_new_n16161__;
  assign new_new_n16163__ = ~new_new_n16058__ & ~new_new_n16069__;
  assign new_new_n16164__ = ~new_new_n16059__ & ~new_new_n16163__;
  assign new_new_n16165__ = new_new_n16162__ & ~new_new_n16164__;
  assign new_new_n16166__ = ~new_new_n16162__ & new_new_n16164__;
  assign new_new_n16167__ = ~new_new_n16165__ & ~new_new_n16166__;
  assign new_new_n16168__ = ~new_new_n16069__ & new_new_n16167__;
  assign new_new_n16169__ = new_new_n16069__ & ~new_new_n16167__;
  assign new_new_n16170__ = ~new_new_n16168__ & ~new_new_n16169__;
  assign new_new_n16171__ = ~new_new_n16060__ & ~new_new_n16170__;
  assign new_new_n16172__ = new_new_n16060__ & new_new_n16162__;
  assign new_new_n16173__ = ~new_new_n16075__ & ~new_new_n16172__;
  assign new_new_n16174__ = ~new_new_n16171__ & new_new_n16173__;
  assign new_new_n16175__ = ~new_new_n16007__ & ~new_new_n16167__;
  assign new_new_n16176__ = new_new_n16007__ & new_new_n16167__;
  assign new_new_n16177__ = new_new_n16075__ & ~new_new_n16175__;
  assign new_new_n16178__ = ~new_new_n16176__ & new_new_n16177__;
  assign new_new_n16179__ = ~new_new_n16174__ & ~new_new_n16178__;
  assign new_new_n16180__ = ~new_new_n16049__ & ~new_new_n16053__;
  assign new_new_n16181__ = ~new_new_n16052__ & ~new_new_n16180__;
  assign new_new_n16182__ = pi63 & new_new_n16181__;
  assign new_new_n16183__ = pi25 & new_new_n16182__;
  assign new_new_n16184__ = ~pi63 & ~new_new_n16181__;
  assign new_new_n16185__ = ~pi25 & ~new_new_n16181__;
  assign new_new_n16186__ = ~new_new_n16184__ & ~new_new_n16185__;
  assign new_new_n16187__ = ~new_new_n16183__ & new_new_n16186__;
  assign new_new_n16188__ = pi43 & ~new_new_n16187__;
  assign new_new_n16189__ = ~pi43 & new_new_n16182__;
  assign new_new_n16190__ = pi25 & new_new_n16184__;
  assign new_new_n16191__ = ~new_new_n16189__ & ~new_new_n16190__;
  assign new_new_n16192__ = pi62 & ~new_new_n16191__;
  assign new_new_n16193__ = ~new_new_n16188__ & ~new_new_n16192__;
  assign new_new_n16194__ = pi44 & ~new_new_n16193__;
  assign new_new_n16195__ = pi43 & pi44;
  assign new_new_n16196__ = pi44 & pi62;
  assign new_new_n16197__ = ~new_new_n16182__ & ~new_new_n16196__;
  assign new_new_n16198__ = pi25 & ~new_new_n16197__;
  assign new_new_n16199__ = new_new_n16186__ & ~new_new_n16195__;
  assign new_new_n16200__ = ~new_new_n16198__ & new_new_n16199__;
  assign new_new_n16201__ = ~new_new_n16194__ & ~new_new_n16200__;
  assign new_new_n16202__ = ~new_new_n15963__ & ~new_new_n15968__;
  assign new_new_n16203__ = ~new_new_n15969__ & ~new_new_n16202__;
  assign new_new_n16204__ = pi40 & pi48;
  assign new_new_n16205__ = pi32 & pi56;
  assign new_new_n16206__ = ~new_new_n8827__ & ~new_new_n16205__;
  assign new_new_n16207__ = new_new_n8827__ & new_new_n16205__;
  assign new_new_n16208__ = ~new_new_n16206__ & ~new_new_n16207__;
  assign new_new_n16209__ = new_new_n16204__ & ~new_new_n16208__;
  assign new_new_n16210__ = ~new_new_n16204__ & new_new_n16208__;
  assign new_new_n16211__ = ~new_new_n16209__ & ~new_new_n16210__;
  assign new_new_n16212__ = pi39 & pi49;
  assign new_new_n16213__ = pi38 & pi50;
  assign new_new_n16214__ = ~new_new_n9333__ & ~new_new_n16213__;
  assign new_new_n16215__ = new_new_n9333__ & new_new_n16213__;
  assign new_new_n16216__ = ~new_new_n16214__ & ~new_new_n16215__;
  assign new_new_n16217__ = new_new_n16212__ & ~new_new_n16216__;
  assign new_new_n16218__ = ~new_new_n16212__ & new_new_n16216__;
  assign new_new_n16219__ = ~new_new_n16217__ & ~new_new_n16218__;
  assign new_new_n16220__ = new_new_n16211__ & new_new_n16219__;
  assign new_new_n16221__ = ~new_new_n16211__ & ~new_new_n16219__;
  assign new_new_n16222__ = ~new_new_n16220__ & ~new_new_n16221__;
  assign new_new_n16223__ = new_new_n16203__ & new_new_n16222__;
  assign new_new_n16224__ = ~new_new_n16203__ & ~new_new_n16222__;
  assign new_new_n16225__ = ~new_new_n16223__ & ~new_new_n16224__;
  assign new_new_n16226__ = ~new_new_n16201__ & new_new_n16225__;
  assign new_new_n16227__ = new_new_n16201__ & ~new_new_n16225__;
  assign new_new_n16228__ = ~new_new_n16226__ & ~new_new_n16227__;
  assign new_new_n16229__ = pi37 & pi51;
  assign new_new_n16230__ = pi36 & pi52;
  assign new_new_n16231__ = pi35 & pi53;
  assign new_new_n16232__ = ~new_new_n16230__ & ~new_new_n16231__;
  assign new_new_n16233__ = new_new_n16230__ & new_new_n16231__;
  assign new_new_n16234__ = ~new_new_n16232__ & ~new_new_n16233__;
  assign new_new_n16235__ = new_new_n16229__ & ~new_new_n16234__;
  assign new_new_n16236__ = ~new_new_n16229__ & new_new_n16234__;
  assign new_new_n16237__ = ~new_new_n16235__ & ~new_new_n16236__;
  assign new_new_n16238__ = pi28 & pi60;
  assign new_new_n16239__ = pi27 & pi61;
  assign new_new_n16240__ = pi26 & pi62;
  assign new_new_n16241__ = ~new_new_n16239__ & ~new_new_n16240__;
  assign new_new_n16242__ = new_new_n16239__ & new_new_n16240__;
  assign new_new_n16243__ = ~new_new_n16241__ & ~new_new_n16242__;
  assign new_new_n16244__ = new_new_n16238__ & ~new_new_n16243__;
  assign new_new_n16245__ = ~new_new_n16238__ & new_new_n16243__;
  assign new_new_n16246__ = ~new_new_n16244__ & ~new_new_n16245__;
  assign new_new_n16247__ = new_new_n16237__ & new_new_n16246__;
  assign new_new_n16248__ = ~new_new_n16237__ & ~new_new_n16246__;
  assign new_new_n16249__ = ~new_new_n16247__ & ~new_new_n16248__;
  assign new_new_n16250__ = pi42 & pi46;
  assign new_new_n16251__ = pi31 & pi57;
  assign new_new_n16252__ = pi41 & pi47;
  assign new_new_n16253__ = ~new_new_n16251__ & ~new_new_n16252__;
  assign new_new_n16254__ = new_new_n16251__ & new_new_n16252__;
  assign new_new_n16255__ = ~new_new_n16253__ & ~new_new_n16254__;
  assign new_new_n16256__ = new_new_n16250__ & ~new_new_n16255__;
  assign new_new_n16257__ = ~new_new_n16250__ & new_new_n16255__;
  assign new_new_n16258__ = ~new_new_n16256__ & ~new_new_n16257__;
  assign new_new_n16259__ = new_new_n16249__ & ~new_new_n16258__;
  assign new_new_n16260__ = ~new_new_n16249__ & new_new_n16258__;
  assign new_new_n16261__ = ~new_new_n16259__ & ~new_new_n16260__;
  assign new_new_n16262__ = new_new_n16228__ & ~new_new_n16261__;
  assign new_new_n16263__ = ~new_new_n16228__ & new_new_n16261__;
  assign new_new_n16264__ = ~new_new_n16262__ & ~new_new_n16263__;
  assign new_new_n16265__ = ~new_new_n15960__ & new_new_n15973__;
  assign new_new_n16266__ = ~new_new_n15959__ & ~new_new_n16265__;
  assign new_new_n16267__ = ~new_new_n16040__ & ~new_new_n16044__;
  assign new_new_n16268__ = ~new_new_n16043__ & ~new_new_n16267__;
  assign new_new_n16269__ = ~new_new_n16017__ & ~new_new_n16021__;
  assign new_new_n16270__ = ~new_new_n16020__ & ~new_new_n16269__;
  assign new_new_n16271__ = ~new_new_n16061__ & ~new_new_n16065__;
  assign new_new_n16272__ = ~new_new_n16064__ & ~new_new_n16271__;
  assign new_new_n16273__ = new_new_n16270__ & new_new_n16272__;
  assign new_new_n16274__ = ~new_new_n16270__ & ~new_new_n16272__;
  assign new_new_n16275__ = ~new_new_n16273__ & ~new_new_n16274__;
  assign new_new_n16276__ = ~new_new_n16268__ & ~new_new_n16275__;
  assign new_new_n16277__ = new_new_n16268__ & new_new_n16275__;
  assign new_new_n16278__ = ~new_new_n16276__ & ~new_new_n16277__;
  assign new_new_n16279__ = ~new_new_n15999__ & ~new_new_n16004__;
  assign new_new_n16280__ = ~new_new_n15998__ & ~new_new_n16279__;
  assign new_new_n16281__ = ~new_new_n15989__ & ~new_new_n15993__;
  assign new_new_n16282__ = ~new_new_n15992__ & ~new_new_n16281__;
  assign new_new_n16283__ = pi43 & pi45;
  assign new_new_n16284__ = pi34 & pi54;
  assign new_new_n16285__ = pi33 & pi55;
  assign new_new_n16286__ = ~new_new_n16284__ & ~new_new_n16285__;
  assign new_new_n16287__ = new_new_n16284__ & new_new_n16285__;
  assign new_new_n16288__ = ~new_new_n16286__ & ~new_new_n16287__;
  assign new_new_n16289__ = new_new_n16283__ & ~new_new_n16288__;
  assign new_new_n16290__ = ~new_new_n16283__ & new_new_n16288__;
  assign new_new_n16291__ = ~new_new_n16289__ & ~new_new_n16290__;
  assign new_new_n16292__ = ~new_new_n16282__ & new_new_n16291__;
  assign new_new_n16293__ = new_new_n16282__ & ~new_new_n16291__;
  assign new_new_n16294__ = ~new_new_n16292__ & ~new_new_n16293__;
  assign new_new_n16295__ = ~new_new_n16008__ & ~new_new_n16012__;
  assign new_new_n16296__ = ~new_new_n16011__ & ~new_new_n16295__;
  assign new_new_n16297__ = new_new_n16294__ & ~new_new_n16296__;
  assign new_new_n16298__ = ~new_new_n16294__ & new_new_n16296__;
  assign new_new_n16299__ = ~new_new_n16297__ & ~new_new_n16298__;
  assign new_new_n16300__ = new_new_n16280__ & ~new_new_n16299__;
  assign new_new_n16301__ = ~new_new_n16280__ & new_new_n16299__;
  assign new_new_n16302__ = ~new_new_n16300__ & ~new_new_n16301__;
  assign new_new_n16303__ = new_new_n16278__ & ~new_new_n16302__;
  assign new_new_n16304__ = ~new_new_n16278__ & new_new_n16302__;
  assign new_new_n16305__ = ~new_new_n16303__ & ~new_new_n16304__;
  assign new_new_n16306__ = new_new_n16266__ & ~new_new_n16305__;
  assign new_new_n16307__ = ~new_new_n16266__ & new_new_n16305__;
  assign new_new_n16308__ = ~new_new_n16306__ & ~new_new_n16307__;
  assign new_new_n16309__ = ~new_new_n16093__ & ~new_new_n16124__;
  assign new_new_n16310__ = ~new_new_n16125__ & ~new_new_n16309__;
  assign new_new_n16311__ = new_new_n16308__ & ~new_new_n16310__;
  assign new_new_n16312__ = ~new_new_n16308__ & new_new_n16310__;
  assign new_new_n16313__ = ~new_new_n16311__ & ~new_new_n16312__;
  assign new_new_n16314__ = new_new_n16264__ & ~new_new_n16313__;
  assign new_new_n16315__ = ~new_new_n16264__ & new_new_n16313__;
  assign new_new_n16316__ = ~new_new_n16314__ & ~new_new_n16315__;
  assign new_new_n16317__ = new_new_n16179__ & new_new_n16316__;
  assign new_new_n16318__ = ~new_new_n16179__ & ~new_new_n16316__;
  assign new_new_n16319__ = ~new_new_n16317__ & ~new_new_n16318__;
  assign new_new_n16320__ = ~new_new_n16080__ & ~new_new_n16083__;
  assign new_new_n16321__ = ~new_new_n16079__ & ~new_new_n16320__;
  assign new_new_n16322__ = new_new_n16319__ & ~new_new_n16321__;
  assign new_new_n16323__ = ~new_new_n16319__ & new_new_n16321__;
  assign new_new_n16324__ = ~new_new_n16322__ & ~new_new_n16323__;
  assign new_new_n16325__ = new_new_n16156__ & new_new_n16324__;
  assign new_new_n16326__ = ~new_new_n16156__ & ~new_new_n16324__;
  assign new_new_n16327__ = ~new_new_n16325__ & ~new_new_n16326__;
  assign new_new_n16328__ = ~new_new_n16137__ & new_new_n16327__;
  assign new_new_n16329__ = new_new_n16137__ & ~new_new_n16327__;
  assign new_new_n16330__ = ~new_new_n16328__ & ~new_new_n16329__;
  assign new_new_n16331__ = ~new_new_n15931__ & ~new_new_n16132__;
  assign new_new_n16332__ = ~new_new_n15932__ & ~new_new_n16331__;
  assign new_new_n16333__ = new_new_n16330__ & ~new_new_n16332__;
  assign new_new_n16334__ = ~new_new_n16330__ & new_new_n16332__;
  assign po089 = ~new_new_n16333__ & ~new_new_n16334__;
  assign new_new_n16336__ = ~new_new_n16328__ & ~new_new_n16332__;
  assign new_new_n16337__ = ~new_new_n16329__ & ~new_new_n16336__;
  assign new_new_n16338__ = ~new_new_n16139__ & ~new_new_n16179__;
  assign new_new_n16339__ = new_new_n16139__ & new_new_n16179__;
  assign new_new_n16340__ = ~new_new_n16338__ & ~new_new_n16339__;
  assign new_new_n16341__ = new_new_n16321__ & new_new_n16340__;
  assign new_new_n16342__ = ~new_new_n16321__ & ~new_new_n16340__;
  assign new_new_n16343__ = new_new_n16153__ & new_new_n16316__;
  assign new_new_n16344__ = ~new_new_n16153__ & ~new_new_n16316__;
  assign new_new_n16345__ = ~new_new_n16342__ & ~new_new_n16343__;
  assign new_new_n16346__ = ~new_new_n16344__ & new_new_n16345__;
  assign new_new_n16347__ = ~new_new_n16341__ & ~new_new_n16346__;
  assign new_new_n16348__ = new_new_n16337__ & ~new_new_n16347__;
  assign new_new_n16349__ = ~new_new_n16337__ & new_new_n16347__;
  assign new_new_n16350__ = ~new_new_n16348__ & ~new_new_n16349__;
  assign new_new_n16351__ = ~new_new_n16167__ & new_new_n16179__;
  assign new_new_n16352__ = ~new_new_n16338__ & ~new_new_n16351__;
  assign new_new_n16353__ = ~new_new_n16238__ & ~new_new_n16242__;
  assign new_new_n16354__ = ~new_new_n16241__ & ~new_new_n16353__;
  assign new_new_n16355__ = ~new_new_n16204__ & ~new_new_n16207__;
  assign new_new_n16356__ = ~new_new_n16206__ & ~new_new_n16355__;
  assign new_new_n16357__ = ~new_new_n16354__ & ~new_new_n16356__;
  assign new_new_n16358__ = new_new_n16354__ & new_new_n16356__;
  assign new_new_n16359__ = ~new_new_n16357__ & ~new_new_n16358__;
  assign new_new_n16360__ = ~new_new_n16229__ & ~new_new_n16233__;
  assign new_new_n16361__ = ~new_new_n16232__ & ~new_new_n16360__;
  assign new_new_n16362__ = ~new_new_n16359__ & new_new_n16361__;
  assign new_new_n16363__ = new_new_n16359__ & ~new_new_n16361__;
  assign new_new_n16364__ = ~new_new_n16362__ & ~new_new_n16363__;
  assign new_new_n16365__ = pi32 & pi57;
  assign new_new_n16366__ = pi31 & pi58;
  assign new_new_n16367__ = pi30 & pi59;
  assign new_new_n16368__ = ~new_new_n16366__ & ~new_new_n16367__;
  assign new_new_n16369__ = new_new_n16366__ & new_new_n16367__;
  assign new_new_n16370__ = ~new_new_n16368__ & ~new_new_n16369__;
  assign new_new_n16371__ = new_new_n16365__ & ~new_new_n16370__;
  assign new_new_n16372__ = ~new_new_n16365__ & new_new_n16370__;
  assign new_new_n16373__ = ~new_new_n16371__ & ~new_new_n16372__;
  assign new_new_n16374__ = pi38 & pi51;
  assign new_new_n16375__ = pi37 & pi52;
  assign new_new_n16376__ = pi36 & pi53;
  assign new_new_n16377__ = ~new_new_n16375__ & ~new_new_n16376__;
  assign new_new_n16378__ = new_new_n16375__ & new_new_n16376__;
  assign new_new_n16379__ = ~new_new_n16377__ & ~new_new_n16378__;
  assign new_new_n16380__ = new_new_n16374__ & ~new_new_n16379__;
  assign new_new_n16381__ = ~new_new_n16374__ & new_new_n16379__;
  assign new_new_n16382__ = ~new_new_n16380__ & ~new_new_n16381__;
  assign new_new_n16383__ = new_new_n16373__ & new_new_n16382__;
  assign new_new_n16384__ = ~new_new_n16373__ & ~new_new_n16382__;
  assign new_new_n16385__ = ~new_new_n16383__ & ~new_new_n16384__;
  assign new_new_n16386__ = pi41 & pi48;
  assign new_new_n16387__ = pi33 & pi56;
  assign new_new_n16388__ = pi35 & pi54;
  assign new_new_n16389__ = ~new_new_n16387__ & ~new_new_n16388__;
  assign new_new_n16390__ = new_new_n16387__ & new_new_n16388__;
  assign new_new_n16391__ = ~new_new_n16389__ & ~new_new_n16390__;
  assign new_new_n16392__ = new_new_n16386__ & ~new_new_n16391__;
  assign new_new_n16393__ = ~new_new_n16386__ & new_new_n16391__;
  assign new_new_n16394__ = ~new_new_n16392__ & ~new_new_n16393__;
  assign new_new_n16395__ = new_new_n16385__ & ~new_new_n16394__;
  assign new_new_n16396__ = ~new_new_n16385__ & new_new_n16394__;
  assign new_new_n16397__ = ~new_new_n16395__ & ~new_new_n16396__;
  assign new_new_n16398__ = ~new_new_n16283__ & ~new_new_n16287__;
  assign new_new_n16399__ = ~new_new_n16286__ & ~new_new_n16398__;
  assign new_new_n16400__ = pi29 & pi60;
  assign new_new_n16401__ = pi28 & pi61;
  assign new_new_n16402__ = ~new_new_n16400__ & ~new_new_n16401__;
  assign new_new_n16403__ = new_new_n16400__ & new_new_n16401__;
  assign new_new_n16404__ = ~new_new_n16402__ & ~new_new_n16403__;
  assign new_new_n16405__ = new_new_n16399__ & ~new_new_n16404__;
  assign new_new_n16406__ = ~new_new_n16399__ & new_new_n16404__;
  assign new_new_n16407__ = ~new_new_n16405__ & ~new_new_n16406__;
  assign new_new_n16408__ = pi43 & pi46;
  assign new_new_n16409__ = pi34 & pi55;
  assign new_new_n16410__ = pi42 & pi47;
  assign new_new_n16411__ = ~new_new_n16409__ & ~new_new_n16410__;
  assign new_new_n16412__ = new_new_n16409__ & new_new_n16410__;
  assign new_new_n16413__ = ~new_new_n16411__ & ~new_new_n16412__;
  assign new_new_n16414__ = new_new_n16408__ & ~new_new_n16413__;
  assign new_new_n16415__ = ~new_new_n16408__ & new_new_n16413__;
  assign new_new_n16416__ = ~new_new_n16414__ & ~new_new_n16415__;
  assign new_new_n16417__ = new_new_n16407__ & new_new_n16416__;
  assign new_new_n16418__ = ~new_new_n16407__ & ~new_new_n16416__;
  assign new_new_n16419__ = ~new_new_n16417__ & ~new_new_n16418__;
  assign new_new_n16420__ = pi27 & pi62;
  assign new_new_n16421__ = ~pi44 & pi45;
  assign new_new_n16422__ = new_new_n16420__ & ~new_new_n16421__;
  assign new_new_n16423__ = ~new_new_n16420__ & new_new_n16421__;
  assign new_new_n16424__ = ~new_new_n16422__ & ~new_new_n16423__;
  assign new_new_n16425__ = ~new_new_n16419__ & new_new_n16424__;
  assign new_new_n16426__ = new_new_n16419__ & ~new_new_n16424__;
  assign new_new_n16427__ = ~new_new_n16425__ & ~new_new_n16426__;
  assign new_new_n16428__ = ~new_new_n16397__ & ~new_new_n16427__;
  assign new_new_n16429__ = new_new_n16397__ & new_new_n16427__;
  assign new_new_n16430__ = ~new_new_n16428__ & ~new_new_n16429__;
  assign new_new_n16431__ = new_new_n16364__ & new_new_n16430__;
  assign new_new_n16432__ = ~new_new_n16364__ & ~new_new_n16430__;
  assign new_new_n16433__ = ~new_new_n16431__ & ~new_new_n16432__;
  assign new_new_n16434__ = new_new_n16352__ & ~new_new_n16433__;
  assign new_new_n16435__ = ~new_new_n16352__ & new_new_n16433__;
  assign new_new_n16436__ = ~new_new_n16434__ & ~new_new_n16435__;
  assign new_new_n16437__ = ~new_new_n16273__ & ~new_new_n16277__;
  assign new_new_n16438__ = ~pi43 & ~new_new_n15739__;
  assign new_new_n16439__ = pi44 & ~new_new_n16438__;
  assign new_new_n16440__ = new_new_n16186__ & new_new_n16439__;
  assign new_new_n16441__ = ~new_new_n16183__ & ~new_new_n16440__;
  assign new_new_n16442__ = ~new_new_n16437__ & ~new_new_n16441__;
  assign new_new_n16443__ = new_new_n16437__ & new_new_n16441__;
  assign new_new_n16444__ = ~new_new_n16442__ & ~new_new_n16443__;
  assign new_new_n16445__ = ~new_new_n16292__ & new_new_n16296__;
  assign new_new_n16446__ = ~new_new_n16293__ & ~new_new_n16445__;
  assign new_new_n16447__ = new_new_n16444__ & ~new_new_n16446__;
  assign new_new_n16448__ = ~new_new_n16444__ & new_new_n16446__;
  assign new_new_n16449__ = ~new_new_n16447__ & ~new_new_n16448__;
  assign new_new_n16450__ = ~new_new_n16161__ & ~new_new_n16164__;
  assign new_new_n16451__ = ~new_new_n16160__ & ~new_new_n16450__;
  assign new_new_n16452__ = new_new_n16449__ & ~new_new_n16451__;
  assign new_new_n16453__ = ~new_new_n16449__ & new_new_n16451__;
  assign new_new_n16454__ = ~new_new_n16452__ & ~new_new_n16453__;
  assign new_new_n16455__ = new_new_n16278__ & ~new_new_n16301__;
  assign new_new_n16456__ = ~new_new_n16300__ & ~new_new_n16455__;
  assign new_new_n16457__ = new_new_n16454__ & ~new_new_n16456__;
  assign new_new_n16458__ = ~new_new_n16454__ & new_new_n16456__;
  assign new_new_n16459__ = ~new_new_n16457__ & ~new_new_n16458__;
  assign new_new_n16460__ = new_new_n16436__ & ~new_new_n16459__;
  assign new_new_n16461__ = ~new_new_n16436__ & new_new_n16459__;
  assign new_new_n16462__ = ~new_new_n16460__ & ~new_new_n16461__;
  assign new_new_n16463__ = ~new_new_n16153__ & ~new_new_n16314__;
  assign new_new_n16464__ = ~new_new_n16315__ & ~new_new_n16463__;
  assign new_new_n16465__ = ~new_new_n16462__ & ~new_new_n16464__;
  assign new_new_n16466__ = new_new_n16462__ & new_new_n16464__;
  assign new_new_n16467__ = ~new_new_n16465__ & ~new_new_n16466__;
  assign new_new_n16468__ = ~new_new_n16212__ & ~new_new_n16215__;
  assign new_new_n16469__ = ~new_new_n16214__ & ~new_new_n16468__;
  assign new_new_n16470__ = ~new_new_n16250__ & ~new_new_n16254__;
  assign new_new_n16471__ = ~new_new_n16253__ & ~new_new_n16470__;
  assign new_new_n16472__ = pi40 & pi49;
  assign new_new_n16473__ = pi26 & pi63;
  assign new_new_n16474__ = pi39 & pi50;
  assign new_new_n16475__ = ~new_new_n16473__ & ~new_new_n16474__;
  assign new_new_n16476__ = new_new_n16473__ & new_new_n16474__;
  assign new_new_n16477__ = ~new_new_n16475__ & ~new_new_n16476__;
  assign new_new_n16478__ = new_new_n16472__ & ~new_new_n16477__;
  assign new_new_n16479__ = ~new_new_n16472__ & new_new_n16477__;
  assign new_new_n16480__ = ~new_new_n16478__ & ~new_new_n16479__;
  assign new_new_n16481__ = ~new_new_n16471__ & ~new_new_n16480__;
  assign new_new_n16482__ = new_new_n16471__ & new_new_n16480__;
  assign new_new_n16483__ = ~new_new_n16481__ & ~new_new_n16482__;
  assign new_new_n16484__ = new_new_n16469__ & new_new_n16483__;
  assign new_new_n16485__ = ~new_new_n16469__ & ~new_new_n16483__;
  assign new_new_n16486__ = ~new_new_n16484__ & ~new_new_n16485__;
  assign new_new_n16487__ = ~new_new_n16307__ & ~new_new_n16310__;
  assign new_new_n16488__ = ~new_new_n16306__ & ~new_new_n16487__;
  assign new_new_n16489__ = ~new_new_n16247__ & ~new_new_n16258__;
  assign new_new_n16490__ = ~new_new_n16248__ & ~new_new_n16489__;
  assign new_new_n16491__ = new_new_n16203__ & ~new_new_n16220__;
  assign new_new_n16492__ = ~new_new_n16221__ & ~new_new_n16491__;
  assign new_new_n16493__ = new_new_n16490__ & new_new_n16492__;
  assign new_new_n16494__ = ~new_new_n16490__ & ~new_new_n16492__;
  assign new_new_n16495__ = ~new_new_n16493__ & ~new_new_n16494__;
  assign new_new_n16496__ = ~new_new_n16227__ & new_new_n16261__;
  assign new_new_n16497__ = ~new_new_n16226__ & ~new_new_n16496__;
  assign new_new_n16498__ = ~new_new_n16495__ & new_new_n16497__;
  assign new_new_n16499__ = new_new_n16495__ & ~new_new_n16497__;
  assign new_new_n16500__ = ~new_new_n16498__ & ~new_new_n16499__;
  assign new_new_n16501__ = new_new_n16488__ & ~new_new_n16500__;
  assign new_new_n16502__ = ~new_new_n16488__ & new_new_n16500__;
  assign new_new_n16503__ = ~new_new_n16501__ & ~new_new_n16502__;
  assign new_new_n16504__ = new_new_n16486__ & new_new_n16503__;
  assign new_new_n16505__ = ~new_new_n16486__ & ~new_new_n16503__;
  assign new_new_n16506__ = ~new_new_n16504__ & ~new_new_n16505__;
  assign new_new_n16507__ = new_new_n16467__ & ~new_new_n16506__;
  assign new_new_n16508__ = ~new_new_n16467__ & new_new_n16506__;
  assign new_new_n16509__ = ~new_new_n16507__ & ~new_new_n16508__;
  assign new_new_n16510__ = new_new_n16350__ & ~new_new_n16509__;
  assign new_new_n16511__ = ~new_new_n16350__ & new_new_n16509__;
  assign po090 = new_new_n16510__ | new_new_n16511__;
  assign new_new_n16513__ = ~new_new_n16466__ & ~new_new_n16506__;
  assign new_new_n16514__ = ~new_new_n16465__ & ~new_new_n16513__;
  assign new_new_n16515__ = ~new_new_n16349__ & ~new_new_n16509__;
  assign new_new_n16516__ = ~new_new_n16348__ & ~new_new_n16515__;
  assign new_new_n16517__ = ~new_new_n16514__ & new_new_n16516__;
  assign new_new_n16518__ = new_new_n16514__ & ~new_new_n16516__;
  assign new_new_n16519__ = ~new_new_n16517__ & ~new_new_n16518__;
  assign new_new_n16520__ = new_new_n16364__ & ~new_new_n16429__;
  assign new_new_n16521__ = ~new_new_n16428__ & ~new_new_n16520__;
  assign new_new_n16522__ = ~pi44 & ~new_new_n16420__;
  assign new_new_n16523__ = pi45 & ~new_new_n16522__;
  assign new_new_n16524__ = ~new_new_n16408__ & ~new_new_n16412__;
  assign new_new_n16525__ = ~new_new_n16411__ & ~new_new_n16524__;
  assign new_new_n16526__ = ~new_new_n16386__ & ~new_new_n16390__;
  assign new_new_n16527__ = ~new_new_n16389__ & ~new_new_n16526__;
  assign new_new_n16528__ = new_new_n16525__ & new_new_n16527__;
  assign new_new_n16529__ = ~new_new_n16525__ & ~new_new_n16527__;
  assign new_new_n16530__ = ~new_new_n16528__ & ~new_new_n16529__;
  assign new_new_n16531__ = new_new_n16523__ & ~new_new_n16530__;
  assign new_new_n16532__ = ~new_new_n16523__ & new_new_n16530__;
  assign new_new_n16533__ = ~new_new_n16531__ & ~new_new_n16532__;
  assign new_new_n16534__ = ~new_new_n16418__ & new_new_n16424__;
  assign new_new_n16535__ = ~new_new_n16417__ & ~new_new_n16534__;
  assign new_new_n16536__ = ~new_new_n16533__ & new_new_n16535__;
  assign new_new_n16537__ = new_new_n16533__ & ~new_new_n16535__;
  assign new_new_n16538__ = ~new_new_n16536__ & ~new_new_n16537__;
  assign new_new_n16539__ = ~new_new_n16383__ & ~new_new_n16394__;
  assign new_new_n16540__ = ~new_new_n16384__ & ~new_new_n16539__;
  assign new_new_n16541__ = new_new_n16538__ & ~new_new_n16540__;
  assign new_new_n16542__ = ~new_new_n16538__ & new_new_n16540__;
  assign new_new_n16543__ = ~new_new_n16541__ & ~new_new_n16542__;
  assign new_new_n16544__ = new_new_n16521__ & new_new_n16543__;
  assign new_new_n16545__ = ~new_new_n16521__ & ~new_new_n16543__;
  assign new_new_n16546__ = ~new_new_n16544__ & ~new_new_n16545__;
  assign new_new_n16547__ = ~new_new_n16453__ & ~new_new_n16456__;
  assign new_new_n16548__ = ~new_new_n16452__ & ~new_new_n16547__;
  assign new_new_n16549__ = new_new_n16546__ & ~new_new_n16548__;
  assign new_new_n16550__ = ~new_new_n16546__ & new_new_n16548__;
  assign new_new_n16551__ = ~new_new_n16549__ & ~new_new_n16550__;
  assign new_new_n16552__ = ~new_new_n16358__ & ~new_new_n16361__;
  assign new_new_n16553__ = ~new_new_n16357__ & ~new_new_n16552__;
  assign new_new_n16554__ = new_new_n16469__ & ~new_new_n16480__;
  assign new_new_n16555__ = ~new_new_n16469__ & new_new_n16480__;
  assign new_new_n16556__ = new_new_n16471__ & ~new_new_n16555__;
  assign new_new_n16557__ = ~new_new_n16554__ & ~new_new_n16556__;
  assign new_new_n16558__ = pi41 & pi49;
  assign new_new_n16559__ = pi40 & pi50;
  assign new_new_n16560__ = pi39 & pi51;
  assign new_new_n16561__ = ~new_new_n16559__ & ~new_new_n16560__;
  assign new_new_n16562__ = new_new_n16559__ & new_new_n16560__;
  assign new_new_n16563__ = ~new_new_n16561__ & ~new_new_n16562__;
  assign new_new_n16564__ = new_new_n16558__ & ~new_new_n16563__;
  assign new_new_n16565__ = ~new_new_n16558__ & new_new_n16563__;
  assign new_new_n16566__ = ~new_new_n16564__ & ~new_new_n16565__;
  assign new_new_n16567__ = ~new_new_n16557__ & ~new_new_n16566__;
  assign new_new_n16568__ = new_new_n16557__ & new_new_n16566__;
  assign new_new_n16569__ = ~new_new_n16567__ & ~new_new_n16568__;
  assign new_new_n16570__ = new_new_n16553__ & new_new_n16569__;
  assign new_new_n16571__ = ~new_new_n16553__ & ~new_new_n16569__;
  assign new_new_n16572__ = ~new_new_n16570__ & ~new_new_n16571__;
  assign new_new_n16573__ = ~new_new_n16486__ & ~new_new_n16493__;
  assign new_new_n16574__ = ~new_new_n16494__ & ~new_new_n16573__;
  assign new_new_n16575__ = ~new_new_n16572__ & new_new_n16574__;
  assign new_new_n16576__ = new_new_n16572__ & ~new_new_n16574__;
  assign new_new_n16577__ = ~new_new_n16575__ & ~new_new_n16576__;
  assign new_new_n16578__ = pi32 & pi58;
  assign new_new_n16579__ = pi31 & pi59;
  assign new_new_n16580__ = pi30 & pi60;
  assign new_new_n16581__ = ~new_new_n16579__ & ~new_new_n16580__;
  assign new_new_n16582__ = new_new_n16579__ & new_new_n16580__;
  assign new_new_n16583__ = ~new_new_n16581__ & ~new_new_n16582__;
  assign new_new_n16584__ = new_new_n16578__ & ~new_new_n16583__;
  assign new_new_n16585__ = ~new_new_n16578__ & new_new_n16583__;
  assign new_new_n16586__ = ~new_new_n16584__ & ~new_new_n16585__;
  assign new_new_n16587__ = ~new_new_n16399__ & ~new_new_n16403__;
  assign new_new_n16588__ = ~new_new_n16402__ & ~new_new_n16587__;
  assign new_new_n16589__ = pi29 & pi61;
  assign new_new_n16590__ = pi27 & pi63;
  assign new_new_n16591__ = pi28 & pi62;
  assign new_new_n16592__ = ~new_new_n16590__ & ~new_new_n16591__;
  assign new_new_n16593__ = new_new_n16590__ & new_new_n16591__;
  assign new_new_n16594__ = ~new_new_n16592__ & ~new_new_n16593__;
  assign new_new_n16595__ = new_new_n16589__ & ~new_new_n16594__;
  assign new_new_n16596__ = ~new_new_n16589__ & new_new_n16594__;
  assign new_new_n16597__ = ~new_new_n16595__ & ~new_new_n16596__;
  assign new_new_n16598__ = ~new_new_n16588__ & new_new_n16597__;
  assign new_new_n16599__ = new_new_n16588__ & ~new_new_n16597__;
  assign new_new_n16600__ = ~new_new_n16586__ & ~new_new_n16598__;
  assign new_new_n16601__ = ~new_new_n16599__ & ~new_new_n16600__;
  assign new_new_n16602__ = ~new_new_n16598__ & new_new_n16601__;
  assign new_new_n16603__ = new_new_n16586__ & ~new_new_n16602__;
  assign new_new_n16604__ = ~new_new_n16599__ & new_new_n16600__;
  assign new_new_n16605__ = ~new_new_n16603__ & ~new_new_n16604__;
  assign new_new_n16606__ = new_new_n16577__ & ~new_new_n16605__;
  assign new_new_n16607__ = ~new_new_n16577__ & new_new_n16605__;
  assign new_new_n16608__ = ~new_new_n16606__ & ~new_new_n16607__;
  assign new_new_n16609__ = ~new_new_n16435__ & new_new_n16459__;
  assign new_new_n16610__ = ~new_new_n16434__ & ~new_new_n16609__;
  assign new_new_n16611__ = new_new_n16608__ & new_new_n16610__;
  assign new_new_n16612__ = ~new_new_n16608__ & ~new_new_n16610__;
  assign new_new_n16613__ = ~new_new_n16611__ & ~new_new_n16612__;
  assign new_new_n16614__ = ~new_new_n16365__ & ~new_new_n16369__;
  assign new_new_n16615__ = ~new_new_n16368__ & ~new_new_n16614__;
  assign new_new_n16616__ = ~new_new_n16472__ & ~new_new_n16476__;
  assign new_new_n16617__ = ~new_new_n16475__ & ~new_new_n16616__;
  assign new_new_n16618__ = ~new_new_n16615__ & ~new_new_n16617__;
  assign new_new_n16619__ = new_new_n16615__ & new_new_n16617__;
  assign new_new_n16620__ = ~new_new_n16618__ & ~new_new_n16619__;
  assign new_new_n16621__ = ~new_new_n16374__ & ~new_new_n16378__;
  assign new_new_n16622__ = ~new_new_n16377__ & ~new_new_n16621__;
  assign new_new_n16623__ = ~new_new_n16620__ & new_new_n16622__;
  assign new_new_n16624__ = ~new_new_n16619__ & ~new_new_n16622__;
  assign new_new_n16625__ = ~new_new_n16618__ & new_new_n16624__;
  assign new_new_n16626__ = ~new_new_n16623__ & ~new_new_n16625__;
  assign new_new_n16627__ = ~new_new_n16442__ & ~new_new_n16447__;
  assign new_new_n16628__ = pi35 & pi55;
  assign new_new_n16629__ = pi33 & pi57;
  assign new_new_n16630__ = pi34 & pi56;
  assign new_new_n16631__ = ~new_new_n16629__ & ~new_new_n16630__;
  assign new_new_n16632__ = new_new_n16629__ & new_new_n16630__;
  assign new_new_n16633__ = ~new_new_n16631__ & ~new_new_n16632__;
  assign new_new_n16634__ = new_new_n16628__ & ~new_new_n16633__;
  assign new_new_n16635__ = ~new_new_n16628__ & new_new_n16633__;
  assign new_new_n16636__ = ~new_new_n16634__ & ~new_new_n16635__;
  assign new_new_n16637__ = pi38 & pi52;
  assign new_new_n16638__ = pi37 & pi53;
  assign new_new_n16639__ = pi36 & pi54;
  assign new_new_n16640__ = ~new_new_n16638__ & ~new_new_n16639__;
  assign new_new_n16641__ = new_new_n16638__ & new_new_n16639__;
  assign new_new_n16642__ = ~new_new_n16640__ & ~new_new_n16641__;
  assign new_new_n16643__ = new_new_n16637__ & ~new_new_n16642__;
  assign new_new_n16644__ = ~new_new_n16637__ & new_new_n16642__;
  assign new_new_n16645__ = ~new_new_n16643__ & ~new_new_n16644__;
  assign new_new_n16646__ = new_new_n16636__ & new_new_n16645__;
  assign new_new_n16647__ = ~new_new_n16636__ & ~new_new_n16645__;
  assign new_new_n16648__ = ~new_new_n16646__ & ~new_new_n16647__;
  assign new_new_n16649__ = pi44 & pi46;
  assign new_new_n16650__ = pi43 & pi47;
  assign new_new_n16651__ = pi42 & pi48;
  assign new_new_n16652__ = ~new_new_n16650__ & ~new_new_n16651__;
  assign new_new_n16653__ = new_new_n16650__ & new_new_n16651__;
  assign new_new_n16654__ = ~new_new_n16652__ & ~new_new_n16653__;
  assign new_new_n16655__ = new_new_n16649__ & ~new_new_n16654__;
  assign new_new_n16656__ = ~new_new_n16649__ & new_new_n16654__;
  assign new_new_n16657__ = ~new_new_n16655__ & ~new_new_n16656__;
  assign new_new_n16658__ = new_new_n16648__ & ~new_new_n16657__;
  assign new_new_n16659__ = ~new_new_n16648__ & new_new_n16657__;
  assign new_new_n16660__ = ~new_new_n16658__ & ~new_new_n16659__;
  assign new_new_n16661__ = ~new_new_n16627__ & new_new_n16660__;
  assign new_new_n16662__ = new_new_n16627__ & ~new_new_n16660__;
  assign new_new_n16663__ = ~new_new_n16661__ & ~new_new_n16662__;
  assign new_new_n16664__ = ~new_new_n16626__ & new_new_n16663__;
  assign new_new_n16665__ = new_new_n16626__ & ~new_new_n16663__;
  assign new_new_n16666__ = ~new_new_n16664__ & ~new_new_n16665__;
  assign new_new_n16667__ = new_new_n16488__ & new_new_n16497__;
  assign new_new_n16668__ = ~new_new_n16488__ & ~new_new_n16497__;
  assign new_new_n16669__ = new_new_n16469__ & ~new_new_n16495__;
  assign new_new_n16670__ = ~new_new_n16469__ & new_new_n16495__;
  assign new_new_n16671__ = ~new_new_n16669__ & ~new_new_n16670__;
  assign new_new_n16672__ = new_new_n16483__ & new_new_n16671__;
  assign new_new_n16673__ = ~new_new_n16483__ & ~new_new_n16671__;
  assign new_new_n16674__ = ~new_new_n16672__ & ~new_new_n16673__;
  assign new_new_n16675__ = ~new_new_n16668__ & ~new_new_n16674__;
  assign new_new_n16676__ = ~new_new_n16667__ & ~new_new_n16675__;
  assign new_new_n16677__ = ~new_new_n16666__ & ~new_new_n16676__;
  assign new_new_n16678__ = new_new_n16666__ & new_new_n16676__;
  assign new_new_n16679__ = ~new_new_n16677__ & ~new_new_n16678__;
  assign new_new_n16680__ = new_new_n16613__ & ~new_new_n16679__;
  assign new_new_n16681__ = ~new_new_n16613__ & new_new_n16679__;
  assign new_new_n16682__ = ~new_new_n16680__ & ~new_new_n16681__;
  assign new_new_n16683__ = new_new_n16551__ & new_new_n16682__;
  assign new_new_n16684__ = ~new_new_n16551__ & ~new_new_n16682__;
  assign new_new_n16685__ = ~new_new_n16683__ & ~new_new_n16684__;
  assign new_new_n16686__ = new_new_n16519__ & new_new_n16685__;
  assign new_new_n16687__ = ~new_new_n16519__ & ~new_new_n16685__;
  assign po091 = new_new_n16686__ | new_new_n16687__;
  assign new_new_n16689__ = ~new_new_n16646__ & ~new_new_n16657__;
  assign new_new_n16690__ = ~new_new_n16647__ & ~new_new_n16689__;
  assign new_new_n16691__ = new_new_n16601__ & new_new_n16690__;
  assign new_new_n16692__ = ~new_new_n16601__ & ~new_new_n16690__;
  assign new_new_n16693__ = ~new_new_n16691__ & ~new_new_n16692__;
  assign new_new_n16694__ = ~new_new_n16628__ & ~new_new_n16632__;
  assign new_new_n16695__ = ~new_new_n16631__ & ~new_new_n16694__;
  assign new_new_n16696__ = ~new_new_n16649__ & ~new_new_n16653__;
  assign new_new_n16697__ = ~new_new_n16652__ & ~new_new_n16696__;
  assign new_new_n16698__ = new_new_n9881__ & new_new_n16697__;
  assign new_new_n16699__ = ~new_new_n9881__ & ~new_new_n16697__;
  assign new_new_n16700__ = ~new_new_n16698__ & ~new_new_n16699__;
  assign new_new_n16701__ = new_new_n16695__ & ~new_new_n16700__;
  assign new_new_n16702__ = ~new_new_n16695__ & new_new_n16700__;
  assign new_new_n16703__ = ~new_new_n16701__ & ~new_new_n16702__;
  assign new_new_n16704__ = new_new_n16693__ & ~new_new_n16703__;
  assign new_new_n16705__ = ~new_new_n16693__ & new_new_n16703__;
  assign new_new_n16706__ = ~new_new_n16704__ & ~new_new_n16705__;
  assign new_new_n16707__ = ~new_new_n16576__ & ~new_new_n16605__;
  assign new_new_n16708__ = ~new_new_n16575__ & ~new_new_n16707__;
  assign new_new_n16709__ = new_new_n16706__ & new_new_n16708__;
  assign new_new_n16710__ = new_new_n16626__ & ~new_new_n16661__;
  assign new_new_n16711__ = ~new_new_n16706__ & ~new_new_n16708__;
  assign new_new_n16712__ = ~new_new_n16662__ & ~new_new_n16710__;
  assign new_new_n16713__ = ~new_new_n16711__ & new_new_n16712__;
  assign new_new_n16714__ = ~new_new_n16709__ & new_new_n16713__;
  assign new_new_n16715__ = new_new_n16626__ & new_new_n16711__;
  assign new_new_n16716__ = ~new_new_n16660__ & new_new_n16709__;
  assign new_new_n16717__ = ~new_new_n16715__ & ~new_new_n16716__;
  assign new_new_n16718__ = new_new_n16627__ & ~new_new_n16717__;
  assign new_new_n16719__ = ~new_new_n16660__ & new_new_n16711__;
  assign new_new_n16720__ = new_new_n16663__ & new_new_n16709__;
  assign new_new_n16721__ = ~new_new_n16719__ & ~new_new_n16720__;
  assign new_new_n16722__ = new_new_n16666__ & ~new_new_n16721__;
  assign new_new_n16723__ = ~new_new_n16714__ & ~new_new_n16718__;
  assign new_new_n16724__ = ~new_new_n16722__ & new_new_n16723__;
  assign new_new_n16725__ = new_new_n16608__ & ~new_new_n16678__;
  assign new_new_n16726__ = ~new_new_n16677__ & ~new_new_n16725__;
  assign new_new_n16727__ = ~new_new_n16589__ & ~new_new_n16593__;
  assign new_new_n16728__ = ~new_new_n16592__ & ~new_new_n16727__;
  assign new_new_n16729__ = ~new_new_n16578__ & ~new_new_n16582__;
  assign new_new_n16730__ = ~new_new_n16581__ & ~new_new_n16729__;
  assign new_new_n16731__ = ~new_new_n16728__ & ~new_new_n16730__;
  assign new_new_n16732__ = new_new_n16728__ & new_new_n16730__;
  assign new_new_n16733__ = ~new_new_n16731__ & ~new_new_n16732__;
  assign new_new_n16734__ = ~new_new_n16637__ & ~new_new_n16641__;
  assign new_new_n16735__ = ~new_new_n16640__ & ~new_new_n16734__;
  assign new_new_n16736__ = ~new_new_n16733__ & new_new_n16735__;
  assign new_new_n16737__ = ~new_new_n16732__ & ~new_new_n16735__;
  assign new_new_n16738__ = ~new_new_n16731__ & new_new_n16737__;
  assign new_new_n16739__ = ~new_new_n16736__ & ~new_new_n16738__;
  assign new_new_n16740__ = new_new_n16553__ & ~new_new_n16568__;
  assign new_new_n16741__ = ~new_new_n16567__ & ~new_new_n16740__;
  assign new_new_n16742__ = pi29 & pi62;
  assign new_new_n16743__ = ~pi45 & pi46;
  assign new_new_n16744__ = ~new_new_n16742__ & new_new_n16743__;
  assign new_new_n16745__ = new_new_n16742__ & ~new_new_n16743__;
  assign new_new_n16746__ = ~new_new_n16744__ & ~new_new_n16745__;
  assign new_new_n16747__ = pi41 & pi50;
  assign new_new_n16748__ = pi28 & pi63;
  assign new_new_n16749__ = pi40 & pi51;
  assign new_new_n16750__ = ~new_new_n16748__ & ~new_new_n16749__;
  assign new_new_n16751__ = new_new_n16748__ & new_new_n16749__;
  assign new_new_n16752__ = ~new_new_n16750__ & ~new_new_n16751__;
  assign new_new_n16753__ = new_new_n16747__ & ~new_new_n16752__;
  assign new_new_n16754__ = ~new_new_n16747__ & new_new_n16752__;
  assign new_new_n16755__ = ~new_new_n16753__ & ~new_new_n16754__;
  assign new_new_n16756__ = pi44 & pi47;
  assign new_new_n16757__ = pi35 & pi56;
  assign new_new_n16758__ = pi43 & pi48;
  assign new_new_n16759__ = ~new_new_n16757__ & ~new_new_n16758__;
  assign new_new_n16760__ = new_new_n16757__ & new_new_n16758__;
  assign new_new_n16761__ = ~new_new_n16759__ & ~new_new_n16760__;
  assign new_new_n16762__ = new_new_n16756__ & ~new_new_n16761__;
  assign new_new_n16763__ = ~new_new_n16756__ & new_new_n16761__;
  assign new_new_n16764__ = ~new_new_n16762__ & ~new_new_n16763__;
  assign new_new_n16765__ = new_new_n16755__ & new_new_n16764__;
  assign new_new_n16766__ = ~new_new_n16755__ & ~new_new_n16764__;
  assign new_new_n16767__ = ~new_new_n16765__ & ~new_new_n16766__;
  assign new_new_n16768__ = new_new_n16746__ & new_new_n16767__;
  assign new_new_n16769__ = ~new_new_n16746__ & ~new_new_n16767__;
  assign new_new_n16770__ = ~new_new_n16768__ & ~new_new_n16769__;
  assign new_new_n16771__ = new_new_n16741__ & new_new_n16770__;
  assign new_new_n16772__ = ~new_new_n16741__ & ~new_new_n16770__;
  assign new_new_n16773__ = ~new_new_n16771__ & ~new_new_n16772__;
  assign new_new_n16774__ = ~new_new_n16739__ & new_new_n16773__;
  assign new_new_n16775__ = new_new_n16739__ & ~new_new_n16773__;
  assign new_new_n16776__ = ~new_new_n16774__ & ~new_new_n16775__;
  assign new_new_n16777__ = ~new_new_n16545__ & ~new_new_n16548__;
  assign new_new_n16778__ = ~new_new_n16544__ & ~new_new_n16777__;
  assign new_new_n16779__ = new_new_n16776__ & ~new_new_n16778__;
  assign new_new_n16780__ = ~new_new_n16776__ & new_new_n16778__;
  assign new_new_n16781__ = ~new_new_n16779__ & ~new_new_n16780__;
  assign new_new_n16782__ = ~new_new_n16536__ & new_new_n16540__;
  assign new_new_n16783__ = ~new_new_n16537__ & ~new_new_n16782__;
  assign new_new_n16784__ = ~new_new_n16523__ & ~new_new_n16528__;
  assign new_new_n16785__ = ~new_new_n16529__ & ~new_new_n16784__;
  assign new_new_n16786__ = pi42 & pi49;
  assign new_new_n16787__ = pi34 & pi57;
  assign new_new_n16788__ = pi36 & pi55;
  assign new_new_n16789__ = ~new_new_n16787__ & ~new_new_n16788__;
  assign new_new_n16790__ = new_new_n16787__ & new_new_n16788__;
  assign new_new_n16791__ = ~new_new_n16789__ & ~new_new_n16790__;
  assign new_new_n16792__ = new_new_n16786__ & ~new_new_n16791__;
  assign new_new_n16793__ = ~new_new_n16786__ & new_new_n16791__;
  assign new_new_n16794__ = ~new_new_n16792__ & ~new_new_n16793__;
  assign new_new_n16795__ = ~new_new_n16785__ & new_new_n16794__;
  assign new_new_n16796__ = new_new_n16785__ & ~new_new_n16794__;
  assign new_new_n16797__ = ~new_new_n16795__ & ~new_new_n16796__;
  assign new_new_n16798__ = ~new_new_n16618__ & ~new_new_n16624__;
  assign new_new_n16799__ = new_new_n16797__ & ~new_new_n16798__;
  assign new_new_n16800__ = ~new_new_n16797__ & new_new_n16798__;
  assign new_new_n16801__ = ~new_new_n16799__ & ~new_new_n16800__;
  assign new_new_n16802__ = new_new_n16783__ & ~new_new_n16801__;
  assign new_new_n16803__ = ~new_new_n16783__ & new_new_n16801__;
  assign new_new_n16804__ = ~new_new_n16802__ & ~new_new_n16803__;
  assign new_new_n16805__ = ~new_new_n16558__ & ~new_new_n16562__;
  assign new_new_n16806__ = ~new_new_n16561__ & ~new_new_n16805__;
  assign new_new_n16807__ = pi33 & pi58;
  assign new_new_n16808__ = pi32 & pi59;
  assign new_new_n16809__ = ~new_new_n9339__ & ~new_new_n16808__;
  assign new_new_n16810__ = new_new_n9339__ & new_new_n16808__;
  assign new_new_n16811__ = ~new_new_n16809__ & ~new_new_n16810__;
  assign new_new_n16812__ = new_new_n16807__ & ~new_new_n16811__;
  assign new_new_n16813__ = ~new_new_n16807__ & new_new_n16811__;
  assign new_new_n16814__ = ~new_new_n16812__ & ~new_new_n16813__;
  assign new_new_n16815__ = pi39 & pi52;
  assign new_new_n16816__ = pi37 & pi54;
  assign new_new_n16817__ = pi38 & pi53;
  assign new_new_n16818__ = ~new_new_n16816__ & ~new_new_n16817__;
  assign new_new_n16819__ = new_new_n16816__ & new_new_n16817__;
  assign new_new_n16820__ = ~new_new_n16818__ & ~new_new_n16819__;
  assign new_new_n16821__ = new_new_n16815__ & ~new_new_n16820__;
  assign new_new_n16822__ = ~new_new_n16815__ & new_new_n16820__;
  assign new_new_n16823__ = ~new_new_n16821__ & ~new_new_n16822__;
  assign new_new_n16824__ = new_new_n16814__ & new_new_n16823__;
  assign new_new_n16825__ = ~new_new_n16814__ & ~new_new_n16823__;
  assign new_new_n16826__ = ~new_new_n16824__ & ~new_new_n16825__;
  assign new_new_n16827__ = new_new_n16806__ & new_new_n16826__;
  assign new_new_n16828__ = ~new_new_n16806__ & ~new_new_n16826__;
  assign new_new_n16829__ = ~new_new_n16827__ & ~new_new_n16828__;
  assign new_new_n16830__ = new_new_n16804__ & ~new_new_n16829__;
  assign new_new_n16831__ = ~new_new_n16804__ & new_new_n16829__;
  assign new_new_n16832__ = ~new_new_n16830__ & ~new_new_n16831__;
  assign new_new_n16833__ = new_new_n16781__ & ~new_new_n16832__;
  assign new_new_n16834__ = ~new_new_n16781__ & new_new_n16832__;
  assign new_new_n16835__ = ~new_new_n16833__ & ~new_new_n16834__;
  assign new_new_n16836__ = new_new_n16726__ & new_new_n16835__;
  assign new_new_n16837__ = ~new_new_n16726__ & ~new_new_n16835__;
  assign new_new_n16838__ = ~new_new_n16836__ & ~new_new_n16837__;
  assign new_new_n16839__ = new_new_n16551__ & ~new_new_n16610__;
  assign new_new_n16840__ = ~new_new_n16551__ & new_new_n16610__;
  assign new_new_n16841__ = ~new_new_n16608__ & new_new_n16679__;
  assign new_new_n16842__ = new_new_n16608__ & ~new_new_n16679__;
  assign new_new_n16843__ = ~new_new_n16841__ & ~new_new_n16842__;
  assign new_new_n16844__ = ~new_new_n16840__ & new_new_n16843__;
  assign new_new_n16845__ = ~new_new_n16839__ & ~new_new_n16844__;
  assign new_new_n16846__ = ~new_new_n16517__ & new_new_n16685__;
  assign new_new_n16847__ = ~new_new_n16518__ & ~new_new_n16846__;
  assign new_new_n16848__ = ~new_new_n16845__ & new_new_n16847__;
  assign new_new_n16849__ = new_new_n16845__ & ~new_new_n16847__;
  assign new_new_n16850__ = ~new_new_n16848__ & ~new_new_n16849__;
  assign new_new_n16851__ = new_new_n16838__ & ~new_new_n16850__;
  assign new_new_n16852__ = ~new_new_n16838__ & new_new_n16850__;
  assign new_new_n16853__ = ~new_new_n16851__ & ~new_new_n16852__;
  assign new_new_n16854__ = new_new_n16724__ & new_new_n16853__;
  assign new_new_n16855__ = ~new_new_n16724__ & ~new_new_n16853__;
  assign po092 = new_new_n16854__ | new_new_n16855__;
  assign new_new_n16857__ = ~new_new_n16709__ & ~new_new_n16713__;
  assign new_new_n16858__ = ~new_new_n16803__ & new_new_n16829__;
  assign new_new_n16859__ = ~new_new_n16802__ & ~new_new_n16858__;
  assign new_new_n16860__ = ~new_new_n16857__ & ~new_new_n16859__;
  assign new_new_n16861__ = new_new_n16857__ & new_new_n16859__;
  assign new_new_n16862__ = ~new_new_n16860__ & ~new_new_n16861__;
  assign new_new_n16863__ = pi31 & pi61;
  assign new_new_n16864__ = ~pi30 & ~new_new_n16863__;
  assign new_new_n16865__ = ~pi62 & ~new_new_n16863__;
  assign new_new_n16866__ = ~new_new_n16864__ & ~new_new_n16865__;
  assign new_new_n16867__ = pi45 & ~new_new_n16866__;
  assign new_new_n16868__ = pi30 & new_new_n16863__;
  assign new_new_n16869__ = ~new_new_n16864__ & ~new_new_n16868__;
  assign new_new_n16870__ = pi29 & ~new_new_n16869__;
  assign new_new_n16871__ = new_new_n9881__ & new_new_n13473__;
  assign new_new_n16872__ = ~new_new_n16870__ & ~new_new_n16871__;
  assign new_new_n16873__ = pi62 & ~new_new_n16872__;
  assign new_new_n16874__ = ~new_new_n16867__ & ~new_new_n16873__;
  assign new_new_n16875__ = pi46 & ~new_new_n16874__;
  assign new_new_n16876__ = pi45 & pi46;
  assign new_new_n16877__ = ~new_new_n13280__ & ~new_new_n16868__;
  assign new_new_n16878__ = pi62 & ~new_new_n16877__;
  assign new_new_n16879__ = new_new_n16866__ & ~new_new_n16876__;
  assign new_new_n16880__ = ~new_new_n16878__ & new_new_n16879__;
  assign new_new_n16881__ = ~new_new_n16875__ & ~new_new_n16880__;
  assign new_new_n16882__ = pi41 & pi51;
  assign new_new_n16883__ = pi39 & pi53;
  assign new_new_n16884__ = pi40 & pi52;
  assign new_new_n16885__ = ~new_new_n16883__ & ~new_new_n16884__;
  assign new_new_n16886__ = new_new_n16883__ & new_new_n16884__;
  assign new_new_n16887__ = ~new_new_n16885__ & ~new_new_n16886__;
  assign new_new_n16888__ = new_new_n16882__ & ~new_new_n16887__;
  assign new_new_n16889__ = ~new_new_n16882__ & new_new_n16887__;
  assign new_new_n16890__ = ~new_new_n16888__ & ~new_new_n16889__;
  assign new_new_n16891__ = new_new_n16881__ & new_new_n16890__;
  assign new_new_n16892__ = ~new_new_n16881__ & ~new_new_n16890__;
  assign new_new_n16893__ = ~new_new_n16891__ & ~new_new_n16892__;
  assign new_new_n16894__ = ~new_new_n16695__ & ~new_new_n16698__;
  assign new_new_n16895__ = ~new_new_n16699__ & ~new_new_n16894__;
  assign new_new_n16896__ = new_new_n16893__ & ~new_new_n16895__;
  assign new_new_n16897__ = ~new_new_n16893__ & new_new_n16895__;
  assign new_new_n16898__ = ~new_new_n16896__ & ~new_new_n16897__;
  assign new_new_n16899__ = ~new_new_n16692__ & new_new_n16703__;
  assign new_new_n16900__ = ~new_new_n16691__ & ~new_new_n16899__;
  assign new_new_n16901__ = ~new_new_n16898__ & new_new_n16900__;
  assign new_new_n16902__ = new_new_n16898__ & ~new_new_n16900__;
  assign new_new_n16903__ = pi42 & pi50;
  assign new_new_n16904__ = pi35 & pi57;
  assign new_new_n16905__ = pi34 & pi58;
  assign new_new_n16906__ = ~new_new_n16904__ & ~new_new_n16905__;
  assign new_new_n16907__ = new_new_n16904__ & new_new_n16905__;
  assign new_new_n16908__ = ~new_new_n16906__ & ~new_new_n16907__;
  assign new_new_n16909__ = new_new_n16903__ & ~new_new_n16908__;
  assign new_new_n16910__ = ~new_new_n16903__ & new_new_n16908__;
  assign new_new_n16911__ = ~new_new_n16909__ & ~new_new_n16910__;
  assign new_new_n16912__ = pi45 & pi47;
  assign new_new_n16913__ = pi44 & pi48;
  assign new_new_n16914__ = pi43 & pi49;
  assign new_new_n16915__ = ~new_new_n16913__ & ~new_new_n16914__;
  assign new_new_n16916__ = new_new_n16913__ & new_new_n16914__;
  assign new_new_n16917__ = ~new_new_n16915__ & ~new_new_n16916__;
  assign new_new_n16918__ = new_new_n16912__ & ~new_new_n16917__;
  assign new_new_n16919__ = ~new_new_n16912__ & new_new_n16917__;
  assign new_new_n16920__ = ~new_new_n16918__ & ~new_new_n16919__;
  assign new_new_n16921__ = new_new_n16911__ & new_new_n16920__;
  assign new_new_n16922__ = ~new_new_n16911__ & ~new_new_n16920__;
  assign new_new_n16923__ = ~new_new_n16921__ & ~new_new_n16922__;
  assign new_new_n16924__ = pi36 & pi56;
  assign new_new_n16925__ = pi29 & pi63;
  assign new_new_n16926__ = pi33 & pi59;
  assign new_new_n16927__ = ~new_new_n16925__ & ~new_new_n16926__;
  assign new_new_n16928__ = new_new_n16925__ & new_new_n16926__;
  assign new_new_n16929__ = ~new_new_n16927__ & ~new_new_n16928__;
  assign new_new_n16930__ = new_new_n16924__ & ~new_new_n16929__;
  assign new_new_n16931__ = ~new_new_n16924__ & new_new_n16929__;
  assign new_new_n16932__ = ~new_new_n16930__ & ~new_new_n16931__;
  assign new_new_n16933__ = ~new_new_n16923__ & new_new_n16932__;
  assign new_new_n16934__ = new_new_n16923__ & ~new_new_n16932__;
  assign new_new_n16935__ = ~new_new_n16933__ & ~new_new_n16934__;
  assign new_new_n16936__ = ~new_new_n16901__ & ~new_new_n16935__;
  assign new_new_n16937__ = ~new_new_n16902__ & ~new_new_n16936__;
  assign new_new_n16938__ = ~new_new_n16901__ & new_new_n16937__;
  assign new_new_n16939__ = ~new_new_n16902__ & new_new_n16936__;
  assign new_new_n16940__ = ~new_new_n16935__ & ~new_new_n16939__;
  assign new_new_n16941__ = ~new_new_n16938__ & ~new_new_n16940__;
  assign new_new_n16942__ = new_new_n16862__ & ~new_new_n16941__;
  assign new_new_n16943__ = ~new_new_n16862__ & new_new_n16941__;
  assign new_new_n16944__ = ~new_new_n16942__ & ~new_new_n16943__;
  assign new_new_n16945__ = ~new_new_n16779__ & new_new_n16832__;
  assign new_new_n16946__ = ~new_new_n16780__ & ~new_new_n16945__;
  assign new_new_n16947__ = new_new_n16944__ & ~new_new_n16946__;
  assign new_new_n16948__ = ~new_new_n16944__ & new_new_n16946__;
  assign new_new_n16949__ = ~new_new_n16947__ & ~new_new_n16948__;
  assign new_new_n16950__ = ~new_new_n16739__ & ~new_new_n16771__;
  assign new_new_n16951__ = ~new_new_n16772__ & ~new_new_n16950__;
  assign new_new_n16952__ = ~new_new_n16731__ & ~new_new_n16737__;
  assign new_new_n16953__ = ~new_new_n16746__ & ~new_new_n16765__;
  assign new_new_n16954__ = ~new_new_n16766__ & ~new_new_n16953__;
  assign new_new_n16955__ = new_new_n16806__ & ~new_new_n16824__;
  assign new_new_n16956__ = ~new_new_n16825__ & ~new_new_n16955__;
  assign new_new_n16957__ = new_new_n16954__ & new_new_n16956__;
  assign new_new_n16958__ = ~new_new_n16954__ & ~new_new_n16956__;
  assign new_new_n16959__ = ~new_new_n16957__ & ~new_new_n16958__;
  assign new_new_n16960__ = new_new_n16952__ & ~new_new_n16959__;
  assign new_new_n16961__ = ~new_new_n16952__ & new_new_n16959__;
  assign new_new_n16962__ = ~new_new_n16960__ & ~new_new_n16961__;
  assign new_new_n16963__ = ~new_new_n16815__ & ~new_new_n16819__;
  assign new_new_n16964__ = ~new_new_n16818__ & ~new_new_n16963__;
  assign new_new_n16965__ = ~new_new_n16747__ & ~new_new_n16751__;
  assign new_new_n16966__ = ~new_new_n16750__ & ~new_new_n16965__;
  assign new_new_n16967__ = ~new_new_n16964__ & ~new_new_n16966__;
  assign new_new_n16968__ = new_new_n16964__ & new_new_n16966__;
  assign new_new_n16969__ = ~new_new_n16967__ & ~new_new_n16968__;
  assign new_new_n16970__ = ~new_new_n16807__ & ~new_new_n16810__;
  assign new_new_n16971__ = ~new_new_n16809__ & ~new_new_n16970__;
  assign new_new_n16972__ = ~new_new_n16969__ & new_new_n16971__;
  assign new_new_n16973__ = ~new_new_n16968__ & ~new_new_n16971__;
  assign new_new_n16974__ = ~new_new_n16967__ & new_new_n16973__;
  assign new_new_n16975__ = ~new_new_n16972__ & ~new_new_n16974__;
  assign new_new_n16976__ = ~new_new_n16795__ & new_new_n16798__;
  assign new_new_n16977__ = ~new_new_n16796__ & ~new_new_n16976__;
  assign new_new_n16978__ = ~new_new_n16975__ & ~new_new_n16977__;
  assign new_new_n16979__ = new_new_n16975__ & new_new_n16977__;
  assign new_new_n16980__ = ~new_new_n16978__ & ~new_new_n16979__;
  assign new_new_n16981__ = ~new_new_n16786__ & ~new_new_n16790__;
  assign new_new_n16982__ = ~new_new_n16789__ & ~new_new_n16981__;
  assign new_new_n16983__ = ~new_new_n16756__ & ~new_new_n16760__;
  assign new_new_n16984__ = ~new_new_n16759__ & ~new_new_n16983__;
  assign new_new_n16985__ = ~new_new_n16982__ & ~new_new_n16984__;
  assign new_new_n16986__ = new_new_n16982__ & new_new_n16984__;
  assign new_new_n16987__ = ~new_new_n16985__ & ~new_new_n16986__;
  assign new_new_n16988__ = pi38 & pi54;
  assign new_new_n16989__ = pi37 & pi55;
  assign new_new_n16990__ = pi32 & pi60;
  assign new_new_n16991__ = ~new_new_n16989__ & ~new_new_n16990__;
  assign new_new_n16992__ = new_new_n16989__ & new_new_n16990__;
  assign new_new_n16993__ = ~new_new_n16991__ & ~new_new_n16992__;
  assign new_new_n16994__ = new_new_n16988__ & ~new_new_n16993__;
  assign new_new_n16995__ = ~new_new_n16988__ & new_new_n16993__;
  assign new_new_n16996__ = ~new_new_n16994__ & ~new_new_n16995__;
  assign new_new_n16997__ = new_new_n16987__ & ~new_new_n16996__;
  assign new_new_n16998__ = ~new_new_n16987__ & new_new_n16996__;
  assign new_new_n16999__ = ~new_new_n16997__ & ~new_new_n16998__;
  assign new_new_n17000__ = new_new_n16980__ & ~new_new_n16999__;
  assign new_new_n17001__ = ~new_new_n16980__ & new_new_n16999__;
  assign new_new_n17002__ = ~new_new_n17000__ & ~new_new_n17001__;
  assign new_new_n17003__ = new_new_n16962__ & new_new_n17002__;
  assign new_new_n17004__ = ~new_new_n16962__ & ~new_new_n17002__;
  assign new_new_n17005__ = ~new_new_n17003__ & ~new_new_n17004__;
  assign new_new_n17006__ = new_new_n16951__ & new_new_n17005__;
  assign new_new_n17007__ = ~new_new_n16951__ & ~new_new_n17005__;
  assign new_new_n17008__ = ~new_new_n17006__ & ~new_new_n17007__;
  assign new_new_n17009__ = new_new_n16949__ & ~new_new_n17008__;
  assign new_new_n17010__ = ~new_new_n16949__ & new_new_n17008__;
  assign new_new_n17011__ = ~new_new_n17009__ & ~new_new_n17010__;
  assign new_new_n17012__ = ~new_new_n16724__ & ~new_new_n16836__;
  assign new_new_n17013__ = ~new_new_n16837__ & ~new_new_n17012__;
  assign new_new_n17014__ = ~new_new_n16849__ & new_new_n17013__;
  assign new_new_n17015__ = ~new_new_n16848__ & ~new_new_n17013__;
  assign new_new_n17016__ = ~new_new_n17014__ & ~new_new_n17015__;
  assign new_new_n17017__ = new_new_n16724__ & new_new_n16836__;
  assign new_new_n17018__ = ~new_new_n16724__ & new_new_n16837__;
  assign new_new_n17019__ = ~new_new_n17017__ & ~new_new_n17018__;
  assign new_new_n17020__ = new_new_n16850__ & new_new_n17019__;
  assign new_new_n17021__ = ~new_new_n17016__ & ~new_new_n17020__;
  assign new_new_n17022__ = ~new_new_n17011__ & ~new_new_n17021__;
  assign new_new_n17023__ = new_new_n16836__ & new_new_n16848__;
  assign new_new_n17024__ = new_new_n16835__ & new_new_n16848__;
  assign new_new_n17025__ = ~new_new_n16835__ & ~new_new_n16848__;
  assign new_new_n17026__ = new_new_n16726__ & ~new_new_n16849__;
  assign new_new_n17027__ = ~new_new_n17025__ & new_new_n17026__;
  assign new_new_n17028__ = ~new_new_n17024__ & ~new_new_n17027__;
  assign new_new_n17029__ = new_new_n16724__ & ~new_new_n17028__;
  assign new_new_n17030__ = ~new_new_n16836__ & new_new_n16849__;
  assign new_new_n17031__ = ~new_new_n16726__ & new_new_n17025__;
  assign new_new_n17032__ = ~new_new_n17030__ & ~new_new_n17031__;
  assign new_new_n17033__ = ~new_new_n16724__ & ~new_new_n17032__;
  assign new_new_n17034__ = new_new_n16837__ & new_new_n16849__;
  assign new_new_n17035__ = ~new_new_n17023__ & ~new_new_n17034__;
  assign new_new_n17036__ = ~new_new_n17029__ & new_new_n17035__;
  assign new_new_n17037__ = ~new_new_n17033__ & new_new_n17036__;
  assign new_new_n17038__ = new_new_n17011__ & ~new_new_n17037__;
  assign po093 = new_new_n17022__ | new_new_n17038__;
  assign new_new_n17040__ = ~new_new_n17011__ & ~new_new_n17014__;
  assign new_new_n17041__ = new_new_n16849__ & ~new_new_n17013__;
  assign new_new_n17042__ = new_new_n17011__ & ~new_new_n17018__;
  assign new_new_n17043__ = ~new_new_n17017__ & ~new_new_n17042__;
  assign new_new_n17044__ = ~new_new_n16848__ & new_new_n17043__;
  assign new_new_n17045__ = ~new_new_n17041__ & ~new_new_n17044__;
  assign new_new_n17046__ = ~new_new_n17040__ & new_new_n17045__;
  assign new_new_n17047__ = ~new_new_n16948__ & new_new_n17008__;
  assign new_new_n17048__ = ~new_new_n16947__ & ~new_new_n17047__;
  assign new_new_n17049__ = new_new_n17046__ & new_new_n17048__;
  assign new_new_n17050__ = ~new_new_n17046__ & ~new_new_n17048__;
  assign new_new_n17051__ = ~new_new_n17049__ & ~new_new_n17050__;
  assign new_new_n17052__ = ~new_new_n16967__ & ~new_new_n16973__;
  assign new_new_n17053__ = ~new_new_n16921__ & ~new_new_n16932__;
  assign new_new_n17054__ = ~new_new_n16922__ & ~new_new_n17053__;
  assign new_new_n17055__ = ~new_new_n17052__ & new_new_n17054__;
  assign new_new_n17056__ = new_new_n17052__ & ~new_new_n17054__;
  assign new_new_n17057__ = ~new_new_n17055__ & ~new_new_n17056__;
  assign new_new_n17058__ = ~new_new_n16986__ & new_new_n16996__;
  assign new_new_n17059__ = ~new_new_n16985__ & ~new_new_n17058__;
  assign new_new_n17060__ = new_new_n17057__ & new_new_n17059__;
  assign new_new_n17061__ = ~new_new_n17057__ & ~new_new_n17059__;
  assign new_new_n17062__ = ~new_new_n17060__ & ~new_new_n17061__;
  assign new_new_n17063__ = ~new_new_n16891__ & new_new_n16895__;
  assign new_new_n17064__ = ~new_new_n16892__ & ~new_new_n17063__;
  assign new_new_n17065__ = ~new_new_n16924__ & ~new_new_n16928__;
  assign new_new_n17066__ = ~new_new_n16927__ & ~new_new_n17065__;
  assign new_new_n17067__ = pi29 & ~new_new_n16864__;
  assign new_new_n17068__ = ~new_new_n13253__ & ~new_new_n17067__;
  assign new_new_n17069__ = pi46 & ~new_new_n17068__;
  assign new_new_n17070__ = ~new_new_n16868__ & ~new_new_n17069__;
  assign new_new_n17071__ = pi62 & ~new_new_n17070__;
  assign new_new_n17072__ = new_new_n16863__ & new_new_n16876__;
  assign new_new_n17073__ = ~new_new_n17071__ & ~new_new_n17072__;
  assign new_new_n17074__ = ~new_new_n16988__ & ~new_new_n16992__;
  assign new_new_n17075__ = ~new_new_n16991__ & ~new_new_n17074__;
  assign new_new_n17076__ = new_new_n17073__ & ~new_new_n17075__;
  assign new_new_n17077__ = ~new_new_n17073__ & new_new_n17075__;
  assign new_new_n17078__ = ~new_new_n17076__ & ~new_new_n17077__;
  assign new_new_n17079__ = new_new_n17066__ & new_new_n17078__;
  assign new_new_n17080__ = ~new_new_n17066__ & ~new_new_n17078__;
  assign new_new_n17081__ = ~new_new_n17079__ & ~new_new_n17080__;
  assign new_new_n17082__ = ~new_new_n17064__ & new_new_n17081__;
  assign new_new_n17083__ = new_new_n17064__ & ~new_new_n17081__;
  assign new_new_n17084__ = ~new_new_n17082__ & ~new_new_n17083__;
  assign new_new_n17085__ = ~new_new_n16912__ & ~new_new_n16916__;
  assign new_new_n17086__ = ~new_new_n16915__ & ~new_new_n17085__;
  assign new_new_n17087__ = ~new_new_n16882__ & ~new_new_n16886__;
  assign new_new_n17088__ = ~new_new_n16885__ & ~new_new_n17087__;
  assign new_new_n17089__ = ~new_new_n16903__ & ~new_new_n16907__;
  assign new_new_n17090__ = ~new_new_n16906__ & ~new_new_n17089__;
  assign new_new_n17091__ = ~new_new_n17088__ & ~new_new_n17090__;
  assign new_new_n17092__ = new_new_n17088__ & new_new_n17090__;
  assign new_new_n17093__ = ~new_new_n17091__ & ~new_new_n17092__;
  assign new_new_n17094__ = new_new_n17086__ & ~new_new_n17093__;
  assign new_new_n17095__ = ~new_new_n17086__ & new_new_n17093__;
  assign new_new_n17096__ = ~new_new_n17094__ & ~new_new_n17095__;
  assign new_new_n17097__ = new_new_n17084__ & new_new_n17096__;
  assign new_new_n17098__ = ~new_new_n17084__ & ~new_new_n17096__;
  assign new_new_n17099__ = ~new_new_n17097__ & ~new_new_n17098__;
  assign new_new_n17100__ = ~new_new_n17062__ & new_new_n17099__;
  assign new_new_n17101__ = new_new_n17062__ & ~new_new_n17099__;
  assign new_new_n17102__ = ~new_new_n17100__ & ~new_new_n17101__;
  assign new_new_n17103__ = ~new_new_n16978__ & ~new_new_n16999__;
  assign new_new_n17104__ = ~new_new_n16979__ & ~new_new_n17103__;
  assign new_new_n17105__ = new_new_n17102__ & new_new_n17104__;
  assign new_new_n17106__ = ~new_new_n17102__ & ~new_new_n17104__;
  assign new_new_n17107__ = ~new_new_n17105__ & ~new_new_n17106__;
  assign new_new_n17108__ = ~new_new_n16860__ & ~new_new_n16941__;
  assign new_new_n17109__ = ~new_new_n16861__ & ~new_new_n17108__;
  assign new_new_n17110__ = new_new_n17107__ & new_new_n17109__;
  assign new_new_n17111__ = ~new_new_n17107__ & ~new_new_n17109__;
  assign new_new_n17112__ = ~new_new_n17110__ & ~new_new_n17111__;
  assign new_new_n17113__ = ~new_new_n16951__ & ~new_new_n17003__;
  assign new_new_n17114__ = ~new_new_n17004__ & ~new_new_n17113__;
  assign new_new_n17115__ = ~new_new_n16937__ & new_new_n17114__;
  assign new_new_n17116__ = new_new_n16937__ & ~new_new_n17114__;
  assign new_new_n17117__ = ~new_new_n17115__ & ~new_new_n17116__;
  assign new_new_n17118__ = new_new_n16952__ & ~new_new_n16957__;
  assign new_new_n17119__ = ~new_new_n16958__ & ~new_new_n17118__;
  assign new_new_n17120__ = pi33 & pi60;
  assign new_new_n17121__ = pi30 & pi63;
  assign new_new_n17122__ = pi32 & pi61;
  assign new_new_n17123__ = ~new_new_n17121__ & ~new_new_n17122__;
  assign new_new_n17124__ = new_new_n17121__ & new_new_n17122__;
  assign new_new_n17125__ = ~new_new_n17123__ & ~new_new_n17124__;
  assign new_new_n17126__ = new_new_n17120__ & ~new_new_n17125__;
  assign new_new_n17127__ = ~new_new_n17120__ & new_new_n17125__;
  assign new_new_n17128__ = ~new_new_n17126__ & ~new_new_n17127__;
  assign new_new_n17129__ = pi39 & pi54;
  assign new_new_n17130__ = pi35 & pi58;
  assign new_new_n17131__ = pi36 & pi57;
  assign new_new_n17132__ = ~new_new_n17130__ & ~new_new_n17131__;
  assign new_new_n17133__ = new_new_n17130__ & new_new_n17131__;
  assign new_new_n17134__ = ~new_new_n17132__ & ~new_new_n17133__;
  assign new_new_n17135__ = new_new_n17129__ & ~new_new_n17134__;
  assign new_new_n17136__ = ~new_new_n17129__ & new_new_n17134__;
  assign new_new_n17137__ = ~new_new_n17135__ & ~new_new_n17136__;
  assign new_new_n17138__ = ~new_new_n17128__ & ~new_new_n17137__;
  assign new_new_n17139__ = new_new_n17128__ & new_new_n17137__;
  assign new_new_n17140__ = ~new_new_n17138__ & ~new_new_n17139__;
  assign new_new_n17141__ = pi41 & pi52;
  assign new_new_n17142__ = pi40 & pi53;
  assign new_new_n17143__ = pi34 & pi59;
  assign new_new_n17144__ = ~new_new_n17142__ & ~new_new_n17143__;
  assign new_new_n17145__ = new_new_n17142__ & new_new_n17143__;
  assign new_new_n17146__ = ~new_new_n17144__ & ~new_new_n17145__;
  assign new_new_n17147__ = new_new_n17141__ & ~new_new_n17146__;
  assign new_new_n17148__ = ~new_new_n17141__ & new_new_n17146__;
  assign new_new_n17149__ = ~new_new_n17147__ & ~new_new_n17148__;
  assign new_new_n17150__ = ~new_new_n17140__ & new_new_n17149__;
  assign new_new_n17151__ = new_new_n17140__ & ~new_new_n17149__;
  assign new_new_n17152__ = ~new_new_n17150__ & ~new_new_n17151__;
  assign new_new_n17153__ = new_new_n17119__ & ~new_new_n17152__;
  assign new_new_n17154__ = ~new_new_n17119__ & new_new_n17152__;
  assign new_new_n17155__ = ~new_new_n17153__ & ~new_new_n17154__;
  assign new_new_n17156__ = pi45 & pi48;
  assign new_new_n17157__ = pi38 & pi55;
  assign new_new_n17158__ = pi37 & pi56;
  assign new_new_n17159__ = ~new_new_n17157__ & ~new_new_n17158__;
  assign new_new_n17160__ = new_new_n17157__ & new_new_n17158__;
  assign new_new_n17161__ = ~new_new_n17159__ & ~new_new_n17160__;
  assign new_new_n17162__ = new_new_n17156__ & ~new_new_n17161__;
  assign new_new_n17163__ = ~new_new_n17156__ & new_new_n17161__;
  assign new_new_n17164__ = ~new_new_n17162__ & ~new_new_n17163__;
  assign new_new_n17165__ = pi44 & pi49;
  assign new_new_n17166__ = pi43 & pi50;
  assign new_new_n17167__ = pi42 & pi51;
  assign new_new_n17168__ = ~new_new_n17166__ & ~new_new_n17167__;
  assign new_new_n17169__ = new_new_n17166__ & new_new_n17167__;
  assign new_new_n17170__ = ~new_new_n17168__ & ~new_new_n17169__;
  assign new_new_n17171__ = new_new_n17165__ & ~new_new_n17170__;
  assign new_new_n17172__ = ~new_new_n17165__ & new_new_n17170__;
  assign new_new_n17173__ = ~new_new_n17171__ & ~new_new_n17172__;
  assign new_new_n17174__ = new_new_n17164__ & new_new_n17173__;
  assign new_new_n17175__ = ~new_new_n17164__ & ~new_new_n17173__;
  assign new_new_n17176__ = ~new_new_n17174__ & ~new_new_n17175__;
  assign new_new_n17177__ = pi31 & pi62;
  assign new_new_n17178__ = ~pi46 & pi47;
  assign new_new_n17179__ = new_new_n17177__ & ~new_new_n17178__;
  assign new_new_n17180__ = ~new_new_n17177__ & new_new_n17178__;
  assign new_new_n17181__ = ~new_new_n17179__ & ~new_new_n17180__;
  assign new_new_n17182__ = new_new_n17176__ & ~new_new_n17181__;
  assign new_new_n17183__ = ~new_new_n17176__ & new_new_n17181__;
  assign new_new_n17184__ = ~new_new_n17182__ & ~new_new_n17183__;
  assign new_new_n17185__ = ~new_new_n17155__ & new_new_n17184__;
  assign new_new_n17186__ = new_new_n17155__ & ~new_new_n17184__;
  assign new_new_n17187__ = ~new_new_n17185__ & ~new_new_n17186__;
  assign new_new_n17188__ = new_new_n17117__ & new_new_n17187__;
  assign new_new_n17189__ = ~new_new_n17117__ & ~new_new_n17187__;
  assign new_new_n17190__ = ~new_new_n17188__ & ~new_new_n17189__;
  assign new_new_n17191__ = new_new_n17112__ & ~new_new_n17190__;
  assign new_new_n17192__ = ~new_new_n17112__ & new_new_n17190__;
  assign new_new_n17193__ = ~new_new_n17191__ & ~new_new_n17192__;
  assign new_new_n17194__ = new_new_n17051__ & ~new_new_n17193__;
  assign new_new_n17195__ = ~new_new_n17051__ & new_new_n17193__;
  assign po094 = new_new_n17194__ | new_new_n17195__;
  assign new_new_n17197__ = ~new_new_n17110__ & new_new_n17190__;
  assign new_new_n17198__ = ~new_new_n17111__ & ~new_new_n17197__;
  assign new_new_n17199__ = ~new_new_n17050__ & new_new_n17193__;
  assign new_new_n17200__ = ~new_new_n17049__ & ~new_new_n17199__;
  assign new_new_n17201__ = new_new_n17198__ & ~new_new_n17200__;
  assign new_new_n17202__ = ~new_new_n17198__ & new_new_n17200__;
  assign new_new_n17203__ = ~new_new_n17201__ & ~new_new_n17202__;
  assign new_new_n17204__ = ~new_new_n17141__ & ~new_new_n17145__;
  assign new_new_n17205__ = ~new_new_n17144__ & ~new_new_n17204__;
  assign new_new_n17206__ = ~new_new_n17120__ & ~new_new_n17124__;
  assign new_new_n17207__ = ~new_new_n17123__ & ~new_new_n17206__;
  assign new_new_n17208__ = ~new_new_n17205__ & ~new_new_n17207__;
  assign new_new_n17209__ = new_new_n17205__ & new_new_n17207__;
  assign new_new_n17210__ = ~new_new_n17208__ & ~new_new_n17209__;
  assign new_new_n17211__ = ~new_new_n17129__ & ~new_new_n17133__;
  assign new_new_n17212__ = ~new_new_n17132__ & ~new_new_n17211__;
  assign new_new_n17213__ = ~new_new_n17210__ & new_new_n17212__;
  assign new_new_n17214__ = new_new_n17210__ & ~new_new_n17212__;
  assign new_new_n17215__ = ~new_new_n17213__ & ~new_new_n17214__;
  assign new_new_n17216__ = ~new_new_n17174__ & ~new_new_n17181__;
  assign new_new_n17217__ = ~new_new_n17175__ & ~new_new_n17216__;
  assign new_new_n17218__ = ~new_new_n17156__ & ~new_new_n17160__;
  assign new_new_n17219__ = ~new_new_n17159__ & ~new_new_n17218__;
  assign new_new_n17220__ = pi63 & new_new_n17219__;
  assign new_new_n17221__ = pi31 & new_new_n17220__;
  assign new_new_n17222__ = ~pi63 & ~new_new_n17219__;
  assign new_new_n17223__ = ~pi31 & ~new_new_n17219__;
  assign new_new_n17224__ = ~new_new_n17222__ & ~new_new_n17223__;
  assign new_new_n17225__ = ~new_new_n17221__ & new_new_n17224__;
  assign new_new_n17226__ = pi46 & ~new_new_n17225__;
  assign new_new_n17227__ = ~pi46 & new_new_n17220__;
  assign new_new_n17228__ = pi31 & new_new_n17222__;
  assign new_new_n17229__ = ~new_new_n17227__ & ~new_new_n17228__;
  assign new_new_n17230__ = pi62 & ~new_new_n17229__;
  assign new_new_n17231__ = ~new_new_n17226__ & ~new_new_n17230__;
  assign new_new_n17232__ = pi47 & ~new_new_n17231__;
  assign new_new_n17233__ = pi46 & pi47;
  assign new_new_n17234__ = pi47 & pi62;
  assign new_new_n17235__ = ~new_new_n17220__ & ~new_new_n17234__;
  assign new_new_n17236__ = pi31 & ~new_new_n17235__;
  assign new_new_n17237__ = new_new_n17224__ & ~new_new_n17233__;
  assign new_new_n17238__ = ~new_new_n17236__ & new_new_n17237__;
  assign new_new_n17239__ = ~new_new_n17232__ & ~new_new_n17238__;
  assign new_new_n17240__ = new_new_n17217__ & new_new_n17239__;
  assign new_new_n17241__ = ~new_new_n17217__ & ~new_new_n17239__;
  assign new_new_n17242__ = ~new_new_n17240__ & ~new_new_n17241__;
  assign new_new_n17243__ = ~new_new_n17215__ & new_new_n17242__;
  assign new_new_n17244__ = new_new_n17215__ & ~new_new_n17242__;
  assign new_new_n17245__ = ~new_new_n17243__ & ~new_new_n17244__;
  assign new_new_n17246__ = ~new_new_n17056__ & ~new_new_n17059__;
  assign new_new_n17247__ = ~new_new_n17055__ & ~new_new_n17246__;
  assign new_new_n17248__ = pi44 & pi50;
  assign new_new_n17249__ = pi36 & pi58;
  assign new_new_n17250__ = pi43 & pi51;
  assign new_new_n17251__ = ~new_new_n17249__ & ~new_new_n17250__;
  assign new_new_n17252__ = new_new_n17249__ & new_new_n17250__;
  assign new_new_n17253__ = ~new_new_n17251__ & ~new_new_n17252__;
  assign new_new_n17254__ = new_new_n17248__ & ~new_new_n17253__;
  assign new_new_n17255__ = ~new_new_n17248__ & new_new_n17253__;
  assign new_new_n17256__ = ~new_new_n17254__ & ~new_new_n17255__;
  assign new_new_n17257__ = pi42 & pi52;
  assign new_new_n17258__ = pi40 & pi54;
  assign new_new_n17259__ = pi41 & pi53;
  assign new_new_n17260__ = ~new_new_n17258__ & ~new_new_n17259__;
  assign new_new_n17261__ = new_new_n17258__ & new_new_n17259__;
  assign new_new_n17262__ = ~new_new_n17260__ & ~new_new_n17261__;
  assign new_new_n17263__ = new_new_n17257__ & ~new_new_n17262__;
  assign new_new_n17264__ = ~new_new_n17257__ & new_new_n17262__;
  assign new_new_n17265__ = ~new_new_n17263__ & ~new_new_n17264__;
  assign new_new_n17266__ = new_new_n17256__ & new_new_n17265__;
  assign new_new_n17267__ = ~new_new_n17256__ & ~new_new_n17265__;
  assign new_new_n17268__ = ~new_new_n17266__ & ~new_new_n17267__;
  assign new_new_n17269__ = pi46 & pi48;
  assign new_new_n17270__ = pi38 & pi56;
  assign new_new_n17271__ = pi45 & pi49;
  assign new_new_n17272__ = ~new_new_n17270__ & ~new_new_n17271__;
  assign new_new_n17273__ = new_new_n17270__ & new_new_n17271__;
  assign new_new_n17274__ = ~new_new_n17272__ & ~new_new_n17273__;
  assign new_new_n17275__ = new_new_n17269__ & ~new_new_n17274__;
  assign new_new_n17276__ = ~new_new_n17269__ & new_new_n17274__;
  assign new_new_n17277__ = ~new_new_n17275__ & ~new_new_n17276__;
  assign new_new_n17278__ = new_new_n17268__ & ~new_new_n17277__;
  assign new_new_n17279__ = ~new_new_n17268__ & new_new_n17277__;
  assign new_new_n17280__ = ~new_new_n17278__ & ~new_new_n17279__;
  assign new_new_n17281__ = new_new_n17247__ & new_new_n17280__;
  assign new_new_n17282__ = ~new_new_n17247__ & ~new_new_n17280__;
  assign new_new_n17283__ = ~new_new_n17281__ & ~new_new_n17282__;
  assign new_new_n17284__ = ~new_new_n17165__ & ~new_new_n17169__;
  assign new_new_n17285__ = ~new_new_n17168__ & ~new_new_n17284__;
  assign new_new_n17286__ = pi39 & pi55;
  assign new_new_n17287__ = pi37 & pi57;
  assign new_new_n17288__ = pi34 & pi60;
  assign new_new_n17289__ = ~new_new_n17287__ & ~new_new_n17288__;
  assign new_new_n17290__ = new_new_n17287__ & new_new_n17288__;
  assign new_new_n17291__ = ~new_new_n17289__ & ~new_new_n17290__;
  assign new_new_n17292__ = new_new_n17286__ & ~new_new_n17291__;
  assign new_new_n17293__ = ~new_new_n17286__ & new_new_n17291__;
  assign new_new_n17294__ = ~new_new_n17292__ & ~new_new_n17293__;
  assign new_new_n17295__ = ~new_new_n17285__ & new_new_n17294__;
  assign new_new_n17296__ = new_new_n17285__ & ~new_new_n17294__;
  assign new_new_n17297__ = ~new_new_n17295__ & ~new_new_n17296__;
  assign new_new_n17298__ = pi35 & pi59;
  assign new_new_n17299__ = pi33 & pi61;
  assign new_new_n17300__ = ~new_new_n10300__ & ~new_new_n17299__;
  assign new_new_n17301__ = new_new_n10300__ & new_new_n17299__;
  assign new_new_n17302__ = ~new_new_n17300__ & ~new_new_n17301__;
  assign new_new_n17303__ = new_new_n17298__ & ~new_new_n17302__;
  assign new_new_n17304__ = ~new_new_n17298__ & new_new_n17302__;
  assign new_new_n17305__ = ~new_new_n17303__ & ~new_new_n17304__;
  assign new_new_n17306__ = ~new_new_n17297__ & new_new_n17305__;
  assign new_new_n17307__ = new_new_n17297__ & ~new_new_n17305__;
  assign new_new_n17308__ = ~new_new_n17306__ & ~new_new_n17307__;
  assign new_new_n17309__ = new_new_n17283__ & ~new_new_n17308__;
  assign new_new_n17310__ = ~new_new_n17283__ & new_new_n17308__;
  assign new_new_n17311__ = ~new_new_n17309__ & ~new_new_n17310__;
  assign new_new_n17312__ = new_new_n17245__ & ~new_new_n17311__;
  assign new_new_n17313__ = ~new_new_n17245__ & new_new_n17311__;
  assign new_new_n17314__ = ~new_new_n17312__ & ~new_new_n17313__;
  assign new_new_n17315__ = ~new_new_n17101__ & ~new_new_n17104__;
  assign new_new_n17316__ = ~new_new_n17100__ & ~new_new_n17315__;
  assign new_new_n17317__ = new_new_n17314__ & new_new_n17316__;
  assign new_new_n17318__ = ~new_new_n17314__ & ~new_new_n17316__;
  assign new_new_n17319__ = ~new_new_n17317__ & ~new_new_n17318__;
  assign new_new_n17320__ = ~new_new_n17082__ & new_new_n17096__;
  assign new_new_n17321__ = ~new_new_n17083__ & ~new_new_n17320__;
  assign new_new_n17322__ = ~new_new_n17086__ & ~new_new_n17092__;
  assign new_new_n17323__ = ~new_new_n17091__ & ~new_new_n17322__;
  assign new_new_n17324__ = ~new_new_n17139__ & ~new_new_n17149__;
  assign new_new_n17325__ = ~new_new_n17138__ & ~new_new_n17324__;
  assign new_new_n17326__ = ~new_new_n17066__ & ~new_new_n17077__;
  assign new_new_n17327__ = ~new_new_n17076__ & ~new_new_n17326__;
  assign new_new_n17328__ = ~new_new_n17325__ & new_new_n17327__;
  assign new_new_n17329__ = new_new_n17325__ & ~new_new_n17327__;
  assign new_new_n17330__ = ~new_new_n17328__ & ~new_new_n17329__;
  assign new_new_n17331__ = new_new_n17323__ & new_new_n17330__;
  assign new_new_n17332__ = ~new_new_n17323__ & ~new_new_n17330__;
  assign new_new_n17333__ = ~new_new_n17331__ & ~new_new_n17332__;
  assign new_new_n17334__ = ~new_new_n17321__ & ~new_new_n17333__;
  assign new_new_n17335__ = new_new_n17321__ & new_new_n17333__;
  assign new_new_n17336__ = ~new_new_n17334__ & ~new_new_n17335__;
  assign new_new_n17337__ = ~new_new_n17154__ & ~new_new_n17336__;
  assign new_new_n17338__ = ~new_new_n17153__ & new_new_n17336__;
  assign new_new_n17339__ = new_new_n17184__ & ~new_new_n17338__;
  assign new_new_n17340__ = ~new_new_n17186__ & ~new_new_n17339__;
  assign new_new_n17341__ = ~new_new_n17115__ & ~new_new_n17337__;
  assign new_new_n17342__ = ~new_new_n17340__ & new_new_n17341__;
  assign new_new_n17343__ = ~new_new_n17154__ & ~new_new_n17184__;
  assign new_new_n17344__ = ~new_new_n17153__ & ~new_new_n17343__;
  assign new_new_n17345__ = ~new_new_n17336__ & ~new_new_n17344__;
  assign new_new_n17346__ = new_new_n17116__ & ~new_new_n17338__;
  assign new_new_n17347__ = ~new_new_n17345__ & new_new_n17346__;
  assign new_new_n17348__ = ~new_new_n17342__ & ~new_new_n17347__;
  assign new_new_n17349__ = new_new_n17319__ & ~new_new_n17348__;
  assign new_new_n17350__ = new_new_n17154__ & new_new_n17336__;
  assign new_new_n17351__ = ~new_new_n17345__ & ~new_new_n17350__;
  assign new_new_n17352__ = new_new_n17115__ & ~new_new_n17351__;
  assign new_new_n17353__ = ~new_new_n17153__ & ~new_new_n17336__;
  assign new_new_n17354__ = new_new_n17336__ & new_new_n17343__;
  assign new_new_n17355__ = ~new_new_n17116__ & ~new_new_n17185__;
  assign new_new_n17356__ = ~new_new_n17353__ & ~new_new_n17354__;
  assign new_new_n17357__ = new_new_n17355__ & new_new_n17356__;
  assign new_new_n17358__ = ~new_new_n17352__ & ~new_new_n17357__;
  assign new_new_n17359__ = ~new_new_n17319__ & ~new_new_n17358__;
  assign new_new_n17360__ = new_new_n17319__ & new_new_n17358__;
  assign new_new_n17361__ = new_new_n17348__ & ~new_new_n17360__;
  assign new_new_n17362__ = ~new_new_n17359__ & new_new_n17361__;
  assign new_new_n17363__ = ~new_new_n17349__ & ~new_new_n17362__;
  assign new_new_n17364__ = new_new_n17203__ & new_new_n17363__;
  assign new_new_n17365__ = ~new_new_n17203__ & ~new_new_n17363__;
  assign po095 = new_new_n17364__ | new_new_n17365__;
  assign new_new_n17367__ = ~new_new_n17312__ & ~new_new_n17316__;
  assign new_new_n17368__ = ~new_new_n17313__ & ~new_new_n17367__;
  assign new_new_n17369__ = ~new_new_n17266__ & ~new_new_n17277__;
  assign new_new_n17370__ = ~new_new_n17267__ & ~new_new_n17369__;
  assign new_new_n17371__ = ~new_new_n17257__ & ~new_new_n17261__;
  assign new_new_n17372__ = ~new_new_n17260__ & ~new_new_n17371__;
  assign new_new_n17373__ = ~new_new_n17298__ & ~new_new_n17301__;
  assign new_new_n17374__ = ~new_new_n17300__ & ~new_new_n17373__;
  assign new_new_n17375__ = ~new_new_n17286__ & ~new_new_n17290__;
  assign new_new_n17376__ = ~new_new_n17289__ & ~new_new_n17375__;
  assign new_new_n17377__ = ~new_new_n17374__ & ~new_new_n17376__;
  assign new_new_n17378__ = new_new_n17374__ & new_new_n17376__;
  assign new_new_n17379__ = ~new_new_n17377__ & ~new_new_n17378__;
  assign new_new_n17380__ = ~new_new_n17296__ & new_new_n17305__;
  assign new_new_n17381__ = ~new_new_n17295__ & ~new_new_n17380__;
  assign new_new_n17382__ = new_new_n17379__ & ~new_new_n17381__;
  assign new_new_n17383__ = ~new_new_n17379__ & new_new_n17381__;
  assign new_new_n17384__ = ~new_new_n17382__ & ~new_new_n17383__;
  assign new_new_n17385__ = new_new_n17372__ & ~new_new_n17384__;
  assign new_new_n17386__ = ~new_new_n17372__ & new_new_n17384__;
  assign new_new_n17387__ = ~new_new_n17385__ & ~new_new_n17386__;
  assign new_new_n17388__ = ~new_new_n17370__ & new_new_n17387__;
  assign new_new_n17389__ = new_new_n17370__ & ~new_new_n17387__;
  assign new_new_n17390__ = ~new_new_n17388__ & ~new_new_n17389__;
  assign new_new_n17391__ = ~new_new_n17335__ & ~new_new_n17344__;
  assign new_new_n17392__ = ~new_new_n17334__ & ~new_new_n17391__;
  assign new_new_n17393__ = ~new_new_n17323__ & ~new_new_n17328__;
  assign new_new_n17394__ = ~new_new_n17329__ & ~new_new_n17393__;
  assign new_new_n17395__ = pi44 & pi51;
  assign new_new_n17396__ = pi43 & pi52;
  assign new_new_n17397__ = pi42 & pi53;
  assign new_new_n17398__ = ~new_new_n17396__ & ~new_new_n17397__;
  assign new_new_n17399__ = new_new_n17396__ & new_new_n17397__;
  assign new_new_n17400__ = ~new_new_n17398__ & ~new_new_n17399__;
  assign new_new_n17401__ = new_new_n17395__ & ~new_new_n17400__;
  assign new_new_n17402__ = ~new_new_n17395__ & new_new_n17400__;
  assign new_new_n17403__ = ~new_new_n17401__ & ~new_new_n17402__;
  assign new_new_n17404__ = pi46 & pi49;
  assign new_new_n17405__ = pi39 & pi56;
  assign new_new_n17406__ = pi45 & pi50;
  assign new_new_n17407__ = ~new_new_n17405__ & ~new_new_n17406__;
  assign new_new_n17408__ = new_new_n17405__ & new_new_n17406__;
  assign new_new_n17409__ = ~new_new_n17407__ & ~new_new_n17408__;
  assign new_new_n17410__ = new_new_n17404__ & ~new_new_n17409__;
  assign new_new_n17411__ = ~new_new_n17404__ & new_new_n17409__;
  assign new_new_n17412__ = ~new_new_n17410__ & ~new_new_n17411__;
  assign new_new_n17413__ = new_new_n17403__ & new_new_n17412__;
  assign new_new_n17414__ = ~new_new_n17403__ & ~new_new_n17412__;
  assign new_new_n17415__ = ~new_new_n17413__ & ~new_new_n17414__;
  assign new_new_n17416__ = pi33 & pi62;
  assign new_new_n17417__ = ~pi47 & pi48;
  assign new_new_n17418__ = new_new_n17416__ & ~new_new_n17417__;
  assign new_new_n17419__ = ~new_new_n17416__ & new_new_n17417__;
  assign new_new_n17420__ = ~new_new_n17418__ & ~new_new_n17419__;
  assign new_new_n17421__ = new_new_n17415__ & ~new_new_n17420__;
  assign new_new_n17422__ = ~new_new_n17415__ & new_new_n17420__;
  assign new_new_n17423__ = ~new_new_n17421__ & ~new_new_n17422__;
  assign new_new_n17424__ = ~new_new_n17394__ & ~new_new_n17423__;
  assign new_new_n17425__ = new_new_n17394__ & new_new_n17423__;
  assign new_new_n17426__ = ~new_new_n17424__ & ~new_new_n17425__;
  assign new_new_n17427__ = ~new_new_n17248__ & ~new_new_n17252__;
  assign new_new_n17428__ = ~new_new_n17251__ & ~new_new_n17427__;
  assign new_new_n17429__ = pi40 & pi55;
  assign new_new_n17430__ = pi38 & pi57;
  assign new_new_n17431__ = pi37 & pi58;
  assign new_new_n17432__ = ~new_new_n17430__ & ~new_new_n17431__;
  assign new_new_n17433__ = new_new_n17430__ & new_new_n17431__;
  assign new_new_n17434__ = ~new_new_n17432__ & ~new_new_n17433__;
  assign new_new_n17435__ = new_new_n17429__ & ~new_new_n17434__;
  assign new_new_n17436__ = ~new_new_n17429__ & new_new_n17434__;
  assign new_new_n17437__ = ~new_new_n17435__ & ~new_new_n17436__;
  assign new_new_n17438__ = ~new_new_n17428__ & new_new_n17437__;
  assign new_new_n17439__ = new_new_n17428__ & ~new_new_n17437__;
  assign new_new_n17440__ = ~new_new_n17438__ & ~new_new_n17439__;
  assign new_new_n17441__ = pi41 & pi54;
  assign new_new_n17442__ = pi32 & pi63;
  assign new_new_n17443__ = pi34 & pi61;
  assign new_new_n17444__ = ~new_new_n17442__ & ~new_new_n17443__;
  assign new_new_n17445__ = new_new_n17442__ & new_new_n17443__;
  assign new_new_n17446__ = ~new_new_n17444__ & ~new_new_n17445__;
  assign new_new_n17447__ = new_new_n17441__ & ~new_new_n17446__;
  assign new_new_n17448__ = ~new_new_n17441__ & new_new_n17446__;
  assign new_new_n17449__ = ~new_new_n17447__ & ~new_new_n17448__;
  assign new_new_n17450__ = ~new_new_n17440__ & new_new_n17449__;
  assign new_new_n17451__ = new_new_n17440__ & ~new_new_n17449__;
  assign new_new_n17452__ = ~new_new_n17450__ & ~new_new_n17451__;
  assign new_new_n17453__ = new_new_n17426__ & new_new_n17452__;
  assign new_new_n17454__ = ~new_new_n17426__ & ~new_new_n17452__;
  assign new_new_n17455__ = ~new_new_n17453__ & ~new_new_n17454__;
  assign new_new_n17456__ = ~new_new_n17392__ & ~new_new_n17455__;
  assign new_new_n17457__ = new_new_n17392__ & new_new_n17455__;
  assign new_new_n17458__ = ~new_new_n17456__ & ~new_new_n17457__;
  assign new_new_n17459__ = new_new_n17390__ & new_new_n17458__;
  assign new_new_n17460__ = ~new_new_n17390__ & ~new_new_n17458__;
  assign new_new_n17461__ = ~new_new_n17459__ & ~new_new_n17460__;
  assign new_new_n17462__ = new_new_n17368__ & new_new_n17461__;
  assign new_new_n17463__ = ~new_new_n17368__ & ~new_new_n17461__;
  assign new_new_n17464__ = ~new_new_n17462__ & ~new_new_n17463__;
  assign new_new_n17465__ = ~new_new_n17215__ & ~new_new_n17240__;
  assign new_new_n17466__ = ~new_new_n17241__ & ~new_new_n17465__;
  assign new_new_n17467__ = ~new_new_n17281__ & ~new_new_n17308__;
  assign new_new_n17468__ = ~new_new_n17282__ & ~new_new_n17467__;
  assign new_new_n17469__ = ~new_new_n17209__ & ~new_new_n17212__;
  assign new_new_n17470__ = ~new_new_n17208__ & ~new_new_n17469__;
  assign new_new_n17471__ = ~new_new_n17269__ & ~new_new_n17273__;
  assign new_new_n17472__ = ~new_new_n17272__ & ~new_new_n17471__;
  assign new_new_n17473__ = pi36 & pi59;
  assign new_new_n17474__ = pi35 & pi60;
  assign new_new_n17475__ = ~new_new_n17473__ & ~new_new_n17474__;
  assign new_new_n17476__ = new_new_n17473__ & new_new_n17474__;
  assign new_new_n17477__ = ~new_new_n17475__ & ~new_new_n17476__;
  assign new_new_n17478__ = new_new_n17472__ & ~new_new_n17477__;
  assign new_new_n17479__ = ~new_new_n17472__ & new_new_n17477__;
  assign new_new_n17480__ = ~new_new_n17478__ & ~new_new_n17479__;
  assign new_new_n17481__ = ~pi46 & ~new_new_n17177__;
  assign new_new_n17482__ = pi47 & ~new_new_n17481__;
  assign new_new_n17483__ = new_new_n17224__ & new_new_n17482__;
  assign new_new_n17484__ = ~new_new_n17221__ & ~new_new_n17483__;
  assign new_new_n17485__ = new_new_n17480__ & new_new_n17484__;
  assign new_new_n17486__ = ~new_new_n17480__ & ~new_new_n17484__;
  assign new_new_n17487__ = ~new_new_n17485__ & ~new_new_n17486__;
  assign new_new_n17488__ = new_new_n17470__ & new_new_n17487__;
  assign new_new_n17489__ = ~new_new_n17470__ & ~new_new_n17487__;
  assign new_new_n17490__ = ~new_new_n17488__ & ~new_new_n17489__;
  assign new_new_n17491__ = ~new_new_n17468__ & ~new_new_n17490__;
  assign new_new_n17492__ = new_new_n17468__ & new_new_n17490__;
  assign new_new_n17493__ = ~new_new_n17491__ & ~new_new_n17492__;
  assign new_new_n17494__ = new_new_n17466__ & ~new_new_n17493__;
  assign new_new_n17495__ = ~new_new_n17466__ & new_new_n17493__;
  assign new_new_n17496__ = ~new_new_n17494__ & ~new_new_n17495__;
  assign new_new_n17497__ = new_new_n17464__ & ~new_new_n17496__;
  assign new_new_n17498__ = ~new_new_n17464__ & new_new_n17496__;
  assign new_new_n17499__ = ~new_new_n17497__ & ~new_new_n17498__;
  assign new_new_n17500__ = new_new_n17359__ & new_new_n17499__;
  assign new_new_n17501__ = new_new_n17319__ & new_new_n17348__;
  assign new_new_n17502__ = ~new_new_n17499__ & new_new_n17501__;
  assign new_new_n17503__ = ~new_new_n17500__ & ~new_new_n17502__;
  assign new_new_n17504__ = new_new_n17203__ & ~new_new_n17503__;
  assign new_new_n17505__ = new_new_n17202__ & new_new_n17499__;
  assign new_new_n17506__ = new_new_n17201__ & ~new_new_n17499__;
  assign new_new_n17507__ = ~new_new_n17505__ & ~new_new_n17506__;
  assign new_new_n17508__ = new_new_n17361__ & ~new_new_n17507__;
  assign new_new_n17509__ = ~new_new_n17319__ & new_new_n17348__;
  assign new_new_n17510__ = new_new_n17201__ & ~new_new_n17509__;
  assign new_new_n17511__ = ~new_new_n17202__ & new_new_n17349__;
  assign new_new_n17512__ = new_new_n17499__ & ~new_new_n17510__;
  assign new_new_n17513__ = ~new_new_n17511__ & new_new_n17512__;
  assign new_new_n17514__ = new_new_n17203__ & ~new_new_n17319__;
  assign new_new_n17515__ = new_new_n17202__ & ~new_new_n17509__;
  assign new_new_n17516__ = ~new_new_n17499__ & ~new_new_n17515__;
  assign new_new_n17517__ = ~new_new_n17514__ & new_new_n17516__;
  assign new_new_n17518__ = new_new_n17358__ & ~new_new_n17513__;
  assign new_new_n17519__ = ~new_new_n17517__ & new_new_n17518__;
  assign new_new_n17520__ = ~new_new_n17504__ & ~new_new_n17508__;
  assign po096 = ~new_new_n17519__ & new_new_n17520__;
  assign new_new_n17522__ = ~new_new_n17201__ & new_new_n17499__;
  assign new_new_n17523__ = ~new_new_n17361__ & ~new_new_n17522__;
  assign new_new_n17524__ = ~new_new_n17349__ & new_new_n17499__;
  assign new_new_n17525__ = ~new_new_n17359__ & ~new_new_n17524__;
  assign new_new_n17526__ = ~new_new_n17202__ & new_new_n17525__;
  assign new_new_n17527__ = ~new_new_n17506__ & ~new_new_n17526__;
  assign new_new_n17528__ = ~new_new_n17523__ & new_new_n17527__;
  assign new_new_n17529__ = ~new_new_n17462__ & ~new_new_n17496__;
  assign new_new_n17530__ = ~new_new_n17463__ & ~new_new_n17529__;
  assign new_new_n17531__ = ~new_new_n17528__ & new_new_n17530__;
  assign new_new_n17532__ = new_new_n17528__ & ~new_new_n17530__;
  assign new_new_n17533__ = ~new_new_n17531__ & ~new_new_n17532__;
  assign new_new_n17534__ = ~new_new_n17390__ & ~new_new_n17457__;
  assign new_new_n17535__ = ~new_new_n17456__ & ~new_new_n17534__;
  assign new_new_n17536__ = ~new_new_n17413__ & ~new_new_n17420__;
  assign new_new_n17537__ = ~new_new_n17414__ & ~new_new_n17536__;
  assign new_new_n17538__ = ~pi47 & ~new_new_n17416__;
  assign new_new_n17539__ = pi48 & ~new_new_n17538__;
  assign new_new_n17540__ = ~new_new_n17395__ & ~new_new_n17399__;
  assign new_new_n17541__ = ~new_new_n17398__ & ~new_new_n17540__;
  assign new_new_n17542__ = ~new_new_n17404__ & ~new_new_n17408__;
  assign new_new_n17543__ = ~new_new_n17407__ & ~new_new_n17542__;
  assign new_new_n17544__ = ~new_new_n17541__ & ~new_new_n17543__;
  assign new_new_n17545__ = new_new_n17541__ & new_new_n17543__;
  assign new_new_n17546__ = ~new_new_n17544__ & ~new_new_n17545__;
  assign new_new_n17547__ = new_new_n17539__ & ~new_new_n17546__;
  assign new_new_n17548__ = ~new_new_n17539__ & new_new_n17546__;
  assign new_new_n17549__ = ~new_new_n17547__ & ~new_new_n17548__;
  assign new_new_n17550__ = new_new_n17537__ & new_new_n17549__;
  assign new_new_n17551__ = ~new_new_n17537__ & ~new_new_n17549__;
  assign new_new_n17552__ = ~new_new_n17550__ & ~new_new_n17551__;
  assign new_new_n17553__ = ~new_new_n17439__ & new_new_n17449__;
  assign new_new_n17554__ = ~new_new_n17438__ & ~new_new_n17553__;
  assign new_new_n17555__ = new_new_n17552__ & new_new_n17554__;
  assign new_new_n17556__ = ~new_new_n17552__ & ~new_new_n17554__;
  assign new_new_n17557__ = ~new_new_n17555__ & ~new_new_n17556__;
  assign new_new_n17558__ = ~new_new_n17429__ & ~new_new_n17433__;
  assign new_new_n17559__ = ~new_new_n17432__ & ~new_new_n17558__;
  assign new_new_n17560__ = ~new_new_n17441__ & ~new_new_n17445__;
  assign new_new_n17561__ = ~new_new_n17444__ & ~new_new_n17560__;
  assign new_new_n17562__ = ~new_new_n17472__ & ~new_new_n17476__;
  assign new_new_n17563__ = ~new_new_n17475__ & ~new_new_n17562__;
  assign new_new_n17564__ = ~new_new_n17561__ & ~new_new_n17563__;
  assign new_new_n17565__ = new_new_n17561__ & new_new_n17563__;
  assign new_new_n17566__ = ~new_new_n17564__ & ~new_new_n17565__;
  assign new_new_n17567__ = new_new_n17559__ & ~new_new_n17566__;
  assign new_new_n17568__ = ~new_new_n17559__ & new_new_n17566__;
  assign new_new_n17569__ = ~new_new_n17567__ & ~new_new_n17568__;
  assign new_new_n17570__ = new_new_n17470__ & ~new_new_n17485__;
  assign new_new_n17571__ = ~new_new_n17486__ & ~new_new_n17570__;
  assign new_new_n17572__ = pi43 & pi53;
  assign new_new_n17573__ = pi41 & pi55;
  assign new_new_n17574__ = pi42 & pi54;
  assign new_new_n17575__ = ~new_new_n17573__ & ~new_new_n17574__;
  assign new_new_n17576__ = new_new_n17573__ & new_new_n17574__;
  assign new_new_n17577__ = ~new_new_n17575__ & ~new_new_n17576__;
  assign new_new_n17578__ = new_new_n17572__ & ~new_new_n17577__;
  assign new_new_n17579__ = ~new_new_n17572__ & new_new_n17577__;
  assign new_new_n17580__ = ~new_new_n17578__ & ~new_new_n17579__;
  assign new_new_n17581__ = pi35 & pi61;
  assign new_new_n17582__ = pi33 & pi63;
  assign new_new_n17583__ = pi34 & pi62;
  assign new_new_n17584__ = ~new_new_n17582__ & ~new_new_n17583__;
  assign new_new_n17585__ = new_new_n17582__ & new_new_n17583__;
  assign new_new_n17586__ = ~new_new_n17584__ & ~new_new_n17585__;
  assign new_new_n17587__ = new_new_n17581__ & ~new_new_n17586__;
  assign new_new_n17588__ = ~new_new_n17581__ & new_new_n17586__;
  assign new_new_n17589__ = ~new_new_n17587__ & ~new_new_n17588__;
  assign new_new_n17590__ = new_new_n17580__ & new_new_n17589__;
  assign new_new_n17591__ = ~new_new_n17580__ & ~new_new_n17589__;
  assign new_new_n17592__ = ~new_new_n17590__ & ~new_new_n17591__;
  assign new_new_n17593__ = ~new_new_n17372__ & ~new_new_n17378__;
  assign new_new_n17594__ = ~new_new_n17377__ & ~new_new_n17593__;
  assign new_new_n17595__ = new_new_n17592__ & new_new_n17594__;
  assign new_new_n17596__ = ~new_new_n17592__ & ~new_new_n17594__;
  assign new_new_n17597__ = ~new_new_n17595__ & ~new_new_n17596__;
  assign new_new_n17598__ = ~new_new_n17571__ & new_new_n17597__;
  assign new_new_n17599__ = new_new_n17571__ & ~new_new_n17597__;
  assign new_new_n17600__ = ~new_new_n17598__ & ~new_new_n17599__;
  assign new_new_n17601__ = new_new_n17569__ & new_new_n17600__;
  assign new_new_n17602__ = ~new_new_n17569__ & ~new_new_n17600__;
  assign new_new_n17603__ = ~new_new_n17601__ & ~new_new_n17602__;
  assign new_new_n17604__ = ~new_new_n17557__ & new_new_n17603__;
  assign new_new_n17605__ = new_new_n17557__ & ~new_new_n17603__;
  assign new_new_n17606__ = ~new_new_n17604__ & ~new_new_n17605__;
  assign new_new_n17607__ = new_new_n17466__ & ~new_new_n17492__;
  assign new_new_n17608__ = ~new_new_n17491__ & ~new_new_n17607__;
  assign new_new_n17609__ = new_new_n17606__ & new_new_n17608__;
  assign new_new_n17610__ = ~new_new_n17606__ & ~new_new_n17608__;
  assign new_new_n17611__ = ~new_new_n17609__ & ~new_new_n17610__;
  assign new_new_n17612__ = new_new_n17535__ & new_new_n17611__;
  assign new_new_n17613__ = ~new_new_n17535__ & ~new_new_n17611__;
  assign new_new_n17614__ = ~new_new_n17612__ & ~new_new_n17613__;
  assign new_new_n17615__ = ~new_new_n17425__ & ~new_new_n17452__;
  assign new_new_n17616__ = ~new_new_n17424__ & ~new_new_n17615__;
  assign new_new_n17617__ = new_new_n17372__ & new_new_n17379__;
  assign new_new_n17618__ = ~new_new_n17372__ & ~new_new_n17379__;
  assign new_new_n17619__ = ~new_new_n17617__ & ~new_new_n17618__;
  assign new_new_n17620__ = new_new_n17381__ & new_new_n17619__;
  assign new_new_n17621__ = ~new_new_n17388__ & ~new_new_n17620__;
  assign new_new_n17622__ = ~new_new_n17616__ & new_new_n17621__;
  assign new_new_n17623__ = new_new_n17616__ & ~new_new_n17621__;
  assign new_new_n17624__ = ~new_new_n17622__ & ~new_new_n17623__;
  assign new_new_n17625__ = pi44 & pi52;
  assign new_new_n17626__ = pi38 & pi58;
  assign new_new_n17627__ = pi39 & pi57;
  assign new_new_n17628__ = ~new_new_n17626__ & ~new_new_n17627__;
  assign new_new_n17629__ = new_new_n17626__ & new_new_n17627__;
  assign new_new_n17630__ = ~new_new_n17628__ & ~new_new_n17629__;
  assign new_new_n17631__ = new_new_n17625__ & ~new_new_n17630__;
  assign new_new_n17632__ = ~new_new_n17625__ & new_new_n17630__;
  assign new_new_n17633__ = ~new_new_n17631__ & ~new_new_n17632__;
  assign new_new_n17634__ = pi47 & pi49;
  assign new_new_n17635__ = pi46 & pi50;
  assign new_new_n17636__ = pi45 & pi51;
  assign new_new_n17637__ = ~new_new_n17635__ & ~new_new_n17636__;
  assign new_new_n17638__ = new_new_n17635__ & new_new_n17636__;
  assign new_new_n17639__ = ~new_new_n17637__ & ~new_new_n17638__;
  assign new_new_n17640__ = new_new_n17634__ & ~new_new_n17639__;
  assign new_new_n17641__ = ~new_new_n17634__ & new_new_n17639__;
  assign new_new_n17642__ = ~new_new_n17640__ & ~new_new_n17641__;
  assign new_new_n17643__ = ~new_new_n17633__ & ~new_new_n17642__;
  assign new_new_n17644__ = new_new_n17633__ & new_new_n17642__;
  assign new_new_n17645__ = ~new_new_n17643__ & ~new_new_n17644__;
  assign new_new_n17646__ = pi40 & pi56;
  assign new_new_n17647__ = pi36 & pi60;
  assign new_new_n17648__ = pi37 & pi59;
  assign new_new_n17649__ = ~new_new_n17647__ & ~new_new_n17648__;
  assign new_new_n17650__ = new_new_n17647__ & new_new_n17648__;
  assign new_new_n17651__ = ~new_new_n17649__ & ~new_new_n17650__;
  assign new_new_n17652__ = new_new_n17646__ & ~new_new_n17651__;
  assign new_new_n17653__ = ~new_new_n17646__ & new_new_n17651__;
  assign new_new_n17654__ = ~new_new_n17652__ & ~new_new_n17653__;
  assign new_new_n17655__ = ~new_new_n17645__ & new_new_n17654__;
  assign new_new_n17656__ = new_new_n17645__ & ~new_new_n17654__;
  assign new_new_n17657__ = ~new_new_n17655__ & ~new_new_n17656__;
  assign new_new_n17658__ = new_new_n17624__ & new_new_n17657__;
  assign new_new_n17659__ = ~new_new_n17624__ & ~new_new_n17657__;
  assign new_new_n17660__ = ~new_new_n17658__ & ~new_new_n17659__;
  assign new_new_n17661__ = new_new_n17614__ & ~new_new_n17660__;
  assign new_new_n17662__ = ~new_new_n17614__ & new_new_n17660__;
  assign new_new_n17663__ = ~new_new_n17661__ & ~new_new_n17662__;
  assign new_new_n17664__ = new_new_n17533__ & new_new_n17663__;
  assign new_new_n17665__ = ~new_new_n17533__ & ~new_new_n17663__;
  assign po097 = new_new_n17664__ | new_new_n17665__;
  assign new_new_n17667__ = ~new_new_n17605__ & ~new_new_n17608__;
  assign new_new_n17668__ = ~new_new_n17604__ & ~new_new_n17667__;
  assign new_new_n17669__ = ~new_new_n17559__ & ~new_new_n17565__;
  assign new_new_n17670__ = ~new_new_n17564__ & ~new_new_n17669__;
  assign new_new_n17671__ = pi36 & pi61;
  assign new_new_n17672__ = ~new_new_n17634__ & ~new_new_n17638__;
  assign new_new_n17673__ = ~new_new_n17637__ & ~new_new_n17672__;
  assign new_new_n17674__ = ~new_new_n17625__ & ~new_new_n17629__;
  assign new_new_n17675__ = ~new_new_n17628__ & ~new_new_n17674__;
  assign new_new_n17676__ = new_new_n17673__ & new_new_n17675__;
  assign new_new_n17677__ = ~new_new_n17673__ & ~new_new_n17675__;
  assign new_new_n17678__ = ~new_new_n17676__ & ~new_new_n17677__;
  assign new_new_n17679__ = new_new_n17671__ & ~new_new_n17678__;
  assign new_new_n17680__ = ~new_new_n17671__ & new_new_n17678__;
  assign new_new_n17681__ = ~new_new_n17679__ & ~new_new_n17680__;
  assign new_new_n17682__ = ~new_new_n17670__ & new_new_n17681__;
  assign new_new_n17683__ = new_new_n17670__ & ~new_new_n17681__;
  assign new_new_n17684__ = ~new_new_n17682__ & ~new_new_n17683__;
  assign new_new_n17685__ = ~new_new_n17644__ & ~new_new_n17654__;
  assign new_new_n17686__ = ~new_new_n17643__ & ~new_new_n17685__;
  assign new_new_n17687__ = new_new_n17684__ & ~new_new_n17686__;
  assign new_new_n17688__ = ~new_new_n17684__ & new_new_n17686__;
  assign new_new_n17689__ = ~new_new_n17687__ & ~new_new_n17688__;
  assign new_new_n17690__ = ~new_new_n17591__ & ~new_new_n17594__;
  assign new_new_n17691__ = ~new_new_n17590__ & ~new_new_n17690__;
  assign new_new_n17692__ = pi35 & pi62;
  assign new_new_n17693__ = ~pi48 & pi49;
  assign new_new_n17694__ = ~new_new_n17692__ & new_new_n17693__;
  assign new_new_n17695__ = new_new_n17692__ & ~new_new_n17693__;
  assign new_new_n17696__ = ~new_new_n17694__ & ~new_new_n17695__;
  assign new_new_n17697__ = ~new_new_n17539__ & ~new_new_n17545__;
  assign new_new_n17698__ = ~new_new_n17544__ & ~new_new_n17697__;
  assign new_new_n17699__ = pi47 & pi50;
  assign new_new_n17700__ = pi46 & pi51;
  assign new_new_n17701__ = pi40 & pi57;
  assign new_new_n17702__ = ~new_new_n17700__ & ~new_new_n17701__;
  assign new_new_n17703__ = new_new_n17700__ & new_new_n17701__;
  assign new_new_n17704__ = ~new_new_n17702__ & ~new_new_n17703__;
  assign new_new_n17705__ = new_new_n17699__ & ~new_new_n17704__;
  assign new_new_n17706__ = ~new_new_n17699__ & new_new_n17704__;
  assign new_new_n17707__ = ~new_new_n17705__ & ~new_new_n17706__;
  assign new_new_n17708__ = ~new_new_n17698__ & new_new_n17707__;
  assign new_new_n17709__ = new_new_n17698__ & ~new_new_n17707__;
  assign new_new_n17710__ = ~new_new_n17708__ & ~new_new_n17709__;
  assign new_new_n17711__ = ~new_new_n17696__ & ~new_new_n17710__;
  assign new_new_n17712__ = new_new_n17696__ & new_new_n17710__;
  assign new_new_n17713__ = ~new_new_n17711__ & ~new_new_n17712__;
  assign new_new_n17714__ = new_new_n17691__ & ~new_new_n17713__;
  assign new_new_n17715__ = ~new_new_n17691__ & new_new_n17713__;
  assign new_new_n17716__ = ~new_new_n17714__ & ~new_new_n17715__;
  assign new_new_n17717__ = ~new_new_n17581__ & ~new_new_n17585__;
  assign new_new_n17718__ = ~new_new_n17584__ & ~new_new_n17717__;
  assign new_new_n17719__ = ~new_new_n17572__ & ~new_new_n17576__;
  assign new_new_n17720__ = ~new_new_n17575__ & ~new_new_n17719__;
  assign new_new_n17721__ = ~new_new_n17646__ & ~new_new_n17650__;
  assign new_new_n17722__ = ~new_new_n17649__ & ~new_new_n17721__;
  assign new_new_n17723__ = ~new_new_n17720__ & ~new_new_n17722__;
  assign new_new_n17724__ = new_new_n17720__ & new_new_n17722__;
  assign new_new_n17725__ = ~new_new_n17723__ & ~new_new_n17724__;
  assign new_new_n17726__ = new_new_n17718__ & ~new_new_n17725__;
  assign new_new_n17727__ = ~new_new_n17718__ & new_new_n17725__;
  assign new_new_n17728__ = ~new_new_n17726__ & ~new_new_n17727__;
  assign new_new_n17729__ = new_new_n17716__ & new_new_n17728__;
  assign new_new_n17730__ = ~new_new_n17716__ & ~new_new_n17728__;
  assign new_new_n17731__ = ~new_new_n17729__ & ~new_new_n17730__;
  assign new_new_n17732__ = ~new_new_n17689__ & new_new_n17731__;
  assign new_new_n17733__ = new_new_n17689__ & ~new_new_n17731__;
  assign new_new_n17734__ = ~new_new_n17732__ & ~new_new_n17733__;
  assign new_new_n17735__ = ~new_new_n17623__ & ~new_new_n17657__;
  assign new_new_n17736__ = ~new_new_n17622__ & ~new_new_n17735__;
  assign new_new_n17737__ = new_new_n17734__ & ~new_new_n17736__;
  assign new_new_n17738__ = ~new_new_n17734__ & new_new_n17736__;
  assign new_new_n17739__ = ~new_new_n17737__ & ~new_new_n17738__;
  assign new_new_n17740__ = new_new_n17668__ & ~new_new_n17739__;
  assign new_new_n17741__ = ~new_new_n17668__ & new_new_n17739__;
  assign new_new_n17742__ = ~new_new_n17740__ & ~new_new_n17741__;
  assign new_new_n17743__ = new_new_n17569__ & ~new_new_n17598__;
  assign new_new_n17744__ = ~new_new_n17599__ & ~new_new_n17743__;
  assign new_new_n17745__ = ~new_new_n17551__ & ~new_new_n17554__;
  assign new_new_n17746__ = ~new_new_n17550__ & ~new_new_n17745__;
  assign new_new_n17747__ = new_new_n17744__ & new_new_n17746__;
  assign new_new_n17748__ = ~new_new_n17744__ & ~new_new_n17746__;
  assign new_new_n17749__ = ~new_new_n17747__ & ~new_new_n17748__;
  assign new_new_n17750__ = pi45 & pi52;
  assign new_new_n17751__ = pi43 & pi54;
  assign new_new_n17752__ = pi44 & pi53;
  assign new_new_n17753__ = ~new_new_n17751__ & ~new_new_n17752__;
  assign new_new_n17754__ = new_new_n17751__ & new_new_n17752__;
  assign new_new_n17755__ = ~new_new_n17753__ & ~new_new_n17754__;
  assign new_new_n17756__ = new_new_n17750__ & ~new_new_n17755__;
  assign new_new_n17757__ = ~new_new_n17750__ & new_new_n17755__;
  assign new_new_n17758__ = ~new_new_n17756__ & ~new_new_n17757__;
  assign new_new_n17759__ = pi39 & pi58;
  assign new_new_n17760__ = pi38 & pi59;
  assign new_new_n17761__ = pi37 & pi60;
  assign new_new_n17762__ = ~new_new_n17760__ & ~new_new_n17761__;
  assign new_new_n17763__ = new_new_n17760__ & new_new_n17761__;
  assign new_new_n17764__ = ~new_new_n17762__ & ~new_new_n17763__;
  assign new_new_n17765__ = new_new_n17759__ & ~new_new_n17764__;
  assign new_new_n17766__ = ~new_new_n17759__ & new_new_n17764__;
  assign new_new_n17767__ = ~new_new_n17765__ & ~new_new_n17766__;
  assign new_new_n17768__ = new_new_n17758__ & new_new_n17767__;
  assign new_new_n17769__ = ~new_new_n17758__ & ~new_new_n17767__;
  assign new_new_n17770__ = ~new_new_n17768__ & ~new_new_n17769__;
  assign new_new_n17771__ = pi42 & pi55;
  assign new_new_n17772__ = pi34 & pi63;
  assign new_new_n17773__ = pi41 & pi56;
  assign new_new_n17774__ = ~new_new_n17772__ & ~new_new_n17773__;
  assign new_new_n17775__ = new_new_n17772__ & new_new_n17773__;
  assign new_new_n17776__ = ~new_new_n17774__ & ~new_new_n17775__;
  assign new_new_n17777__ = new_new_n17771__ & ~new_new_n17776__;
  assign new_new_n17778__ = ~new_new_n17771__ & new_new_n17776__;
  assign new_new_n17779__ = ~new_new_n17777__ & ~new_new_n17778__;
  assign new_new_n17780__ = ~new_new_n17770__ & new_new_n17779__;
  assign new_new_n17781__ = new_new_n17770__ & ~new_new_n17779__;
  assign new_new_n17782__ = ~new_new_n17780__ & ~new_new_n17781__;
  assign new_new_n17783__ = ~new_new_n17749__ & new_new_n17782__;
  assign new_new_n17784__ = new_new_n17749__ & ~new_new_n17782__;
  assign new_new_n17785__ = ~new_new_n17783__ & ~new_new_n17784__;
  assign new_new_n17786__ = new_new_n17742__ & ~new_new_n17785__;
  assign new_new_n17787__ = ~new_new_n17742__ & new_new_n17785__;
  assign new_new_n17788__ = ~new_new_n17786__ & ~new_new_n17787__;
  assign new_new_n17789__ = new_new_n17612__ & new_new_n17660__;
  assign new_new_n17790__ = new_new_n17613__ & ~new_new_n17660__;
  assign new_new_n17791__ = ~new_new_n17789__ & ~new_new_n17790__;
  assign new_new_n17792__ = new_new_n17533__ & new_new_n17791__;
  assign new_new_n17793__ = ~new_new_n17612__ & ~new_new_n17660__;
  assign new_new_n17794__ = ~new_new_n17613__ & ~new_new_n17793__;
  assign new_new_n17795__ = new_new_n17531__ & ~new_new_n17794__;
  assign new_new_n17796__ = new_new_n17532__ & new_new_n17794__;
  assign new_new_n17797__ = ~new_new_n17795__ & ~new_new_n17796__;
  assign new_new_n17798__ = ~new_new_n17792__ & new_new_n17797__;
  assign new_new_n17799__ = ~new_new_n17788__ & ~new_new_n17798__;
  assign new_new_n17800__ = new_new_n17531__ & new_new_n17612__;
  assign new_new_n17801__ = new_new_n17531__ & new_new_n17611__;
  assign new_new_n17802__ = ~new_new_n17531__ & ~new_new_n17611__;
  assign new_new_n17803__ = ~new_new_n17532__ & new_new_n17535__;
  assign new_new_n17804__ = ~new_new_n17802__ & new_new_n17803__;
  assign new_new_n17805__ = ~new_new_n17801__ & ~new_new_n17804__;
  assign new_new_n17806__ = new_new_n17660__ & ~new_new_n17805__;
  assign new_new_n17807__ = new_new_n17532__ & ~new_new_n17612__;
  assign new_new_n17808__ = ~new_new_n17535__ & new_new_n17802__;
  assign new_new_n17809__ = ~new_new_n17807__ & ~new_new_n17808__;
  assign new_new_n17810__ = ~new_new_n17660__ & ~new_new_n17809__;
  assign new_new_n17811__ = new_new_n17532__ & new_new_n17613__;
  assign new_new_n17812__ = ~new_new_n17800__ & ~new_new_n17811__;
  assign new_new_n17813__ = ~new_new_n17806__ & new_new_n17812__;
  assign new_new_n17814__ = ~new_new_n17810__ & new_new_n17813__;
  assign new_new_n17815__ = new_new_n17788__ & ~new_new_n17814__;
  assign po098 = new_new_n17799__ | new_new_n17815__;
  assign new_new_n17817__ = new_new_n17613__ & ~new_new_n17788__;
  assign new_new_n17818__ = ~new_new_n17613__ & new_new_n17788__;
  assign new_new_n17819__ = ~new_new_n17531__ & ~new_new_n17660__;
  assign new_new_n17820__ = ~new_new_n17532__ & ~new_new_n17819__;
  assign new_new_n17821__ = ~new_new_n17818__ & ~new_new_n17820__;
  assign new_new_n17822__ = ~new_new_n17532__ & new_new_n17788__;
  assign new_new_n17823__ = ~new_new_n17531__ & ~new_new_n17788__;
  assign new_new_n17824__ = new_new_n17660__ & ~new_new_n17823__;
  assign new_new_n17825__ = ~new_new_n17612__ & ~new_new_n17822__;
  assign new_new_n17826__ = ~new_new_n17824__ & new_new_n17825__;
  assign new_new_n17827__ = ~new_new_n17817__ & ~new_new_n17821__;
  assign new_new_n17828__ = ~new_new_n17826__ & new_new_n17827__;
  assign new_new_n17829__ = ~new_new_n17740__ & new_new_n17785__;
  assign new_new_n17830__ = ~new_new_n17741__ & ~new_new_n17829__;
  assign new_new_n17831__ = new_new_n17828__ & new_new_n17830__;
  assign new_new_n17832__ = ~new_new_n17828__ & ~new_new_n17830__;
  assign new_new_n17833__ = ~new_new_n17831__ & ~new_new_n17832__;
  assign new_new_n17834__ = ~new_new_n17771__ & ~new_new_n17775__;
  assign new_new_n17835__ = ~new_new_n17774__ & ~new_new_n17834__;
  assign new_new_n17836__ = ~new_new_n17750__ & ~new_new_n17754__;
  assign new_new_n17837__ = ~new_new_n17753__ & ~new_new_n17836__;
  assign new_new_n17838__ = ~new_new_n17759__ & ~new_new_n17763__;
  assign new_new_n17839__ = ~new_new_n17762__ & ~new_new_n17838__;
  assign new_new_n17840__ = ~new_new_n17837__ & ~new_new_n17839__;
  assign new_new_n17841__ = new_new_n17837__ & new_new_n17839__;
  assign new_new_n17842__ = ~new_new_n17840__ & ~new_new_n17841__;
  assign new_new_n17843__ = new_new_n17835__ & ~new_new_n17842__;
  assign new_new_n17844__ = ~new_new_n17835__ & new_new_n17842__;
  assign new_new_n17845__ = ~new_new_n17843__ & ~new_new_n17844__;
  assign new_new_n17846__ = pi37 & pi62;
  assign new_new_n17847__ = new_new_n17671__ & new_new_n17846__;
  assign new_new_n17848__ = pi37 & pi61;
  assign new_new_n17849__ = pi48 & new_new_n17848__;
  assign new_new_n17850__ = ~pi62 & ~new_new_n17849__;
  assign new_new_n17851__ = ~pi36 & ~new_new_n17848__;
  assign new_new_n17852__ = ~pi35 & ~pi48;
  assign new_new_n17853__ = pi49 & ~new_new_n17852__;
  assign new_new_n17854__ = ~new_new_n17847__ & new_new_n17853__;
  assign new_new_n17855__ = ~new_new_n17851__ & new_new_n17854__;
  assign new_new_n17856__ = ~new_new_n17850__ & new_new_n17855__;
  assign new_new_n17857__ = pi48 & pi49;
  assign new_new_n17858__ = pi36 & ~new_new_n17848__;
  assign new_new_n17859__ = ~new_new_n15362__ & ~new_new_n17858__;
  assign new_new_n17860__ = pi62 & ~new_new_n17859__;
  assign new_new_n17861__ = pi36 & pi62;
  assign new_new_n17862__ = new_new_n17848__ & ~new_new_n17861__;
  assign new_new_n17863__ = ~new_new_n17857__ & ~new_new_n17862__;
  assign new_new_n17864__ = ~new_new_n17860__ & new_new_n17863__;
  assign new_new_n17865__ = ~new_new_n17856__ & ~new_new_n17864__;
  assign new_new_n17866__ = pi48 & pi50;
  assign new_new_n17867__ = pi47 & pi51;
  assign new_new_n17868__ = pi46 & pi52;
  assign new_new_n17869__ = ~new_new_n17867__ & ~new_new_n17868__;
  assign new_new_n17870__ = new_new_n17867__ & new_new_n17868__;
  assign new_new_n17871__ = ~new_new_n17869__ & ~new_new_n17870__;
  assign new_new_n17872__ = new_new_n17866__ & ~new_new_n17871__;
  assign new_new_n17873__ = ~new_new_n17866__ & new_new_n17871__;
  assign new_new_n17874__ = ~new_new_n17872__ & ~new_new_n17873__;
  assign new_new_n17875__ = new_new_n17865__ & ~new_new_n17874__;
  assign new_new_n17876__ = ~new_new_n17865__ & new_new_n17874__;
  assign new_new_n17877__ = ~new_new_n17875__ & ~new_new_n17876__;
  assign new_new_n17878__ = pi45 & pi53;
  assign new_new_n17879__ = pi40 & pi58;
  assign new_new_n17880__ = pi39 & pi59;
  assign new_new_n17881__ = ~new_new_n17879__ & ~new_new_n17880__;
  assign new_new_n17882__ = new_new_n17879__ & new_new_n17880__;
  assign new_new_n17883__ = ~new_new_n17881__ & ~new_new_n17882__;
  assign new_new_n17884__ = new_new_n17878__ & ~new_new_n17883__;
  assign new_new_n17885__ = ~new_new_n17878__ & new_new_n17883__;
  assign new_new_n17886__ = ~new_new_n17884__ & ~new_new_n17885__;
  assign new_new_n17887__ = ~new_new_n17877__ & new_new_n17886__;
  assign new_new_n17888__ = new_new_n17877__ & ~new_new_n17886__;
  assign new_new_n17889__ = ~new_new_n17887__ & ~new_new_n17888__;
  assign new_new_n17890__ = ~new_new_n17696__ & ~new_new_n17708__;
  assign new_new_n17891__ = ~new_new_n17709__ & ~new_new_n17890__;
  assign new_new_n17892__ = new_new_n17889__ & ~new_new_n17891__;
  assign new_new_n17893__ = ~new_new_n17889__ & new_new_n17891__;
  assign new_new_n17894__ = ~new_new_n17892__ & ~new_new_n17893__;
  assign new_new_n17895__ = new_new_n17845__ & new_new_n17894__;
  assign new_new_n17896__ = ~new_new_n17845__ & ~new_new_n17894__;
  assign new_new_n17897__ = ~new_new_n17895__ & ~new_new_n17896__;
  assign new_new_n17898__ = ~new_new_n17718__ & ~new_new_n17724__;
  assign new_new_n17899__ = ~new_new_n17723__ & ~new_new_n17898__;
  assign new_new_n17900__ = ~new_new_n17768__ & ~new_new_n17779__;
  assign new_new_n17901__ = ~new_new_n17769__ & ~new_new_n17900__;
  assign new_new_n17902__ = ~new_new_n17671__ & ~new_new_n17676__;
  assign new_new_n17903__ = ~new_new_n17677__ & ~new_new_n17902__;
  assign new_new_n17904__ = ~new_new_n17901__ & new_new_n17903__;
  assign new_new_n17905__ = new_new_n17901__ & ~new_new_n17903__;
  assign new_new_n17906__ = ~new_new_n17904__ & ~new_new_n17905__;
  assign new_new_n17907__ = ~new_new_n17899__ & ~new_new_n17906__;
  assign new_new_n17908__ = new_new_n17899__ & new_new_n17906__;
  assign new_new_n17909__ = ~new_new_n17907__ & ~new_new_n17908__;
  assign new_new_n17910__ = ~new_new_n17897__ & new_new_n17909__;
  assign new_new_n17911__ = new_new_n17897__ & ~new_new_n17909__;
  assign new_new_n17912__ = ~new_new_n17910__ & ~new_new_n17911__;
  assign new_new_n17913__ = ~new_new_n17748__ & new_new_n17782__;
  assign new_new_n17914__ = ~new_new_n17747__ & ~new_new_n17913__;
  assign new_new_n17915__ = new_new_n17912__ & ~new_new_n17914__;
  assign new_new_n17916__ = ~new_new_n17912__ & new_new_n17914__;
  assign new_new_n17917__ = ~new_new_n17915__ & ~new_new_n17916__;
  assign new_new_n17918__ = ~new_new_n17733__ & ~new_new_n17736__;
  assign new_new_n17919__ = ~new_new_n17732__ & ~new_new_n17918__;
  assign new_new_n17920__ = new_new_n17917__ & new_new_n17919__;
  assign new_new_n17921__ = ~new_new_n17917__ & ~new_new_n17919__;
  assign new_new_n17922__ = ~new_new_n17920__ & ~new_new_n17921__;
  assign new_new_n17923__ = ~new_new_n17714__ & new_new_n17728__;
  assign new_new_n17924__ = ~new_new_n17715__ & ~new_new_n17923__;
  assign new_new_n17925__ = ~new_new_n17683__ & new_new_n17686__;
  assign new_new_n17926__ = ~new_new_n17682__ & ~new_new_n17925__;
  assign new_new_n17927__ = ~new_new_n17924__ & ~new_new_n17926__;
  assign new_new_n17928__ = new_new_n17924__ & new_new_n17926__;
  assign new_new_n17929__ = ~new_new_n17927__ & ~new_new_n17928__;
  assign new_new_n17930__ = pi42 & pi56;
  assign new_new_n17931__ = pi41 & pi57;
  assign new_new_n17932__ = pi38 & pi60;
  assign new_new_n17933__ = ~new_new_n17931__ & ~new_new_n17932__;
  assign new_new_n17934__ = new_new_n17931__ & new_new_n17932__;
  assign new_new_n17935__ = ~new_new_n17933__ & ~new_new_n17934__;
  assign new_new_n17936__ = new_new_n17930__ & ~new_new_n17935__;
  assign new_new_n17937__ = ~new_new_n17930__ & new_new_n17935__;
  assign new_new_n17938__ = ~new_new_n17936__ & ~new_new_n17937__;
  assign new_new_n17939__ = ~new_new_n17699__ & ~new_new_n17703__;
  assign new_new_n17940__ = ~new_new_n17702__ & ~new_new_n17939__;
  assign new_new_n17941__ = pi44 & pi54;
  assign new_new_n17942__ = pi43 & pi55;
  assign new_new_n17943__ = pi35 & pi63;
  assign new_new_n17944__ = ~new_new_n17942__ & ~new_new_n17943__;
  assign new_new_n17945__ = new_new_n17942__ & new_new_n17943__;
  assign new_new_n17946__ = ~new_new_n17944__ & ~new_new_n17945__;
  assign new_new_n17947__ = new_new_n17941__ & ~new_new_n17946__;
  assign new_new_n17948__ = ~new_new_n17941__ & new_new_n17946__;
  assign new_new_n17949__ = ~new_new_n17947__ & ~new_new_n17948__;
  assign new_new_n17950__ = ~new_new_n17940__ & new_new_n17949__;
  assign new_new_n17951__ = new_new_n17940__ & ~new_new_n17949__;
  assign new_new_n17952__ = ~new_new_n17950__ & ~new_new_n17951__;
  assign new_new_n17953__ = new_new_n17938__ & new_new_n17952__;
  assign new_new_n17954__ = ~new_new_n17938__ & ~new_new_n17952__;
  assign new_new_n17955__ = ~new_new_n17953__ & ~new_new_n17954__;
  assign new_new_n17956__ = new_new_n17929__ & new_new_n17955__;
  assign new_new_n17957__ = ~new_new_n17929__ & ~new_new_n17955__;
  assign new_new_n17958__ = ~new_new_n17956__ & ~new_new_n17957__;
  assign new_new_n17959__ = new_new_n17922__ & ~new_new_n17958__;
  assign new_new_n17960__ = ~new_new_n17922__ & new_new_n17958__;
  assign new_new_n17961__ = ~new_new_n17959__ & ~new_new_n17960__;
  assign new_new_n17962__ = ~new_new_n17833__ & new_new_n17961__;
  assign new_new_n17963__ = new_new_n17833__ & ~new_new_n17961__;
  assign po099 = new_new_n17962__ | new_new_n17963__;
  assign new_new_n17965__ = ~new_new_n17921__ & ~new_new_n17958__;
  assign new_new_n17966__ = ~new_new_n17920__ & ~new_new_n17965__;
  assign new_new_n17967__ = ~new_new_n17832__ & new_new_n17961__;
  assign new_new_n17968__ = ~new_new_n17831__ & ~new_new_n17967__;
  assign new_new_n17969__ = new_new_n17966__ & new_new_n17968__;
  assign new_new_n17970__ = ~new_new_n17966__ & ~new_new_n17968__;
  assign new_new_n17971__ = ~new_new_n17969__ & ~new_new_n17970__;
  assign new_new_n17972__ = ~new_new_n17911__ & ~new_new_n17914__;
  assign new_new_n17973__ = ~new_new_n17910__ & ~new_new_n17972__;
  assign new_new_n17974__ = ~new_new_n17835__ & ~new_new_n17841__;
  assign new_new_n17975__ = ~new_new_n17840__ & ~new_new_n17974__;
  assign new_new_n17976__ = ~new_new_n17938__ & ~new_new_n17950__;
  assign new_new_n17977__ = ~new_new_n17951__ & ~new_new_n17976__;
  assign new_new_n17978__ = ~pi49 & pi50;
  assign new_new_n17979__ = new_new_n17846__ & ~new_new_n17978__;
  assign new_new_n17980__ = ~new_new_n17846__ & new_new_n17978__;
  assign new_new_n17981__ = ~new_new_n17979__ & ~new_new_n17980__;
  assign new_new_n17982__ = ~new_new_n17977__ & ~new_new_n17981__;
  assign new_new_n17983__ = new_new_n17977__ & new_new_n17981__;
  assign new_new_n17984__ = ~new_new_n17982__ & ~new_new_n17983__;
  assign new_new_n17985__ = new_new_n17975__ & new_new_n17984__;
  assign new_new_n17986__ = ~new_new_n17975__ & ~new_new_n17984__;
  assign new_new_n17987__ = ~new_new_n17985__ & ~new_new_n17986__;
  assign new_new_n17988__ = ~new_new_n17927__ & ~new_new_n17955__;
  assign new_new_n17989__ = ~new_new_n17928__ & ~new_new_n17988__;
  assign new_new_n17990__ = new_new_n17987__ & ~new_new_n17989__;
  assign new_new_n17991__ = ~new_new_n17987__ & new_new_n17989__;
  assign new_new_n17992__ = ~new_new_n17990__ & ~new_new_n17991__;
  assign new_new_n17993__ = ~new_new_n17878__ & ~new_new_n17882__;
  assign new_new_n17994__ = ~new_new_n17881__ & ~new_new_n17993__;
  assign new_new_n17995__ = ~new_new_n17866__ & ~new_new_n17870__;
  assign new_new_n17996__ = ~new_new_n17869__ & ~new_new_n17995__;
  assign new_new_n17997__ = ~new_new_n17941__ & ~new_new_n17945__;
  assign new_new_n17998__ = ~new_new_n17944__ & ~new_new_n17997__;
  assign new_new_n17999__ = new_new_n17996__ & new_new_n17998__;
  assign new_new_n18000__ = ~new_new_n17996__ & ~new_new_n17998__;
  assign new_new_n18001__ = ~new_new_n17999__ & ~new_new_n18000__;
  assign new_new_n18002__ = new_new_n17994__ & ~new_new_n18001__;
  assign new_new_n18003__ = ~new_new_n17994__ & new_new_n18001__;
  assign new_new_n18004__ = ~new_new_n18002__ & ~new_new_n18003__;
  assign new_new_n18005__ = ~new_new_n17875__ & new_new_n17886__;
  assign new_new_n18006__ = ~new_new_n17876__ & ~new_new_n18005__;
  assign new_new_n18007__ = new_new_n18004__ & ~new_new_n18006__;
  assign new_new_n18008__ = ~new_new_n18004__ & new_new_n18006__;
  assign new_new_n18009__ = ~new_new_n18007__ & ~new_new_n18008__;
  assign new_new_n18010__ = ~new_new_n17930__ & ~new_new_n17934__;
  assign new_new_n18011__ = ~new_new_n17933__ & ~new_new_n18010__;
  assign new_new_n18012__ = pi39 & pi60;
  assign new_new_n18013__ = pi36 & pi63;
  assign new_new_n18014__ = pi38 & pi61;
  assign new_new_n18015__ = ~new_new_n18013__ & ~new_new_n18014__;
  assign new_new_n18016__ = new_new_n18013__ & new_new_n18014__;
  assign new_new_n18017__ = ~new_new_n18015__ & ~new_new_n18016__;
  assign new_new_n18018__ = new_new_n18012__ & ~new_new_n18017__;
  assign new_new_n18019__ = ~new_new_n18012__ & new_new_n18017__;
  assign new_new_n18020__ = ~new_new_n18018__ & ~new_new_n18019__;
  assign new_new_n18021__ = ~new_new_n18011__ & new_new_n18020__;
  assign new_new_n18022__ = new_new_n18011__ & ~new_new_n18020__;
  assign new_new_n18023__ = ~new_new_n18021__ & ~new_new_n18022__;
  assign new_new_n18024__ = pi35 & ~new_new_n17851__;
  assign new_new_n18025__ = ~new_new_n15360__ & ~new_new_n18024__;
  assign new_new_n18026__ = pi49 & ~new_new_n18025__;
  assign new_new_n18027__ = pi37 & new_new_n17671__;
  assign new_new_n18028__ = ~new_new_n18026__ & ~new_new_n18027__;
  assign new_new_n18029__ = pi62 & ~new_new_n18028__;
  assign new_new_n18030__ = pi49 & new_new_n17849__;
  assign new_new_n18031__ = ~new_new_n18029__ & ~new_new_n18030__;
  assign new_new_n18032__ = new_new_n18023__ & new_new_n18031__;
  assign new_new_n18033__ = ~new_new_n18023__ & ~new_new_n18031__;
  assign new_new_n18034__ = ~new_new_n18032__ & ~new_new_n18033__;
  assign new_new_n18035__ = new_new_n18009__ & ~new_new_n18034__;
  assign new_new_n18036__ = ~new_new_n18009__ & new_new_n18034__;
  assign new_new_n18037__ = ~new_new_n18035__ & ~new_new_n18036__;
  assign new_new_n18038__ = new_new_n17992__ & ~new_new_n18037__;
  assign new_new_n18039__ = ~new_new_n17992__ & new_new_n18037__;
  assign new_new_n18040__ = ~new_new_n18038__ & ~new_new_n18039__;
  assign new_new_n18041__ = new_new_n17973__ & new_new_n18040__;
  assign new_new_n18042__ = ~new_new_n17973__ & ~new_new_n18040__;
  assign new_new_n18043__ = ~new_new_n18041__ & ~new_new_n18042__;
  assign new_new_n18044__ = ~new_new_n17899__ & ~new_new_n17904__;
  assign new_new_n18045__ = ~new_new_n17905__ & ~new_new_n18044__;
  assign new_new_n18046__ = new_new_n17845__ & ~new_new_n17892__;
  assign new_new_n18047__ = ~new_new_n17893__ & ~new_new_n18046__;
  assign new_new_n18048__ = ~new_new_n18045__ & ~new_new_n18047__;
  assign new_new_n18049__ = new_new_n18045__ & new_new_n18047__;
  assign new_new_n18050__ = ~new_new_n18048__ & ~new_new_n18049__;
  assign new_new_n18051__ = pi44 & pi55;
  assign new_new_n18052__ = pi40 & pi59;
  assign new_new_n18053__ = pi41 & pi58;
  assign new_new_n18054__ = ~new_new_n18052__ & ~new_new_n18053__;
  assign new_new_n18055__ = new_new_n18052__ & new_new_n18053__;
  assign new_new_n18056__ = ~new_new_n18054__ & ~new_new_n18055__;
  assign new_new_n18057__ = new_new_n18051__ & ~new_new_n18056__;
  assign new_new_n18058__ = ~new_new_n18051__ & new_new_n18056__;
  assign new_new_n18059__ = ~new_new_n18057__ & ~new_new_n18058__;
  assign new_new_n18060__ = pi48 & pi51;
  assign new_new_n18061__ = pi43 & pi56;
  assign new_new_n18062__ = pi42 & pi57;
  assign new_new_n18063__ = ~new_new_n18061__ & ~new_new_n18062__;
  assign new_new_n18064__ = new_new_n18061__ & new_new_n18062__;
  assign new_new_n18065__ = ~new_new_n18063__ & ~new_new_n18064__;
  assign new_new_n18066__ = new_new_n18060__ & ~new_new_n18065__;
  assign new_new_n18067__ = ~new_new_n18060__ & new_new_n18065__;
  assign new_new_n18068__ = ~new_new_n18066__ & ~new_new_n18067__;
  assign new_new_n18069__ = pi47 & pi52;
  assign new_new_n18070__ = pi45 & pi54;
  assign new_new_n18071__ = pi46 & pi53;
  assign new_new_n18072__ = ~new_new_n18070__ & ~new_new_n18071__;
  assign new_new_n18073__ = new_new_n18070__ & new_new_n18071__;
  assign new_new_n18074__ = ~new_new_n18072__ & ~new_new_n18073__;
  assign new_new_n18075__ = new_new_n18069__ & ~new_new_n18074__;
  assign new_new_n18076__ = ~new_new_n18069__ & new_new_n18074__;
  assign new_new_n18077__ = ~new_new_n18075__ & ~new_new_n18076__;
  assign new_new_n18078__ = new_new_n18068__ & new_new_n18077__;
  assign new_new_n18079__ = ~new_new_n18068__ & ~new_new_n18077__;
  assign new_new_n18080__ = ~new_new_n18078__ & ~new_new_n18079__;
  assign new_new_n18081__ = new_new_n18059__ & new_new_n18080__;
  assign new_new_n18082__ = ~new_new_n18059__ & ~new_new_n18080__;
  assign new_new_n18083__ = ~new_new_n18081__ & ~new_new_n18082__;
  assign new_new_n18084__ = new_new_n18050__ & new_new_n18083__;
  assign new_new_n18085__ = ~new_new_n18050__ & ~new_new_n18083__;
  assign new_new_n18086__ = ~new_new_n18084__ & ~new_new_n18085__;
  assign new_new_n18087__ = new_new_n18043__ & ~new_new_n18086__;
  assign new_new_n18088__ = ~new_new_n18043__ & new_new_n18086__;
  assign new_new_n18089__ = ~new_new_n18087__ & ~new_new_n18088__;
  assign new_new_n18090__ = new_new_n17971__ & new_new_n18089__;
  assign new_new_n18091__ = ~new_new_n17971__ & ~new_new_n18089__;
  assign po100 = ~new_new_n18090__ & ~new_new_n18091__;
  assign new_new_n18093__ = ~new_new_n17991__ & new_new_n18037__;
  assign new_new_n18094__ = ~new_new_n17990__ & ~new_new_n18093__;
  assign new_new_n18095__ = ~new_new_n18012__ & ~new_new_n18016__;
  assign new_new_n18096__ = ~new_new_n18015__ & ~new_new_n18095__;
  assign new_new_n18097__ = ~new_new_n18069__ & ~new_new_n18073__;
  assign new_new_n18098__ = ~new_new_n18072__ & ~new_new_n18097__;
  assign new_new_n18099__ = ~new_new_n18096__ & ~new_new_n18098__;
  assign new_new_n18100__ = new_new_n18096__ & new_new_n18098__;
  assign new_new_n18101__ = ~new_new_n18099__ & ~new_new_n18100__;
  assign new_new_n18102__ = ~new_new_n18051__ & ~new_new_n18055__;
  assign new_new_n18103__ = ~new_new_n18054__ & ~new_new_n18102__;
  assign new_new_n18104__ = ~new_new_n18101__ & new_new_n18103__;
  assign new_new_n18105__ = new_new_n18101__ & ~new_new_n18103__;
  assign new_new_n18106__ = ~new_new_n18104__ & ~new_new_n18105__;
  assign new_new_n18107__ = ~new_new_n18059__ & ~new_new_n18078__;
  assign new_new_n18108__ = ~new_new_n18079__ & ~new_new_n18107__;
  assign new_new_n18109__ = ~new_new_n18060__ & ~new_new_n18064__;
  assign new_new_n18110__ = ~new_new_n18063__ & ~new_new_n18109__;
  assign new_new_n18111__ = pi37 & pi63;
  assign new_new_n18112__ = new_new_n18110__ & ~new_new_n18111__;
  assign new_new_n18113__ = ~pi37 & pi49;
  assign new_new_n18114__ = pi63 & ~new_new_n18110__;
  assign new_new_n18115__ = ~new_new_n18113__ & new_new_n18114__;
  assign new_new_n18116__ = ~new_new_n18112__ & ~new_new_n18115__;
  assign new_new_n18117__ = ~pi37 & new_new_n18110__;
  assign new_new_n18118__ = pi62 & ~new_new_n18117__;
  assign new_new_n18119__ = ~pi49 & ~new_new_n18118__;
  assign new_new_n18120__ = pi50 & ~new_new_n18116__;
  assign new_new_n18121__ = ~new_new_n18119__ & new_new_n18120__;
  assign new_new_n18122__ = pi50 & pi62;
  assign new_new_n18123__ = ~new_new_n18114__ & ~new_new_n18122__;
  assign new_new_n18124__ = pi37 & ~new_new_n18123__;
  assign new_new_n18125__ = pi49 & pi50;
  assign new_new_n18126__ = ~new_new_n18112__ & ~new_new_n18125__;
  assign new_new_n18127__ = ~new_new_n18124__ & new_new_n18126__;
  assign new_new_n18128__ = ~new_new_n18121__ & ~new_new_n18127__;
  assign new_new_n18129__ = new_new_n18108__ & ~new_new_n18128__;
  assign new_new_n18130__ = ~new_new_n18108__ & new_new_n18128__;
  assign new_new_n18131__ = ~new_new_n18129__ & ~new_new_n18130__;
  assign new_new_n18132__ = new_new_n18106__ & new_new_n18131__;
  assign new_new_n18133__ = ~new_new_n18106__ & ~new_new_n18131__;
  assign new_new_n18134__ = ~new_new_n18132__ & ~new_new_n18133__;
  assign new_new_n18135__ = ~new_new_n18048__ & ~new_new_n18083__;
  assign new_new_n18136__ = ~new_new_n18049__ & ~new_new_n18135__;
  assign new_new_n18137__ = ~new_new_n18134__ & ~new_new_n18136__;
  assign new_new_n18138__ = new_new_n18134__ & new_new_n18136__;
  assign new_new_n18139__ = ~new_new_n18137__ & ~new_new_n18138__;
  assign new_new_n18140__ = ~new_new_n17994__ & ~new_new_n17999__;
  assign new_new_n18141__ = ~new_new_n18000__ & ~new_new_n18140__;
  assign new_new_n18142__ = pi49 & pi51;
  assign new_new_n18143__ = pi48 & pi52;
  assign new_new_n18144__ = pi47 & pi53;
  assign new_new_n18145__ = ~new_new_n18143__ & ~new_new_n18144__;
  assign new_new_n18146__ = new_new_n18143__ & new_new_n18144__;
  assign new_new_n18147__ = ~new_new_n18145__ & ~new_new_n18146__;
  assign new_new_n18148__ = new_new_n18142__ & ~new_new_n18147__;
  assign new_new_n18149__ = ~new_new_n18142__ & new_new_n18147__;
  assign new_new_n18150__ = ~new_new_n18148__ & ~new_new_n18149__;
  assign new_new_n18151__ = ~new_new_n18141__ & new_new_n18150__;
  assign new_new_n18152__ = new_new_n18141__ & ~new_new_n18150__;
  assign new_new_n18153__ = ~new_new_n18151__ & ~new_new_n18152__;
  assign new_new_n18154__ = ~new_new_n18021__ & ~new_new_n18031__;
  assign new_new_n18155__ = ~new_new_n18022__ & ~new_new_n18154__;
  assign new_new_n18156__ = new_new_n18153__ & ~new_new_n18155__;
  assign new_new_n18157__ = ~new_new_n18153__ & new_new_n18155__;
  assign new_new_n18158__ = ~new_new_n18156__ & ~new_new_n18157__;
  assign new_new_n18159__ = new_new_n18139__ & ~new_new_n18158__;
  assign new_new_n18160__ = ~new_new_n18139__ & new_new_n18158__;
  assign new_new_n18161__ = ~new_new_n18159__ & ~new_new_n18160__;
  assign new_new_n18162__ = ~new_new_n18094__ & ~new_new_n18161__;
  assign new_new_n18163__ = new_new_n18094__ & new_new_n18161__;
  assign new_new_n18164__ = ~new_new_n18162__ & ~new_new_n18163__;
  assign new_new_n18165__ = ~new_new_n17975__ & ~new_new_n17982__;
  assign new_new_n18166__ = ~new_new_n17983__ & ~new_new_n18165__;
  assign new_new_n18167__ = ~new_new_n18007__ & ~new_new_n18034__;
  assign new_new_n18168__ = ~new_new_n18008__ & ~new_new_n18167__;
  assign new_new_n18169__ = new_new_n18166__ & ~new_new_n18168__;
  assign new_new_n18170__ = ~new_new_n18166__ & new_new_n18168__;
  assign new_new_n18171__ = ~new_new_n18169__ & ~new_new_n18170__;
  assign new_new_n18172__ = pi45 & pi55;
  assign new_new_n18173__ = pi43 & pi57;
  assign new_new_n18174__ = pi44 & pi56;
  assign new_new_n18175__ = ~new_new_n18173__ & ~new_new_n18174__;
  assign new_new_n18176__ = new_new_n18173__ & new_new_n18174__;
  assign new_new_n18177__ = ~new_new_n18175__ & ~new_new_n18176__;
  assign new_new_n18178__ = new_new_n18172__ & ~new_new_n18177__;
  assign new_new_n18179__ = ~new_new_n18172__ & new_new_n18177__;
  assign new_new_n18180__ = ~new_new_n18178__ & ~new_new_n18179__;
  assign new_new_n18181__ = pi46 & pi54;
  assign new_new_n18182__ = pi41 & pi59;
  assign new_new_n18183__ = pi42 & pi58;
  assign new_new_n18184__ = ~new_new_n18182__ & ~new_new_n18183__;
  assign new_new_n18185__ = new_new_n18182__ & new_new_n18183__;
  assign new_new_n18186__ = ~new_new_n18184__ & ~new_new_n18185__;
  assign new_new_n18187__ = new_new_n18181__ & ~new_new_n18186__;
  assign new_new_n18188__ = ~new_new_n18181__ & new_new_n18186__;
  assign new_new_n18189__ = ~new_new_n18187__ & ~new_new_n18188__;
  assign new_new_n18190__ = new_new_n18180__ & new_new_n18189__;
  assign new_new_n18191__ = ~new_new_n18180__ & ~new_new_n18189__;
  assign new_new_n18192__ = ~new_new_n18190__ & ~new_new_n18191__;
  assign new_new_n18193__ = pi40 & pi60;
  assign new_new_n18194__ = pi38 & pi62;
  assign new_new_n18195__ = pi39 & pi61;
  assign new_new_n18196__ = ~new_new_n18194__ & ~new_new_n18195__;
  assign new_new_n18197__ = new_new_n18194__ & new_new_n18195__;
  assign new_new_n18198__ = ~new_new_n18196__ & ~new_new_n18197__;
  assign new_new_n18199__ = new_new_n18193__ & ~new_new_n18198__;
  assign new_new_n18200__ = ~new_new_n18193__ & new_new_n18198__;
  assign new_new_n18201__ = ~new_new_n18199__ & ~new_new_n18200__;
  assign new_new_n18202__ = ~new_new_n18192__ & new_new_n18201__;
  assign new_new_n18203__ = new_new_n18192__ & ~new_new_n18201__;
  assign new_new_n18204__ = ~new_new_n18202__ & ~new_new_n18203__;
  assign new_new_n18205__ = new_new_n18171__ & new_new_n18204__;
  assign new_new_n18206__ = ~new_new_n18171__ & ~new_new_n18204__;
  assign new_new_n18207__ = ~new_new_n18205__ & ~new_new_n18206__;
  assign new_new_n18208__ = new_new_n18164__ & ~new_new_n18207__;
  assign new_new_n18209__ = ~new_new_n18164__ & new_new_n18207__;
  assign new_new_n18210__ = ~new_new_n18208__ & ~new_new_n18209__;
  assign new_new_n18211__ = ~new_new_n18041__ & ~new_new_n18086__;
  assign new_new_n18212__ = ~new_new_n18042__ & ~new_new_n18211__;
  assign new_new_n18213__ = ~new_new_n17970__ & new_new_n18212__;
  assign new_new_n18214__ = ~new_new_n17969__ & ~new_new_n18212__;
  assign new_new_n18215__ = ~new_new_n18213__ & ~new_new_n18214__;
  assign new_new_n18216__ = new_new_n18042__ & ~new_new_n18086__;
  assign new_new_n18217__ = new_new_n18041__ & new_new_n18086__;
  assign new_new_n18218__ = ~new_new_n18216__ & ~new_new_n18217__;
  assign new_new_n18219__ = new_new_n17971__ & new_new_n18218__;
  assign new_new_n18220__ = new_new_n18210__ & ~new_new_n18215__;
  assign new_new_n18221__ = ~new_new_n18219__ & new_new_n18220__;
  assign new_new_n18222__ = new_new_n17970__ & ~new_new_n17973__;
  assign new_new_n18223__ = ~new_new_n18040__ & new_new_n18222__;
  assign new_new_n18224__ = new_new_n18040__ & ~new_new_n18222__;
  assign new_new_n18225__ = ~new_new_n17969__ & ~new_new_n17973__;
  assign new_new_n18226__ = ~new_new_n17970__ & ~new_new_n18225__;
  assign new_new_n18227__ = ~new_new_n18086__ & ~new_new_n18224__;
  assign new_new_n18228__ = ~new_new_n18226__ & new_new_n18227__;
  assign new_new_n18229__ = new_new_n17969__ & new_new_n17973__;
  assign new_new_n18230__ = new_new_n18040__ & new_new_n18226__;
  assign new_new_n18231__ = ~new_new_n18229__ & ~new_new_n18230__;
  assign new_new_n18232__ = new_new_n18086__ & ~new_new_n18231__;
  assign new_new_n18233__ = new_new_n17969__ & new_new_n18041__;
  assign new_new_n18234__ = ~new_new_n18210__ & ~new_new_n18233__;
  assign new_new_n18235__ = ~new_new_n18223__ & new_new_n18234__;
  assign new_new_n18236__ = ~new_new_n18228__ & new_new_n18235__;
  assign new_new_n18237__ = ~new_new_n18232__ & new_new_n18236__;
  assign po101 = ~new_new_n18221__ & ~new_new_n18237__;
  assign new_new_n18239__ = ~new_new_n18210__ & ~new_new_n18213__;
  assign new_new_n18240__ = new_new_n17970__ & ~new_new_n18212__;
  assign new_new_n18241__ = new_new_n18210__ & ~new_new_n18216__;
  assign new_new_n18242__ = ~new_new_n18217__ & ~new_new_n18241__;
  assign new_new_n18243__ = ~new_new_n17969__ & new_new_n18242__;
  assign new_new_n18244__ = ~new_new_n18240__ & ~new_new_n18243__;
  assign new_new_n18245__ = ~new_new_n18239__ & new_new_n18244__;
  assign new_new_n18246__ = ~new_new_n18163__ & new_new_n18207__;
  assign new_new_n18247__ = ~new_new_n18162__ & ~new_new_n18246__;
  assign new_new_n18248__ = ~new_new_n18245__ & ~new_new_n18247__;
  assign new_new_n18249__ = new_new_n18245__ & new_new_n18247__;
  assign new_new_n18250__ = ~new_new_n18248__ & ~new_new_n18249__;
  assign new_new_n18251__ = ~new_new_n18138__ & new_new_n18158__;
  assign new_new_n18252__ = ~new_new_n18137__ & ~new_new_n18251__;
  assign new_new_n18253__ = ~new_new_n18106__ & ~new_new_n18129__;
  assign new_new_n18254__ = ~new_new_n18130__ & ~new_new_n18253__;
  assign new_new_n18255__ = ~new_new_n18100__ & ~new_new_n18103__;
  assign new_new_n18256__ = ~new_new_n18099__ & ~new_new_n18255__;
  assign new_new_n18257__ = ~new_new_n18190__ & ~new_new_n18201__;
  assign new_new_n18258__ = ~new_new_n18191__ & ~new_new_n18257__;
  assign new_new_n18259__ = ~new_new_n18172__ & ~new_new_n18176__;
  assign new_new_n18260__ = ~new_new_n18175__ & ~new_new_n18259__;
  assign new_new_n18261__ = ~new_new_n18181__ & ~new_new_n18185__;
  assign new_new_n18262__ = ~new_new_n18184__ & ~new_new_n18261__;
  assign new_new_n18263__ = ~new_new_n18193__ & ~new_new_n18197__;
  assign new_new_n18264__ = ~new_new_n18196__ & ~new_new_n18263__;
  assign new_new_n18265__ = new_new_n18262__ & new_new_n18264__;
  assign new_new_n18266__ = ~new_new_n18262__ & ~new_new_n18264__;
  assign new_new_n18267__ = ~new_new_n18265__ & ~new_new_n18266__;
  assign new_new_n18268__ = new_new_n18260__ & ~new_new_n18267__;
  assign new_new_n18269__ = ~new_new_n18260__ & new_new_n18267__;
  assign new_new_n18270__ = ~new_new_n18268__ & ~new_new_n18269__;
  assign new_new_n18271__ = ~new_new_n18258__ & ~new_new_n18270__;
  assign new_new_n18272__ = new_new_n18258__ & new_new_n18270__;
  assign new_new_n18273__ = ~new_new_n18271__ & ~new_new_n18272__;
  assign new_new_n18274__ = new_new_n18256__ & ~new_new_n18273__;
  assign new_new_n18275__ = ~new_new_n18256__ & new_new_n18273__;
  assign new_new_n18276__ = ~new_new_n18274__ & ~new_new_n18275__;
  assign new_new_n18277__ = ~new_new_n18254__ & ~new_new_n18276__;
  assign new_new_n18278__ = new_new_n18254__ & new_new_n18276__;
  assign new_new_n18279__ = ~new_new_n18277__ & ~new_new_n18278__;
  assign new_new_n18280__ = ~new_new_n18169__ & ~new_new_n18204__;
  assign new_new_n18281__ = ~new_new_n18170__ & ~new_new_n18280__;
  assign new_new_n18282__ = new_new_n18279__ & ~new_new_n18281__;
  assign new_new_n18283__ = ~new_new_n18279__ & new_new_n18281__;
  assign new_new_n18284__ = ~new_new_n18282__ & ~new_new_n18283__;
  assign new_new_n18285__ = new_new_n18252__ & new_new_n18284__;
  assign new_new_n18286__ = ~new_new_n18252__ & ~new_new_n18284__;
  assign new_new_n18287__ = ~new_new_n18285__ & ~new_new_n18286__;
  assign new_new_n18288__ = ~new_new_n18151__ & ~new_new_n18155__;
  assign new_new_n18289__ = ~new_new_n18152__ & ~new_new_n18288__;
  assign new_new_n18290__ = ~new_new_n18142__ & ~new_new_n18146__;
  assign new_new_n18291__ = ~new_new_n18145__ & ~new_new_n18290__;
  assign new_new_n18292__ = pi41 & pi60;
  assign new_new_n18293__ = pi40 & pi61;
  assign new_new_n18294__ = ~new_new_n18292__ & ~new_new_n18293__;
  assign new_new_n18295__ = new_new_n18292__ & new_new_n18293__;
  assign new_new_n18296__ = ~new_new_n18294__ & ~new_new_n18295__;
  assign new_new_n18297__ = new_new_n18291__ & ~new_new_n18296__;
  assign new_new_n18298__ = ~new_new_n18291__ & new_new_n18296__;
  assign new_new_n18299__ = ~new_new_n18297__ & ~new_new_n18298__;
  assign new_new_n18300__ = ~pi49 & ~new_new_n17846__;
  assign new_new_n18301__ = pi50 & ~new_new_n18300__;
  assign new_new_n18302__ = new_new_n18110__ & new_new_n18301__;
  assign new_new_n18303__ = ~new_new_n18111__ & ~new_new_n18302__;
  assign new_new_n18304__ = ~new_new_n18110__ & ~new_new_n18301__;
  assign new_new_n18305__ = ~new_new_n18303__ & ~new_new_n18304__;
  assign new_new_n18306__ = ~new_new_n18299__ & new_new_n18305__;
  assign new_new_n18307__ = new_new_n18299__ & ~new_new_n18305__;
  assign new_new_n18308__ = ~new_new_n18306__ & ~new_new_n18307__;
  assign new_new_n18309__ = pi39 & pi62;
  assign new_new_n18310__ = ~pi50 & pi51;
  assign new_new_n18311__ = new_new_n18309__ & ~new_new_n18310__;
  assign new_new_n18312__ = ~new_new_n18309__ & new_new_n18310__;
  assign new_new_n18313__ = ~new_new_n18311__ & ~new_new_n18312__;
  assign new_new_n18314__ = ~new_new_n18308__ & new_new_n18313__;
  assign new_new_n18315__ = new_new_n18308__ & ~new_new_n18313__;
  assign new_new_n18316__ = ~new_new_n18314__ & ~new_new_n18315__;
  assign new_new_n18317__ = ~new_new_n18289__ & new_new_n18316__;
  assign new_new_n18318__ = new_new_n18289__ & ~new_new_n18316__;
  assign new_new_n18319__ = ~new_new_n18317__ & ~new_new_n18318__;
  assign new_new_n18320__ = pi47 & pi54;
  assign new_new_n18321__ = pi38 & pi63;
  assign new_new_n18322__ = pi46 & pi55;
  assign new_new_n18323__ = ~new_new_n18321__ & ~new_new_n18322__;
  assign new_new_n18324__ = new_new_n18321__ & new_new_n18322__;
  assign new_new_n18325__ = ~new_new_n18323__ & ~new_new_n18324__;
  assign new_new_n18326__ = new_new_n18320__ & ~new_new_n18325__;
  assign new_new_n18327__ = ~new_new_n18320__ & new_new_n18325__;
  assign new_new_n18328__ = ~new_new_n18326__ & ~new_new_n18327__;
  assign new_new_n18329__ = pi49 & pi52;
  assign new_new_n18330__ = pi44 & pi57;
  assign new_new_n18331__ = pi48 & pi53;
  assign new_new_n18332__ = ~new_new_n18330__ & ~new_new_n18331__;
  assign new_new_n18333__ = new_new_n18330__ & new_new_n18331__;
  assign new_new_n18334__ = ~new_new_n18332__ & ~new_new_n18333__;
  assign new_new_n18335__ = new_new_n18329__ & ~new_new_n18334__;
  assign new_new_n18336__ = ~new_new_n18329__ & new_new_n18334__;
  assign new_new_n18337__ = ~new_new_n18335__ & ~new_new_n18336__;
  assign new_new_n18338__ = pi45 & pi56;
  assign new_new_n18339__ = pi43 & pi58;
  assign new_new_n18340__ = pi42 & pi59;
  assign new_new_n18341__ = ~new_new_n18339__ & ~new_new_n18340__;
  assign new_new_n18342__ = new_new_n18339__ & new_new_n18340__;
  assign new_new_n18343__ = ~new_new_n18341__ & ~new_new_n18342__;
  assign new_new_n18344__ = new_new_n18338__ & ~new_new_n18343__;
  assign new_new_n18345__ = ~new_new_n18338__ & new_new_n18343__;
  assign new_new_n18346__ = ~new_new_n18344__ & ~new_new_n18345__;
  assign new_new_n18347__ = new_new_n18337__ & new_new_n18346__;
  assign new_new_n18348__ = ~new_new_n18337__ & ~new_new_n18346__;
  assign new_new_n18349__ = ~new_new_n18347__ & ~new_new_n18348__;
  assign new_new_n18350__ = ~new_new_n18328__ & new_new_n18349__;
  assign new_new_n18351__ = new_new_n18328__ & ~new_new_n18349__;
  assign new_new_n18352__ = ~new_new_n18350__ & ~new_new_n18351__;
  assign new_new_n18353__ = new_new_n18319__ & ~new_new_n18352__;
  assign new_new_n18354__ = ~new_new_n18319__ & new_new_n18352__;
  assign new_new_n18355__ = ~new_new_n18353__ & ~new_new_n18354__;
  assign new_new_n18356__ = new_new_n18287__ & ~new_new_n18355__;
  assign new_new_n18357__ = ~new_new_n18287__ & new_new_n18355__;
  assign new_new_n18358__ = ~new_new_n18356__ & ~new_new_n18357__;
  assign new_new_n18359__ = new_new_n18250__ & new_new_n18358__;
  assign new_new_n18360__ = ~new_new_n18250__ & ~new_new_n18358__;
  assign po102 = ~new_new_n18359__ & ~new_new_n18360__;
  assign new_new_n18362__ = ~new_new_n18306__ & new_new_n18313__;
  assign new_new_n18363__ = ~new_new_n18307__ & ~new_new_n18362__;
  assign new_new_n18364__ = ~new_new_n18338__ & ~new_new_n18342__;
  assign new_new_n18365__ = ~new_new_n18341__ & ~new_new_n18364__;
  assign new_new_n18366__ = ~new_new_n18291__ & ~new_new_n18295__;
  assign new_new_n18367__ = ~new_new_n18294__ & ~new_new_n18366__;
  assign new_new_n18368__ = pi42 & pi60;
  assign new_new_n18369__ = pi39 & pi63;
  assign new_new_n18370__ = pi41 & pi61;
  assign new_new_n18371__ = ~new_new_n18369__ & ~new_new_n18370__;
  assign new_new_n18372__ = new_new_n18369__ & new_new_n18370__;
  assign new_new_n18373__ = ~new_new_n18371__ & ~new_new_n18372__;
  assign new_new_n18374__ = new_new_n18368__ & ~new_new_n18373__;
  assign new_new_n18375__ = ~new_new_n18368__ & new_new_n18373__;
  assign new_new_n18376__ = ~new_new_n18374__ & ~new_new_n18375__;
  assign new_new_n18377__ = new_new_n18367__ & ~new_new_n18376__;
  assign new_new_n18378__ = ~new_new_n18367__ & new_new_n18376__;
  assign new_new_n18379__ = ~new_new_n18377__ & ~new_new_n18378__;
  assign new_new_n18380__ = new_new_n18365__ & ~new_new_n18379__;
  assign new_new_n18381__ = ~new_new_n18365__ & new_new_n18379__;
  assign new_new_n18382__ = ~new_new_n18380__ & ~new_new_n18381__;
  assign new_new_n18383__ = new_new_n18363__ & ~new_new_n18382__;
  assign new_new_n18384__ = ~new_new_n18363__ & new_new_n18382__;
  assign new_new_n18385__ = ~new_new_n18383__ & ~new_new_n18384__;
  assign new_new_n18386__ = pi50 & pi52;
  assign new_new_n18387__ = pi49 & pi53;
  assign new_new_n18388__ = pi48 & pi54;
  assign new_new_n18389__ = ~new_new_n18387__ & ~new_new_n18388__;
  assign new_new_n18390__ = new_new_n18387__ & new_new_n18388__;
  assign new_new_n18391__ = ~new_new_n18389__ & ~new_new_n18390__;
  assign new_new_n18392__ = new_new_n18386__ & ~new_new_n18391__;
  assign new_new_n18393__ = ~new_new_n18386__ & new_new_n18391__;
  assign new_new_n18394__ = ~new_new_n18392__ & ~new_new_n18393__;
  assign new_new_n18395__ = pi44 & pi58;
  assign new_new_n18396__ = pi43 & pi59;
  assign new_new_n18397__ = pi40 & pi62;
  assign new_new_n18398__ = ~new_new_n18396__ & ~new_new_n18397__;
  assign new_new_n18399__ = new_new_n18396__ & new_new_n18397__;
  assign new_new_n18400__ = ~new_new_n18398__ & ~new_new_n18399__;
  assign new_new_n18401__ = new_new_n18395__ & ~new_new_n18400__;
  assign new_new_n18402__ = ~new_new_n18395__ & new_new_n18400__;
  assign new_new_n18403__ = ~new_new_n18401__ & ~new_new_n18402__;
  assign new_new_n18404__ = new_new_n18394__ & new_new_n18403__;
  assign new_new_n18405__ = ~new_new_n18394__ & ~new_new_n18403__;
  assign new_new_n18406__ = ~new_new_n18404__ & ~new_new_n18405__;
  assign new_new_n18407__ = pi47 & pi55;
  assign new_new_n18408__ = pi45 & pi57;
  assign new_new_n18409__ = pi46 & pi56;
  assign new_new_n18410__ = ~new_new_n18408__ & ~new_new_n18409__;
  assign new_new_n18411__ = new_new_n18408__ & new_new_n18409__;
  assign new_new_n18412__ = ~new_new_n18410__ & ~new_new_n18411__;
  assign new_new_n18413__ = new_new_n18407__ & ~new_new_n18412__;
  assign new_new_n18414__ = ~new_new_n18407__ & new_new_n18412__;
  assign new_new_n18415__ = ~new_new_n18413__ & ~new_new_n18414__;
  assign new_new_n18416__ = new_new_n18406__ & ~new_new_n18415__;
  assign new_new_n18417__ = ~new_new_n18406__ & new_new_n18415__;
  assign new_new_n18418__ = ~new_new_n18416__ & ~new_new_n18417__;
  assign new_new_n18419__ = new_new_n18385__ & ~new_new_n18418__;
  assign new_new_n18420__ = ~new_new_n18385__ & new_new_n18418__;
  assign new_new_n18421__ = ~new_new_n18419__ & ~new_new_n18420__;
  assign new_new_n18422__ = ~new_new_n18260__ & ~new_new_n18265__;
  assign new_new_n18423__ = ~new_new_n18266__ & ~new_new_n18422__;
  assign new_new_n18424__ = ~pi50 & ~new_new_n18309__;
  assign new_new_n18425__ = pi51 & ~new_new_n18424__;
  assign new_new_n18426__ = ~new_new_n18320__ & ~new_new_n18324__;
  assign new_new_n18427__ = ~new_new_n18323__ & ~new_new_n18426__;
  assign new_new_n18428__ = ~new_new_n18329__ & ~new_new_n18333__;
  assign new_new_n18429__ = ~new_new_n18332__ & ~new_new_n18428__;
  assign new_new_n18430__ = new_new_n18427__ & new_new_n18429__;
  assign new_new_n18431__ = ~new_new_n18427__ & ~new_new_n18429__;
  assign new_new_n18432__ = ~new_new_n18430__ & ~new_new_n18431__;
  assign new_new_n18433__ = new_new_n18425__ & ~new_new_n18432__;
  assign new_new_n18434__ = ~new_new_n18425__ & new_new_n18432__;
  assign new_new_n18435__ = ~new_new_n18433__ & ~new_new_n18434__;
  assign new_new_n18436__ = ~new_new_n18423__ & ~new_new_n18435__;
  assign new_new_n18437__ = new_new_n18423__ & new_new_n18435__;
  assign new_new_n18438__ = ~new_new_n18436__ & ~new_new_n18437__;
  assign new_new_n18439__ = ~new_new_n18328__ & ~new_new_n18347__;
  assign new_new_n18440__ = ~new_new_n18348__ & ~new_new_n18439__;
  assign new_new_n18441__ = new_new_n18256__ & ~new_new_n18272__;
  assign new_new_n18442__ = ~new_new_n18271__ & ~new_new_n18441__;
  assign new_new_n18443__ = ~new_new_n18318__ & new_new_n18352__;
  assign new_new_n18444__ = ~new_new_n18317__ & ~new_new_n18443__;
  assign new_new_n18445__ = new_new_n18442__ & new_new_n18444__;
  assign new_new_n18446__ = ~new_new_n18442__ & ~new_new_n18444__;
  assign new_new_n18447__ = ~new_new_n18445__ & ~new_new_n18446__;
  assign new_new_n18448__ = new_new_n18440__ & ~new_new_n18447__;
  assign new_new_n18449__ = ~new_new_n18440__ & new_new_n18447__;
  assign new_new_n18450__ = ~new_new_n18448__ & ~new_new_n18449__;
  assign new_new_n18451__ = new_new_n18438__ & new_new_n18450__;
  assign new_new_n18452__ = ~new_new_n18438__ & ~new_new_n18450__;
  assign new_new_n18453__ = ~new_new_n18451__ & ~new_new_n18452__;
  assign new_new_n18454__ = ~new_new_n18421__ & ~new_new_n18453__;
  assign new_new_n18455__ = new_new_n18421__ & new_new_n18453__;
  assign new_new_n18456__ = ~new_new_n18454__ & ~new_new_n18455__;
  assign new_new_n18457__ = ~new_new_n18278__ & new_new_n18281__;
  assign new_new_n18458__ = ~new_new_n18277__ & ~new_new_n18457__;
  assign new_new_n18459__ = new_new_n18456__ & ~new_new_n18458__;
  assign new_new_n18460__ = ~new_new_n18456__ & new_new_n18458__;
  assign new_new_n18461__ = ~new_new_n18459__ & ~new_new_n18460__;
  assign new_new_n18462__ = new_new_n18285__ & new_new_n18355__;
  assign new_new_n18463__ = new_new_n18286__ & ~new_new_n18355__;
  assign new_new_n18464__ = ~new_new_n18462__ & ~new_new_n18463__;
  assign new_new_n18465__ = new_new_n18250__ & new_new_n18464__;
  assign new_new_n18466__ = ~new_new_n18285__ & ~new_new_n18355__;
  assign new_new_n18467__ = ~new_new_n18286__ & ~new_new_n18466__;
  assign new_new_n18468__ = new_new_n18249__ & ~new_new_n18467__;
  assign new_new_n18469__ = new_new_n18248__ & new_new_n18467__;
  assign new_new_n18470__ = ~new_new_n18461__ & ~new_new_n18468__;
  assign new_new_n18471__ = ~new_new_n18469__ & new_new_n18470__;
  assign new_new_n18472__ = ~new_new_n18465__ & new_new_n18471__;
  assign new_new_n18473__ = ~new_new_n18247__ & ~new_new_n18252__;
  assign new_new_n18474__ = ~new_new_n18245__ & ~new_new_n18284__;
  assign new_new_n18475__ = new_new_n18473__ & new_new_n18474__;
  assign new_new_n18476__ = new_new_n18245__ & new_new_n18284__;
  assign new_new_n18477__ = new_new_n18247__ & new_new_n18252__;
  assign new_new_n18478__ = new_new_n18476__ & new_new_n18477__;
  assign new_new_n18479__ = new_new_n18249__ & new_new_n18284__;
  assign new_new_n18480__ = ~new_new_n18249__ & ~new_new_n18284__;
  assign new_new_n18481__ = ~new_new_n18248__ & ~new_new_n18480__;
  assign new_new_n18482__ = new_new_n18252__ & new_new_n18481__;
  assign new_new_n18483__ = new_new_n18355__ & ~new_new_n18479__;
  assign new_new_n18484__ = ~new_new_n18482__ & new_new_n18483__;
  assign new_new_n18485__ = new_new_n18248__ & ~new_new_n18284__;
  assign new_new_n18486__ = ~new_new_n18252__ & ~new_new_n18481__;
  assign new_new_n18487__ = ~new_new_n18355__ & ~new_new_n18485__;
  assign new_new_n18488__ = ~new_new_n18486__ & new_new_n18487__;
  assign new_new_n18489__ = ~new_new_n18484__ & ~new_new_n18488__;
  assign new_new_n18490__ = new_new_n18461__ & ~new_new_n18475__;
  assign new_new_n18491__ = ~new_new_n18478__ & new_new_n18490__;
  assign new_new_n18492__ = ~new_new_n18489__ & new_new_n18491__;
  assign po103 = ~new_new_n18472__ & ~new_new_n18492__;
  assign new_new_n18494__ = ~pi51 & pi52;
  assign new_new_n18495__ = ~new_new_n14927__ & new_new_n18494__;
  assign new_new_n18496__ = new_new_n14927__ & ~new_new_n18494__;
  assign new_new_n18497__ = ~new_new_n18495__ & ~new_new_n18496__;
  assign new_new_n18498__ = pi50 & pi53;
  assign new_new_n18499__ = pi49 & pi54;
  assign new_new_n18500__ = pi48 & pi55;
  assign new_new_n18501__ = ~new_new_n18499__ & ~new_new_n18500__;
  assign new_new_n18502__ = new_new_n18499__ & new_new_n18500__;
  assign new_new_n18503__ = ~new_new_n18501__ & ~new_new_n18502__;
  assign new_new_n18504__ = new_new_n18498__ & ~new_new_n18503__;
  assign new_new_n18505__ = ~new_new_n18498__ & new_new_n18503__;
  assign new_new_n18506__ = ~new_new_n18504__ & ~new_new_n18505__;
  assign new_new_n18507__ = pi47 & pi56;
  assign new_new_n18508__ = pi46 & pi57;
  assign new_new_n18509__ = pi43 & pi60;
  assign new_new_n18510__ = ~new_new_n18508__ & ~new_new_n18509__;
  assign new_new_n18511__ = new_new_n18508__ & new_new_n18509__;
  assign new_new_n18512__ = ~new_new_n18510__ & ~new_new_n18511__;
  assign new_new_n18513__ = new_new_n18507__ & ~new_new_n18512__;
  assign new_new_n18514__ = ~new_new_n18507__ & new_new_n18512__;
  assign new_new_n18515__ = ~new_new_n18513__ & ~new_new_n18514__;
  assign new_new_n18516__ = new_new_n18506__ & new_new_n18515__;
  assign new_new_n18517__ = ~new_new_n18506__ & ~new_new_n18515__;
  assign new_new_n18518__ = ~new_new_n18516__ & ~new_new_n18517__;
  assign new_new_n18519__ = new_new_n18497__ & new_new_n18518__;
  assign new_new_n18520__ = ~new_new_n18497__ & ~new_new_n18518__;
  assign new_new_n18521__ = ~new_new_n18519__ & ~new_new_n18520__;
  assign new_new_n18522__ = pi40 & pi63;
  assign new_new_n18523__ = ~new_new_n18386__ & ~new_new_n18390__;
  assign new_new_n18524__ = ~new_new_n18389__ & ~new_new_n18523__;
  assign new_new_n18525__ = ~new_new_n18407__ & ~new_new_n18411__;
  assign new_new_n18526__ = ~new_new_n18410__ & ~new_new_n18525__;
  assign new_new_n18527__ = new_new_n18524__ & new_new_n18526__;
  assign new_new_n18528__ = ~new_new_n18524__ & ~new_new_n18526__;
  assign new_new_n18529__ = ~new_new_n18527__ & ~new_new_n18528__;
  assign new_new_n18530__ = new_new_n18522__ & ~new_new_n18529__;
  assign new_new_n18531__ = ~new_new_n18522__ & new_new_n18529__;
  assign new_new_n18532__ = ~new_new_n18530__ & ~new_new_n18531__;
  assign new_new_n18533__ = ~new_new_n18521__ & ~new_new_n18532__;
  assign new_new_n18534__ = new_new_n18521__ & new_new_n18532__;
  assign new_new_n18535__ = ~new_new_n18533__ & ~new_new_n18534__;
  assign new_new_n18536__ = ~new_new_n18368__ & ~new_new_n18372__;
  assign new_new_n18537__ = ~new_new_n18371__ & ~new_new_n18536__;
  assign new_new_n18538__ = ~new_new_n18395__ & ~new_new_n18399__;
  assign new_new_n18539__ = ~new_new_n18398__ & ~new_new_n18538__;
  assign new_new_n18540__ = new_new_n18537__ & new_new_n18539__;
  assign new_new_n18541__ = ~new_new_n18537__ & ~new_new_n18539__;
  assign new_new_n18542__ = ~new_new_n18540__ & ~new_new_n18541__;
  assign new_new_n18543__ = pi45 & pi58;
  assign new_new_n18544__ = pi42 & pi61;
  assign new_new_n18545__ = pi44 & pi59;
  assign new_new_n18546__ = ~new_new_n18544__ & ~new_new_n18545__;
  assign new_new_n18547__ = new_new_n18544__ & new_new_n18545__;
  assign new_new_n18548__ = ~new_new_n18546__ & ~new_new_n18547__;
  assign new_new_n18549__ = new_new_n18543__ & ~new_new_n18548__;
  assign new_new_n18550__ = ~new_new_n18543__ & new_new_n18548__;
  assign new_new_n18551__ = ~new_new_n18549__ & ~new_new_n18550__;
  assign new_new_n18552__ = new_new_n18542__ & ~new_new_n18551__;
  assign new_new_n18553__ = ~new_new_n18542__ & new_new_n18551__;
  assign new_new_n18554__ = ~new_new_n18552__ & ~new_new_n18553__;
  assign new_new_n18555__ = new_new_n18535__ & ~new_new_n18554__;
  assign new_new_n18556__ = ~new_new_n18535__ & new_new_n18554__;
  assign new_new_n18557__ = ~new_new_n18555__ & ~new_new_n18556__;
  assign new_new_n18558__ = ~new_new_n18438__ & new_new_n18440__;
  assign new_new_n18559__ = new_new_n18438__ & ~new_new_n18440__;
  assign new_new_n18560__ = ~new_new_n18558__ & ~new_new_n18559__;
  assign new_new_n18561__ = ~new_new_n18446__ & new_new_n18560__;
  assign new_new_n18562__ = ~new_new_n18445__ & ~new_new_n18561__;
  assign new_new_n18563__ = ~new_new_n18557__ & new_new_n18562__;
  assign new_new_n18564__ = new_new_n18557__ & ~new_new_n18562__;
  assign new_new_n18565__ = ~new_new_n18563__ & ~new_new_n18564__;
  assign new_new_n18566__ = new_new_n18423__ & ~new_new_n18440__;
  assign new_new_n18567__ = new_new_n18435__ & ~new_new_n18566__;
  assign new_new_n18568__ = ~new_new_n18423__ & new_new_n18440__;
  assign new_new_n18569__ = ~new_new_n18567__ & ~new_new_n18568__;
  assign new_new_n18570__ = ~new_new_n18404__ & ~new_new_n18415__;
  assign new_new_n18571__ = ~new_new_n18405__ & ~new_new_n18570__;
  assign new_new_n18572__ = ~new_new_n18425__ & ~new_new_n18430__;
  assign new_new_n18573__ = ~new_new_n18431__ & ~new_new_n18572__;
  assign new_new_n18574__ = ~new_new_n18571__ & new_new_n18573__;
  assign new_new_n18575__ = new_new_n18571__ & ~new_new_n18573__;
  assign new_new_n18576__ = ~new_new_n18574__ & ~new_new_n18575__;
  assign new_new_n18577__ = new_new_n18365__ & ~new_new_n18378__;
  assign new_new_n18578__ = ~new_new_n18377__ & ~new_new_n18577__;
  assign new_new_n18579__ = new_new_n18576__ & new_new_n18578__;
  assign new_new_n18580__ = ~new_new_n18576__ & ~new_new_n18578__;
  assign new_new_n18581__ = ~new_new_n18579__ & ~new_new_n18580__;
  assign new_new_n18582__ = ~new_new_n18384__ & new_new_n18418__;
  assign new_new_n18583__ = ~new_new_n18383__ & ~new_new_n18582__;
  assign new_new_n18584__ = new_new_n18581__ & new_new_n18583__;
  assign new_new_n18585__ = ~new_new_n18581__ & ~new_new_n18583__;
  assign new_new_n18586__ = ~new_new_n18584__ & ~new_new_n18585__;
  assign new_new_n18587__ = ~new_new_n18569__ & new_new_n18586__;
  assign new_new_n18588__ = new_new_n18569__ & ~new_new_n18586__;
  assign new_new_n18589__ = ~new_new_n18587__ & ~new_new_n18588__;
  assign new_new_n18590__ = new_new_n18565__ & new_new_n18589__;
  assign new_new_n18591__ = ~new_new_n18565__ & ~new_new_n18589__;
  assign new_new_n18592__ = ~new_new_n18590__ & ~new_new_n18591__;
  assign new_new_n18593__ = ~new_new_n18355__ & ~new_new_n18477__;
  assign new_new_n18594__ = new_new_n18461__ & ~new_new_n18476__;
  assign new_new_n18595__ = ~new_new_n18473__ & ~new_new_n18593__;
  assign new_new_n18596__ = ~new_new_n18594__ & new_new_n18595__;
  assign new_new_n18597__ = ~new_new_n18355__ & new_new_n18473__;
  assign new_new_n18598__ = ~new_new_n18461__ & ~new_new_n18597__;
  assign new_new_n18599__ = new_new_n18355__ & new_new_n18477__;
  assign new_new_n18600__ = ~new_new_n18598__ & ~new_new_n18599__;
  assign new_new_n18601__ = ~new_new_n18474__ & ~new_new_n18600__;
  assign new_new_n18602__ = ~new_new_n18461__ & new_new_n18476__;
  assign new_new_n18603__ = ~new_new_n18601__ & ~new_new_n18602__;
  assign new_new_n18604__ = ~new_new_n18596__ & new_new_n18603__;
  assign new_new_n18605__ = new_new_n18592__ & ~new_new_n18604__;
  assign new_new_n18606__ = ~new_new_n18592__ & new_new_n18604__;
  assign new_new_n18607__ = ~new_new_n18605__ & ~new_new_n18606__;
  assign new_new_n18608__ = ~new_new_n18455__ & ~new_new_n18458__;
  assign new_new_n18609__ = ~new_new_n18454__ & ~new_new_n18608__;
  assign new_new_n18610__ = new_new_n18607__ & ~new_new_n18609__;
  assign new_new_n18611__ = ~new_new_n18607__ & new_new_n18609__;
  assign po104 = ~new_new_n18610__ & ~new_new_n18611__;
  assign new_new_n18613__ = ~new_new_n18605__ & ~new_new_n18609__;
  assign new_new_n18614__ = ~new_new_n18606__ & ~new_new_n18613__;
  assign new_new_n18615__ = ~new_new_n18564__ & ~new_new_n18589__;
  assign new_new_n18616__ = ~new_new_n18563__ & ~new_new_n18615__;
  assign new_new_n18617__ = new_new_n18614__ & new_new_n18616__;
  assign new_new_n18618__ = ~new_new_n18614__ & ~new_new_n18616__;
  assign new_new_n18619__ = ~new_new_n18617__ & ~new_new_n18618__;
  assign new_new_n18620__ = ~new_new_n18569__ & ~new_new_n18585__;
  assign new_new_n18621__ = ~new_new_n18584__ & ~new_new_n18620__;
  assign new_new_n18622__ = ~new_new_n18534__ & new_new_n18554__;
  assign new_new_n18623__ = ~new_new_n18533__ & ~new_new_n18622__;
  assign new_new_n18624__ = ~pi42 & ~pi63;
  assign new_new_n18625__ = pi42 & pi63;
  assign new_new_n18626__ = ~new_new_n18624__ & ~new_new_n18625__;
  assign new_new_n18627__ = pi42 & ~pi52;
  assign new_new_n18628__ = new_new_n18626__ & ~new_new_n18627__;
  assign new_new_n18629__ = ~new_new_n17141__ & ~new_new_n18626__;
  assign new_new_n18630__ = pi62 & ~new_new_n18628__;
  assign new_new_n18631__ = ~new_new_n18629__ & new_new_n18630__;
  assign new_new_n18632__ = pi51 & pi52;
  assign new_new_n18633__ = pi41 & pi63;
  assign new_new_n18634__ = ~new_new_n18632__ & ~new_new_n18633__;
  assign new_new_n18635__ = ~pi62 & ~new_new_n18633__;
  assign new_new_n18636__ = ~pi42 & ~new_new_n17141__;
  assign new_new_n18637__ = ~new_new_n18635__ & ~new_new_n18636__;
  assign new_new_n18638__ = ~new_new_n18634__ & ~new_new_n18637__;
  assign new_new_n18639__ = ~pi42 & ~new_new_n18633__;
  assign new_new_n18640__ = ~new_new_n18635__ & ~new_new_n18639__;
  assign new_new_n18641__ = ~new_new_n14927__ & ~new_new_n18632__;
  assign new_new_n18642__ = new_new_n18640__ & new_new_n18641__;
  assign new_new_n18643__ = ~new_new_n18638__ & ~new_new_n18642__;
  assign new_new_n18644__ = ~new_new_n18631__ & new_new_n18643__;
  assign new_new_n18645__ = ~new_new_n18522__ & ~new_new_n18527__;
  assign new_new_n18646__ = ~new_new_n18528__ & ~new_new_n18645__;
  assign new_new_n18647__ = new_new_n18644__ & ~new_new_n18646__;
  assign new_new_n18648__ = ~new_new_n18644__ & new_new_n18646__;
  assign new_new_n18649__ = ~new_new_n18647__ & ~new_new_n18648__;
  assign new_new_n18650__ = ~new_new_n18541__ & ~new_new_n18551__;
  assign new_new_n18651__ = ~new_new_n18540__ & ~new_new_n18650__;
  assign new_new_n18652__ = new_new_n18649__ & new_new_n18651__;
  assign new_new_n18653__ = ~new_new_n18649__ & ~new_new_n18651__;
  assign new_new_n18654__ = ~new_new_n18652__ & ~new_new_n18653__;
  assign new_new_n18655__ = ~new_new_n18623__ & ~new_new_n18654__;
  assign new_new_n18656__ = new_new_n18623__ & new_new_n18654__;
  assign new_new_n18657__ = ~new_new_n18655__ & ~new_new_n18656__;
  assign new_new_n18658__ = ~new_new_n18575__ & ~new_new_n18578__;
  assign new_new_n18659__ = ~new_new_n18574__ & ~new_new_n18658__;
  assign new_new_n18660__ = new_new_n18657__ & ~new_new_n18659__;
  assign new_new_n18661__ = ~new_new_n18657__ & new_new_n18659__;
  assign new_new_n18662__ = ~new_new_n18660__ & ~new_new_n18661__;
  assign new_new_n18663__ = ~new_new_n18621__ & ~new_new_n18662__;
  assign new_new_n18664__ = new_new_n18621__ & new_new_n18662__;
  assign new_new_n18665__ = ~new_new_n18663__ & ~new_new_n18664__;
  assign new_new_n18666__ = ~new_new_n18543__ & ~new_new_n18547__;
  assign new_new_n18667__ = ~new_new_n18546__ & ~new_new_n18666__;
  assign new_new_n18668__ = ~new_new_n18498__ & ~new_new_n18502__;
  assign new_new_n18669__ = ~new_new_n18501__ & ~new_new_n18668__;
  assign new_new_n18670__ = ~new_new_n18507__ & ~new_new_n18511__;
  assign new_new_n18671__ = ~new_new_n18510__ & ~new_new_n18670__;
  assign new_new_n18672__ = ~new_new_n18669__ & ~new_new_n18671__;
  assign new_new_n18673__ = new_new_n18669__ & new_new_n18671__;
  assign new_new_n18674__ = ~new_new_n18672__ & ~new_new_n18673__;
  assign new_new_n18675__ = new_new_n18667__ & ~new_new_n18674__;
  assign new_new_n18676__ = ~new_new_n18667__ & new_new_n18674__;
  assign new_new_n18677__ = ~new_new_n18675__ & ~new_new_n18676__;
  assign new_new_n18678__ = ~new_new_n18497__ & ~new_new_n18516__;
  assign new_new_n18679__ = ~new_new_n18517__ & ~new_new_n18678__;
  assign new_new_n18680__ = pi45 & pi59;
  assign new_new_n18681__ = pi44 & pi60;
  assign new_new_n18682__ = pi43 & pi61;
  assign new_new_n18683__ = ~new_new_n18681__ & ~new_new_n18682__;
  assign new_new_n18684__ = new_new_n18681__ & new_new_n18682__;
  assign new_new_n18685__ = ~new_new_n18683__ & ~new_new_n18684__;
  assign new_new_n18686__ = new_new_n18680__ & ~new_new_n18685__;
  assign new_new_n18687__ = ~new_new_n18680__ & new_new_n18685__;
  assign new_new_n18688__ = ~new_new_n18686__ & ~new_new_n18687__;
  assign new_new_n18689__ = pi51 & pi53;
  assign new_new_n18690__ = pi49 & pi55;
  assign new_new_n18691__ = pi50 & pi54;
  assign new_new_n18692__ = ~new_new_n18690__ & ~new_new_n18691__;
  assign new_new_n18693__ = new_new_n18690__ & new_new_n18691__;
  assign new_new_n18694__ = ~new_new_n18692__ & ~new_new_n18693__;
  assign new_new_n18695__ = new_new_n18689__ & ~new_new_n18694__;
  assign new_new_n18696__ = ~new_new_n18689__ & new_new_n18694__;
  assign new_new_n18697__ = ~new_new_n18695__ & ~new_new_n18696__;
  assign new_new_n18698__ = ~new_new_n18688__ & ~new_new_n18697__;
  assign new_new_n18699__ = new_new_n18688__ & new_new_n18697__;
  assign new_new_n18700__ = ~new_new_n18698__ & ~new_new_n18699__;
  assign new_new_n18701__ = pi48 & pi56;
  assign new_new_n18702__ = pi47 & pi57;
  assign new_new_n18703__ = pi46 & pi58;
  assign new_new_n18704__ = ~new_new_n18702__ & ~new_new_n18703__;
  assign new_new_n18705__ = new_new_n18702__ & new_new_n18703__;
  assign new_new_n18706__ = ~new_new_n18704__ & ~new_new_n18705__;
  assign new_new_n18707__ = new_new_n18701__ & ~new_new_n18706__;
  assign new_new_n18708__ = ~new_new_n18701__ & new_new_n18706__;
  assign new_new_n18709__ = ~new_new_n18707__ & ~new_new_n18708__;
  assign new_new_n18710__ = ~new_new_n18700__ & new_new_n18709__;
  assign new_new_n18711__ = new_new_n18700__ & ~new_new_n18709__;
  assign new_new_n18712__ = ~new_new_n18710__ & ~new_new_n18711__;
  assign new_new_n18713__ = new_new_n18679__ & ~new_new_n18712__;
  assign new_new_n18714__ = ~new_new_n18679__ & new_new_n18712__;
  assign new_new_n18715__ = ~new_new_n18713__ & ~new_new_n18714__;
  assign new_new_n18716__ = new_new_n18677__ & new_new_n18715__;
  assign new_new_n18717__ = ~new_new_n18677__ & ~new_new_n18715__;
  assign new_new_n18718__ = ~new_new_n18716__ & ~new_new_n18717__;
  assign new_new_n18719__ = new_new_n18665__ & ~new_new_n18718__;
  assign new_new_n18720__ = ~new_new_n18665__ & new_new_n18718__;
  assign new_new_n18721__ = ~new_new_n18719__ & ~new_new_n18720__;
  assign new_new_n18722__ = new_new_n18619__ & new_new_n18721__;
  assign new_new_n18723__ = ~new_new_n18619__ & ~new_new_n18721__;
  assign po105 = ~new_new_n18722__ & ~new_new_n18723__;
  assign new_new_n18725__ = ~new_new_n18699__ & ~new_new_n18709__;
  assign new_new_n18726__ = ~new_new_n18698__ & ~new_new_n18725__;
  assign new_new_n18727__ = ~new_new_n18647__ & ~new_new_n18651__;
  assign new_new_n18728__ = ~new_new_n18648__ & ~new_new_n18727__;
  assign new_new_n18729__ = ~new_new_n18726__ & ~new_new_n18728__;
  assign new_new_n18730__ = new_new_n18726__ & new_new_n18728__;
  assign new_new_n18731__ = ~new_new_n18729__ & ~new_new_n18730__;
  assign new_new_n18732__ = ~new_new_n18689__ & ~new_new_n18693__;
  assign new_new_n18733__ = ~new_new_n18692__ & ~new_new_n18732__;
  assign new_new_n18734__ = ~new_new_n18680__ & ~new_new_n18684__;
  assign new_new_n18735__ = ~new_new_n18683__ & ~new_new_n18734__;
  assign new_new_n18736__ = ~new_new_n18701__ & ~new_new_n18705__;
  assign new_new_n18737__ = ~new_new_n18704__ & ~new_new_n18736__;
  assign new_new_n18738__ = new_new_n18735__ & new_new_n18737__;
  assign new_new_n18739__ = ~new_new_n18735__ & ~new_new_n18737__;
  assign new_new_n18740__ = ~new_new_n18738__ & ~new_new_n18739__;
  assign new_new_n18741__ = new_new_n18733__ & ~new_new_n18740__;
  assign new_new_n18742__ = ~new_new_n18733__ & new_new_n18740__;
  assign new_new_n18743__ = ~new_new_n18741__ & ~new_new_n18742__;
  assign new_new_n18744__ = new_new_n18731__ & new_new_n18743__;
  assign new_new_n18745__ = ~new_new_n18731__ & ~new_new_n18743__;
  assign new_new_n18746__ = ~new_new_n18744__ & ~new_new_n18745__;
  assign new_new_n18747__ = ~new_new_n18667__ & ~new_new_n18673__;
  assign new_new_n18748__ = ~new_new_n18672__ & ~new_new_n18747__;
  assign new_new_n18749__ = pi51 & pi54;
  assign new_new_n18750__ = pi50 & pi55;
  assign new_new_n18751__ = pi49 & pi56;
  assign new_new_n18752__ = ~new_new_n18750__ & ~new_new_n18751__;
  assign new_new_n18753__ = new_new_n18750__ & new_new_n18751__;
  assign new_new_n18754__ = ~new_new_n18752__ & ~new_new_n18753__;
  assign new_new_n18755__ = new_new_n18749__ & ~new_new_n18754__;
  assign new_new_n18756__ = ~new_new_n18749__ & new_new_n18754__;
  assign new_new_n18757__ = ~new_new_n18755__ & ~new_new_n18756__;
  assign new_new_n18758__ = ~new_new_n18748__ & new_new_n18757__;
  assign new_new_n18759__ = new_new_n18748__ & ~new_new_n18757__;
  assign new_new_n18760__ = ~new_new_n18758__ & ~new_new_n18759__;
  assign new_new_n18761__ = pi43 & pi62;
  assign new_new_n18762__ = ~pi52 & pi53;
  assign new_new_n18763__ = new_new_n18761__ & ~new_new_n18762__;
  assign new_new_n18764__ = ~new_new_n18761__ & new_new_n18762__;
  assign new_new_n18765__ = ~new_new_n18763__ & ~new_new_n18764__;
  assign new_new_n18766__ = new_new_n18760__ & ~new_new_n18765__;
  assign new_new_n18767__ = ~new_new_n18760__ & new_new_n18765__;
  assign new_new_n18768__ = ~new_new_n18766__ & ~new_new_n18767__;
  assign new_new_n18769__ = ~new_new_n18677__ & ~new_new_n18713__;
  assign new_new_n18770__ = ~new_new_n18714__ & ~new_new_n18769__;
  assign new_new_n18771__ = ~new_new_n18768__ & new_new_n18770__;
  assign new_new_n18772__ = new_new_n18768__ & ~new_new_n18770__;
  assign new_new_n18773__ = ~new_new_n18771__ & ~new_new_n18772__;
  assign new_new_n18774__ = new_new_n14927__ & new_new_n18625__;
  assign new_new_n18775__ = new_new_n14927__ & ~new_new_n18624__;
  assign new_new_n18776__ = pi51 & new_new_n18640__;
  assign new_new_n18777__ = ~new_new_n18775__ & ~new_new_n18776__;
  assign new_new_n18778__ = pi52 & ~new_new_n18777__;
  assign new_new_n18779__ = ~new_new_n18774__ & ~new_new_n18778__;
  assign new_new_n18780__ = pi48 & pi57;
  assign new_new_n18781__ = pi47 & pi58;
  assign new_new_n18782__ = pi46 & pi59;
  assign new_new_n18783__ = ~new_new_n18781__ & ~new_new_n18782__;
  assign new_new_n18784__ = new_new_n18781__ & new_new_n18782__;
  assign new_new_n18785__ = ~new_new_n18783__ & ~new_new_n18784__;
  assign new_new_n18786__ = new_new_n18780__ & ~new_new_n18785__;
  assign new_new_n18787__ = ~new_new_n18780__ & new_new_n18785__;
  assign new_new_n18788__ = ~new_new_n18786__ & ~new_new_n18787__;
  assign new_new_n18789__ = new_new_n18779__ & new_new_n18788__;
  assign new_new_n18790__ = ~new_new_n18779__ & ~new_new_n18788__;
  assign new_new_n18791__ = ~new_new_n18789__ & ~new_new_n18790__;
  assign new_new_n18792__ = pi45 & pi60;
  assign new_new_n18793__ = pi44 & pi61;
  assign new_new_n18794__ = ~new_new_n18625__ & ~new_new_n18793__;
  assign new_new_n18795__ = new_new_n18625__ & new_new_n18793__;
  assign new_new_n18796__ = ~new_new_n18794__ & ~new_new_n18795__;
  assign new_new_n18797__ = new_new_n18792__ & ~new_new_n18796__;
  assign new_new_n18798__ = ~new_new_n18792__ & new_new_n18796__;
  assign new_new_n18799__ = ~new_new_n18797__ & ~new_new_n18798__;
  assign new_new_n18800__ = ~new_new_n18791__ & new_new_n18799__;
  assign new_new_n18801__ = new_new_n18791__ & ~new_new_n18799__;
  assign new_new_n18802__ = ~new_new_n18800__ & ~new_new_n18801__;
  assign new_new_n18803__ = new_new_n18773__ & new_new_n18802__;
  assign new_new_n18804__ = ~new_new_n18773__ & ~new_new_n18802__;
  assign new_new_n18805__ = ~new_new_n18803__ & ~new_new_n18804__;
  assign new_new_n18806__ = ~new_new_n18746__ & new_new_n18805__;
  assign new_new_n18807__ = ~new_new_n18655__ & new_new_n18659__;
  assign new_new_n18808__ = new_new_n18746__ & ~new_new_n18805__;
  assign new_new_n18809__ = ~new_new_n18656__ & ~new_new_n18807__;
  assign new_new_n18810__ = ~new_new_n18808__ & new_new_n18809__;
  assign new_new_n18811__ = ~new_new_n18806__ & new_new_n18810__;
  assign new_new_n18812__ = new_new_n18623__ & new_new_n18808__;
  assign new_new_n18813__ = new_new_n18659__ & new_new_n18806__;
  assign new_new_n18814__ = ~new_new_n18812__ & ~new_new_n18813__;
  assign new_new_n18815__ = new_new_n18654__ & ~new_new_n18814__;
  assign new_new_n18816__ = new_new_n18623__ & new_new_n18806__;
  assign new_new_n18817__ = new_new_n18659__ & new_new_n18808__;
  assign new_new_n18818__ = ~new_new_n18816__ & ~new_new_n18817__;
  assign new_new_n18819__ = new_new_n18662__ & ~new_new_n18818__;
  assign new_new_n18820__ = ~new_new_n18811__ & ~new_new_n18815__;
  assign new_new_n18821__ = ~new_new_n18819__ & new_new_n18820__;
  assign new_new_n18822__ = new_new_n18663__ & new_new_n18718__;
  assign new_new_n18823__ = new_new_n18664__ & ~new_new_n18718__;
  assign new_new_n18824__ = ~new_new_n18822__ & ~new_new_n18823__;
  assign new_new_n18825__ = new_new_n18619__ & new_new_n18824__;
  assign new_new_n18826__ = ~new_new_n18663__ & ~new_new_n18718__;
  assign new_new_n18827__ = ~new_new_n18664__ & ~new_new_n18826__;
  assign new_new_n18828__ = new_new_n18617__ & ~new_new_n18827__;
  assign new_new_n18829__ = new_new_n18618__ & new_new_n18827__;
  assign new_new_n18830__ = ~new_new_n18828__ & ~new_new_n18829__;
  assign new_new_n18831__ = ~new_new_n18825__ & new_new_n18830__;
  assign new_new_n18832__ = ~new_new_n18821__ & ~new_new_n18831__;
  assign new_new_n18833__ = ~new_new_n18617__ & new_new_n18621__;
  assign new_new_n18834__ = ~new_new_n18618__ & ~new_new_n18833__;
  assign new_new_n18835__ = new_new_n18662__ & ~new_new_n18834__;
  assign new_new_n18836__ = new_new_n18618__ & new_new_n18621__;
  assign new_new_n18837__ = ~new_new_n18835__ & ~new_new_n18836__;
  assign new_new_n18838__ = ~new_new_n18718__ & ~new_new_n18837__;
  assign new_new_n18839__ = ~new_new_n18662__ & new_new_n18834__;
  assign new_new_n18840__ = new_new_n18617__ & ~new_new_n18621__;
  assign new_new_n18841__ = ~new_new_n18839__ & ~new_new_n18840__;
  assign new_new_n18842__ = new_new_n18718__ & ~new_new_n18841__;
  assign new_new_n18843__ = ~new_new_n18616__ & new_new_n18662__;
  assign new_new_n18844__ = ~new_new_n18663__ & ~new_new_n18843__;
  assign new_new_n18845__ = ~new_new_n18614__ & new_new_n18621__;
  assign new_new_n18846__ = ~new_new_n18617__ & ~new_new_n18845__;
  assign new_new_n18847__ = ~new_new_n18844__ & ~new_new_n18846__;
  assign new_new_n18848__ = ~new_new_n18838__ & ~new_new_n18847__;
  assign new_new_n18849__ = ~new_new_n18842__ & new_new_n18848__;
  assign new_new_n18850__ = new_new_n18821__ & ~new_new_n18849__;
  assign po106 = new_new_n18832__ | new_new_n18850__;
  assign new_new_n18852__ = ~new_new_n18806__ & ~new_new_n18810__;
  assign new_new_n18853__ = new_new_n18616__ & ~new_new_n18662__;
  assign new_new_n18854__ = new_new_n18718__ & ~new_new_n18843__;
  assign new_new_n18855__ = ~new_new_n18853__ & ~new_new_n18854__;
  assign new_new_n18856__ = ~new_new_n18821__ & ~new_new_n18855__;
  assign new_new_n18857__ = new_new_n18821__ & new_new_n18855__;
  assign new_new_n18858__ = ~new_new_n18621__ & ~new_new_n18857__;
  assign new_new_n18859__ = new_new_n18614__ & new_new_n18858__;
  assign new_new_n18860__ = new_new_n18821__ & ~new_new_n18853__;
  assign new_new_n18861__ = ~new_new_n18821__ & ~new_new_n18843__;
  assign new_new_n18862__ = ~new_new_n18718__ & ~new_new_n18861__;
  assign new_new_n18863__ = ~new_new_n18860__ & ~new_new_n18862__;
  assign new_new_n18864__ = ~new_new_n18845__ & new_new_n18863__;
  assign new_new_n18865__ = ~new_new_n18856__ & ~new_new_n18859__;
  assign new_new_n18866__ = ~new_new_n18864__ & new_new_n18865__;
  assign new_new_n18867__ = ~new_new_n18852__ & new_new_n18866__;
  assign new_new_n18868__ = new_new_n18852__ & ~new_new_n18866__;
  assign new_new_n18869__ = ~new_new_n18867__ & ~new_new_n18868__;
  assign new_new_n18870__ = ~new_new_n18730__ & ~new_new_n18743__;
  assign new_new_n18871__ = ~new_new_n18729__ & ~new_new_n18870__;
  assign new_new_n18872__ = ~new_new_n18733__ & ~new_new_n18738__;
  assign new_new_n18873__ = ~new_new_n18739__ & ~new_new_n18872__;
  assign new_new_n18874__ = pi52 & pi54;
  assign new_new_n18875__ = pi50 & pi56;
  assign new_new_n18876__ = pi51 & pi55;
  assign new_new_n18877__ = ~new_new_n18875__ & ~new_new_n18876__;
  assign new_new_n18878__ = new_new_n18875__ & new_new_n18876__;
  assign new_new_n18879__ = ~new_new_n18877__ & ~new_new_n18878__;
  assign new_new_n18880__ = new_new_n18874__ & ~new_new_n18879__;
  assign new_new_n18881__ = ~new_new_n18874__ & new_new_n18879__;
  assign new_new_n18882__ = ~new_new_n18880__ & ~new_new_n18881__;
  assign new_new_n18883__ = pi49 & pi57;
  assign new_new_n18884__ = pi47 & pi59;
  assign new_new_n18885__ = pi48 & pi58;
  assign new_new_n18886__ = ~new_new_n18884__ & ~new_new_n18885__;
  assign new_new_n18887__ = new_new_n18884__ & new_new_n18885__;
  assign new_new_n18888__ = ~new_new_n18886__ & ~new_new_n18887__;
  assign new_new_n18889__ = new_new_n18883__ & ~new_new_n18888__;
  assign new_new_n18890__ = ~new_new_n18883__ & new_new_n18888__;
  assign new_new_n18891__ = ~new_new_n18889__ & ~new_new_n18890__;
  assign new_new_n18892__ = new_new_n18882__ & new_new_n18891__;
  assign new_new_n18893__ = ~new_new_n18882__ & ~new_new_n18891__;
  assign new_new_n18894__ = ~new_new_n18892__ & ~new_new_n18893__;
  assign new_new_n18895__ = new_new_n18873__ & ~new_new_n18894__;
  assign new_new_n18896__ = ~new_new_n18873__ & new_new_n18894__;
  assign new_new_n18897__ = ~new_new_n18895__ & ~new_new_n18896__;
  assign new_new_n18898__ = ~new_new_n18871__ & ~new_new_n18897__;
  assign new_new_n18899__ = new_new_n18871__ & new_new_n18897__;
  assign new_new_n18900__ = ~new_new_n18898__ & ~new_new_n18899__;
  assign new_new_n18901__ = ~new_new_n18780__ & ~new_new_n18784__;
  assign new_new_n18902__ = ~new_new_n18783__ & ~new_new_n18901__;
  assign new_new_n18903__ = pi46 & pi60;
  assign new_new_n18904__ = pi45 & pi61;
  assign new_new_n18905__ = ~new_new_n16196__ & ~new_new_n18904__;
  assign new_new_n18906__ = new_new_n16196__ & new_new_n18904__;
  assign new_new_n18907__ = ~new_new_n18905__ & ~new_new_n18906__;
  assign new_new_n18908__ = new_new_n18903__ & ~new_new_n18907__;
  assign new_new_n18909__ = ~new_new_n18903__ & new_new_n18907__;
  assign new_new_n18910__ = ~new_new_n18908__ & ~new_new_n18909__;
  assign new_new_n18911__ = ~new_new_n18792__ & ~new_new_n18795__;
  assign new_new_n18912__ = ~new_new_n18794__ & ~new_new_n18911__;
  assign new_new_n18913__ = new_new_n18910__ & ~new_new_n18912__;
  assign new_new_n18914__ = ~new_new_n18910__ & new_new_n18912__;
  assign new_new_n18915__ = new_new_n18902__ & ~new_new_n18913__;
  assign new_new_n18916__ = ~new_new_n18914__ & ~new_new_n18915__;
  assign new_new_n18917__ = ~new_new_n18913__ & new_new_n18916__;
  assign new_new_n18918__ = ~new_new_n18902__ & ~new_new_n18917__;
  assign new_new_n18919__ = ~new_new_n18914__ & new_new_n18915__;
  assign new_new_n18920__ = ~new_new_n18918__ & ~new_new_n18919__;
  assign new_new_n18921__ = new_new_n18900__ & ~new_new_n18920__;
  assign new_new_n18922__ = ~new_new_n18900__ & new_new_n18920__;
  assign new_new_n18923__ = ~new_new_n18921__ & ~new_new_n18922__;
  assign new_new_n18924__ = pi43 & pi63;
  assign new_new_n18925__ = ~new_new_n18749__ & ~new_new_n18753__;
  assign new_new_n18926__ = ~new_new_n18752__ & ~new_new_n18925__;
  assign new_new_n18927__ = ~new_new_n18924__ & new_new_n18926__;
  assign new_new_n18928__ = ~pi43 & pi52;
  assign new_new_n18929__ = pi63 & ~new_new_n18926__;
  assign new_new_n18930__ = ~new_new_n18928__ & new_new_n18929__;
  assign new_new_n18931__ = ~new_new_n18927__ & ~new_new_n18930__;
  assign new_new_n18932__ = ~pi43 & new_new_n18926__;
  assign new_new_n18933__ = pi62 & ~new_new_n18932__;
  assign new_new_n18934__ = ~pi52 & ~new_new_n18933__;
  assign new_new_n18935__ = pi53 & ~new_new_n18931__;
  assign new_new_n18936__ = ~new_new_n18934__ & new_new_n18935__;
  assign new_new_n18937__ = pi53 & pi62;
  assign new_new_n18938__ = ~new_new_n18929__ & ~new_new_n18937__;
  assign new_new_n18939__ = pi43 & ~new_new_n18938__;
  assign new_new_n18940__ = pi52 & pi53;
  assign new_new_n18941__ = ~new_new_n18927__ & ~new_new_n18940__;
  assign new_new_n18942__ = ~new_new_n18939__ & new_new_n18941__;
  assign new_new_n18943__ = ~new_new_n18936__ & ~new_new_n18942__;
  assign new_new_n18944__ = ~new_new_n18758__ & ~new_new_n18765__;
  assign new_new_n18945__ = ~new_new_n18759__ & ~new_new_n18944__;
  assign new_new_n18946__ = ~new_new_n18943__ & new_new_n18945__;
  assign new_new_n18947__ = new_new_n18943__ & ~new_new_n18945__;
  assign new_new_n18948__ = ~new_new_n18946__ & ~new_new_n18947__;
  assign new_new_n18949__ = ~new_new_n18790__ & new_new_n18799__;
  assign new_new_n18950__ = ~new_new_n18789__ & ~new_new_n18949__;
  assign new_new_n18951__ = new_new_n18948__ & new_new_n18950__;
  assign new_new_n18952__ = ~new_new_n18948__ & ~new_new_n18950__;
  assign new_new_n18953__ = ~new_new_n18951__ & ~new_new_n18952__;
  assign new_new_n18954__ = new_new_n18923__ & ~new_new_n18953__;
  assign new_new_n18955__ = ~new_new_n18923__ & new_new_n18953__;
  assign new_new_n18956__ = ~new_new_n18954__ & ~new_new_n18955__;
  assign new_new_n18957__ = ~new_new_n18772__ & ~new_new_n18802__;
  assign new_new_n18958__ = ~new_new_n18771__ & ~new_new_n18957__;
  assign new_new_n18959__ = new_new_n18956__ & new_new_n18958__;
  assign new_new_n18960__ = ~new_new_n18956__ & ~new_new_n18958__;
  assign new_new_n18961__ = ~new_new_n18959__ & ~new_new_n18960__;
  assign new_new_n18962__ = new_new_n18869__ & new_new_n18961__;
  assign new_new_n18963__ = ~new_new_n18869__ & ~new_new_n18961__;
  assign po107 = ~new_new_n18962__ & ~new_new_n18963__;
  assign new_new_n18965__ = new_new_n18873__ & ~new_new_n18892__;
  assign new_new_n18966__ = ~new_new_n18893__ & ~new_new_n18965__;
  assign new_new_n18967__ = ~pi52 & ~new_new_n18761__;
  assign new_new_n18968__ = pi53 & ~new_new_n18967__;
  assign new_new_n18969__ = new_new_n18924__ & new_new_n18968__;
  assign new_new_n18970__ = ~new_new_n18926__ & ~new_new_n18969__;
  assign new_new_n18971__ = ~new_new_n18924__ & ~new_new_n18968__;
  assign new_new_n18972__ = ~new_new_n18970__ & ~new_new_n18971__;
  assign new_new_n18973__ = ~new_new_n18966__ & new_new_n18972__;
  assign new_new_n18974__ = new_new_n18966__ & ~new_new_n18972__;
  assign new_new_n18975__ = ~new_new_n18973__ & ~new_new_n18974__;
  assign new_new_n18976__ = ~new_new_n18916__ & ~new_new_n18975__;
  assign new_new_n18977__ = new_new_n18916__ & new_new_n18975__;
  assign new_new_n18978__ = ~new_new_n18976__ & ~new_new_n18977__;
  assign new_new_n18979__ = ~new_new_n18947__ & ~new_new_n18950__;
  assign new_new_n18980__ = ~new_new_n18946__ & ~new_new_n18979__;
  assign new_new_n18981__ = ~new_new_n18874__ & ~new_new_n18878__;
  assign new_new_n18982__ = ~new_new_n18877__ & ~new_new_n18981__;
  assign new_new_n18983__ = pi47 & pi60;
  assign new_new_n18984__ = pi46 & pi61;
  assign new_new_n18985__ = ~new_new_n18983__ & ~new_new_n18984__;
  assign new_new_n18986__ = new_new_n18983__ & new_new_n18984__;
  assign new_new_n18987__ = ~new_new_n18985__ & ~new_new_n18986__;
  assign new_new_n18988__ = new_new_n18982__ & ~new_new_n18987__;
  assign new_new_n18989__ = ~new_new_n18982__ & new_new_n18987__;
  assign new_new_n18990__ = ~new_new_n18988__ & ~new_new_n18989__;
  assign new_new_n18991__ = pi52 & pi55;
  assign new_new_n18992__ = pi51 & pi56;
  assign new_new_n18993__ = pi50 & pi57;
  assign new_new_n18994__ = ~new_new_n18992__ & ~new_new_n18993__;
  assign new_new_n18995__ = new_new_n18992__ & new_new_n18993__;
  assign new_new_n18996__ = ~new_new_n18994__ & ~new_new_n18995__;
  assign new_new_n18997__ = new_new_n18991__ & ~new_new_n18996__;
  assign new_new_n18998__ = ~new_new_n18991__ & new_new_n18996__;
  assign new_new_n18999__ = ~new_new_n18997__ & ~new_new_n18998__;
  assign new_new_n19000__ = new_new_n18990__ & new_new_n18999__;
  assign new_new_n19001__ = ~new_new_n18990__ & ~new_new_n18999__;
  assign new_new_n19002__ = ~new_new_n19000__ & ~new_new_n19001__;
  assign new_new_n19003__ = pi45 & pi62;
  assign new_new_n19004__ = ~pi53 & pi54;
  assign new_new_n19005__ = new_new_n19003__ & ~new_new_n19004__;
  assign new_new_n19006__ = ~new_new_n19003__ & new_new_n19004__;
  assign new_new_n19007__ = ~new_new_n19005__ & ~new_new_n19006__;
  assign new_new_n19008__ = ~new_new_n19002__ & new_new_n19007__;
  assign new_new_n19009__ = new_new_n19002__ & ~new_new_n19007__;
  assign new_new_n19010__ = ~new_new_n19008__ & ~new_new_n19009__;
  assign new_new_n19011__ = new_new_n18980__ & new_new_n19010__;
  assign new_new_n19012__ = ~new_new_n18980__ & ~new_new_n19010__;
  assign new_new_n19013__ = ~new_new_n19011__ & ~new_new_n19012__;
  assign new_new_n19014__ = ~new_new_n18903__ & ~new_new_n18906__;
  assign new_new_n19015__ = ~new_new_n18905__ & ~new_new_n19014__;
  assign new_new_n19016__ = ~new_new_n18883__ & ~new_new_n18887__;
  assign new_new_n19017__ = ~new_new_n18886__ & ~new_new_n19016__;
  assign new_new_n19018__ = ~new_new_n19015__ & ~new_new_n19017__;
  assign new_new_n19019__ = new_new_n19015__ & new_new_n19017__;
  assign new_new_n19020__ = ~new_new_n19018__ & ~new_new_n19019__;
  assign new_new_n19021__ = pi49 & pi58;
  assign new_new_n19022__ = pi44 & pi63;
  assign new_new_n19023__ = pi48 & pi59;
  assign new_new_n19024__ = ~new_new_n19022__ & ~new_new_n19023__;
  assign new_new_n19025__ = new_new_n19022__ & new_new_n19023__;
  assign new_new_n19026__ = ~new_new_n19024__ & ~new_new_n19025__;
  assign new_new_n19027__ = new_new_n19021__ & ~new_new_n19026__;
  assign new_new_n19028__ = ~new_new_n19021__ & new_new_n19026__;
  assign new_new_n19029__ = ~new_new_n19027__ & ~new_new_n19028__;
  assign new_new_n19030__ = new_new_n19020__ & ~new_new_n19029__;
  assign new_new_n19031__ = ~new_new_n19020__ & new_new_n19029__;
  assign new_new_n19032__ = ~new_new_n19030__ & ~new_new_n19031__;
  assign new_new_n19033__ = new_new_n19013__ & ~new_new_n19032__;
  assign new_new_n19034__ = ~new_new_n19013__ & new_new_n19032__;
  assign new_new_n19035__ = ~new_new_n19033__ & ~new_new_n19034__;
  assign new_new_n19036__ = new_new_n18978__ & new_new_n19035__;
  assign new_new_n19037__ = ~new_new_n18978__ & ~new_new_n19035__;
  assign new_new_n19038__ = ~new_new_n19036__ & ~new_new_n19037__;
  assign new_new_n19039__ = ~new_new_n18955__ & ~new_new_n18958__;
  assign new_new_n19040__ = ~new_new_n18954__ & ~new_new_n19039__;
  assign new_new_n19041__ = ~new_new_n18867__ & ~new_new_n18961__;
  assign new_new_n19042__ = ~new_new_n18868__ & ~new_new_n19041__;
  assign new_new_n19043__ = new_new_n19040__ & new_new_n19042__;
  assign new_new_n19044__ = ~new_new_n19040__ & ~new_new_n19042__;
  assign new_new_n19045__ = ~new_new_n19043__ & ~new_new_n19044__;
  assign new_new_n19046__ = ~new_new_n18899__ & new_new_n18920__;
  assign new_new_n19047__ = ~new_new_n18898__ & ~new_new_n19046__;
  assign new_new_n19048__ = new_new_n19045__ & ~new_new_n19047__;
  assign new_new_n19049__ = ~new_new_n19045__ & new_new_n19047__;
  assign new_new_n19050__ = ~new_new_n19048__ & ~new_new_n19049__;
  assign new_new_n19051__ = new_new_n19038__ & ~new_new_n19050__;
  assign new_new_n19052__ = ~new_new_n19038__ & new_new_n19050__;
  assign po108 = new_new_n19051__ | new_new_n19052__;
  assign new_new_n19054__ = ~new_new_n19012__ & new_new_n19032__;
  assign new_new_n19055__ = ~new_new_n19011__ & ~new_new_n19054__;
  assign new_new_n19056__ = ~pi53 & ~new_new_n19003__;
  assign new_new_n19057__ = pi54 & ~new_new_n19056__;
  assign new_new_n19058__ = ~new_new_n19021__ & ~new_new_n19025__;
  assign new_new_n19059__ = ~new_new_n19024__ & ~new_new_n19058__;
  assign new_new_n19060__ = ~new_new_n18991__ & ~new_new_n18995__;
  assign new_new_n19061__ = ~new_new_n18994__ & ~new_new_n19060__;
  assign new_new_n19062__ = ~new_new_n19059__ & ~new_new_n19061__;
  assign new_new_n19063__ = new_new_n19059__ & new_new_n19061__;
  assign new_new_n19064__ = ~new_new_n19062__ & ~new_new_n19063__;
  assign new_new_n19065__ = new_new_n19057__ & ~new_new_n19064__;
  assign new_new_n19066__ = ~new_new_n19057__ & new_new_n19064__;
  assign new_new_n19067__ = ~new_new_n19065__ & ~new_new_n19066__;
  assign new_new_n19068__ = ~new_new_n18916__ & ~new_new_n18974__;
  assign new_new_n19069__ = ~new_new_n18973__ & ~new_new_n19068__;
  assign new_new_n19070__ = new_new_n19067__ & new_new_n19069__;
  assign new_new_n19071__ = ~new_new_n19067__ & ~new_new_n19069__;
  assign new_new_n19072__ = ~new_new_n19070__ & ~new_new_n19071__;
  assign new_new_n19073__ = pi50 & pi58;
  assign new_new_n19074__ = pi48 & pi60;
  assign new_new_n19075__ = pi49 & pi59;
  assign new_new_n19076__ = ~new_new_n19074__ & ~new_new_n19075__;
  assign new_new_n19077__ = new_new_n19074__ & new_new_n19075__;
  assign new_new_n19078__ = ~new_new_n19076__ & ~new_new_n19077__;
  assign new_new_n19079__ = new_new_n19073__ & ~new_new_n19078__;
  assign new_new_n19080__ = ~new_new_n19073__ & new_new_n19078__;
  assign new_new_n19081__ = ~new_new_n19079__ & ~new_new_n19080__;
  assign new_new_n19082__ = ~new_new_n18982__ & ~new_new_n18986__;
  assign new_new_n19083__ = ~new_new_n18985__ & ~new_new_n19082__;
  assign new_new_n19084__ = pi47 & pi61;
  assign new_new_n19085__ = pi45 & pi63;
  assign new_new_n19086__ = pi46 & pi62;
  assign new_new_n19087__ = ~new_new_n19085__ & ~new_new_n19086__;
  assign new_new_n19088__ = new_new_n19085__ & new_new_n19086__;
  assign new_new_n19089__ = ~new_new_n19087__ & ~new_new_n19088__;
  assign new_new_n19090__ = new_new_n19084__ & ~new_new_n19089__;
  assign new_new_n19091__ = ~new_new_n19084__ & new_new_n19089__;
  assign new_new_n19092__ = ~new_new_n19090__ & ~new_new_n19091__;
  assign new_new_n19093__ = ~new_new_n19083__ & new_new_n19092__;
  assign new_new_n19094__ = new_new_n19083__ & ~new_new_n19092__;
  assign new_new_n19095__ = ~new_new_n19093__ & ~new_new_n19094__;
  assign new_new_n19096__ = new_new_n19081__ & new_new_n19095__;
  assign new_new_n19097__ = ~new_new_n19081__ & ~new_new_n19095__;
  assign new_new_n19098__ = ~new_new_n19096__ & ~new_new_n19097__;
  assign new_new_n19099__ = new_new_n19072__ & new_new_n19098__;
  assign new_new_n19100__ = ~new_new_n19072__ & ~new_new_n19098__;
  assign new_new_n19101__ = ~new_new_n19099__ & ~new_new_n19100__;
  assign new_new_n19102__ = ~new_new_n19055__ & ~new_new_n19101__;
  assign new_new_n19103__ = new_new_n19055__ & new_new_n19101__;
  assign new_new_n19104__ = ~new_new_n19102__ & ~new_new_n19103__;
  assign new_new_n19105__ = pi53 & pi55;
  assign new_new_n19106__ = pi51 & pi57;
  assign new_new_n19107__ = pi52 & pi56;
  assign new_new_n19108__ = ~new_new_n19106__ & ~new_new_n19107__;
  assign new_new_n19109__ = new_new_n19106__ & new_new_n19107__;
  assign new_new_n19110__ = ~new_new_n19108__ & ~new_new_n19109__;
  assign new_new_n19111__ = new_new_n19105__ & ~new_new_n19110__;
  assign new_new_n19112__ = ~new_new_n19105__ & new_new_n19110__;
  assign new_new_n19113__ = ~new_new_n19111__ & ~new_new_n19112__;
  assign new_new_n19114__ = ~new_new_n19001__ & new_new_n19007__;
  assign new_new_n19115__ = ~new_new_n19000__ & ~new_new_n19114__;
  assign new_new_n19116__ = ~new_new_n19019__ & new_new_n19029__;
  assign new_new_n19117__ = ~new_new_n19018__ & ~new_new_n19116__;
  assign new_new_n19118__ = ~new_new_n19115__ & ~new_new_n19117__;
  assign new_new_n19119__ = new_new_n19115__ & new_new_n19117__;
  assign new_new_n19120__ = ~new_new_n19118__ & ~new_new_n19119__;
  assign new_new_n19121__ = new_new_n19113__ & new_new_n19120__;
  assign new_new_n19122__ = ~new_new_n19113__ & ~new_new_n19120__;
  assign new_new_n19123__ = ~new_new_n19121__ & ~new_new_n19122__;
  assign new_new_n19124__ = new_new_n19104__ & new_new_n19123__;
  assign new_new_n19125__ = ~new_new_n19104__ & ~new_new_n19123__;
  assign new_new_n19126__ = ~new_new_n19124__ & ~new_new_n19125__;
  assign new_new_n19127__ = ~new_new_n19037__ & ~new_new_n19043__;
  assign new_new_n19128__ = ~new_new_n19044__ & ~new_new_n19047__;
  assign new_new_n19129__ = ~new_new_n19127__ & new_new_n19128__;
  assign new_new_n19130__ = new_new_n19126__ & ~new_new_n19129__;
  assign new_new_n19131__ = new_new_n19045__ & new_new_n19047__;
  assign new_new_n19132__ = ~new_new_n19037__ & new_new_n19047__;
  assign new_new_n19133__ = new_new_n19044__ & ~new_new_n19132__;
  assign new_new_n19134__ = ~new_new_n19126__ & ~new_new_n19133__;
  assign new_new_n19135__ = ~new_new_n19131__ & new_new_n19134__;
  assign new_new_n19136__ = ~new_new_n19036__ & ~new_new_n19130__;
  assign new_new_n19137__ = ~new_new_n19135__ & new_new_n19136__;
  assign new_new_n19138__ = ~new_new_n19036__ & ~new_new_n19047__;
  assign new_new_n19139__ = new_new_n19043__ & ~new_new_n19138__;
  assign new_new_n19140__ = ~new_new_n19126__ & ~new_new_n19139__;
  assign new_new_n19141__ = ~new_new_n19048__ & new_new_n19140__;
  assign new_new_n19142__ = new_new_n19036__ & new_new_n19047__;
  assign new_new_n19143__ = ~new_new_n19043__ & new_new_n19142__;
  assign new_new_n19144__ = new_new_n19044__ & ~new_new_n19138__;
  assign new_new_n19145__ = new_new_n19126__ & ~new_new_n19143__;
  assign new_new_n19146__ = ~new_new_n19144__ & new_new_n19145__;
  assign new_new_n19147__ = ~new_new_n19037__ & ~new_new_n19141__;
  assign new_new_n19148__ = ~new_new_n19146__ & new_new_n19147__;
  assign new_new_n19149__ = new_new_n19037__ & new_new_n19047__;
  assign new_new_n19150__ = new_new_n19126__ & new_new_n19149__;
  assign new_new_n19151__ = new_new_n19043__ & new_new_n19150__;
  assign new_new_n19152__ = ~new_new_n19137__ & ~new_new_n19151__;
  assign po109 = ~new_new_n19148__ & new_new_n19152__;
  assign new_new_n19154__ = ~pi54 & pi55;
  assign new_new_n19155__ = ~new_new_n17234__ & new_new_n19154__;
  assign new_new_n19156__ = new_new_n17234__ & ~new_new_n19154__;
  assign new_new_n19157__ = ~new_new_n19155__ & ~new_new_n19156__;
  assign new_new_n19158__ = new_new_n19081__ & ~new_new_n19094__;
  assign new_new_n19159__ = ~new_new_n19093__ & ~new_new_n19158__;
  assign new_new_n19160__ = ~new_new_n19057__ & ~new_new_n19063__;
  assign new_new_n19161__ = ~new_new_n19062__ & ~new_new_n19160__;
  assign new_new_n19162__ = ~new_new_n19159__ & ~new_new_n19161__;
  assign new_new_n19163__ = new_new_n19159__ & new_new_n19161__;
  assign new_new_n19164__ = ~new_new_n19162__ & ~new_new_n19163__;
  assign new_new_n19165__ = new_new_n19157__ & new_new_n19164__;
  assign new_new_n19166__ = ~new_new_n19157__ & ~new_new_n19164__;
  assign new_new_n19167__ = ~new_new_n19165__ & ~new_new_n19166__;
  assign new_new_n19168__ = ~new_new_n19103__ & ~new_new_n19123__;
  assign new_new_n19169__ = ~new_new_n19102__ & ~new_new_n19168__;
  assign new_new_n19170__ = ~new_new_n19167__ & ~new_new_n19169__;
  assign new_new_n19171__ = new_new_n19167__ & new_new_n19169__;
  assign new_new_n19172__ = ~new_new_n19170__ & ~new_new_n19171__;
  assign new_new_n19173__ = ~new_new_n19113__ & ~new_new_n19118__;
  assign new_new_n19174__ = ~new_new_n19119__ & ~new_new_n19173__;
  assign new_new_n19175__ = pi50 & pi59;
  assign new_new_n19176__ = pi48 & pi61;
  assign new_new_n19177__ = pi49 & pi60;
  assign new_new_n19178__ = ~new_new_n19176__ & ~new_new_n19177__;
  assign new_new_n19179__ = new_new_n19176__ & new_new_n19177__;
  assign new_new_n19180__ = ~new_new_n19178__ & ~new_new_n19179__;
  assign new_new_n19181__ = new_new_n19175__ & ~new_new_n19180__;
  assign new_new_n19182__ = ~new_new_n19175__ & new_new_n19180__;
  assign new_new_n19183__ = ~new_new_n19181__ & ~new_new_n19182__;
  assign new_new_n19184__ = pi53 & pi56;
  assign new_new_n19185__ = pi52 & pi57;
  assign new_new_n19186__ = pi51 & pi58;
  assign new_new_n19187__ = ~new_new_n19185__ & ~new_new_n19186__;
  assign new_new_n19188__ = new_new_n19185__ & new_new_n19186__;
  assign new_new_n19189__ = ~new_new_n19187__ & ~new_new_n19188__;
  assign new_new_n19190__ = new_new_n19184__ & ~new_new_n19189__;
  assign new_new_n19191__ = ~new_new_n19184__ & new_new_n19189__;
  assign new_new_n19192__ = ~new_new_n19190__ & ~new_new_n19191__;
  assign new_new_n19193__ = new_new_n19183__ & new_new_n19192__;
  assign new_new_n19194__ = ~new_new_n19183__ & ~new_new_n19192__;
  assign new_new_n19195__ = ~new_new_n19193__ & ~new_new_n19194__;
  assign new_new_n19196__ = ~new_new_n19084__ & ~new_new_n19088__;
  assign new_new_n19197__ = ~new_new_n19087__ & ~new_new_n19196__;
  assign new_new_n19198__ = new_new_n19195__ & ~new_new_n19197__;
  assign new_new_n19199__ = ~new_new_n19195__ & new_new_n19197__;
  assign new_new_n19200__ = ~new_new_n19198__ & ~new_new_n19199__;
  assign new_new_n19201__ = ~new_new_n19174__ & ~new_new_n19200__;
  assign new_new_n19202__ = new_new_n19174__ & new_new_n19200__;
  assign new_new_n19203__ = ~new_new_n19201__ & ~new_new_n19202__;
  assign new_new_n19204__ = ~new_new_n19105__ & ~new_new_n19109__;
  assign new_new_n19205__ = ~new_new_n19108__ & ~new_new_n19204__;
  assign new_new_n19206__ = pi46 & pi63;
  assign new_new_n19207__ = ~new_new_n19073__ & ~new_new_n19077__;
  assign new_new_n19208__ = ~new_new_n19076__ & ~new_new_n19207__;
  assign new_new_n19209__ = new_new_n19206__ & ~new_new_n19208__;
  assign new_new_n19210__ = ~new_new_n19206__ & new_new_n19208__;
  assign new_new_n19211__ = ~new_new_n19209__ & ~new_new_n19210__;
  assign new_new_n19212__ = new_new_n19205__ & new_new_n19211__;
  assign new_new_n19213__ = ~new_new_n19205__ & ~new_new_n19211__;
  assign new_new_n19214__ = ~new_new_n19212__ & ~new_new_n19213__;
  assign new_new_n19215__ = new_new_n19203__ & new_new_n19214__;
  assign new_new_n19216__ = ~new_new_n19203__ & ~new_new_n19214__;
  assign new_new_n19217__ = ~new_new_n19215__ & ~new_new_n19216__;
  assign new_new_n19218__ = ~new_new_n19037__ & ~new_new_n19138__;
  assign new_new_n19219__ = new_new_n19126__ & new_new_n19218__;
  assign new_new_n19220__ = new_new_n19043__ & ~new_new_n19219__;
  assign new_new_n19221__ = new_new_n19037__ & ~new_new_n19047__;
  assign new_new_n19222__ = new_new_n19126__ & ~new_new_n19221__;
  assign new_new_n19223__ = ~new_new_n19142__ & ~new_new_n19222__;
  assign new_new_n19224__ = ~new_new_n19044__ & new_new_n19223__;
  assign new_new_n19225__ = ~new_new_n19126__ & ~new_new_n19218__;
  assign new_new_n19226__ = ~new_new_n19220__ & ~new_new_n19225__;
  assign new_new_n19227__ = ~new_new_n19224__ & new_new_n19226__;
  assign new_new_n19228__ = new_new_n19217__ & new_new_n19227__;
  assign new_new_n19229__ = ~new_new_n19217__ & ~new_new_n19227__;
  assign new_new_n19230__ = ~new_new_n19228__ & ~new_new_n19229__;
  assign new_new_n19231__ = new_new_n19172__ & ~new_new_n19230__;
  assign new_new_n19232__ = ~new_new_n19172__ & new_new_n19230__;
  assign new_new_n19233__ = ~new_new_n19231__ & ~new_new_n19232__;
  assign new_new_n19234__ = ~new_new_n19070__ & ~new_new_n19098__;
  assign new_new_n19235__ = ~new_new_n19071__ & ~new_new_n19234__;
  assign new_new_n19236__ = new_new_n19233__ & new_new_n19235__;
  assign new_new_n19237__ = ~new_new_n19233__ & ~new_new_n19235__;
  assign po110 = ~new_new_n19236__ & ~new_new_n19237__;
  assign new_new_n19239__ = ~new_new_n19169__ & new_new_n19229__;
  assign new_new_n19240__ = ~new_new_n19167__ & new_new_n19239__;
  assign new_new_n19241__ = ~new_new_n19194__ & ~new_new_n19197__;
  assign new_new_n19242__ = ~new_new_n19193__ & ~new_new_n19241__;
  assign new_new_n19243__ = ~new_new_n19157__ & ~new_new_n19162__;
  assign new_new_n19244__ = ~new_new_n19163__ & ~new_new_n19243__;
  assign new_new_n19245__ = ~new_new_n19242__ & new_new_n19244__;
  assign new_new_n19246__ = new_new_n19242__ & ~new_new_n19244__;
  assign new_new_n19247__ = ~new_new_n19245__ & ~new_new_n19246__;
  assign new_new_n19248__ = ~new_new_n19184__ & ~new_new_n19188__;
  assign new_new_n19249__ = ~new_new_n19187__ & ~new_new_n19248__;
  assign new_new_n19250__ = ~new_new_n19175__ & ~new_new_n19179__;
  assign new_new_n19251__ = ~new_new_n19178__ & ~new_new_n19250__;
  assign new_new_n19252__ = new_new_n19249__ & new_new_n19251__;
  assign new_new_n19253__ = ~new_new_n19249__ & ~new_new_n19251__;
  assign new_new_n19254__ = ~new_new_n19252__ & ~new_new_n19253__;
  assign new_new_n19255__ = pi51 & pi59;
  assign new_new_n19256__ = pi49 & pi61;
  assign new_new_n19257__ = pi50 & pi60;
  assign new_new_n19258__ = ~new_new_n19256__ & ~new_new_n19257__;
  assign new_new_n19259__ = new_new_n19256__ & new_new_n19257__;
  assign new_new_n19260__ = ~new_new_n19258__ & ~new_new_n19259__;
  assign new_new_n19261__ = new_new_n19255__ & ~new_new_n19260__;
  assign new_new_n19262__ = ~new_new_n19255__ & new_new_n19260__;
  assign new_new_n19263__ = ~new_new_n19261__ & ~new_new_n19262__;
  assign new_new_n19264__ = new_new_n19254__ & new_new_n19263__;
  assign new_new_n19265__ = ~new_new_n19254__ & ~new_new_n19263__;
  assign new_new_n19266__ = ~new_new_n19264__ & ~new_new_n19265__;
  assign new_new_n19267__ = new_new_n19247__ & ~new_new_n19266__;
  assign new_new_n19268__ = ~new_new_n19247__ & new_new_n19266__;
  assign new_new_n19269__ = ~new_new_n19267__ & ~new_new_n19268__;
  assign new_new_n19270__ = ~new_new_n19202__ & ~new_new_n19214__;
  assign new_new_n19271__ = ~new_new_n19201__ & ~new_new_n19270__;
  assign new_new_n19272__ = new_new_n19269__ & ~new_new_n19271__;
  assign new_new_n19273__ = ~new_new_n19269__ & new_new_n19271__;
  assign new_new_n19274__ = ~new_new_n19272__ & ~new_new_n19273__;
  assign new_new_n19275__ = pi54 & pi56;
  assign new_new_n19276__ = pi52 & pi58;
  assign new_new_n19277__ = pi53 & pi57;
  assign new_new_n19278__ = ~new_new_n19276__ & ~new_new_n19277__;
  assign new_new_n19279__ = new_new_n19276__ & new_new_n19277__;
  assign new_new_n19280__ = ~new_new_n19278__ & ~new_new_n19279__;
  assign new_new_n19281__ = new_new_n19275__ & ~new_new_n19280__;
  assign new_new_n19282__ = ~new_new_n19275__ & new_new_n19280__;
  assign new_new_n19283__ = ~new_new_n19281__ & ~new_new_n19282__;
  assign new_new_n19284__ = pi48 & pi63;
  assign new_new_n19285__ = ~pi48 & ~pi63;
  assign new_new_n19286__ = ~new_new_n19284__ & ~new_new_n19285__;
  assign new_new_n19287__ = pi48 & ~pi55;
  assign new_new_n19288__ = new_new_n19286__ & ~new_new_n19287__;
  assign new_new_n19289__ = ~new_new_n18407__ & ~new_new_n19286__;
  assign new_new_n19290__ = pi62 & ~new_new_n19288__;
  assign new_new_n19291__ = ~new_new_n19289__ & new_new_n19290__;
  assign new_new_n19292__ = pi54 & pi55;
  assign new_new_n19293__ = pi47 & pi63;
  assign new_new_n19294__ = ~new_new_n19292__ & ~new_new_n19293__;
  assign new_new_n19295__ = ~pi62 & ~new_new_n19293__;
  assign new_new_n19296__ = ~pi48 & ~new_new_n18407__;
  assign new_new_n19297__ = ~new_new_n19295__ & ~new_new_n19296__;
  assign new_new_n19298__ = ~new_new_n19294__ & ~new_new_n19297__;
  assign new_new_n19299__ = ~pi48 & ~new_new_n19293__;
  assign new_new_n19300__ = ~new_new_n19295__ & ~new_new_n19299__;
  assign new_new_n19301__ = ~new_new_n17234__ & ~new_new_n19292__;
  assign new_new_n19302__ = new_new_n19300__ & new_new_n19301__;
  assign new_new_n19303__ = ~new_new_n19298__ & ~new_new_n19302__;
  assign new_new_n19304__ = ~new_new_n19291__ & new_new_n19303__;
  assign new_new_n19305__ = ~new_new_n19206__ & ~new_new_n19208__;
  assign new_new_n19306__ = new_new_n19206__ & new_new_n19208__;
  assign new_new_n19307__ = ~new_new_n19205__ & ~new_new_n19306__;
  assign new_new_n19308__ = ~new_new_n19305__ & ~new_new_n19307__;
  assign new_new_n19309__ = ~new_new_n19304__ & new_new_n19308__;
  assign new_new_n19310__ = new_new_n19304__ & ~new_new_n19308__;
  assign new_new_n19311__ = new_new_n19283__ & ~new_new_n19309__;
  assign new_new_n19312__ = ~new_new_n19310__ & ~new_new_n19311__;
  assign new_new_n19313__ = ~new_new_n19309__ & new_new_n19312__;
  assign new_new_n19314__ = ~new_new_n19283__ & ~new_new_n19313__;
  assign new_new_n19315__ = ~new_new_n19310__ & new_new_n19311__;
  assign new_new_n19316__ = ~new_new_n19314__ & ~new_new_n19315__;
  assign new_new_n19317__ = new_new_n19274__ & ~new_new_n19316__;
  assign new_new_n19318__ = ~new_new_n19274__ & new_new_n19316__;
  assign new_new_n19319__ = ~new_new_n19317__ & ~new_new_n19318__;
  assign new_new_n19320__ = ~new_new_n19169__ & ~new_new_n19217__;
  assign new_new_n19321__ = new_new_n19169__ & new_new_n19217__;
  assign new_new_n19322__ = ~new_new_n19227__ & ~new_new_n19321__;
  assign new_new_n19323__ = ~new_new_n19320__ & ~new_new_n19322__;
  assign new_new_n19324__ = ~new_new_n19167__ & ~new_new_n19323__;
  assign new_new_n19325__ = ~new_new_n19235__ & ~new_new_n19239__;
  assign new_new_n19326__ = ~new_new_n19324__ & new_new_n19325__;
  assign new_new_n19327__ = new_new_n19169__ & new_new_n19228__;
  assign new_new_n19328__ = new_new_n19167__ & new_new_n19323__;
  assign new_new_n19329__ = new_new_n19235__ & ~new_new_n19327__;
  assign new_new_n19330__ = ~new_new_n19328__ & new_new_n19329__;
  assign new_new_n19331__ = ~new_new_n19326__ & ~new_new_n19330__;
  assign new_new_n19332__ = new_new_n19171__ & new_new_n19228__;
  assign new_new_n19333__ = new_new_n19319__ & ~new_new_n19332__;
  assign new_new_n19334__ = ~new_new_n19240__ & new_new_n19333__;
  assign new_new_n19335__ = ~new_new_n19331__ & new_new_n19334__;
  assign new_new_n19336__ = ~new_new_n19171__ & ~new_new_n19235__;
  assign new_new_n19337__ = ~new_new_n19170__ & ~new_new_n19336__;
  assign new_new_n19338__ = new_new_n19229__ & new_new_n19337__;
  assign new_new_n19339__ = new_new_n19171__ & new_new_n19235__;
  assign new_new_n19340__ = new_new_n19170__ & ~new_new_n19235__;
  assign new_new_n19341__ = ~new_new_n19339__ & ~new_new_n19340__;
  assign new_new_n19342__ = new_new_n19230__ & new_new_n19341__;
  assign new_new_n19343__ = new_new_n19228__ & ~new_new_n19337__;
  assign new_new_n19344__ = ~new_new_n19319__ & ~new_new_n19338__;
  assign new_new_n19345__ = ~new_new_n19343__ & new_new_n19344__;
  assign new_new_n19346__ = ~new_new_n19342__ & new_new_n19345__;
  assign po111 = ~new_new_n19335__ & ~new_new_n19346__;
  assign new_new_n19348__ = pi49 & pi62;
  assign new_new_n19349__ = ~pi55 & pi56;
  assign new_new_n19350__ = ~new_new_n19348__ & new_new_n19349__;
  assign new_new_n19351__ = new_new_n19348__ & ~new_new_n19349__;
  assign new_new_n19352__ = ~new_new_n19350__ & ~new_new_n19351__;
  assign new_new_n19353__ = pi54 & pi57;
  assign new_new_n19354__ = pi53 & pi58;
  assign new_new_n19355__ = pi52 & pi59;
  assign new_new_n19356__ = ~new_new_n19354__ & ~new_new_n19355__;
  assign new_new_n19357__ = new_new_n19354__ & new_new_n19355__;
  assign new_new_n19358__ = ~new_new_n19356__ & ~new_new_n19357__;
  assign new_new_n19359__ = new_new_n19353__ & ~new_new_n19358__;
  assign new_new_n19360__ = ~new_new_n19353__ & new_new_n19358__;
  assign new_new_n19361__ = ~new_new_n19359__ & ~new_new_n19360__;
  assign new_new_n19362__ = pi51 & pi60;
  assign new_new_n19363__ = pi50 & pi61;
  assign new_new_n19364__ = ~new_new_n19284__ & ~new_new_n19363__;
  assign new_new_n19365__ = new_new_n19284__ & new_new_n19363__;
  assign new_new_n19366__ = ~new_new_n19364__ & ~new_new_n19365__;
  assign new_new_n19367__ = new_new_n19362__ & ~new_new_n19366__;
  assign new_new_n19368__ = ~new_new_n19362__ & new_new_n19366__;
  assign new_new_n19369__ = ~new_new_n19367__ & ~new_new_n19368__;
  assign new_new_n19370__ = new_new_n19361__ & new_new_n19369__;
  assign new_new_n19371__ = ~new_new_n19361__ & ~new_new_n19369__;
  assign new_new_n19372__ = ~new_new_n19370__ & ~new_new_n19371__;
  assign new_new_n19373__ = new_new_n19352__ & ~new_new_n19372__;
  assign new_new_n19374__ = ~new_new_n19352__ & new_new_n19372__;
  assign new_new_n19375__ = ~new_new_n19373__ & ~new_new_n19374__;
  assign new_new_n19376__ = ~new_new_n19245__ & ~new_new_n19266__;
  assign new_new_n19377__ = ~new_new_n19246__ & ~new_new_n19376__;
  assign new_new_n19378__ = new_new_n19375__ & ~new_new_n19377__;
  assign new_new_n19379__ = ~new_new_n19375__ & new_new_n19377__;
  assign new_new_n19380__ = ~new_new_n19378__ & ~new_new_n19379__;
  assign new_new_n19381__ = ~new_new_n19273__ & ~new_new_n19316__;
  assign new_new_n19382__ = ~new_new_n19272__ & ~new_new_n19381__;
  assign new_new_n19383__ = ~new_new_n19235__ & ~new_new_n19321__;
  assign new_new_n19384__ = new_new_n19167__ & new_new_n19227__;
  assign new_new_n19385__ = new_new_n19319__ & ~new_new_n19384__;
  assign new_new_n19386__ = ~new_new_n19320__ & ~new_new_n19383__;
  assign new_new_n19387__ = ~new_new_n19385__ & new_new_n19386__;
  assign new_new_n19388__ = ~new_new_n19167__ & ~new_new_n19227__;
  assign new_new_n19389__ = ~new_new_n19235__ & new_new_n19320__;
  assign new_new_n19390__ = ~new_new_n19319__ & ~new_new_n19389__;
  assign new_new_n19391__ = new_new_n19235__ & new_new_n19321__;
  assign new_new_n19392__ = ~new_new_n19390__ & ~new_new_n19391__;
  assign new_new_n19393__ = ~new_new_n19388__ & ~new_new_n19392__;
  assign new_new_n19394__ = ~new_new_n19319__ & new_new_n19384__;
  assign new_new_n19395__ = ~new_new_n19393__ & ~new_new_n19394__;
  assign new_new_n19396__ = ~new_new_n19387__ & new_new_n19395__;
  assign new_new_n19397__ = ~new_new_n19382__ & new_new_n19396__;
  assign new_new_n19398__ = new_new_n19382__ & ~new_new_n19396__;
  assign new_new_n19399__ = ~new_new_n19397__ & ~new_new_n19398__;
  assign new_new_n19400__ = ~new_new_n19253__ & ~new_new_n19263__;
  assign new_new_n19401__ = ~new_new_n19252__ & ~new_new_n19400__;
  assign new_new_n19402__ = ~new_new_n19312__ & new_new_n19401__;
  assign new_new_n19403__ = new_new_n19312__ & ~new_new_n19401__;
  assign new_new_n19404__ = ~new_new_n19402__ & ~new_new_n19403__;
  assign new_new_n19405__ = new_new_n17234__ & new_new_n19284__;
  assign new_new_n19406__ = new_new_n17234__ & ~new_new_n19285__;
  assign new_new_n19407__ = pi54 & new_new_n19300__;
  assign new_new_n19408__ = ~new_new_n19406__ & ~new_new_n19407__;
  assign new_new_n19409__ = pi55 & ~new_new_n19408__;
  assign new_new_n19410__ = ~new_new_n19405__ & ~new_new_n19409__;
  assign new_new_n19411__ = ~new_new_n19255__ & ~new_new_n19259__;
  assign new_new_n19412__ = ~new_new_n19258__ & ~new_new_n19411__;
  assign new_new_n19413__ = new_new_n19410__ & ~new_new_n19412__;
  assign new_new_n19414__ = ~new_new_n19410__ & new_new_n19412__;
  assign new_new_n19415__ = ~new_new_n19413__ & ~new_new_n19414__;
  assign new_new_n19416__ = ~new_new_n19275__ & ~new_new_n19279__;
  assign new_new_n19417__ = ~new_new_n19278__ & ~new_new_n19416__;
  assign new_new_n19418__ = new_new_n19415__ & ~new_new_n19417__;
  assign new_new_n19419__ = ~new_new_n19415__ & new_new_n19417__;
  assign new_new_n19420__ = ~new_new_n19418__ & ~new_new_n19419__;
  assign new_new_n19421__ = new_new_n19404__ & ~new_new_n19420__;
  assign new_new_n19422__ = ~new_new_n19404__ & new_new_n19420__;
  assign new_new_n19423__ = ~new_new_n19421__ & ~new_new_n19422__;
  assign new_new_n19424__ = new_new_n19399__ & ~new_new_n19423__;
  assign new_new_n19425__ = ~new_new_n19399__ & new_new_n19423__;
  assign new_new_n19426__ = ~new_new_n19424__ & ~new_new_n19425__;
  assign new_new_n19427__ = new_new_n19380__ & new_new_n19426__;
  assign new_new_n19428__ = ~new_new_n19380__ & ~new_new_n19426__;
  assign po112 = new_new_n19427__ | new_new_n19428__;
  assign new_new_n19430__ = new_new_n19377__ & ~new_new_n19423__;
  assign new_new_n19431__ = ~new_new_n19377__ & new_new_n19423__;
  assign new_new_n19432__ = ~new_new_n19375__ & ~new_new_n19431__;
  assign new_new_n19433__ = ~new_new_n19430__ & ~new_new_n19432__;
  assign new_new_n19434__ = new_new_n19398__ & new_new_n19433__;
  assign new_new_n19435__ = ~new_new_n19430__ & ~new_new_n19431__;
  assign new_new_n19436__ = ~new_new_n19380__ & ~new_new_n19435__;
  assign new_new_n19437__ = new_new_n19399__ & ~new_new_n19436__;
  assign new_new_n19438__ = ~new_new_n19414__ & ~new_new_n19417__;
  assign new_new_n19439__ = ~new_new_n19413__ & ~new_new_n19438__;
  assign new_new_n19440__ = ~new_new_n19352__ & ~new_new_n19370__;
  assign new_new_n19441__ = ~new_new_n19371__ & ~new_new_n19440__;
  assign new_new_n19442__ = ~new_new_n19353__ & ~new_new_n19357__;
  assign new_new_n19443__ = ~new_new_n19356__ & ~new_new_n19442__;
  assign new_new_n19444__ = pi50 & new_new_n19443__;
  assign new_new_n19445__ = ~pi50 & ~new_new_n19443__;
  assign new_new_n19446__ = ~new_new_n19444__ & ~new_new_n19445__;
  assign new_new_n19447__ = pi49 & ~new_new_n19446__;
  assign new_new_n19448__ = pi55 & new_new_n19444__;
  assign new_new_n19449__ = ~new_new_n19447__ & ~new_new_n19448__;
  assign new_new_n19450__ = pi62 & ~new_new_n19449__;
  assign new_new_n19451__ = ~new_new_n18122__ & ~new_new_n19443__;
  assign new_new_n19452__ = pi55 & new_new_n19451__;
  assign new_new_n19453__ = ~new_new_n19450__ & ~new_new_n19452__;
  assign new_new_n19454__ = pi56 & ~new_new_n19453__;
  assign new_new_n19455__ = ~new_new_n18751__ & ~new_new_n19444__;
  assign new_new_n19456__ = pi62 & ~new_new_n19455__;
  assign new_new_n19457__ = pi55 & pi56;
  assign new_new_n19458__ = ~new_new_n19451__ & ~new_new_n19457__;
  assign new_new_n19459__ = ~new_new_n19456__ & new_new_n19458__;
  assign new_new_n19460__ = ~new_new_n19454__ & ~new_new_n19459__;
  assign new_new_n19461__ = new_new_n19441__ & new_new_n19460__;
  assign new_new_n19462__ = ~new_new_n19441__ & ~new_new_n19460__;
  assign new_new_n19463__ = ~new_new_n19461__ & ~new_new_n19462__;
  assign new_new_n19464__ = new_new_n19439__ & ~new_new_n19463__;
  assign new_new_n19465__ = ~new_new_n19439__ & new_new_n19463__;
  assign new_new_n19466__ = ~new_new_n19464__ & ~new_new_n19465__;
  assign new_new_n19467__ = ~new_new_n19402__ & ~new_new_n19420__;
  assign new_new_n19468__ = ~new_new_n19403__ & ~new_new_n19467__;
  assign new_new_n19469__ = new_new_n19466__ & new_new_n19468__;
  assign new_new_n19470__ = ~new_new_n19466__ & ~new_new_n19468__;
  assign new_new_n19471__ = ~new_new_n19469__ & ~new_new_n19470__;
  assign new_new_n19472__ = pi55 & pi57;
  assign new_new_n19473__ = pi53 & pi59;
  assign new_new_n19474__ = pi54 & pi58;
  assign new_new_n19475__ = ~new_new_n19473__ & ~new_new_n19474__;
  assign new_new_n19476__ = new_new_n19473__ & new_new_n19474__;
  assign new_new_n19477__ = ~new_new_n19475__ & ~new_new_n19476__;
  assign new_new_n19478__ = new_new_n19472__ & ~new_new_n19477__;
  assign new_new_n19479__ = ~new_new_n19472__ & new_new_n19477__;
  assign new_new_n19480__ = ~new_new_n19478__ & ~new_new_n19479__;
  assign new_new_n19481__ = pi52 & pi60;
  assign new_new_n19482__ = pi51 & pi61;
  assign new_new_n19483__ = pi49 & pi63;
  assign new_new_n19484__ = ~new_new_n19482__ & ~new_new_n19483__;
  assign new_new_n19485__ = new_new_n19482__ & new_new_n19483__;
  assign new_new_n19486__ = ~new_new_n19484__ & ~new_new_n19485__;
  assign new_new_n19487__ = new_new_n19481__ & ~new_new_n19486__;
  assign new_new_n19488__ = ~new_new_n19481__ & new_new_n19486__;
  assign new_new_n19489__ = ~new_new_n19487__ & ~new_new_n19488__;
  assign new_new_n19490__ = new_new_n19480__ & new_new_n19489__;
  assign new_new_n19491__ = ~new_new_n19480__ & ~new_new_n19489__;
  assign new_new_n19492__ = ~new_new_n19490__ & ~new_new_n19491__;
  assign new_new_n19493__ = ~new_new_n19362__ & ~new_new_n19365__;
  assign new_new_n19494__ = ~new_new_n19364__ & ~new_new_n19493__;
  assign new_new_n19495__ = new_new_n19492__ & ~new_new_n19494__;
  assign new_new_n19496__ = ~new_new_n19492__ & new_new_n19494__;
  assign new_new_n19497__ = ~new_new_n19495__ & ~new_new_n19496__;
  assign new_new_n19498__ = new_new_n19471__ & ~new_new_n19497__;
  assign new_new_n19499__ = ~new_new_n19471__ & new_new_n19497__;
  assign new_new_n19500__ = ~new_new_n19498__ & ~new_new_n19499__;
  assign new_new_n19501__ = new_new_n19397__ & ~new_new_n19433__;
  assign new_new_n19502__ = ~new_new_n19434__ & ~new_new_n19500__;
  assign new_new_n19503__ = ~new_new_n19501__ & new_new_n19502__;
  assign new_new_n19504__ = ~new_new_n19437__ & new_new_n19503__;
  assign new_new_n19505__ = new_new_n19397__ & new_new_n19431__;
  assign new_new_n19506__ = new_new_n19397__ & new_new_n19423__;
  assign new_new_n19507__ = ~new_new_n19397__ & ~new_new_n19423__;
  assign new_new_n19508__ = ~new_new_n19377__ & ~new_new_n19398__;
  assign new_new_n19509__ = ~new_new_n19507__ & new_new_n19508__;
  assign new_new_n19510__ = ~new_new_n19506__ & ~new_new_n19509__;
  assign new_new_n19511__ = new_new_n19375__ & ~new_new_n19510__;
  assign new_new_n19512__ = new_new_n19398__ & ~new_new_n19431__;
  assign new_new_n19513__ = ~new_new_n19397__ & new_new_n19430__;
  assign new_new_n19514__ = ~new_new_n19512__ & ~new_new_n19513__;
  assign new_new_n19515__ = ~new_new_n19375__ & ~new_new_n19514__;
  assign new_new_n19516__ = new_new_n19398__ & new_new_n19430__;
  assign new_new_n19517__ = new_new_n19500__ & ~new_new_n19505__;
  assign new_new_n19518__ = ~new_new_n19516__ & new_new_n19517__;
  assign new_new_n19519__ = ~new_new_n19515__ & new_new_n19518__;
  assign new_new_n19520__ = ~new_new_n19511__ & new_new_n19519__;
  assign po113 = ~new_new_n19504__ & ~new_new_n19520__;
  assign new_new_n19522__ = new_new_n19439__ & ~new_new_n19461__;
  assign new_new_n19523__ = ~new_new_n19462__ & ~new_new_n19522__;
  assign new_new_n19524__ = ~new_new_n19469__ & ~new_new_n19497__;
  assign new_new_n19525__ = ~new_new_n19470__ & ~new_new_n19524__;
  assign new_new_n19526__ = ~new_new_n19523__ & ~new_new_n19525__;
  assign new_new_n19527__ = new_new_n19523__ & new_new_n19525__;
  assign new_new_n19528__ = ~new_new_n19526__ & ~new_new_n19527__;
  assign new_new_n19529__ = ~new_new_n19490__ & new_new_n19494__;
  assign new_new_n19530__ = ~new_new_n19491__ & ~new_new_n19529__;
  assign new_new_n19531__ = pi49 & ~new_new_n19445__;
  assign new_new_n19532__ = ~new_new_n18750__ & ~new_new_n19531__;
  assign new_new_n19533__ = pi56 & ~new_new_n19532__;
  assign new_new_n19534__ = ~new_new_n19444__ & ~new_new_n19533__;
  assign new_new_n19535__ = pi62 & ~new_new_n19534__;
  assign new_new_n19536__ = new_new_n19443__ & new_new_n19457__;
  assign new_new_n19537__ = ~new_new_n19535__ & ~new_new_n19536__;
  assign new_new_n19538__ = ~new_new_n19472__ & ~new_new_n19476__;
  assign new_new_n19539__ = ~new_new_n19475__ & ~new_new_n19538__;
  assign new_new_n19540__ = pi53 & pi60;
  assign new_new_n19541__ = pi52 & pi61;
  assign new_new_n19542__ = ~new_new_n19540__ & ~new_new_n19541__;
  assign new_new_n19543__ = new_new_n19540__ & new_new_n19541__;
  assign new_new_n19544__ = ~new_new_n19542__ & ~new_new_n19543__;
  assign new_new_n19545__ = new_new_n19539__ & ~new_new_n19544__;
  assign new_new_n19546__ = ~new_new_n19539__ & new_new_n19544__;
  assign new_new_n19547__ = ~new_new_n19545__ & ~new_new_n19546__;
  assign new_new_n19548__ = new_new_n19537__ & new_new_n19547__;
  assign new_new_n19549__ = ~new_new_n19537__ & ~new_new_n19547__;
  assign new_new_n19550__ = ~new_new_n19548__ & ~new_new_n19549__;
  assign new_new_n19551__ = new_new_n19530__ & new_new_n19550__;
  assign new_new_n19552__ = ~new_new_n19530__ & ~new_new_n19550__;
  assign new_new_n19553__ = ~new_new_n19551__ & ~new_new_n19552__;
  assign new_new_n19554__ = new_new_n19433__ & new_new_n19500__;
  assign new_new_n19555__ = ~new_new_n19433__ & ~new_new_n19500__;
  assign new_new_n19556__ = new_new_n19397__ & ~new_new_n19555__;
  assign new_new_n19557__ = ~new_new_n19375__ & new_new_n19430__;
  assign new_new_n19558__ = new_new_n19500__ & ~new_new_n19557__;
  assign new_new_n19559__ = new_new_n19375__ & new_new_n19431__;
  assign new_new_n19560__ = ~new_new_n19558__ & ~new_new_n19559__;
  assign new_new_n19561__ = ~new_new_n19398__ & ~new_new_n19560__;
  assign new_new_n19562__ = ~new_new_n19554__ & ~new_new_n19556__;
  assign new_new_n19563__ = ~new_new_n19561__ & new_new_n19562__;
  assign new_new_n19564__ = ~new_new_n19553__ & ~new_new_n19563__;
  assign new_new_n19565__ = new_new_n19553__ & new_new_n19563__;
  assign new_new_n19566__ = ~new_new_n19564__ & ~new_new_n19565__;
  assign new_new_n19567__ = new_new_n19528__ & ~new_new_n19566__;
  assign new_new_n19568__ = ~new_new_n19528__ & new_new_n19566__;
  assign new_new_n19569__ = ~new_new_n19567__ & ~new_new_n19568__;
  assign new_new_n19570__ = ~new_new_n19481__ & ~new_new_n19485__;
  assign new_new_n19571__ = ~new_new_n19484__ & ~new_new_n19570__;
  assign new_new_n19572__ = pi55 & pi58;
  assign new_new_n19573__ = pi50 & pi63;
  assign new_new_n19574__ = pi54 & pi59;
  assign new_new_n19575__ = ~new_new_n19573__ & ~new_new_n19574__;
  assign new_new_n19576__ = new_new_n19573__ & new_new_n19574__;
  assign new_new_n19577__ = ~new_new_n19575__ & ~new_new_n19576__;
  assign new_new_n19578__ = new_new_n19572__ & ~new_new_n19577__;
  assign new_new_n19579__ = ~new_new_n19572__ & new_new_n19577__;
  assign new_new_n19580__ = ~new_new_n19578__ & ~new_new_n19579__;
  assign new_new_n19581__ = ~new_new_n19571__ & new_new_n19580__;
  assign new_new_n19582__ = new_new_n19571__ & ~new_new_n19580__;
  assign new_new_n19583__ = ~new_new_n19581__ & ~new_new_n19582__;
  assign new_new_n19584__ = pi51 & pi62;
  assign new_new_n19585__ = ~pi56 & pi57;
  assign new_new_n19586__ = new_new_n19584__ & ~new_new_n19585__;
  assign new_new_n19587__ = ~new_new_n19584__ & new_new_n19585__;
  assign new_new_n19588__ = ~new_new_n19586__ & ~new_new_n19587__;
  assign new_new_n19589__ = new_new_n19583__ & ~new_new_n19588__;
  assign new_new_n19590__ = ~new_new_n19583__ & new_new_n19588__;
  assign new_new_n19591__ = ~new_new_n19589__ & ~new_new_n19590__;
  assign new_new_n19592__ = new_new_n19569__ & new_new_n19591__;
  assign new_new_n19593__ = ~new_new_n19569__ & ~new_new_n19591__;
  assign po114 = new_new_n19592__ | new_new_n19593__;
  assign new_new_n19595__ = ~new_new_n19525__ & ~new_new_n19565__;
  assign new_new_n19596__ = ~new_new_n19564__ & ~new_new_n19595__;
  assign new_new_n19597__ = new_new_n19523__ & new_new_n19596__;
  assign new_new_n19598__ = new_new_n19525__ & new_new_n19565__;
  assign new_new_n19599__ = ~new_new_n19597__ & ~new_new_n19598__;
  assign new_new_n19600__ = ~new_new_n19591__ & ~new_new_n19599__;
  assign new_new_n19601__ = ~new_new_n19523__ & ~new_new_n19596__;
  assign new_new_n19602__ = ~new_new_n19525__ & new_new_n19564__;
  assign new_new_n19603__ = ~new_new_n19601__ & ~new_new_n19602__;
  assign new_new_n19604__ = new_new_n19591__ & ~new_new_n19603__;
  assign new_new_n19605__ = new_new_n19525__ & new_new_n19563__;
  assign new_new_n19606__ = ~new_new_n19523__ & ~new_new_n19553__;
  assign new_new_n19607__ = ~new_new_n19605__ & ~new_new_n19606__;
  assign new_new_n19608__ = new_new_n19523__ & new_new_n19553__;
  assign new_new_n19609__ = ~new_new_n19525__ & ~new_new_n19563__;
  assign new_new_n19610__ = ~new_new_n19608__ & ~new_new_n19609__;
  assign new_new_n19611__ = ~new_new_n19607__ & ~new_new_n19610__;
  assign new_new_n19612__ = ~new_new_n19530__ & ~new_new_n19548__;
  assign new_new_n19613__ = ~new_new_n19549__ & ~new_new_n19612__;
  assign new_new_n19614__ = ~pi56 & ~new_new_n19584__;
  assign new_new_n19615__ = pi57 & ~new_new_n19614__;
  assign new_new_n19616__ = ~new_new_n19572__ & ~new_new_n19576__;
  assign new_new_n19617__ = ~new_new_n19575__ & ~new_new_n19616__;
  assign new_new_n19618__ = ~new_new_n19539__ & ~new_new_n19543__;
  assign new_new_n19619__ = ~new_new_n19542__ & ~new_new_n19618__;
  assign new_new_n19620__ = ~new_new_n19617__ & ~new_new_n19619__;
  assign new_new_n19621__ = new_new_n19617__ & new_new_n19619__;
  assign new_new_n19622__ = ~new_new_n19620__ & ~new_new_n19621__;
  assign new_new_n19623__ = ~new_new_n19615__ & new_new_n19622__;
  assign new_new_n19624__ = new_new_n19615__ & ~new_new_n19622__;
  assign new_new_n19625__ = ~new_new_n19623__ & ~new_new_n19624__;
  assign new_new_n19626__ = ~new_new_n19613__ & ~new_new_n19625__;
  assign new_new_n19627__ = new_new_n19613__ & new_new_n19625__;
  assign new_new_n19628__ = ~new_new_n19626__ & ~new_new_n19627__;
  assign new_new_n19629__ = pi53 & pi61;
  assign new_new_n19630__ = pi51 & pi63;
  assign new_new_n19631__ = pi52 & pi62;
  assign new_new_n19632__ = ~new_new_n19630__ & ~new_new_n19631__;
  assign new_new_n19633__ = new_new_n19630__ & new_new_n19631__;
  assign new_new_n19634__ = ~new_new_n19632__ & ~new_new_n19633__;
  assign new_new_n19635__ = new_new_n19629__ & ~new_new_n19634__;
  assign new_new_n19636__ = ~new_new_n19629__ & new_new_n19634__;
  assign new_new_n19637__ = ~new_new_n19635__ & ~new_new_n19636__;
  assign new_new_n19638__ = ~new_new_n19581__ & ~new_new_n19588__;
  assign new_new_n19639__ = ~new_new_n19582__ & ~new_new_n19638__;
  assign new_new_n19640__ = new_new_n19637__ & new_new_n19639__;
  assign new_new_n19641__ = ~new_new_n19637__ & ~new_new_n19639__;
  assign new_new_n19642__ = pi56 & pi58;
  assign new_new_n19643__ = pi55 & pi59;
  assign new_new_n19644__ = pi54 & pi60;
  assign new_new_n19645__ = ~new_new_n19643__ & ~new_new_n19644__;
  assign new_new_n19646__ = new_new_n19643__ & new_new_n19644__;
  assign new_new_n19647__ = ~new_new_n19645__ & ~new_new_n19646__;
  assign new_new_n19648__ = new_new_n19642__ & ~new_new_n19647__;
  assign new_new_n19649__ = ~new_new_n19642__ & new_new_n19647__;
  assign new_new_n19650__ = ~new_new_n19648__ & ~new_new_n19649__;
  assign new_new_n19651__ = ~new_new_n19640__ & ~new_new_n19650__;
  assign new_new_n19652__ = ~new_new_n19641__ & ~new_new_n19651__;
  assign new_new_n19653__ = ~new_new_n19640__ & new_new_n19652__;
  assign new_new_n19654__ = ~new_new_n19641__ & new_new_n19651__;
  assign new_new_n19655__ = ~new_new_n19650__ & ~new_new_n19654__;
  assign new_new_n19656__ = ~new_new_n19653__ & ~new_new_n19655__;
  assign new_new_n19657__ = new_new_n19628__ & ~new_new_n19656__;
  assign new_new_n19658__ = ~new_new_n19628__ & new_new_n19656__;
  assign new_new_n19659__ = ~new_new_n19657__ & ~new_new_n19658__;
  assign new_new_n19660__ = ~new_new_n19611__ & new_new_n19659__;
  assign new_new_n19661__ = ~new_new_n19600__ & new_new_n19660__;
  assign new_new_n19662__ = ~new_new_n19604__ & new_new_n19661__;
  assign new_new_n19663__ = new_new_n19526__ & new_new_n19591__;
  assign new_new_n19664__ = new_new_n19527__ & ~new_new_n19591__;
  assign new_new_n19665__ = ~new_new_n19663__ & ~new_new_n19664__;
  assign new_new_n19666__ = new_new_n19566__ & new_new_n19665__;
  assign new_new_n19667__ = ~new_new_n19527__ & new_new_n19591__;
  assign new_new_n19668__ = ~new_new_n19526__ & ~new_new_n19667__;
  assign new_new_n19669__ = new_new_n19565__ & ~new_new_n19668__;
  assign new_new_n19670__ = new_new_n19564__ & new_new_n19668__;
  assign new_new_n19671__ = ~new_new_n19659__ & ~new_new_n19669__;
  assign new_new_n19672__ = ~new_new_n19670__ & new_new_n19671__;
  assign new_new_n19673__ = ~new_new_n19666__ & new_new_n19672__;
  assign po115 = ~new_new_n19662__ & ~new_new_n19673__;
  assign new_new_n19675__ = ~new_new_n19615__ & ~new_new_n19621__;
  assign new_new_n19676__ = ~new_new_n19620__ & ~new_new_n19675__;
  assign new_new_n19677__ = ~pi57 & pi58;
  assign new_new_n19678__ = ~new_new_n19676__ & ~new_new_n19677__;
  assign new_new_n19679__ = ~pi53 & ~new_new_n19678__;
  assign new_new_n19680__ = pi62 & ~new_new_n19676__;
  assign new_new_n19681__ = ~pi62 & new_new_n19676__;
  assign new_new_n19682__ = new_new_n19677__ & ~new_new_n19681__;
  assign new_new_n19683__ = ~new_new_n19680__ & new_new_n19682__;
  assign new_new_n19684__ = ~new_new_n19679__ & ~new_new_n19683__;
  assign new_new_n19685__ = pi56 & pi59;
  assign new_new_n19686__ = pi55 & pi60;
  assign new_new_n19687__ = pi54 & pi61;
  assign new_new_n19688__ = ~new_new_n19686__ & ~new_new_n19687__;
  assign new_new_n19689__ = new_new_n19686__ & new_new_n19687__;
  assign new_new_n19690__ = ~new_new_n19688__ & ~new_new_n19689__;
  assign new_new_n19691__ = new_new_n19685__ & ~new_new_n19690__;
  assign new_new_n19692__ = ~new_new_n19685__ & new_new_n19690__;
  assign new_new_n19693__ = ~new_new_n19691__ & ~new_new_n19692__;
  assign new_new_n19694__ = ~new_new_n19684__ & ~new_new_n19693__;
  assign new_new_n19695__ = ~new_new_n19676__ & new_new_n19693__;
  assign new_new_n19696__ = new_new_n19676__ & ~new_new_n19693__;
  assign new_new_n19697__ = ~new_new_n19695__ & ~new_new_n19696__;
  assign new_new_n19698__ = new_new_n18937__ & ~new_new_n19697__;
  assign new_new_n19699__ = pi62 & ~new_new_n19695__;
  assign new_new_n19700__ = ~new_new_n19697__ & ~new_new_n19699__;
  assign new_new_n19701__ = ~new_new_n18937__ & ~new_new_n19700__;
  assign new_new_n19702__ = ~new_new_n19677__ & ~new_new_n19698__;
  assign new_new_n19703__ = ~new_new_n19701__ & new_new_n19702__;
  assign new_new_n19704__ = pi53 & new_new_n19680__;
  assign new_new_n19705__ = ~new_new_n19681__ & ~new_new_n19704__;
  assign new_new_n19706__ = new_new_n19677__ & new_new_n19693__;
  assign new_new_n19707__ = ~new_new_n19705__ & new_new_n19706__;
  assign new_new_n19708__ = ~new_new_n19694__ & ~new_new_n19707__;
  assign new_new_n19709__ = ~new_new_n19703__ & new_new_n19708__;
  assign new_new_n19710__ = new_new_n19652__ & ~new_new_n19709__;
  assign new_new_n19711__ = ~new_new_n19652__ & new_new_n19709__;
  assign new_new_n19712__ = ~new_new_n19710__ & ~new_new_n19711__;
  assign new_new_n19713__ = ~new_new_n19642__ & ~new_new_n19646__;
  assign new_new_n19714__ = ~new_new_n19645__ & ~new_new_n19713__;
  assign new_new_n19715__ = pi52 & pi63;
  assign new_new_n19716__ = ~new_new_n19629__ & ~new_new_n19633__;
  assign new_new_n19717__ = ~new_new_n19632__ & ~new_new_n19716__;
  assign new_new_n19718__ = new_new_n19715__ & ~new_new_n19717__;
  assign new_new_n19719__ = ~new_new_n19715__ & new_new_n19717__;
  assign new_new_n19720__ = ~new_new_n19718__ & ~new_new_n19719__;
  assign new_new_n19721__ = new_new_n19714__ & new_new_n19720__;
  assign new_new_n19722__ = ~new_new_n19714__ & ~new_new_n19720__;
  assign new_new_n19723__ = ~new_new_n19721__ & ~new_new_n19722__;
  assign new_new_n19724__ = ~new_new_n19712__ & ~new_new_n19723__;
  assign new_new_n19725__ = ~new_new_n19608__ & new_new_n19659__;
  assign new_new_n19726__ = ~new_new_n19591__ & ~new_new_n19609__;
  assign new_new_n19727__ = new_new_n19608__ & ~new_new_n19659__;
  assign new_new_n19728__ = ~new_new_n19605__ & ~new_new_n19727__;
  assign new_new_n19729__ = ~new_new_n19726__ & new_new_n19728__;
  assign new_new_n19730__ = ~new_new_n19725__ & ~new_new_n19729__;
  assign new_new_n19731__ = ~new_new_n19609__ & ~new_new_n19659__;
  assign new_new_n19732__ = new_new_n19591__ & ~new_new_n19731__;
  assign new_new_n19733__ = ~new_new_n19605__ & new_new_n19659__;
  assign new_new_n19734__ = ~new_new_n19606__ & ~new_new_n19733__;
  assign new_new_n19735__ = ~new_new_n19732__ & new_new_n19734__;
  assign new_new_n19736__ = ~new_new_n19730__ & ~new_new_n19735__;
  assign new_new_n19737__ = ~new_new_n19627__ & ~new_new_n19656__;
  assign new_new_n19738__ = ~new_new_n19626__ & ~new_new_n19737__;
  assign new_new_n19739__ = ~new_new_n19736__ & new_new_n19738__;
  assign new_new_n19740__ = new_new_n19724__ & new_new_n19739__;
  assign new_new_n19741__ = new_new_n19710__ & ~new_new_n19736__;
  assign new_new_n19742__ = ~new_new_n19710__ & new_new_n19736__;
  assign new_new_n19743__ = ~new_new_n19711__ & new_new_n19738__;
  assign new_new_n19744__ = ~new_new_n19742__ & new_new_n19743__;
  assign new_new_n19745__ = ~new_new_n19741__ & ~new_new_n19744__;
  assign new_new_n19746__ = new_new_n19723__ & ~new_new_n19745__;
  assign new_new_n19747__ = new_new_n19738__ & new_new_n19741__;
  assign new_new_n19748__ = ~new_new_n19746__ & ~new_new_n19747__;
  assign new_new_n19749__ = new_new_n19712__ & ~new_new_n19723__;
  assign new_new_n19750__ = ~new_new_n19712__ & new_new_n19723__;
  assign new_new_n19751__ = ~new_new_n19738__ & ~new_new_n19749__;
  assign new_new_n19752__ = ~new_new_n19750__ & new_new_n19751__;
  assign new_new_n19753__ = new_new_n19748__ & ~new_new_n19752__;
  assign new_new_n19754__ = new_new_n19736__ & ~new_new_n19753__;
  assign new_new_n19755__ = new_new_n19710__ & new_new_n19738__;
  assign new_new_n19756__ = new_new_n19746__ & ~new_new_n19755__;
  assign new_new_n19757__ = new_new_n19736__ & ~new_new_n19738__;
  assign new_new_n19758__ = ~new_new_n19711__ & new_new_n19723__;
  assign new_new_n19759__ = ~new_new_n19724__ & ~new_new_n19758__;
  assign new_new_n19760__ = ~new_new_n19739__ & new_new_n19759__;
  assign new_new_n19761__ = ~new_new_n19757__ & new_new_n19760__;
  assign new_new_n19762__ = ~new_new_n19740__ & ~new_new_n19761__;
  assign new_new_n19763__ = ~new_new_n19756__ & new_new_n19762__;
  assign po116 = new_new_n19754__ | ~new_new_n19763__;
  assign new_new_n19765__ = pi54 & pi63;
  assign new_new_n19766__ = ~pi54 & ~pi63;
  assign new_new_n19767__ = ~new_new_n19765__ & ~new_new_n19766__;
  assign new_new_n19768__ = pi54 & ~pi58;
  assign new_new_n19769__ = new_new_n19767__ & ~new_new_n19768__;
  assign new_new_n19770__ = ~new_new_n19354__ & ~new_new_n19767__;
  assign new_new_n19771__ = pi62 & ~new_new_n19769__;
  assign new_new_n19772__ = ~new_new_n19770__ & new_new_n19771__;
  assign new_new_n19773__ = pi57 & pi58;
  assign new_new_n19774__ = pi53 & pi63;
  assign new_new_n19775__ = ~new_new_n19773__ & ~new_new_n19774__;
  assign new_new_n19776__ = ~pi62 & ~new_new_n19774__;
  assign new_new_n19777__ = ~pi54 & ~new_new_n19354__;
  assign new_new_n19778__ = ~new_new_n19776__ & ~new_new_n19777__;
  assign new_new_n19779__ = ~new_new_n19775__ & ~new_new_n19778__;
  assign new_new_n19780__ = ~pi54 & ~new_new_n19774__;
  assign new_new_n19781__ = ~new_new_n19776__ & ~new_new_n19780__;
  assign new_new_n19782__ = ~new_new_n18937__ & ~new_new_n19773__;
  assign new_new_n19783__ = new_new_n19781__ & new_new_n19782__;
  assign new_new_n19784__ = ~new_new_n19779__ & ~new_new_n19783__;
  assign new_new_n19785__ = ~new_new_n19772__ & new_new_n19784__;
  assign new_new_n19786__ = ~new_new_n19685__ & ~new_new_n19689__;
  assign new_new_n19787__ = ~new_new_n19688__ & ~new_new_n19786__;
  assign new_new_n19788__ = new_new_n19785__ & ~new_new_n19787__;
  assign new_new_n19789__ = ~new_new_n19785__ & new_new_n19787__;
  assign new_new_n19790__ = ~new_new_n19788__ & ~new_new_n19789__;
  assign new_new_n19791__ = pi57 & pi59;
  assign new_new_n19792__ = pi55 & pi61;
  assign new_new_n19793__ = pi56 & pi60;
  assign new_new_n19794__ = ~new_new_n19792__ & ~new_new_n19793__;
  assign new_new_n19795__ = new_new_n19792__ & new_new_n19793__;
  assign new_new_n19796__ = ~new_new_n19794__ & ~new_new_n19795__;
  assign new_new_n19797__ = new_new_n19791__ & ~new_new_n19796__;
  assign new_new_n19798__ = ~new_new_n19791__ & new_new_n19796__;
  assign new_new_n19799__ = ~new_new_n19797__ & ~new_new_n19798__;
  assign new_new_n19800__ = new_new_n19790__ & new_new_n19799__;
  assign new_new_n19801__ = ~new_new_n19790__ & ~new_new_n19799__;
  assign new_new_n19802__ = ~new_new_n19800__ & ~new_new_n19801__;
  assign new_new_n19803__ = ~new_new_n19677__ & ~new_new_n19699__;
  assign new_new_n19804__ = pi53 & ~new_new_n19682__;
  assign new_new_n19805__ = ~new_new_n19803__ & new_new_n19804__;
  assign new_new_n19806__ = new_new_n18937__ & ~new_new_n19676__;
  assign new_new_n19807__ = ~new_new_n19678__ & ~new_new_n19693__;
  assign new_new_n19808__ = ~new_new_n19806__ & new_new_n19807__;
  assign new_new_n19809__ = ~new_new_n19805__ & ~new_new_n19808__;
  assign new_new_n19810__ = new_new_n19802__ & new_new_n19809__;
  assign new_new_n19811__ = ~new_new_n19802__ & ~new_new_n19809__;
  assign new_new_n19812__ = ~new_new_n19810__ & ~new_new_n19811__;
  assign new_new_n19813__ = new_new_n19711__ & new_new_n19757__;
  assign new_new_n19814__ = new_new_n19711__ & ~new_new_n19739__;
  assign new_new_n19815__ = ~new_new_n19710__ & new_new_n19757__;
  assign new_new_n19816__ = ~new_new_n19814__ & ~new_new_n19815__;
  assign new_new_n19817__ = ~new_new_n19723__ & ~new_new_n19816__;
  assign new_new_n19818__ = ~new_new_n19813__ & ~new_new_n19817__;
  assign new_new_n19819__ = new_new_n19748__ & new_new_n19818__;
  assign new_new_n19820__ = new_new_n19812__ & ~new_new_n19819__;
  assign new_new_n19821__ = ~new_new_n19812__ & new_new_n19819__;
  assign new_new_n19822__ = ~new_new_n19820__ & ~new_new_n19821__;
  assign new_new_n19823__ = ~new_new_n19715__ & ~new_new_n19717__;
  assign new_new_n19824__ = new_new_n19715__ & new_new_n19717__;
  assign new_new_n19825__ = ~new_new_n19714__ & ~new_new_n19824__;
  assign new_new_n19826__ = ~new_new_n19823__ & ~new_new_n19825__;
  assign new_new_n19827__ = new_new_n19822__ & ~new_new_n19826__;
  assign new_new_n19828__ = ~new_new_n19822__ & new_new_n19826__;
  assign po117 = ~new_new_n19827__ & ~new_new_n19828__;
  assign new_new_n19830__ = pi55 & pi62;
  assign new_new_n19831__ = ~pi58 & pi59;
  assign new_new_n19832__ = new_new_n19830__ & ~new_new_n19831__;
  assign new_new_n19833__ = ~new_new_n19830__ & new_new_n19831__;
  assign new_new_n19834__ = ~new_new_n19832__ & ~new_new_n19833__;
  assign new_new_n19835__ = ~new_new_n19788__ & ~new_new_n19799__;
  assign new_new_n19836__ = ~new_new_n19789__ & ~new_new_n19835__;
  assign new_new_n19837__ = new_new_n19834__ & new_new_n19836__;
  assign new_new_n19838__ = ~new_new_n19834__ & ~new_new_n19836__;
  assign new_new_n19839__ = ~new_new_n19837__ & ~new_new_n19838__;
  assign new_new_n19840__ = new_new_n18937__ & new_new_n19765__;
  assign new_new_n19841__ = new_new_n18937__ & ~new_new_n19766__;
  assign new_new_n19842__ = pi57 & new_new_n19781__;
  assign new_new_n19843__ = ~new_new_n19841__ & ~new_new_n19842__;
  assign new_new_n19844__ = pi58 & ~new_new_n19843__;
  assign new_new_n19845__ = ~new_new_n19840__ & ~new_new_n19844__;
  assign new_new_n19846__ = ~new_new_n19791__ & ~new_new_n19795__;
  assign new_new_n19847__ = ~new_new_n19794__ & ~new_new_n19846__;
  assign new_new_n19848__ = ~new_new_n19845__ & new_new_n19847__;
  assign new_new_n19849__ = new_new_n19845__ & ~new_new_n19847__;
  assign new_new_n19850__ = pi57 & pi60;
  assign new_new_n19851__ = pi56 & pi61;
  assign new_new_n19852__ = ~new_new_n19765__ & ~new_new_n19851__;
  assign new_new_n19853__ = new_new_n19765__ & new_new_n19851__;
  assign new_new_n19854__ = ~new_new_n19852__ & ~new_new_n19853__;
  assign new_new_n19855__ = new_new_n19850__ & ~new_new_n19854__;
  assign new_new_n19856__ = ~new_new_n19850__ & new_new_n19854__;
  assign new_new_n19857__ = ~new_new_n19855__ & ~new_new_n19856__;
  assign new_new_n19858__ = ~new_new_n19848__ & new_new_n19857__;
  assign new_new_n19859__ = ~new_new_n19849__ & ~new_new_n19858__;
  assign new_new_n19860__ = ~new_new_n19848__ & new_new_n19859__;
  assign new_new_n19861__ = ~new_new_n19849__ & new_new_n19858__;
  assign new_new_n19862__ = new_new_n19857__ & ~new_new_n19861__;
  assign new_new_n19863__ = ~new_new_n19860__ & ~new_new_n19862__;
  assign new_new_n19864__ = new_new_n19839__ & ~new_new_n19863__;
  assign new_new_n19865__ = ~new_new_n19839__ & new_new_n19863__;
  assign new_new_n19866__ = ~new_new_n19864__ & ~new_new_n19865__;
  assign new_new_n19867__ = new_new_n19810__ & ~new_new_n19866__;
  assign new_new_n19868__ = new_new_n19748__ & new_new_n19866__;
  assign new_new_n19869__ = ~new_new_n19809__ & new_new_n19868__;
  assign new_new_n19870__ = ~new_new_n19867__ & ~new_new_n19869__;
  assign new_new_n19871__ = new_new_n19818__ & ~new_new_n19870__;
  assign new_new_n19872__ = ~new_new_n19748__ & ~new_new_n19809__;
  assign new_new_n19873__ = ~new_new_n19818__ & ~new_new_n19872__;
  assign new_new_n19874__ = new_new_n19866__ & ~new_new_n19873__;
  assign new_new_n19875__ = new_new_n19748__ & ~new_new_n19866__;
  assign new_new_n19876__ = ~new_new_n19811__ & ~new_new_n19875__;
  assign new_new_n19877__ = ~new_new_n19874__ & new_new_n19876__;
  assign new_new_n19878__ = ~new_new_n19871__ & ~new_new_n19877__;
  assign new_new_n19879__ = ~new_new_n19826__ & ~new_new_n19878__;
  assign new_new_n19880__ = new_new_n19818__ & new_new_n19869__;
  assign new_new_n19881__ = new_new_n19818__ & new_new_n19866__;
  assign new_new_n19882__ = new_new_n19809__ & ~new_new_n19875__;
  assign new_new_n19883__ = ~new_new_n19881__ & new_new_n19882__;
  assign new_new_n19884__ = ~new_new_n19880__ & ~new_new_n19883__;
  assign new_new_n19885__ = new_new_n19802__ & ~new_new_n19884__;
  assign new_new_n19886__ = new_new_n19802__ & ~new_new_n19826__;
  assign new_new_n19887__ = new_new_n19818__ & ~new_new_n19866__;
  assign new_new_n19888__ = new_new_n19809__ & ~new_new_n19819__;
  assign new_new_n19889__ = ~new_new_n19886__ & ~new_new_n19887__;
  assign new_new_n19890__ = ~new_new_n19869__ & new_new_n19889__;
  assign new_new_n19891__ = ~new_new_n19888__ & new_new_n19890__;
  assign new_new_n19892__ = new_new_n19748__ & ~new_new_n19809__;
  assign new_new_n19893__ = new_new_n19887__ & ~new_new_n19892__;
  assign new_new_n19894__ = ~new_new_n19802__ & new_new_n19826__;
  assign new_new_n19895__ = ~new_new_n19868__ & new_new_n19894__;
  assign new_new_n19896__ = ~new_new_n19893__ & new_new_n19895__;
  assign new_new_n19897__ = ~new_new_n19891__ & ~new_new_n19896__;
  assign new_new_n19898__ = ~new_new_n19885__ & new_new_n19897__;
  assign po118 = new_new_n19879__ | ~new_new_n19898__;
  assign new_new_n19900__ = ~new_new_n19837__ & new_new_n19863__;
  assign new_new_n19901__ = ~new_new_n19838__ & ~new_new_n19900__;
  assign new_new_n19902__ = ~new_new_n19811__ & new_new_n19866__;
  assign new_new_n19903__ = new_new_n19811__ & ~new_new_n19866__;
  assign new_new_n19904__ = new_new_n19748__ & new_new_n19826__;
  assign new_new_n19905__ = new_new_n19818__ & ~new_new_n19903__;
  assign new_new_n19906__ = ~new_new_n19904__ & new_new_n19905__;
  assign new_new_n19907__ = ~new_new_n19902__ & ~new_new_n19906__;
  assign new_new_n19908__ = ~new_new_n19826__ & ~new_new_n19875__;
  assign new_new_n19909__ = ~new_new_n19810__ & ~new_new_n19881__;
  assign new_new_n19910__ = ~new_new_n19908__ & new_new_n19909__;
  assign new_new_n19911__ = ~new_new_n19907__ & ~new_new_n19910__;
  assign new_new_n19912__ = ~new_new_n19901__ & ~new_new_n19911__;
  assign new_new_n19913__ = new_new_n19901__ & new_new_n19911__;
  assign new_new_n19914__ = ~new_new_n19912__ & ~new_new_n19913__;
  assign new_new_n19915__ = ~new_new_n19850__ & ~new_new_n19853__;
  assign new_new_n19916__ = ~new_new_n19852__ & ~new_new_n19915__;
  assign new_new_n19917__ = pi63 & new_new_n19916__;
  assign new_new_n19918__ = pi55 & new_new_n19917__;
  assign new_new_n19919__ = ~pi63 & ~new_new_n19916__;
  assign new_new_n19920__ = ~pi55 & ~new_new_n19916__;
  assign new_new_n19921__ = ~new_new_n19919__ & ~new_new_n19920__;
  assign new_new_n19922__ = ~new_new_n19918__ & new_new_n19921__;
  assign new_new_n19923__ = pi58 & ~new_new_n19922__;
  assign new_new_n19924__ = ~pi58 & new_new_n19917__;
  assign new_new_n19925__ = pi55 & new_new_n19919__;
  assign new_new_n19926__ = ~new_new_n19924__ & ~new_new_n19925__;
  assign new_new_n19927__ = pi62 & ~new_new_n19926__;
  assign new_new_n19928__ = ~new_new_n19923__ & ~new_new_n19927__;
  assign new_new_n19929__ = pi59 & ~new_new_n19928__;
  assign new_new_n19930__ = pi58 & pi59;
  assign new_new_n19931__ = pi59 & pi62;
  assign new_new_n19932__ = ~new_new_n19917__ & ~new_new_n19931__;
  assign new_new_n19933__ = pi55 & ~new_new_n19932__;
  assign new_new_n19934__ = new_new_n19921__ & ~new_new_n19930__;
  assign new_new_n19935__ = ~new_new_n19933__ & new_new_n19934__;
  assign new_new_n19936__ = ~new_new_n19929__ & ~new_new_n19935__;
  assign new_new_n19937__ = ~new_new_n19859__ & new_new_n19936__;
  assign new_new_n19938__ = new_new_n19859__ & ~new_new_n19936__;
  assign new_new_n19939__ = ~new_new_n19937__ & ~new_new_n19938__;
  assign new_new_n19940__ = pi58 & pi60;
  assign new_new_n19941__ = pi56 & pi62;
  assign new_new_n19942__ = pi57 & pi61;
  assign new_new_n19943__ = ~new_new_n19941__ & ~new_new_n19942__;
  assign new_new_n19944__ = new_new_n19941__ & new_new_n19942__;
  assign new_new_n19945__ = ~new_new_n19943__ & ~new_new_n19944__;
  assign new_new_n19946__ = new_new_n19940__ & ~new_new_n19945__;
  assign new_new_n19947__ = ~new_new_n19940__ & new_new_n19945__;
  assign new_new_n19948__ = ~new_new_n19946__ & ~new_new_n19947__;
  assign new_new_n19949__ = new_new_n19939__ & ~new_new_n19948__;
  assign new_new_n19950__ = ~new_new_n19939__ & new_new_n19948__;
  assign new_new_n19951__ = ~new_new_n19949__ & ~new_new_n19950__;
  assign new_new_n19952__ = new_new_n19914__ & new_new_n19951__;
  assign new_new_n19953__ = ~new_new_n19914__ & ~new_new_n19951__;
  assign po119 = ~new_new_n19952__ & ~new_new_n19953__;
  assign new_new_n19955__ = new_new_n19937__ & new_new_n19948__;
  assign new_new_n19956__ = new_new_n19938__ & ~new_new_n19948__;
  assign new_new_n19957__ = ~new_new_n19955__ & ~new_new_n19956__;
  assign new_new_n19958__ = new_new_n19914__ & new_new_n19957__;
  assign new_new_n19959__ = ~new_new_n19937__ & ~new_new_n19948__;
  assign new_new_n19960__ = ~new_new_n19938__ & ~new_new_n19959__;
  assign new_new_n19961__ = new_new_n19913__ & ~new_new_n19960__;
  assign new_new_n19962__ = new_new_n19912__ & new_new_n19960__;
  assign new_new_n19963__ = ~new_new_n19961__ & ~new_new_n19962__;
  assign new_new_n19964__ = ~new_new_n19958__ & new_new_n19963__;
  assign new_new_n19965__ = pi58 & pi61;
  assign new_new_n19966__ = pi56 & pi63;
  assign new_new_n19967__ = ~new_new_n19940__ & ~new_new_n19944__;
  assign new_new_n19968__ = ~new_new_n19943__ & ~new_new_n19967__;
  assign new_new_n19969__ = ~new_new_n19966__ & ~new_new_n19968__;
  assign new_new_n19970__ = pi63 & new_new_n19968__;
  assign new_new_n19971__ = ~new_new_n19969__ & ~new_new_n19970__;
  assign new_new_n19972__ = ~new_new_n19965__ & ~new_new_n19971__;
  assign new_new_n19973__ = new_new_n19965__ & ~new_new_n19969__;
  assign new_new_n19974__ = pi56 & new_new_n19970__;
  assign new_new_n19975__ = new_new_n19973__ & ~new_new_n19974__;
  assign new_new_n19976__ = ~new_new_n19972__ & ~new_new_n19975__;
  assign new_new_n19977__ = ~pi58 & ~new_new_n19830__;
  assign new_new_n19978__ = pi59 & ~new_new_n19977__;
  assign new_new_n19979__ = new_new_n19921__ & new_new_n19978__;
  assign new_new_n19980__ = ~new_new_n19918__ & ~new_new_n19979__;
  assign new_new_n19981__ = ~new_new_n19976__ & ~new_new_n19980__;
  assign new_new_n19982__ = new_new_n19976__ & new_new_n19980__;
  assign new_new_n19983__ = ~new_new_n19981__ & ~new_new_n19982__;
  assign new_new_n19984__ = ~pi59 & pi60;
  assign new_new_n19985__ = ~pi62 & new_new_n19984__;
  assign new_new_n19986__ = pi57 & pi62;
  assign new_new_n19987__ = ~new_new_n19984__ & new_new_n19986__;
  assign new_new_n19988__ = ~new_new_n19985__ & ~new_new_n19987__;
  assign new_new_n19989__ = ~new_new_n19983__ & ~new_new_n19988__;
  assign new_new_n19990__ = ~pi57 & new_new_n19984__;
  assign new_new_n19991__ = new_new_n19982__ & new_new_n19990__;
  assign new_new_n19992__ = new_new_n19984__ & ~new_new_n19986__;
  assign new_new_n19993__ = ~new_new_n19987__ & ~new_new_n19992__;
  assign new_new_n19994__ = new_new_n19983__ & new_new_n19993__;
  assign new_new_n19995__ = ~new_new_n19989__ & ~new_new_n19991__;
  assign new_new_n19996__ = ~new_new_n19994__ & new_new_n19995__;
  assign new_new_n19997__ = ~new_new_n19964__ & ~new_new_n19996__;
  assign new_new_n19998__ = ~new_new_n19911__ & ~new_new_n19936__;
  assign new_new_n19999__ = new_new_n19911__ & new_new_n19936__;
  assign new_new_n20000__ = ~new_new_n19901__ & ~new_new_n19999__;
  assign new_new_n20001__ = ~new_new_n19998__ & ~new_new_n20000__;
  assign new_new_n20002__ = ~new_new_n19859__ & new_new_n20001__;
  assign new_new_n20003__ = new_new_n19913__ & new_new_n19936__;
  assign new_new_n20004__ = ~new_new_n20002__ & ~new_new_n20003__;
  assign new_new_n20005__ = new_new_n19948__ & ~new_new_n20004__;
  assign new_new_n20006__ = new_new_n19859__ & ~new_new_n20001__;
  assign new_new_n20007__ = new_new_n19912__ & ~new_new_n19936__;
  assign new_new_n20008__ = ~new_new_n20006__ & ~new_new_n20007__;
  assign new_new_n20009__ = ~new_new_n19948__ & ~new_new_n20008__;
  assign new_new_n20010__ = ~new_new_n19859__ & new_new_n19901__;
  assign new_new_n20011__ = ~new_new_n19912__ & ~new_new_n20010__;
  assign new_new_n20012__ = ~new_new_n19938__ & ~new_new_n19999__;
  assign new_new_n20013__ = ~new_new_n20011__ & ~new_new_n20012__;
  assign new_new_n20014__ = ~new_new_n20005__ & ~new_new_n20013__;
  assign new_new_n20015__ = ~new_new_n20009__ & new_new_n20014__;
  assign new_new_n20016__ = new_new_n19996__ & ~new_new_n20015__;
  assign po120 = new_new_n19997__ | new_new_n20016__;
  assign new_new_n20018__ = new_new_n19859__ & ~new_new_n19901__;
  assign new_new_n20019__ = ~new_new_n19948__ & ~new_new_n20010__;
  assign new_new_n20020__ = ~new_new_n20018__ & ~new_new_n20019__;
  assign new_new_n20021__ = ~new_new_n19996__ & new_new_n20020__;
  assign new_new_n20022__ = new_new_n19996__ & ~new_new_n20020__;
  assign new_new_n20023__ = ~new_new_n19998__ & ~new_new_n20022__;
  assign new_new_n20024__ = ~new_new_n20021__ & ~new_new_n20023__;
  assign new_new_n20025__ = ~new_new_n19996__ & ~new_new_n20018__;
  assign new_new_n20026__ = new_new_n19996__ & ~new_new_n20010__;
  assign new_new_n20027__ = new_new_n19948__ & ~new_new_n20026__;
  assign new_new_n20028__ = ~new_new_n20025__ & ~new_new_n20027__;
  assign new_new_n20029__ = ~new_new_n19999__ & new_new_n20028__;
  assign new_new_n20030__ = ~new_new_n20024__ & ~new_new_n20029__;
  assign new_new_n20031__ = ~new_new_n19970__ & ~new_new_n19973__;
  assign new_new_n20032__ = pi59 & pi61;
  assign new_new_n20033__ = pi57 & pi63;
  assign new_new_n20034__ = pi58 & pi62;
  assign new_new_n20035__ = ~new_new_n20033__ & ~new_new_n20034__;
  assign new_new_n20036__ = new_new_n20033__ & new_new_n20034__;
  assign new_new_n20037__ = ~new_new_n20035__ & ~new_new_n20036__;
  assign new_new_n20038__ = new_new_n20032__ & ~new_new_n20037__;
  assign new_new_n20039__ = ~new_new_n20032__ & new_new_n20037__;
  assign new_new_n20040__ = ~new_new_n20038__ & ~new_new_n20039__;
  assign new_new_n20041__ = ~new_new_n20031__ & ~new_new_n20040__;
  assign new_new_n20042__ = new_new_n20031__ & new_new_n20040__;
  assign new_new_n20043__ = ~new_new_n20041__ & ~new_new_n20042__;
  assign new_new_n20044__ = ~pi59 & ~pi62;
  assign new_new_n20045__ = pi60 & ~new_new_n20044__;
  assign new_new_n20046__ = new_new_n20043__ & ~new_new_n20045__;
  assign new_new_n20047__ = ~pi57 & new_new_n20031__;
  assign new_new_n20048__ = ~pi59 & new_new_n20037__;
  assign new_new_n20049__ = new_new_n20047__ & new_new_n20048__;
  assign new_new_n20050__ = ~pi59 & ~new_new_n19986__;
  assign new_new_n20051__ = pi60 & ~new_new_n20050__;
  assign new_new_n20052__ = ~new_new_n20043__ & new_new_n20051__;
  assign new_new_n20053__ = ~new_new_n20046__ & ~new_new_n20049__;
  assign new_new_n20054__ = ~new_new_n20052__ & new_new_n20053__;
  assign new_new_n20055__ = ~new_new_n20030__ & ~new_new_n20054__;
  assign new_new_n20056__ = new_new_n20030__ & new_new_n20054__;
  assign new_new_n20057__ = ~new_new_n20055__ & ~new_new_n20056__;
  assign new_new_n20058__ = ~new_new_n19976__ & new_new_n19980__;
  assign new_new_n20059__ = new_new_n19980__ & ~new_new_n19990__;
  assign new_new_n20060__ = new_new_n19976__ & ~new_new_n20059__;
  assign new_new_n20061__ = new_new_n19988__ & ~new_new_n20060__;
  assign new_new_n20062__ = ~new_new_n20058__ & ~new_new_n20061__;
  assign new_new_n20063__ = ~new_new_n20057__ & new_new_n20062__;
  assign new_new_n20064__ = new_new_n20057__ & ~new_new_n20062__;
  assign po121 = new_new_n20063__ | new_new_n20064__;
  assign new_new_n20066__ = pi58 & pi63;
  assign new_new_n20067__ = ~pi60 & pi61;
  assign new_new_n20068__ = ~new_new_n19931__ & new_new_n20067__;
  assign new_new_n20069__ = new_new_n19931__ & ~new_new_n20067__;
  assign new_new_n20070__ = ~new_new_n20068__ & ~new_new_n20069__;
  assign new_new_n20071__ = ~new_new_n20032__ & ~new_new_n20036__;
  assign new_new_n20072__ = ~new_new_n20035__ & ~new_new_n20071__;
  assign new_new_n20073__ = pi62 & ~new_new_n20047__;
  assign new_new_n20074__ = ~pi59 & ~new_new_n20073__;
  assign new_new_n20075__ = pi60 & ~new_new_n20042__;
  assign new_new_n20076__ = ~new_new_n20074__ & new_new_n20075__;
  assign new_new_n20077__ = ~new_new_n20041__ & ~new_new_n20076__;
  assign new_new_n20078__ = ~new_new_n20055__ & ~new_new_n20062__;
  assign new_new_n20079__ = ~new_new_n20056__ & ~new_new_n20078__;
  assign new_new_n20080__ = new_new_n20077__ & ~new_new_n20079__;
  assign new_new_n20081__ = ~new_new_n20077__ & new_new_n20079__;
  assign new_new_n20082__ = ~new_new_n20080__ & ~new_new_n20081__;
  assign new_new_n20083__ = ~new_new_n20072__ & new_new_n20082__;
  assign new_new_n20084__ = new_new_n20072__ & ~new_new_n20082__;
  assign new_new_n20085__ = ~new_new_n20083__ & ~new_new_n20084__;
  assign new_new_n20086__ = ~new_new_n20070__ & new_new_n20085__;
  assign new_new_n20087__ = new_new_n20070__ & ~new_new_n20085__;
  assign new_new_n20088__ = new_new_n20066__ & ~new_new_n20086__;
  assign new_new_n20089__ = ~new_new_n20087__ & new_new_n20088__;
  assign new_new_n20090__ = new_new_n20070__ & ~new_new_n20072__;
  assign new_new_n20091__ = new_new_n20080__ & new_new_n20090__;
  assign new_new_n20092__ = new_new_n20072__ & new_new_n20080__;
  assign new_new_n20093__ = ~new_new_n20083__ & ~new_new_n20092__;
  assign new_new_n20094__ = ~new_new_n20070__ & ~new_new_n20093__;
  assign new_new_n20095__ = new_new_n20072__ & ~new_new_n20077__;
  assign new_new_n20096__ = ~new_new_n20072__ & new_new_n20077__;
  assign new_new_n20097__ = new_new_n20070__ & ~new_new_n20096__;
  assign new_new_n20098__ = ~new_new_n20095__ & ~new_new_n20097__;
  assign new_new_n20099__ = new_new_n20079__ & ~new_new_n20098__;
  assign new_new_n20100__ = ~new_new_n20066__ & ~new_new_n20099__;
  assign new_new_n20101__ = ~new_new_n20091__ & new_new_n20100__;
  assign new_new_n20102__ = ~new_new_n20094__ & new_new_n20101__;
  assign po122 = new_new_n20089__ | new_new_n20102__;
  assign new_new_n20104__ = ~pi61 & ~pi62;
  assign new_new_n20105__ = pi60 & ~new_new_n20104__;
  assign new_new_n20106__ = ~pi59 & ~new_new_n20105__;
  assign new_new_n20107__ = pi60 & ~pi61;
  assign new_new_n20108__ = pi63 & ~new_new_n20107__;
  assign new_new_n20109__ = ~pi63 & new_new_n20107__;
  assign new_new_n20110__ = ~new_new_n20108__ & ~new_new_n20109__;
  assign new_new_n20111__ = ~new_new_n20070__ & new_new_n20110__;
  assign new_new_n20112__ = ~new_new_n20106__ & ~new_new_n20111__;
  assign new_new_n20113__ = ~new_new_n20070__ & new_new_n20095__;
  assign new_new_n20114__ = new_new_n20112__ & new_new_n20113__;
  assign new_new_n20115__ = pi60 & pi61;
  assign new_new_n20116__ = pi62 & new_new_n20115__;
  assign new_new_n20117__ = ~pi61 & pi63;
  assign new_new_n20118__ = pi61 & ~pi63;
  assign new_new_n20119__ = pi59 & ~new_new_n20117__;
  assign new_new_n20120__ = ~new_new_n20118__ & new_new_n20119__;
  assign new_new_n20121__ = ~new_new_n20116__ & ~new_new_n20120__;
  assign new_new_n20122__ = new_new_n20070__ & ~new_new_n20121__;
  assign new_new_n20123__ = new_new_n20112__ & ~new_new_n20122__;
  assign new_new_n20124__ = ~new_new_n20070__ & new_new_n20077__;
  assign new_new_n20125__ = ~new_new_n20097__ & ~new_new_n20124__;
  assign new_new_n20126__ = ~new_new_n20123__ & ~new_new_n20125__;
  assign new_new_n20127__ = ~new_new_n20079__ & new_new_n20126__;
  assign new_new_n20128__ = ~new_new_n20114__ & ~new_new_n20127__;
  assign new_new_n20129__ = new_new_n20066__ & ~new_new_n20128__;
  assign new_new_n20130__ = new_new_n20066__ & ~new_new_n20070__;
  assign new_new_n20131__ = new_new_n20123__ & ~new_new_n20130__;
  assign new_new_n20132__ = ~new_new_n20066__ & new_new_n20090__;
  assign new_new_n20133__ = ~new_new_n20131__ & ~new_new_n20132__;
  assign new_new_n20134__ = new_new_n20077__ & ~new_new_n20133__;
  assign new_new_n20135__ = new_new_n20072__ & new_new_n20123__;
  assign new_new_n20136__ = new_new_n20070__ & ~new_new_n20095__;
  assign new_new_n20137__ = new_new_n20066__ & ~new_new_n20096__;
  assign new_new_n20138__ = ~new_new_n20136__ & new_new_n20137__;
  assign new_new_n20139__ = ~new_new_n20113__ & ~new_new_n20123__;
  assign new_new_n20140__ = ~new_new_n20138__ & new_new_n20139__;
  assign new_new_n20141__ = ~new_new_n20135__ & ~new_new_n20140__;
  assign new_new_n20142__ = ~new_new_n20134__ & ~new_new_n20141__;
  assign new_new_n20143__ = new_new_n20079__ & new_new_n20142__;
  assign new_new_n20144__ = ~new_new_n20066__ & new_new_n20070__;
  assign new_new_n20145__ = ~new_new_n20096__ & ~new_new_n20144__;
  assign new_new_n20146__ = new_new_n20131__ & ~new_new_n20145__;
  assign new_new_n20147__ = new_new_n20066__ & ~new_new_n20077__;
  assign new_new_n20148__ = new_new_n20072__ & new_new_n20147__;
  assign new_new_n20149__ = ~new_new_n20070__ & ~new_new_n20112__;
  assign new_new_n20150__ = ~new_new_n20096__ & new_new_n20149__;
  assign new_new_n20151__ = ~new_new_n20148__ & new_new_n20150__;
  assign new_new_n20152__ = ~new_new_n20146__ & ~new_new_n20151__;
  assign new_new_n20153__ = ~new_new_n20079__ & ~new_new_n20152__;
  assign new_new_n20154__ = new_new_n20123__ & new_new_n20144__;
  assign new_new_n20155__ = new_new_n20096__ & new_new_n20154__;
  assign new_new_n20156__ = ~new_new_n20143__ & ~new_new_n20155__;
  assign new_new_n20157__ = ~new_new_n20153__ & new_new_n20156__;
  assign po123 = new_new_n20129__ | ~new_new_n20157__;
  assign new_new_n20159__ = new_new_n20123__ & ~new_new_n20144__;
  assign new_new_n20160__ = ~new_new_n20123__ & ~new_new_n20130__;
  assign new_new_n20161__ = new_new_n20079__ & ~new_new_n20160__;
  assign new_new_n20162__ = ~new_new_n20079__ & ~new_new_n20130__;
  assign new_new_n20163__ = ~new_new_n20077__ & ~new_new_n20162__;
  assign new_new_n20164__ = ~new_new_n20159__ & ~new_new_n20161__;
  assign new_new_n20165__ = ~new_new_n20163__ & new_new_n20164__;
  assign new_new_n20166__ = new_new_n20072__ & ~new_new_n20165__;
  assign new_new_n20167__ = ~new_new_n20080__ & new_new_n20159__;
  assign new_new_n20168__ = new_new_n20066__ & new_new_n20123__;
  assign new_new_n20169__ = new_new_n20079__ & new_new_n20147__;
  assign new_new_n20170__ = ~new_new_n20168__ & ~new_new_n20169__;
  assign new_new_n20171__ = ~new_new_n20070__ & ~new_new_n20170__;
  assign new_new_n20172__ = ~new_new_n20167__ & ~new_new_n20171__;
  assign new_new_n20173__ = ~new_new_n20166__ & new_new_n20172__;
  assign new_new_n20174__ = pi60 & pi63;
  assign new_new_n20175__ = ~pi62 & ~new_new_n20174__;
  assign new_new_n20176__ = ~pi60 & ~pi63;
  assign new_new_n20177__ = pi59 & ~pi62;
  assign new_new_n20178__ = ~new_new_n20176__ & ~new_new_n20177__;
  assign new_new_n20179__ = pi61 & ~new_new_n20178__;
  assign new_new_n20180__ = pi62 & pi63;
  assign new_new_n20181__ = ~pi60 & ~pi61;
  assign new_new_n20182__ = ~pi59 & new_new_n20180__;
  assign new_new_n20183__ = ~new_new_n20181__ & new_new_n20182__;
  assign new_new_n20184__ = ~new_new_n20175__ & ~new_new_n20179__;
  assign new_new_n20185__ = ~new_new_n20183__ & new_new_n20184__;
  assign new_new_n20186__ = new_new_n20173__ & ~new_new_n20185__;
  assign new_new_n20187__ = pi62 & ~new_new_n20174__;
  assign new_new_n20188__ = ~new_new_n20176__ & new_new_n20187__;
  assign new_new_n20189__ = ~new_new_n20107__ & ~new_new_n20188__;
  assign new_new_n20190__ = pi59 & ~new_new_n20189__;
  assign new_new_n20191__ = ~new_new_n19985__ & ~new_new_n20190__;
  assign new_new_n20192__ = ~new_new_n20173__ & ~new_new_n20191__;
  assign po124 = ~new_new_n20186__ & ~new_new_n20192__;
  assign new_new_n20194__ = ~pi61 & ~new_new_n20173__;
  assign new_new_n20195__ = pi62 & ~new_new_n20194__;
  assign new_new_n20196__ = ~new_new_n20173__ & ~new_new_n20180__;
  assign new_new_n20197__ = pi60 & ~new_new_n20196__;
  assign new_new_n20198__ = ~new_new_n20195__ & new_new_n20197__;
  assign new_new_n20199__ = ~pi60 & pi63;
  assign new_new_n20200__ = new_new_n20104__ & new_new_n20199__;
  assign new_new_n20201__ = ~new_new_n20198__ & ~new_new_n20200__;
  assign new_new_n20202__ = pi59 & ~new_new_n20201__;
  assign new_new_n20203__ = pi62 & ~new_new_n20199__;
  assign new_new_n20204__ = ~pi62 & pi63;
  assign new_new_n20205__ = pi59 & ~new_new_n20173__;
  assign new_new_n20206__ = ~new_new_n20203__ & ~new_new_n20204__;
  assign new_new_n20207__ = ~new_new_n20194__ & new_new_n20206__;
  assign new_new_n20208__ = ~new_new_n20205__ & new_new_n20207__;
  assign new_new_n20209__ = pi61 & new_new_n20173__;
  assign new_new_n20210__ = ~new_new_n20115__ & ~new_new_n20173__;
  assign new_new_n20211__ = ~new_new_n20180__ & ~new_new_n20209__;
  assign new_new_n20212__ = ~new_new_n20210__ & new_new_n20211__;
  assign new_new_n20213__ = ~new_new_n20208__ & ~new_new_n20212__;
  assign po125 = ~new_new_n20202__ & new_new_n20213__;
  assign new_new_n20215__ = pi60 & new_new_n20205__;
  assign new_new_n20216__ = ~pi61 & ~new_new_n20215__;
  assign new_new_n20217__ = pi62 & ~new_new_n20216__;
  assign new_new_n20218__ = ~pi59 & new_new_n20173__;
  assign new_new_n20219__ = new_new_n20115__ & ~new_new_n20218__;
  assign new_new_n20220__ = ~pi62 & ~new_new_n20219__;
  assign new_new_n20221__ = ~new_new_n20217__ & ~new_new_n20220__;
  assign po126 = pi63 & ~new_new_n20221__;
  assign po127 = pi63 & ~new_new_n20220__;
  assign po000 = pi00;
  assign po001 = 1'b0;
endmodule


