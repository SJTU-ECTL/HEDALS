// Benchmark "div" written by ABC on Wed Jul 13 18:49:02 2022

module div ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127;
  wire new_new_n257__, new_new_n258__, new_new_n259__, new_new_n260__,
    new_new_n261__, new_new_n262__, new_new_n263__, new_new_n264__,
    new_new_n265__, new_new_n266__, new_new_n267__, new_new_n268__,
    new_new_n269__, new_new_n270__, new_new_n271__, new_new_n272__,
    new_new_n273__, new_new_n274__, new_new_n275__, new_new_n276__,
    new_new_n277__, new_new_n278__, new_new_n279__, new_new_n280__,
    new_new_n281__, new_new_n282__, new_new_n283__, new_new_n284__,
    new_new_n285__, new_new_n286__, new_new_n287__, new_new_n288__,
    new_new_n289__, new_new_n290__, new_new_n291__, new_new_n292__,
    new_new_n293__, new_new_n294__, new_new_n295__, new_new_n296__,
    new_new_n297__, new_new_n298__, new_new_n299__, new_new_n300__,
    new_new_n301__, new_new_n302__, new_new_n303__, new_new_n304__,
    new_new_n305__, new_new_n306__, new_new_n307__, new_new_n308__,
    new_new_n309__, new_new_n310__, new_new_n311__, new_new_n312__,
    new_new_n313__, new_new_n314__, new_new_n315__, new_new_n316__,
    new_new_n317__, new_new_n318__, new_new_n319__, new_new_n320__,
    new_new_n321__, new_new_n322__, new_new_n323__, new_new_n324__,
    new_new_n325__, new_new_n326__, new_new_n327__, new_new_n328__,
    new_new_n329__, new_new_n330__, new_new_n331__, new_new_n332__,
    new_new_n333__, new_new_n334__, new_new_n335__, new_new_n336__,
    new_new_n337__, new_new_n338__, new_new_n339__, new_new_n340__,
    new_new_n342__, new_new_n343__, new_new_n344__, new_new_n345__,
    new_new_n346__, new_new_n347__, new_new_n348__, new_new_n349__,
    new_new_n350__, new_new_n351__, new_new_n352__, new_new_n353__,
    new_new_n354__, new_new_n355__, new_new_n356__, new_new_n357__,
    new_new_n358__, new_new_n359__, new_new_n360__, new_new_n361__,
    new_new_n362__, new_new_n363__, new_new_n364__, new_new_n365__,
    new_new_n366__, new_new_n367__, new_new_n368__, new_new_n369__,
    new_new_n370__, new_new_n371__, new_new_n372__, new_new_n373__,
    new_new_n374__, new_new_n375__, new_new_n376__, new_new_n377__,
    new_new_n378__, new_new_n379__, new_new_n380__, new_new_n381__,
    new_new_n383__, new_new_n384__, new_new_n385__, new_new_n386__,
    new_new_n387__, new_new_n388__, new_new_n389__, new_new_n390__,
    new_new_n391__, new_new_n392__, new_new_n393__, new_new_n394__,
    new_new_n395__, new_new_n396__, new_new_n397__, new_new_n398__,
    new_new_n399__, new_new_n400__, new_new_n401__, new_new_n402__,
    new_new_n403__, new_new_n404__, new_new_n405__, new_new_n406__,
    new_new_n407__, new_new_n408__, new_new_n409__, new_new_n410__,
    new_new_n411__, new_new_n412__, new_new_n413__, new_new_n414__,
    new_new_n415__, new_new_n416__, new_new_n417__, new_new_n418__,
    new_new_n419__, new_new_n420__, new_new_n421__, new_new_n422__,
    new_new_n423__, new_new_n424__, new_new_n426__, new_new_n427__,
    new_new_n428__, new_new_n429__, new_new_n430__, new_new_n431__,
    new_new_n432__, new_new_n433__, new_new_n434__, new_new_n435__,
    new_new_n436__, new_new_n437__, new_new_n438__, new_new_n439__,
    new_new_n440__, new_new_n441__, new_new_n442__, new_new_n443__,
    new_new_n444__, new_new_n445__, new_new_n446__, new_new_n447__,
    new_new_n448__, new_new_n449__, new_new_n450__, new_new_n451__,
    new_new_n452__, new_new_n453__, new_new_n454__, new_new_n455__,
    new_new_n456__, new_new_n457__, new_new_n458__, new_new_n459__,
    new_new_n460__, new_new_n461__, new_new_n462__, new_new_n463__,
    new_new_n464__, new_new_n465__, new_new_n466__, new_new_n467__,
    new_new_n468__, new_new_n469__, new_new_n470__, new_new_n471__,
    new_new_n472__, new_new_n473__, new_new_n474__, new_new_n475__,
    new_new_n476__, new_new_n477__, new_new_n478__, new_new_n479__,
    new_new_n480__, new_new_n481__, new_new_n482__, new_new_n483__,
    new_new_n484__, new_new_n485__, new_new_n486__, new_new_n487__,
    new_new_n488__, new_new_n489__, new_new_n490__, new_new_n491__,
    new_new_n492__, new_new_n493__, new_new_n494__, new_new_n495__,
    new_new_n496__, new_new_n497__, new_new_n498__, new_new_n499__,
    new_new_n501__, new_new_n502__, new_new_n503__, new_new_n504__,
    new_new_n505__, new_new_n506__, new_new_n507__, new_new_n508__,
    new_new_n509__, new_new_n510__, new_new_n511__, new_new_n512__,
    new_new_n513__, new_new_n514__, new_new_n515__, new_new_n516__,
    new_new_n517__, new_new_n518__, new_new_n519__, new_new_n520__,
    new_new_n521__, new_new_n522__, new_new_n523__, new_new_n524__,
    new_new_n525__, new_new_n526__, new_new_n527__, new_new_n528__,
    new_new_n529__, new_new_n530__, new_new_n531__, new_new_n532__,
    new_new_n533__, new_new_n534__, new_new_n535__, new_new_n536__,
    new_new_n537__, new_new_n538__, new_new_n539__, new_new_n540__,
    new_new_n541__, new_new_n542__, new_new_n543__, new_new_n544__,
    new_new_n545__, new_new_n546__, new_new_n547__, new_new_n548__,
    new_new_n549__, new_new_n550__, new_new_n551__, new_new_n552__,
    new_new_n553__, new_new_n554__, new_new_n555__, new_new_n556__,
    new_new_n557__, new_new_n558__, new_new_n559__, new_new_n560__,
    new_new_n561__, new_new_n562__, new_new_n563__, new_new_n564__,
    new_new_n565__, new_new_n566__, new_new_n567__, new_new_n568__,
    new_new_n569__, new_new_n570__, new_new_n571__, new_new_n572__,
    new_new_n573__, new_new_n574__, new_new_n575__, new_new_n576__,
    new_new_n577__, new_new_n578__, new_new_n579__, new_new_n581__,
    new_new_n582__, new_new_n583__, new_new_n584__, new_new_n585__,
    new_new_n586__, new_new_n587__, new_new_n588__, new_new_n589__,
    new_new_n590__, new_new_n591__, new_new_n592__, new_new_n593__,
    new_new_n594__, new_new_n595__, new_new_n596__, new_new_n597__,
    new_new_n598__, new_new_n599__, new_new_n600__, new_new_n601__,
    new_new_n602__, new_new_n603__, new_new_n604__, new_new_n605__,
    new_new_n606__, new_new_n607__, new_new_n608__, new_new_n609__,
    new_new_n610__, new_new_n611__, new_new_n612__, new_new_n613__,
    new_new_n614__, new_new_n615__, new_new_n616__, new_new_n617__,
    new_new_n618__, new_new_n619__, new_new_n620__, new_new_n621__,
    new_new_n622__, new_new_n623__, new_new_n624__, new_new_n625__,
    new_new_n626__, new_new_n627__, new_new_n628__, new_new_n629__,
    new_new_n630__, new_new_n631__, new_new_n632__, new_new_n633__,
    new_new_n634__, new_new_n635__, new_new_n636__, new_new_n637__,
    new_new_n638__, new_new_n639__, new_new_n640__, new_new_n641__,
    new_new_n642__, new_new_n643__, new_new_n644__, new_new_n645__,
    new_new_n646__, new_new_n647__, new_new_n648__, new_new_n649__,
    new_new_n650__, new_new_n651__, new_new_n652__, new_new_n653__,
    new_new_n654__, new_new_n655__, new_new_n656__, new_new_n657__,
    new_new_n658__, new_new_n659__, new_new_n660__, new_new_n661__,
    new_new_n662__, new_new_n663__, new_new_n664__, new_new_n665__,
    new_new_n666__, new_new_n667__, new_new_n668__, new_new_n669__,
    new_new_n670__, new_new_n671__, new_new_n672__, new_new_n673__,
    new_new_n674__, new_new_n676__, new_new_n677__, new_new_n678__,
    new_new_n679__, new_new_n680__, new_new_n681__, new_new_n682__,
    new_new_n683__, new_new_n684__, new_new_n685__, new_new_n686__,
    new_new_n687__, new_new_n688__, new_new_n689__, new_new_n690__,
    new_new_n691__, new_new_n692__, new_new_n693__, new_new_n694__,
    new_new_n695__, new_new_n696__, new_new_n697__, new_new_n698__,
    new_new_n699__, new_new_n700__, new_new_n701__, new_new_n702__,
    new_new_n703__, new_new_n704__, new_new_n705__, new_new_n706__,
    new_new_n707__, new_new_n708__, new_new_n709__, new_new_n710__,
    new_new_n711__, new_new_n712__, new_new_n713__, new_new_n714__,
    new_new_n715__, new_new_n716__, new_new_n717__, new_new_n718__,
    new_new_n719__, new_new_n720__, new_new_n721__, new_new_n722__,
    new_new_n723__, new_new_n724__, new_new_n725__, new_new_n726__,
    new_new_n727__, new_new_n728__, new_new_n729__, new_new_n730__,
    new_new_n731__, new_new_n732__, new_new_n733__, new_new_n734__,
    new_new_n735__, new_new_n736__, new_new_n737__, new_new_n738__,
    new_new_n739__, new_new_n740__, new_new_n741__, new_new_n742__,
    new_new_n743__, new_new_n744__, new_new_n745__, new_new_n746__,
    new_new_n747__, new_new_n748__, new_new_n749__, new_new_n750__,
    new_new_n751__, new_new_n752__, new_new_n753__, new_new_n754__,
    new_new_n755__, new_new_n756__, new_new_n757__, new_new_n758__,
    new_new_n759__, new_new_n760__, new_new_n761__, new_new_n762__,
    new_new_n764__, new_new_n765__, new_new_n766__, new_new_n767__,
    new_new_n768__, new_new_n769__, new_new_n770__, new_new_n771__,
    new_new_n772__, new_new_n773__, new_new_n774__, new_new_n775__,
    new_new_n776__, new_new_n777__, new_new_n778__, new_new_n779__,
    new_new_n780__, new_new_n781__, new_new_n782__, new_new_n783__,
    new_new_n784__, new_new_n785__, new_new_n786__, new_new_n787__,
    new_new_n788__, new_new_n789__, new_new_n790__, new_new_n791__,
    new_new_n792__, new_new_n793__, new_new_n794__, new_new_n795__,
    new_new_n796__, new_new_n797__, new_new_n798__, new_new_n799__,
    new_new_n800__, new_new_n801__, new_new_n802__, new_new_n803__,
    new_new_n804__, new_new_n805__, new_new_n806__, new_new_n807__,
    new_new_n808__, new_new_n809__, new_new_n810__, new_new_n811__,
    new_new_n812__, new_new_n813__, new_new_n814__, new_new_n815__,
    new_new_n816__, new_new_n817__, new_new_n818__, new_new_n819__,
    new_new_n820__, new_new_n821__, new_new_n822__, new_new_n823__,
    new_new_n824__, new_new_n825__, new_new_n826__, new_new_n827__,
    new_new_n828__, new_new_n829__, new_new_n830__, new_new_n831__,
    new_new_n832__, new_new_n833__, new_new_n834__, new_new_n835__,
    new_new_n836__, new_new_n837__, new_new_n838__, new_new_n839__,
    new_new_n840__, new_new_n841__, new_new_n842__, new_new_n843__,
    new_new_n844__, new_new_n845__, new_new_n846__, new_new_n847__,
    new_new_n848__, new_new_n849__, new_new_n850__, new_new_n851__,
    new_new_n852__, new_new_n853__, new_new_n854__, new_new_n855__,
    new_new_n856__, new_new_n857__, new_new_n858__, new_new_n859__,
    new_new_n860__, new_new_n861__, new_new_n862__, new_new_n863__,
    new_new_n864__, new_new_n865__, new_new_n866__, new_new_n867__,
    new_new_n868__, new_new_n869__, new_new_n870__, new_new_n871__,
    new_new_n872__, new_new_n873__, new_new_n875__, new_new_n876__,
    new_new_n877__, new_new_n878__, new_new_n879__, new_new_n880__,
    new_new_n881__, new_new_n882__, new_new_n883__, new_new_n884__,
    new_new_n885__, new_new_n886__, new_new_n887__, new_new_n888__,
    new_new_n889__, new_new_n890__, new_new_n891__, new_new_n892__,
    new_new_n893__, new_new_n894__, new_new_n895__, new_new_n896__,
    new_new_n897__, new_new_n898__, new_new_n899__, new_new_n900__,
    new_new_n901__, new_new_n902__, new_new_n903__, new_new_n904__,
    new_new_n905__, new_new_n906__, new_new_n907__, new_new_n908__,
    new_new_n909__, new_new_n910__, new_new_n911__, new_new_n912__,
    new_new_n913__, new_new_n914__, new_new_n915__, new_new_n916__,
    new_new_n917__, new_new_n918__, new_new_n919__, new_new_n920__,
    new_new_n921__, new_new_n922__, new_new_n923__, new_new_n924__,
    new_new_n925__, new_new_n926__, new_new_n927__, new_new_n928__,
    new_new_n929__, new_new_n930__, new_new_n931__, new_new_n932__,
    new_new_n933__, new_new_n934__, new_new_n935__, new_new_n936__,
    new_new_n937__, new_new_n938__, new_new_n939__, new_new_n940__,
    new_new_n941__, new_new_n942__, new_new_n943__, new_new_n944__,
    new_new_n945__, new_new_n946__, new_new_n947__, new_new_n948__,
    new_new_n949__, new_new_n950__, new_new_n951__, new_new_n952__,
    new_new_n953__, new_new_n954__, new_new_n955__, new_new_n956__,
    new_new_n957__, new_new_n958__, new_new_n959__, new_new_n960__,
    new_new_n961__, new_new_n962__, new_new_n963__, new_new_n964__,
    new_new_n965__, new_new_n966__, new_new_n967__, new_new_n968__,
    new_new_n969__, new_new_n970__, new_new_n971__, new_new_n972__,
    new_new_n973__, new_new_n974__, new_new_n975__, new_new_n976__,
    new_new_n977__, new_new_n978__, new_new_n979__, new_new_n980__,
    new_new_n981__, new_new_n982__, new_new_n983__, new_new_n984__,
    new_new_n985__, new_new_n986__, new_new_n987__, new_new_n988__,
    new_new_n989__, new_new_n990__, new_new_n991__, new_new_n992__,
    new_new_n993__, new_new_n994__, new_new_n995__, new_new_n996__,
    new_new_n997__, new_new_n998__, new_new_n1000__, new_new_n1001__,
    new_new_n1002__, new_new_n1003__, new_new_n1004__, new_new_n1005__,
    new_new_n1006__, new_new_n1007__, new_new_n1008__, new_new_n1009__,
    new_new_n1010__, new_new_n1011__, new_new_n1012__, new_new_n1013__,
    new_new_n1014__, new_new_n1015__, new_new_n1016__, new_new_n1017__,
    new_new_n1018__, new_new_n1019__, new_new_n1020__, new_new_n1021__,
    new_new_n1022__, new_new_n1023__, new_new_n1024__, new_new_n1025__,
    new_new_n1026__, new_new_n1027__, new_new_n1028__, new_new_n1029__,
    new_new_n1030__, new_new_n1031__, new_new_n1032__, new_new_n1033__,
    new_new_n1034__, new_new_n1035__, new_new_n1036__, new_new_n1037__,
    new_new_n1038__, new_new_n1039__, new_new_n1040__, new_new_n1041__,
    new_new_n1042__, new_new_n1043__, new_new_n1044__, new_new_n1045__,
    new_new_n1046__, new_new_n1047__, new_new_n1048__, new_new_n1049__,
    new_new_n1050__, new_new_n1051__, new_new_n1052__, new_new_n1053__,
    new_new_n1054__, new_new_n1055__, new_new_n1056__, new_new_n1057__,
    new_new_n1058__, new_new_n1059__, new_new_n1060__, new_new_n1061__,
    new_new_n1062__, new_new_n1063__, new_new_n1064__, new_new_n1065__,
    new_new_n1066__, new_new_n1067__, new_new_n1068__, new_new_n1069__,
    new_new_n1070__, new_new_n1071__, new_new_n1072__, new_new_n1073__,
    new_new_n1074__, new_new_n1075__, new_new_n1076__, new_new_n1077__,
    new_new_n1078__, new_new_n1079__, new_new_n1080__, new_new_n1081__,
    new_new_n1082__, new_new_n1083__, new_new_n1084__, new_new_n1085__,
    new_new_n1086__, new_new_n1087__, new_new_n1088__, new_new_n1089__,
    new_new_n1090__, new_new_n1091__, new_new_n1092__, new_new_n1093__,
    new_new_n1094__, new_new_n1095__, new_new_n1096__, new_new_n1097__,
    new_new_n1098__, new_new_n1099__, new_new_n1100__, new_new_n1101__,
    new_new_n1102__, new_new_n1103__, new_new_n1104__, new_new_n1105__,
    new_new_n1106__, new_new_n1107__, new_new_n1108__, new_new_n1109__,
    new_new_n1110__, new_new_n1111__, new_new_n1112__, new_new_n1113__,
    new_new_n1114__, new_new_n1115__, new_new_n1116__, new_new_n1117__,
    new_new_n1118__, new_new_n1119__, new_new_n1120__, new_new_n1121__,
    new_new_n1122__, new_new_n1123__, new_new_n1124__, new_new_n1125__,
    new_new_n1126__, new_new_n1127__, new_new_n1128__, new_new_n1129__,
    new_new_n1130__, new_new_n1131__, new_new_n1132__, new_new_n1133__,
    new_new_n1135__, new_new_n1136__, new_new_n1137__, new_new_n1138__,
    new_new_n1139__, new_new_n1140__, new_new_n1141__, new_new_n1142__,
    new_new_n1143__, new_new_n1144__, new_new_n1145__, new_new_n1146__,
    new_new_n1147__, new_new_n1148__, new_new_n1149__, new_new_n1150__,
    new_new_n1151__, new_new_n1152__, new_new_n1153__, new_new_n1154__,
    new_new_n1155__, new_new_n1156__, new_new_n1157__, new_new_n1158__,
    new_new_n1159__, new_new_n1160__, new_new_n1161__, new_new_n1162__,
    new_new_n1163__, new_new_n1164__, new_new_n1165__, new_new_n1166__,
    new_new_n1167__, new_new_n1168__, new_new_n1169__, new_new_n1170__,
    new_new_n1171__, new_new_n1172__, new_new_n1173__, new_new_n1174__,
    new_new_n1175__, new_new_n1176__, new_new_n1177__, new_new_n1178__,
    new_new_n1179__, new_new_n1180__, new_new_n1181__, new_new_n1182__,
    new_new_n1183__, new_new_n1184__, new_new_n1185__, new_new_n1186__,
    new_new_n1187__, new_new_n1188__, new_new_n1189__, new_new_n1190__,
    new_new_n1191__, new_new_n1192__, new_new_n1193__, new_new_n1194__,
    new_new_n1195__, new_new_n1196__, new_new_n1197__, new_new_n1198__,
    new_new_n1199__, new_new_n1200__, new_new_n1201__, new_new_n1202__,
    new_new_n1203__, new_new_n1204__, new_new_n1205__, new_new_n1206__,
    new_new_n1207__, new_new_n1208__, new_new_n1209__, new_new_n1210__,
    new_new_n1211__, new_new_n1212__, new_new_n1213__, new_new_n1214__,
    new_new_n1215__, new_new_n1216__, new_new_n1217__, new_new_n1218__,
    new_new_n1219__, new_new_n1220__, new_new_n1221__, new_new_n1222__,
    new_new_n1223__, new_new_n1224__, new_new_n1225__, new_new_n1226__,
    new_new_n1227__, new_new_n1228__, new_new_n1229__, new_new_n1230__,
    new_new_n1231__, new_new_n1232__, new_new_n1233__, new_new_n1234__,
    new_new_n1235__, new_new_n1236__, new_new_n1237__, new_new_n1238__,
    new_new_n1239__, new_new_n1240__, new_new_n1241__, new_new_n1242__,
    new_new_n1243__, new_new_n1244__, new_new_n1245__, new_new_n1246__,
    new_new_n1247__, new_new_n1248__, new_new_n1249__, new_new_n1250__,
    new_new_n1251__, new_new_n1252__, new_new_n1253__, new_new_n1254__,
    new_new_n1255__, new_new_n1256__, new_new_n1257__, new_new_n1258__,
    new_new_n1259__, new_new_n1260__, new_new_n1261__, new_new_n1262__,
    new_new_n1263__, new_new_n1264__, new_new_n1265__, new_new_n1266__,
    new_new_n1267__, new_new_n1268__, new_new_n1269__, new_new_n1270__,
    new_new_n1271__, new_new_n1272__, new_new_n1273__, new_new_n1274__,
    new_new_n1275__, new_new_n1276__, new_new_n1277__, new_new_n1279__,
    new_new_n1280__, new_new_n1281__, new_new_n1282__, new_new_n1283__,
    new_new_n1284__, new_new_n1285__, new_new_n1286__, new_new_n1287__,
    new_new_n1288__, new_new_n1289__, new_new_n1290__, new_new_n1291__,
    new_new_n1292__, new_new_n1293__, new_new_n1294__, new_new_n1295__,
    new_new_n1296__, new_new_n1297__, new_new_n1298__, new_new_n1299__,
    new_new_n1300__, new_new_n1301__, new_new_n1302__, new_new_n1303__,
    new_new_n1304__, new_new_n1305__, new_new_n1306__, new_new_n1307__,
    new_new_n1308__, new_new_n1309__, new_new_n1310__, new_new_n1311__,
    new_new_n1312__, new_new_n1313__, new_new_n1314__, new_new_n1315__,
    new_new_n1316__, new_new_n1317__, new_new_n1318__, new_new_n1319__,
    new_new_n1320__, new_new_n1321__, new_new_n1322__, new_new_n1323__,
    new_new_n1324__, new_new_n1325__, new_new_n1326__, new_new_n1327__,
    new_new_n1328__, new_new_n1329__, new_new_n1330__, new_new_n1331__,
    new_new_n1332__, new_new_n1333__, new_new_n1334__, new_new_n1335__,
    new_new_n1336__, new_new_n1337__, new_new_n1338__, new_new_n1339__,
    new_new_n1340__, new_new_n1341__, new_new_n1342__, new_new_n1343__,
    new_new_n1344__, new_new_n1345__, new_new_n1346__, new_new_n1347__,
    new_new_n1348__, new_new_n1349__, new_new_n1350__, new_new_n1351__,
    new_new_n1352__, new_new_n1353__, new_new_n1354__, new_new_n1355__,
    new_new_n1356__, new_new_n1357__, new_new_n1358__, new_new_n1359__,
    new_new_n1360__, new_new_n1361__, new_new_n1362__, new_new_n1363__,
    new_new_n1364__, new_new_n1365__, new_new_n1366__, new_new_n1367__,
    new_new_n1368__, new_new_n1369__, new_new_n1370__, new_new_n1371__,
    new_new_n1372__, new_new_n1373__, new_new_n1374__, new_new_n1375__,
    new_new_n1376__, new_new_n1377__, new_new_n1378__, new_new_n1379__,
    new_new_n1380__, new_new_n1381__, new_new_n1382__, new_new_n1383__,
    new_new_n1384__, new_new_n1385__, new_new_n1386__, new_new_n1387__,
    new_new_n1388__, new_new_n1389__, new_new_n1390__, new_new_n1391__,
    new_new_n1392__, new_new_n1393__, new_new_n1394__, new_new_n1395__,
    new_new_n1396__, new_new_n1397__, new_new_n1398__, new_new_n1399__,
    new_new_n1400__, new_new_n1401__, new_new_n1402__, new_new_n1403__,
    new_new_n1404__, new_new_n1405__, new_new_n1406__, new_new_n1407__,
    new_new_n1408__, new_new_n1409__, new_new_n1410__, new_new_n1411__,
    new_new_n1412__, new_new_n1413__, new_new_n1414__, new_new_n1415__,
    new_new_n1416__, new_new_n1417__, new_new_n1418__, new_new_n1419__,
    new_new_n1420__, new_new_n1421__, new_new_n1422__, new_new_n1423__,
    new_new_n1424__, new_new_n1425__, new_new_n1426__, new_new_n1427__,
    new_new_n1428__, new_new_n1429__, new_new_n1430__, new_new_n1431__,
    new_new_n1433__, new_new_n1434__, new_new_n1435__, new_new_n1436__,
    new_new_n1437__, new_new_n1438__, new_new_n1439__, new_new_n1440__,
    new_new_n1441__, new_new_n1442__, new_new_n1443__, new_new_n1444__,
    new_new_n1445__, new_new_n1446__, new_new_n1447__, new_new_n1448__,
    new_new_n1449__, new_new_n1450__, new_new_n1451__, new_new_n1452__,
    new_new_n1453__, new_new_n1454__, new_new_n1455__, new_new_n1456__,
    new_new_n1457__, new_new_n1458__, new_new_n1459__, new_new_n1460__,
    new_new_n1461__, new_new_n1462__, new_new_n1463__, new_new_n1464__,
    new_new_n1465__, new_new_n1466__, new_new_n1467__, new_new_n1468__,
    new_new_n1469__, new_new_n1470__, new_new_n1471__, new_new_n1472__,
    new_new_n1473__, new_new_n1474__, new_new_n1475__, new_new_n1476__,
    new_new_n1477__, new_new_n1478__, new_new_n1479__, new_new_n1480__,
    new_new_n1481__, new_new_n1482__, new_new_n1483__, new_new_n1484__,
    new_new_n1485__, new_new_n1486__, new_new_n1487__, new_new_n1488__,
    new_new_n1489__, new_new_n1490__, new_new_n1491__, new_new_n1492__,
    new_new_n1493__, new_new_n1494__, new_new_n1495__, new_new_n1496__,
    new_new_n1497__, new_new_n1498__, new_new_n1499__, new_new_n1500__,
    new_new_n1501__, new_new_n1502__, new_new_n1503__, new_new_n1504__,
    new_new_n1505__, new_new_n1506__, new_new_n1507__, new_new_n1508__,
    new_new_n1509__, new_new_n1510__, new_new_n1511__, new_new_n1512__,
    new_new_n1513__, new_new_n1514__, new_new_n1515__, new_new_n1516__,
    new_new_n1517__, new_new_n1518__, new_new_n1519__, new_new_n1520__,
    new_new_n1521__, new_new_n1522__, new_new_n1523__, new_new_n1524__,
    new_new_n1525__, new_new_n1526__, new_new_n1527__, new_new_n1528__,
    new_new_n1529__, new_new_n1530__, new_new_n1531__, new_new_n1532__,
    new_new_n1533__, new_new_n1534__, new_new_n1535__, new_new_n1536__,
    new_new_n1537__, new_new_n1538__, new_new_n1539__, new_new_n1540__,
    new_new_n1541__, new_new_n1542__, new_new_n1543__, new_new_n1544__,
    new_new_n1545__, new_new_n1546__, new_new_n1547__, new_new_n1548__,
    new_new_n1549__, new_new_n1550__, new_new_n1551__, new_new_n1552__,
    new_new_n1553__, new_new_n1554__, new_new_n1555__, new_new_n1556__,
    new_new_n1557__, new_new_n1558__, new_new_n1559__, new_new_n1560__,
    new_new_n1561__, new_new_n1562__, new_new_n1563__, new_new_n1564__,
    new_new_n1565__, new_new_n1566__, new_new_n1567__, new_new_n1568__,
    new_new_n1569__, new_new_n1570__, new_new_n1571__, new_new_n1572__,
    new_new_n1573__, new_new_n1574__, new_new_n1575__, new_new_n1576__,
    new_new_n1577__, new_new_n1578__, new_new_n1579__, new_new_n1580__,
    new_new_n1581__, new_new_n1582__, new_new_n1583__, new_new_n1584__,
    new_new_n1585__, new_new_n1586__, new_new_n1587__, new_new_n1588__,
    new_new_n1589__, new_new_n1590__, new_new_n1591__, new_new_n1592__,
    new_new_n1593__, new_new_n1594__, new_new_n1595__, new_new_n1596__,
    new_new_n1597__, new_new_n1598__, new_new_n1599__, new_new_n1600__,
    new_new_n1601__, new_new_n1602__, new_new_n1603__, new_new_n1604__,
    new_new_n1605__, new_new_n1607__, new_new_n1608__, new_new_n1609__,
    new_new_n1610__, new_new_n1611__, new_new_n1612__, new_new_n1613__,
    new_new_n1614__, new_new_n1615__, new_new_n1616__, new_new_n1617__,
    new_new_n1618__, new_new_n1619__, new_new_n1620__, new_new_n1621__,
    new_new_n1622__, new_new_n1623__, new_new_n1624__, new_new_n1625__,
    new_new_n1626__, new_new_n1627__, new_new_n1628__, new_new_n1629__,
    new_new_n1630__, new_new_n1631__, new_new_n1632__, new_new_n1633__,
    new_new_n1634__, new_new_n1635__, new_new_n1636__, new_new_n1637__,
    new_new_n1638__, new_new_n1639__, new_new_n1640__, new_new_n1641__,
    new_new_n1642__, new_new_n1643__, new_new_n1644__, new_new_n1645__,
    new_new_n1646__, new_new_n1647__, new_new_n1648__, new_new_n1649__,
    new_new_n1650__, new_new_n1651__, new_new_n1652__, new_new_n1653__,
    new_new_n1654__, new_new_n1655__, new_new_n1656__, new_new_n1657__,
    new_new_n1658__, new_new_n1659__, new_new_n1660__, new_new_n1661__,
    new_new_n1662__, new_new_n1663__, new_new_n1664__, new_new_n1665__,
    new_new_n1666__, new_new_n1667__, new_new_n1668__, new_new_n1669__,
    new_new_n1670__, new_new_n1671__, new_new_n1672__, new_new_n1673__,
    new_new_n1674__, new_new_n1675__, new_new_n1676__, new_new_n1677__,
    new_new_n1678__, new_new_n1679__, new_new_n1680__, new_new_n1681__,
    new_new_n1682__, new_new_n1683__, new_new_n1684__, new_new_n1685__,
    new_new_n1686__, new_new_n1687__, new_new_n1688__, new_new_n1689__,
    new_new_n1690__, new_new_n1691__, new_new_n1692__, new_new_n1693__,
    new_new_n1694__, new_new_n1695__, new_new_n1696__, new_new_n1697__,
    new_new_n1698__, new_new_n1699__, new_new_n1700__, new_new_n1701__,
    new_new_n1702__, new_new_n1703__, new_new_n1704__, new_new_n1705__,
    new_new_n1706__, new_new_n1707__, new_new_n1708__, new_new_n1709__,
    new_new_n1710__, new_new_n1711__, new_new_n1712__, new_new_n1713__,
    new_new_n1714__, new_new_n1715__, new_new_n1716__, new_new_n1717__,
    new_new_n1718__, new_new_n1719__, new_new_n1720__, new_new_n1721__,
    new_new_n1722__, new_new_n1723__, new_new_n1724__, new_new_n1725__,
    new_new_n1726__, new_new_n1727__, new_new_n1728__, new_new_n1729__,
    new_new_n1730__, new_new_n1731__, new_new_n1732__, new_new_n1733__,
    new_new_n1734__, new_new_n1735__, new_new_n1736__, new_new_n1737__,
    new_new_n1738__, new_new_n1739__, new_new_n1740__, new_new_n1741__,
    new_new_n1742__, new_new_n1743__, new_new_n1744__, new_new_n1745__,
    new_new_n1746__, new_new_n1747__, new_new_n1748__, new_new_n1749__,
    new_new_n1750__, new_new_n1751__, new_new_n1752__, new_new_n1753__,
    new_new_n1754__, new_new_n1755__, new_new_n1756__, new_new_n1757__,
    new_new_n1758__, new_new_n1759__, new_new_n1760__, new_new_n1761__,
    new_new_n1762__, new_new_n1763__, new_new_n1764__, new_new_n1765__,
    new_new_n1766__, new_new_n1767__, new_new_n1768__, new_new_n1769__,
    new_new_n1770__, new_new_n1771__, new_new_n1772__, new_new_n1773__,
    new_new_n1774__, new_new_n1775__, new_new_n1776__, new_new_n1777__,
    new_new_n1778__, new_new_n1779__, new_new_n1780__, new_new_n1782__,
    new_new_n1783__, new_new_n1784__, new_new_n1785__, new_new_n1786__,
    new_new_n1787__, new_new_n1788__, new_new_n1789__, new_new_n1790__,
    new_new_n1791__, new_new_n1792__, new_new_n1793__, new_new_n1794__,
    new_new_n1795__, new_new_n1796__, new_new_n1797__, new_new_n1798__,
    new_new_n1799__, new_new_n1800__, new_new_n1801__, new_new_n1802__,
    new_new_n1803__, new_new_n1804__, new_new_n1805__, new_new_n1806__,
    new_new_n1807__, new_new_n1808__, new_new_n1809__, new_new_n1810__,
    new_new_n1811__, new_new_n1812__, new_new_n1813__, new_new_n1814__,
    new_new_n1815__, new_new_n1816__, new_new_n1817__, new_new_n1818__,
    new_new_n1819__, new_new_n1820__, new_new_n1821__, new_new_n1822__,
    new_new_n1823__, new_new_n1824__, new_new_n1825__, new_new_n1826__,
    new_new_n1827__, new_new_n1828__, new_new_n1829__, new_new_n1830__,
    new_new_n1831__, new_new_n1832__, new_new_n1833__, new_new_n1834__,
    new_new_n1835__, new_new_n1836__, new_new_n1837__, new_new_n1838__,
    new_new_n1839__, new_new_n1840__, new_new_n1841__, new_new_n1842__,
    new_new_n1843__, new_new_n1844__, new_new_n1845__, new_new_n1846__,
    new_new_n1847__, new_new_n1848__, new_new_n1849__, new_new_n1850__,
    new_new_n1851__, new_new_n1852__, new_new_n1853__, new_new_n1854__,
    new_new_n1855__, new_new_n1856__, new_new_n1857__, new_new_n1858__,
    new_new_n1859__, new_new_n1860__, new_new_n1861__, new_new_n1862__,
    new_new_n1863__, new_new_n1864__, new_new_n1865__, new_new_n1866__,
    new_new_n1867__, new_new_n1868__, new_new_n1869__, new_new_n1870__,
    new_new_n1871__, new_new_n1872__, new_new_n1873__, new_new_n1874__,
    new_new_n1875__, new_new_n1876__, new_new_n1877__, new_new_n1878__,
    new_new_n1879__, new_new_n1880__, new_new_n1881__, new_new_n1882__,
    new_new_n1883__, new_new_n1884__, new_new_n1885__, new_new_n1886__,
    new_new_n1887__, new_new_n1888__, new_new_n1889__, new_new_n1890__,
    new_new_n1891__, new_new_n1892__, new_new_n1893__, new_new_n1894__,
    new_new_n1895__, new_new_n1896__, new_new_n1897__, new_new_n1898__,
    new_new_n1899__, new_new_n1900__, new_new_n1901__, new_new_n1902__,
    new_new_n1903__, new_new_n1904__, new_new_n1905__, new_new_n1906__,
    new_new_n1907__, new_new_n1908__, new_new_n1909__, new_new_n1910__,
    new_new_n1911__, new_new_n1912__, new_new_n1913__, new_new_n1914__,
    new_new_n1915__, new_new_n1916__, new_new_n1917__, new_new_n1918__,
    new_new_n1919__, new_new_n1920__, new_new_n1921__, new_new_n1922__,
    new_new_n1923__, new_new_n1924__, new_new_n1925__, new_new_n1926__,
    new_new_n1927__, new_new_n1928__, new_new_n1929__, new_new_n1930__,
    new_new_n1931__, new_new_n1932__, new_new_n1933__, new_new_n1934__,
    new_new_n1935__, new_new_n1936__, new_new_n1937__, new_new_n1938__,
    new_new_n1939__, new_new_n1940__, new_new_n1941__, new_new_n1942__,
    new_new_n1943__, new_new_n1944__, new_new_n1945__, new_new_n1946__,
    new_new_n1947__, new_new_n1948__, new_new_n1949__, new_new_n1950__,
    new_new_n1951__, new_new_n1952__, new_new_n1953__, new_new_n1954__,
    new_new_n1955__, new_new_n1956__, new_new_n1957__, new_new_n1958__,
    new_new_n1959__, new_new_n1960__, new_new_n1961__, new_new_n1962__,
    new_new_n1963__, new_new_n1964__, new_new_n1965__, new_new_n1966__,
    new_new_n1967__, new_new_n1968__, new_new_n1970__, new_new_n1971__,
    new_new_n1972__, new_new_n1973__, new_new_n1974__, new_new_n1975__,
    new_new_n1976__, new_new_n1977__, new_new_n1978__, new_new_n1979__,
    new_new_n1980__, new_new_n1981__, new_new_n1982__, new_new_n1983__,
    new_new_n1984__, new_new_n1985__, new_new_n1986__, new_new_n1987__,
    new_new_n1988__, new_new_n1989__, new_new_n1990__, new_new_n1991__,
    new_new_n1992__, new_new_n1993__, new_new_n1994__, new_new_n1995__,
    new_new_n1996__, new_new_n1997__, new_new_n1998__, new_new_n1999__,
    new_new_n2000__, new_new_n2001__, new_new_n2002__, new_new_n2003__,
    new_new_n2004__, new_new_n2005__, new_new_n2006__, new_new_n2007__,
    new_new_n2008__, new_new_n2009__, new_new_n2010__, new_new_n2011__,
    new_new_n2012__, new_new_n2013__, new_new_n2014__, new_new_n2015__,
    new_new_n2016__, new_new_n2017__, new_new_n2018__, new_new_n2019__,
    new_new_n2020__, new_new_n2021__, new_new_n2022__, new_new_n2023__,
    new_new_n2024__, new_new_n2025__, new_new_n2026__, new_new_n2027__,
    new_new_n2028__, new_new_n2029__, new_new_n2030__, new_new_n2031__,
    new_new_n2032__, new_new_n2033__, new_new_n2034__, new_new_n2035__,
    new_new_n2036__, new_new_n2037__, new_new_n2038__, new_new_n2039__,
    new_new_n2040__, new_new_n2041__, new_new_n2042__, new_new_n2043__,
    new_new_n2044__, new_new_n2045__, new_new_n2046__, new_new_n2047__,
    new_new_n2048__, new_new_n2049__, new_new_n2050__, new_new_n2051__,
    new_new_n2052__, new_new_n2053__, new_new_n2054__, new_new_n2055__,
    new_new_n2056__, new_new_n2057__, new_new_n2058__, new_new_n2059__,
    new_new_n2060__, new_new_n2061__, new_new_n2062__, new_new_n2063__,
    new_new_n2064__, new_new_n2065__, new_new_n2066__, new_new_n2067__,
    new_new_n2068__, new_new_n2069__, new_new_n2070__, new_new_n2071__,
    new_new_n2072__, new_new_n2073__, new_new_n2074__, new_new_n2075__,
    new_new_n2076__, new_new_n2077__, new_new_n2078__, new_new_n2079__,
    new_new_n2080__, new_new_n2081__, new_new_n2082__, new_new_n2083__,
    new_new_n2084__, new_new_n2085__, new_new_n2086__, new_new_n2087__,
    new_new_n2088__, new_new_n2089__, new_new_n2090__, new_new_n2091__,
    new_new_n2092__, new_new_n2093__, new_new_n2094__, new_new_n2095__,
    new_new_n2096__, new_new_n2097__, new_new_n2098__, new_new_n2099__,
    new_new_n2100__, new_new_n2101__, new_new_n2102__, new_new_n2103__,
    new_new_n2104__, new_new_n2105__, new_new_n2106__, new_new_n2107__,
    new_new_n2108__, new_new_n2109__, new_new_n2110__, new_new_n2111__,
    new_new_n2112__, new_new_n2113__, new_new_n2114__, new_new_n2115__,
    new_new_n2116__, new_new_n2117__, new_new_n2118__, new_new_n2119__,
    new_new_n2120__, new_new_n2121__, new_new_n2122__, new_new_n2123__,
    new_new_n2124__, new_new_n2125__, new_new_n2126__, new_new_n2127__,
    new_new_n2128__, new_new_n2129__, new_new_n2130__, new_new_n2131__,
    new_new_n2132__, new_new_n2133__, new_new_n2134__, new_new_n2135__,
    new_new_n2136__, new_new_n2137__, new_new_n2138__, new_new_n2139__,
    new_new_n2140__, new_new_n2141__, new_new_n2142__, new_new_n2143__,
    new_new_n2144__, new_new_n2145__, new_new_n2146__, new_new_n2147__,
    new_new_n2148__, new_new_n2149__, new_new_n2150__, new_new_n2151__,
    new_new_n2152__, new_new_n2153__, new_new_n2154__, new_new_n2155__,
    new_new_n2156__, new_new_n2157__, new_new_n2158__, new_new_n2159__,
    new_new_n2160__, new_new_n2161__, new_new_n2162__, new_new_n2163__,
    new_new_n2164__, new_new_n2165__, new_new_n2166__, new_new_n2167__,
    new_new_n2168__, new_new_n2169__, new_new_n2170__, new_new_n2171__,
    new_new_n2173__, new_new_n2174__, new_new_n2175__, new_new_n2176__,
    new_new_n2177__, new_new_n2178__, new_new_n2179__, new_new_n2180__,
    new_new_n2181__, new_new_n2182__, new_new_n2183__, new_new_n2184__,
    new_new_n2185__, new_new_n2186__, new_new_n2187__, new_new_n2188__,
    new_new_n2189__, new_new_n2190__, new_new_n2191__, new_new_n2192__,
    new_new_n2193__, new_new_n2194__, new_new_n2195__, new_new_n2196__,
    new_new_n2197__, new_new_n2198__, new_new_n2199__, new_new_n2200__,
    new_new_n2201__, new_new_n2202__, new_new_n2203__, new_new_n2204__,
    new_new_n2205__, new_new_n2206__, new_new_n2207__, new_new_n2208__,
    new_new_n2209__, new_new_n2210__, new_new_n2211__, new_new_n2212__,
    new_new_n2213__, new_new_n2214__, new_new_n2215__, new_new_n2216__,
    new_new_n2217__, new_new_n2218__, new_new_n2219__, new_new_n2220__,
    new_new_n2221__, new_new_n2222__, new_new_n2223__, new_new_n2224__,
    new_new_n2225__, new_new_n2226__, new_new_n2227__, new_new_n2228__,
    new_new_n2229__, new_new_n2230__, new_new_n2231__, new_new_n2232__,
    new_new_n2233__, new_new_n2234__, new_new_n2235__, new_new_n2236__,
    new_new_n2237__, new_new_n2238__, new_new_n2239__, new_new_n2240__,
    new_new_n2241__, new_new_n2242__, new_new_n2243__, new_new_n2244__,
    new_new_n2245__, new_new_n2246__, new_new_n2247__, new_new_n2248__,
    new_new_n2249__, new_new_n2250__, new_new_n2251__, new_new_n2252__,
    new_new_n2253__, new_new_n2254__, new_new_n2255__, new_new_n2256__,
    new_new_n2257__, new_new_n2258__, new_new_n2259__, new_new_n2260__,
    new_new_n2261__, new_new_n2262__, new_new_n2263__, new_new_n2264__,
    new_new_n2265__, new_new_n2266__, new_new_n2267__, new_new_n2268__,
    new_new_n2269__, new_new_n2270__, new_new_n2271__, new_new_n2272__,
    new_new_n2273__, new_new_n2274__, new_new_n2275__, new_new_n2276__,
    new_new_n2277__, new_new_n2278__, new_new_n2279__, new_new_n2280__,
    new_new_n2281__, new_new_n2282__, new_new_n2283__, new_new_n2284__,
    new_new_n2285__, new_new_n2286__, new_new_n2287__, new_new_n2288__,
    new_new_n2289__, new_new_n2290__, new_new_n2291__, new_new_n2292__,
    new_new_n2293__, new_new_n2294__, new_new_n2295__, new_new_n2296__,
    new_new_n2297__, new_new_n2298__, new_new_n2299__, new_new_n2300__,
    new_new_n2301__, new_new_n2302__, new_new_n2303__, new_new_n2304__,
    new_new_n2305__, new_new_n2306__, new_new_n2307__, new_new_n2308__,
    new_new_n2309__, new_new_n2310__, new_new_n2311__, new_new_n2312__,
    new_new_n2313__, new_new_n2314__, new_new_n2315__, new_new_n2316__,
    new_new_n2317__, new_new_n2318__, new_new_n2319__, new_new_n2320__,
    new_new_n2321__, new_new_n2322__, new_new_n2323__, new_new_n2324__,
    new_new_n2325__, new_new_n2326__, new_new_n2327__, new_new_n2328__,
    new_new_n2329__, new_new_n2330__, new_new_n2331__, new_new_n2332__,
    new_new_n2333__, new_new_n2334__, new_new_n2335__, new_new_n2336__,
    new_new_n2337__, new_new_n2338__, new_new_n2339__, new_new_n2340__,
    new_new_n2341__, new_new_n2342__, new_new_n2343__, new_new_n2344__,
    new_new_n2345__, new_new_n2346__, new_new_n2347__, new_new_n2348__,
    new_new_n2349__, new_new_n2350__, new_new_n2351__, new_new_n2352__,
    new_new_n2353__, new_new_n2354__, new_new_n2355__, new_new_n2356__,
    new_new_n2357__, new_new_n2358__, new_new_n2359__, new_new_n2360__,
    new_new_n2361__, new_new_n2362__, new_new_n2363__, new_new_n2364__,
    new_new_n2365__, new_new_n2366__, new_new_n2367__, new_new_n2368__,
    new_new_n2369__, new_new_n2370__, new_new_n2371__, new_new_n2372__,
    new_new_n2373__, new_new_n2374__, new_new_n2375__, new_new_n2376__,
    new_new_n2377__, new_new_n2378__, new_new_n2379__, new_new_n2380__,
    new_new_n2382__, new_new_n2383__, new_new_n2384__, new_new_n2385__,
    new_new_n2386__, new_new_n2387__, new_new_n2388__, new_new_n2389__,
    new_new_n2390__, new_new_n2391__, new_new_n2392__, new_new_n2393__,
    new_new_n2394__, new_new_n2395__, new_new_n2396__, new_new_n2397__,
    new_new_n2398__, new_new_n2399__, new_new_n2400__, new_new_n2401__,
    new_new_n2402__, new_new_n2403__, new_new_n2404__, new_new_n2405__,
    new_new_n2406__, new_new_n2407__, new_new_n2408__, new_new_n2409__,
    new_new_n2410__, new_new_n2411__, new_new_n2412__, new_new_n2413__,
    new_new_n2414__, new_new_n2415__, new_new_n2416__, new_new_n2417__,
    new_new_n2418__, new_new_n2419__, new_new_n2420__, new_new_n2421__,
    new_new_n2422__, new_new_n2423__, new_new_n2424__, new_new_n2425__,
    new_new_n2426__, new_new_n2427__, new_new_n2428__, new_new_n2429__,
    new_new_n2430__, new_new_n2431__, new_new_n2432__, new_new_n2433__,
    new_new_n2434__, new_new_n2435__, new_new_n2436__, new_new_n2437__,
    new_new_n2438__, new_new_n2439__, new_new_n2440__, new_new_n2441__,
    new_new_n2442__, new_new_n2443__, new_new_n2444__, new_new_n2445__,
    new_new_n2446__, new_new_n2447__, new_new_n2448__, new_new_n2449__,
    new_new_n2450__, new_new_n2451__, new_new_n2452__, new_new_n2453__,
    new_new_n2454__, new_new_n2455__, new_new_n2456__, new_new_n2457__,
    new_new_n2458__, new_new_n2459__, new_new_n2460__, new_new_n2461__,
    new_new_n2462__, new_new_n2463__, new_new_n2464__, new_new_n2465__,
    new_new_n2466__, new_new_n2467__, new_new_n2468__, new_new_n2469__,
    new_new_n2470__, new_new_n2471__, new_new_n2472__, new_new_n2473__,
    new_new_n2474__, new_new_n2475__, new_new_n2476__, new_new_n2477__,
    new_new_n2478__, new_new_n2479__, new_new_n2480__, new_new_n2481__,
    new_new_n2482__, new_new_n2483__, new_new_n2484__, new_new_n2485__,
    new_new_n2486__, new_new_n2487__, new_new_n2488__, new_new_n2489__,
    new_new_n2490__, new_new_n2491__, new_new_n2492__, new_new_n2493__,
    new_new_n2494__, new_new_n2495__, new_new_n2496__, new_new_n2497__,
    new_new_n2498__, new_new_n2499__, new_new_n2500__, new_new_n2501__,
    new_new_n2502__, new_new_n2503__, new_new_n2504__, new_new_n2505__,
    new_new_n2506__, new_new_n2507__, new_new_n2508__, new_new_n2509__,
    new_new_n2510__, new_new_n2511__, new_new_n2512__, new_new_n2513__,
    new_new_n2514__, new_new_n2515__, new_new_n2516__, new_new_n2517__,
    new_new_n2518__, new_new_n2519__, new_new_n2520__, new_new_n2521__,
    new_new_n2522__, new_new_n2523__, new_new_n2524__, new_new_n2525__,
    new_new_n2526__, new_new_n2527__, new_new_n2528__, new_new_n2529__,
    new_new_n2530__, new_new_n2531__, new_new_n2532__, new_new_n2533__,
    new_new_n2534__, new_new_n2535__, new_new_n2536__, new_new_n2537__,
    new_new_n2538__, new_new_n2539__, new_new_n2540__, new_new_n2541__,
    new_new_n2542__, new_new_n2543__, new_new_n2544__, new_new_n2545__,
    new_new_n2546__, new_new_n2547__, new_new_n2548__, new_new_n2549__,
    new_new_n2550__, new_new_n2551__, new_new_n2552__, new_new_n2553__,
    new_new_n2554__, new_new_n2555__, new_new_n2556__, new_new_n2557__,
    new_new_n2558__, new_new_n2559__, new_new_n2560__, new_new_n2561__,
    new_new_n2562__, new_new_n2563__, new_new_n2564__, new_new_n2565__,
    new_new_n2566__, new_new_n2567__, new_new_n2568__, new_new_n2569__,
    new_new_n2570__, new_new_n2571__, new_new_n2572__, new_new_n2573__,
    new_new_n2574__, new_new_n2575__, new_new_n2576__, new_new_n2577__,
    new_new_n2578__, new_new_n2579__, new_new_n2580__, new_new_n2581__,
    new_new_n2582__, new_new_n2583__, new_new_n2584__, new_new_n2585__,
    new_new_n2586__, new_new_n2587__, new_new_n2588__, new_new_n2589__,
    new_new_n2590__, new_new_n2591__, new_new_n2592__, new_new_n2593__,
    new_new_n2594__, new_new_n2595__, new_new_n2596__, new_new_n2597__,
    new_new_n2598__, new_new_n2599__, new_new_n2600__, new_new_n2601__,
    new_new_n2602__, new_new_n2603__, new_new_n2604__, new_new_n2605__,
    new_new_n2607__, new_new_n2608__, new_new_n2609__, new_new_n2610__,
    new_new_n2611__, new_new_n2612__, new_new_n2613__, new_new_n2614__,
    new_new_n2615__, new_new_n2616__, new_new_n2617__, new_new_n2618__,
    new_new_n2619__, new_new_n2620__, new_new_n2621__, new_new_n2622__,
    new_new_n2623__, new_new_n2624__, new_new_n2625__, new_new_n2626__,
    new_new_n2627__, new_new_n2628__, new_new_n2629__, new_new_n2630__,
    new_new_n2631__, new_new_n2632__, new_new_n2633__, new_new_n2634__,
    new_new_n2635__, new_new_n2636__, new_new_n2637__, new_new_n2638__,
    new_new_n2639__, new_new_n2640__, new_new_n2641__, new_new_n2642__,
    new_new_n2643__, new_new_n2644__, new_new_n2645__, new_new_n2646__,
    new_new_n2647__, new_new_n2648__, new_new_n2649__, new_new_n2650__,
    new_new_n2651__, new_new_n2652__, new_new_n2653__, new_new_n2654__,
    new_new_n2655__, new_new_n2656__, new_new_n2657__, new_new_n2658__,
    new_new_n2659__, new_new_n2660__, new_new_n2661__, new_new_n2662__,
    new_new_n2663__, new_new_n2664__, new_new_n2665__, new_new_n2666__,
    new_new_n2667__, new_new_n2668__, new_new_n2669__, new_new_n2670__,
    new_new_n2671__, new_new_n2672__, new_new_n2673__, new_new_n2674__,
    new_new_n2675__, new_new_n2676__, new_new_n2677__, new_new_n2678__,
    new_new_n2679__, new_new_n2680__, new_new_n2681__, new_new_n2682__,
    new_new_n2683__, new_new_n2684__, new_new_n2685__, new_new_n2686__,
    new_new_n2687__, new_new_n2688__, new_new_n2689__, new_new_n2690__,
    new_new_n2691__, new_new_n2692__, new_new_n2693__, new_new_n2694__,
    new_new_n2695__, new_new_n2696__, new_new_n2697__, new_new_n2698__,
    new_new_n2699__, new_new_n2700__, new_new_n2701__, new_new_n2702__,
    new_new_n2703__, new_new_n2704__, new_new_n2705__, new_new_n2706__,
    new_new_n2707__, new_new_n2708__, new_new_n2709__, new_new_n2710__,
    new_new_n2711__, new_new_n2712__, new_new_n2713__, new_new_n2714__,
    new_new_n2715__, new_new_n2716__, new_new_n2717__, new_new_n2718__,
    new_new_n2719__, new_new_n2720__, new_new_n2721__, new_new_n2722__,
    new_new_n2723__, new_new_n2724__, new_new_n2725__, new_new_n2726__,
    new_new_n2727__, new_new_n2728__, new_new_n2729__, new_new_n2730__,
    new_new_n2731__, new_new_n2732__, new_new_n2733__, new_new_n2734__,
    new_new_n2735__, new_new_n2736__, new_new_n2737__, new_new_n2738__,
    new_new_n2739__, new_new_n2740__, new_new_n2741__, new_new_n2742__,
    new_new_n2743__, new_new_n2744__, new_new_n2745__, new_new_n2746__,
    new_new_n2747__, new_new_n2748__, new_new_n2749__, new_new_n2750__,
    new_new_n2751__, new_new_n2752__, new_new_n2753__, new_new_n2754__,
    new_new_n2755__, new_new_n2756__, new_new_n2757__, new_new_n2758__,
    new_new_n2759__, new_new_n2760__, new_new_n2761__, new_new_n2762__,
    new_new_n2763__, new_new_n2764__, new_new_n2765__, new_new_n2766__,
    new_new_n2767__, new_new_n2768__, new_new_n2769__, new_new_n2770__,
    new_new_n2771__, new_new_n2772__, new_new_n2773__, new_new_n2774__,
    new_new_n2775__, new_new_n2776__, new_new_n2777__, new_new_n2778__,
    new_new_n2779__, new_new_n2780__, new_new_n2781__, new_new_n2782__,
    new_new_n2783__, new_new_n2784__, new_new_n2785__, new_new_n2786__,
    new_new_n2787__, new_new_n2788__, new_new_n2789__, new_new_n2790__,
    new_new_n2791__, new_new_n2792__, new_new_n2793__, new_new_n2794__,
    new_new_n2795__, new_new_n2796__, new_new_n2797__, new_new_n2798__,
    new_new_n2799__, new_new_n2800__, new_new_n2801__, new_new_n2802__,
    new_new_n2803__, new_new_n2804__, new_new_n2805__, new_new_n2806__,
    new_new_n2807__, new_new_n2808__, new_new_n2809__, new_new_n2810__,
    new_new_n2811__, new_new_n2812__, new_new_n2813__, new_new_n2814__,
    new_new_n2815__, new_new_n2816__, new_new_n2817__, new_new_n2818__,
    new_new_n2819__, new_new_n2820__, new_new_n2821__, new_new_n2822__,
    new_new_n2823__, new_new_n2824__, new_new_n2825__, new_new_n2826__,
    new_new_n2827__, new_new_n2828__, new_new_n2829__, new_new_n2830__,
    new_new_n2831__, new_new_n2832__, new_new_n2833__, new_new_n2834__,
    new_new_n2835__, new_new_n2836__, new_new_n2837__, new_new_n2838__,
    new_new_n2839__, new_new_n2841__, new_new_n2842__, new_new_n2843__,
    new_new_n2844__, new_new_n2845__, new_new_n2846__, new_new_n2847__,
    new_new_n2848__, new_new_n2849__, new_new_n2850__, new_new_n2851__,
    new_new_n2852__, new_new_n2853__, new_new_n2854__, new_new_n2855__,
    new_new_n2856__, new_new_n2857__, new_new_n2858__, new_new_n2859__,
    new_new_n2860__, new_new_n2861__, new_new_n2862__, new_new_n2863__,
    new_new_n2864__, new_new_n2865__, new_new_n2866__, new_new_n2867__,
    new_new_n2868__, new_new_n2869__, new_new_n2870__, new_new_n2871__,
    new_new_n2872__, new_new_n2873__, new_new_n2874__, new_new_n2875__,
    new_new_n2876__, new_new_n2877__, new_new_n2878__, new_new_n2879__,
    new_new_n2880__, new_new_n2881__, new_new_n2882__, new_new_n2883__,
    new_new_n2884__, new_new_n2885__, new_new_n2886__, new_new_n2887__,
    new_new_n2888__, new_new_n2889__, new_new_n2890__, new_new_n2891__,
    new_new_n2892__, new_new_n2893__, new_new_n2894__, new_new_n2895__,
    new_new_n2896__, new_new_n2897__, new_new_n2898__, new_new_n2899__,
    new_new_n2900__, new_new_n2901__, new_new_n2902__, new_new_n2903__,
    new_new_n2904__, new_new_n2905__, new_new_n2906__, new_new_n2907__,
    new_new_n2908__, new_new_n2909__, new_new_n2910__, new_new_n2911__,
    new_new_n2912__, new_new_n2913__, new_new_n2914__, new_new_n2915__,
    new_new_n2916__, new_new_n2917__, new_new_n2918__, new_new_n2919__,
    new_new_n2920__, new_new_n2921__, new_new_n2922__, new_new_n2923__,
    new_new_n2924__, new_new_n2925__, new_new_n2926__, new_new_n2927__,
    new_new_n2928__, new_new_n2929__, new_new_n2930__, new_new_n2931__,
    new_new_n2932__, new_new_n2933__, new_new_n2934__, new_new_n2935__,
    new_new_n2936__, new_new_n2937__, new_new_n2938__, new_new_n2939__,
    new_new_n2940__, new_new_n2941__, new_new_n2942__, new_new_n2943__,
    new_new_n2944__, new_new_n2945__, new_new_n2946__, new_new_n2947__,
    new_new_n2948__, new_new_n2949__, new_new_n2950__, new_new_n2951__,
    new_new_n2952__, new_new_n2953__, new_new_n2954__, new_new_n2955__,
    new_new_n2956__, new_new_n2957__, new_new_n2958__, new_new_n2959__,
    new_new_n2960__, new_new_n2961__, new_new_n2962__, new_new_n2963__,
    new_new_n2964__, new_new_n2965__, new_new_n2966__, new_new_n2967__,
    new_new_n2968__, new_new_n2969__, new_new_n2970__, new_new_n2971__,
    new_new_n2972__, new_new_n2973__, new_new_n2974__, new_new_n2975__,
    new_new_n2976__, new_new_n2977__, new_new_n2978__, new_new_n2979__,
    new_new_n2980__, new_new_n2981__, new_new_n2982__, new_new_n2983__,
    new_new_n2984__, new_new_n2985__, new_new_n2986__, new_new_n2987__,
    new_new_n2988__, new_new_n2989__, new_new_n2990__, new_new_n2991__,
    new_new_n2992__, new_new_n2993__, new_new_n2994__, new_new_n2995__,
    new_new_n2996__, new_new_n2997__, new_new_n2998__, new_new_n2999__,
    new_new_n3000__, new_new_n3001__, new_new_n3002__, new_new_n3003__,
    new_new_n3004__, new_new_n3005__, new_new_n3006__, new_new_n3007__,
    new_new_n3008__, new_new_n3009__, new_new_n3010__, new_new_n3011__,
    new_new_n3012__, new_new_n3013__, new_new_n3014__, new_new_n3015__,
    new_new_n3016__, new_new_n3017__, new_new_n3018__, new_new_n3019__,
    new_new_n3020__, new_new_n3021__, new_new_n3022__, new_new_n3023__,
    new_new_n3024__, new_new_n3025__, new_new_n3026__, new_new_n3027__,
    new_new_n3028__, new_new_n3029__, new_new_n3030__, new_new_n3031__,
    new_new_n3032__, new_new_n3033__, new_new_n3034__, new_new_n3035__,
    new_new_n3036__, new_new_n3037__, new_new_n3038__, new_new_n3039__,
    new_new_n3040__, new_new_n3041__, new_new_n3042__, new_new_n3043__,
    new_new_n3044__, new_new_n3045__, new_new_n3046__, new_new_n3047__,
    new_new_n3048__, new_new_n3049__, new_new_n3050__, new_new_n3051__,
    new_new_n3052__, new_new_n3053__, new_new_n3054__, new_new_n3055__,
    new_new_n3056__, new_new_n3057__, new_new_n3058__, new_new_n3059__,
    new_new_n3060__, new_new_n3061__, new_new_n3062__, new_new_n3063__,
    new_new_n3064__, new_new_n3065__, new_new_n3066__, new_new_n3067__,
    new_new_n3068__, new_new_n3069__, new_new_n3070__, new_new_n3071__,
    new_new_n3072__, new_new_n3073__, new_new_n3074__, new_new_n3075__,
    new_new_n3076__, new_new_n3077__, new_new_n3078__, new_new_n3080__,
    new_new_n3081__, new_new_n3082__, new_new_n3083__, new_new_n3084__,
    new_new_n3085__, new_new_n3086__, new_new_n3087__, new_new_n3088__,
    new_new_n3089__, new_new_n3090__, new_new_n3091__, new_new_n3092__,
    new_new_n3093__, new_new_n3094__, new_new_n3095__, new_new_n3096__,
    new_new_n3097__, new_new_n3098__, new_new_n3099__, new_new_n3100__,
    new_new_n3101__, new_new_n3102__, new_new_n3103__, new_new_n3104__,
    new_new_n3105__, new_new_n3106__, new_new_n3107__, new_new_n3108__,
    new_new_n3109__, new_new_n3110__, new_new_n3111__, new_new_n3112__,
    new_new_n3113__, new_new_n3114__, new_new_n3115__, new_new_n3116__,
    new_new_n3117__, new_new_n3118__, new_new_n3119__, new_new_n3120__,
    new_new_n3121__, new_new_n3122__, new_new_n3123__, new_new_n3124__,
    new_new_n3125__, new_new_n3126__, new_new_n3127__, new_new_n3128__,
    new_new_n3129__, new_new_n3130__, new_new_n3131__, new_new_n3132__,
    new_new_n3133__, new_new_n3134__, new_new_n3135__, new_new_n3136__,
    new_new_n3137__, new_new_n3138__, new_new_n3139__, new_new_n3140__,
    new_new_n3141__, new_new_n3142__, new_new_n3143__, new_new_n3144__,
    new_new_n3145__, new_new_n3146__, new_new_n3147__, new_new_n3148__,
    new_new_n3149__, new_new_n3150__, new_new_n3151__, new_new_n3152__,
    new_new_n3153__, new_new_n3154__, new_new_n3155__, new_new_n3156__,
    new_new_n3157__, new_new_n3158__, new_new_n3159__, new_new_n3160__,
    new_new_n3161__, new_new_n3162__, new_new_n3163__, new_new_n3164__,
    new_new_n3165__, new_new_n3166__, new_new_n3167__, new_new_n3168__,
    new_new_n3169__, new_new_n3170__, new_new_n3171__, new_new_n3172__,
    new_new_n3173__, new_new_n3174__, new_new_n3175__, new_new_n3176__,
    new_new_n3177__, new_new_n3178__, new_new_n3179__, new_new_n3180__,
    new_new_n3181__, new_new_n3182__, new_new_n3183__, new_new_n3184__,
    new_new_n3185__, new_new_n3186__, new_new_n3187__, new_new_n3188__,
    new_new_n3189__, new_new_n3190__, new_new_n3191__, new_new_n3192__,
    new_new_n3193__, new_new_n3194__, new_new_n3195__, new_new_n3196__,
    new_new_n3197__, new_new_n3198__, new_new_n3199__, new_new_n3200__,
    new_new_n3201__, new_new_n3202__, new_new_n3203__, new_new_n3204__,
    new_new_n3205__, new_new_n3206__, new_new_n3207__, new_new_n3208__,
    new_new_n3209__, new_new_n3210__, new_new_n3211__, new_new_n3212__,
    new_new_n3213__, new_new_n3214__, new_new_n3215__, new_new_n3216__,
    new_new_n3217__, new_new_n3218__, new_new_n3219__, new_new_n3220__,
    new_new_n3221__, new_new_n3222__, new_new_n3223__, new_new_n3224__,
    new_new_n3225__, new_new_n3226__, new_new_n3227__, new_new_n3228__,
    new_new_n3229__, new_new_n3230__, new_new_n3231__, new_new_n3232__,
    new_new_n3233__, new_new_n3234__, new_new_n3235__, new_new_n3236__,
    new_new_n3237__, new_new_n3238__, new_new_n3239__, new_new_n3240__,
    new_new_n3241__, new_new_n3242__, new_new_n3243__, new_new_n3244__,
    new_new_n3245__, new_new_n3246__, new_new_n3247__, new_new_n3248__,
    new_new_n3249__, new_new_n3250__, new_new_n3251__, new_new_n3252__,
    new_new_n3253__, new_new_n3254__, new_new_n3255__, new_new_n3256__,
    new_new_n3257__, new_new_n3258__, new_new_n3259__, new_new_n3260__,
    new_new_n3261__, new_new_n3262__, new_new_n3263__, new_new_n3264__,
    new_new_n3265__, new_new_n3266__, new_new_n3267__, new_new_n3268__,
    new_new_n3269__, new_new_n3270__, new_new_n3271__, new_new_n3272__,
    new_new_n3273__, new_new_n3274__, new_new_n3275__, new_new_n3276__,
    new_new_n3277__, new_new_n3278__, new_new_n3279__, new_new_n3280__,
    new_new_n3281__, new_new_n3282__, new_new_n3283__, new_new_n3284__,
    new_new_n3285__, new_new_n3286__, new_new_n3287__, new_new_n3288__,
    new_new_n3289__, new_new_n3290__, new_new_n3291__, new_new_n3292__,
    new_new_n3293__, new_new_n3294__, new_new_n3295__, new_new_n3296__,
    new_new_n3297__, new_new_n3298__, new_new_n3299__, new_new_n3300__,
    new_new_n3301__, new_new_n3302__, new_new_n3303__, new_new_n3304__,
    new_new_n3305__, new_new_n3306__, new_new_n3307__, new_new_n3308__,
    new_new_n3309__, new_new_n3310__, new_new_n3311__, new_new_n3312__,
    new_new_n3313__, new_new_n3314__, new_new_n3315__, new_new_n3316__,
    new_new_n3317__, new_new_n3318__, new_new_n3319__, new_new_n3320__,
    new_new_n3321__, new_new_n3322__, new_new_n3323__, new_new_n3324__,
    new_new_n3325__, new_new_n3326__, new_new_n3327__, new_new_n3328__,
    new_new_n3329__, new_new_n3330__, new_new_n3331__, new_new_n3332__,
    new_new_n3333__, new_new_n3334__, new_new_n3335__, new_new_n3336__,
    new_new_n3337__, new_new_n3338__, new_new_n3339__, new_new_n3340__,
    new_new_n3342__, new_new_n3343__, new_new_n3344__, new_new_n3345__,
    new_new_n3346__, new_new_n3347__, new_new_n3348__, new_new_n3349__,
    new_new_n3350__, new_new_n3351__, new_new_n3352__, new_new_n3353__,
    new_new_n3354__, new_new_n3355__, new_new_n3356__, new_new_n3357__,
    new_new_n3358__, new_new_n3359__, new_new_n3360__, new_new_n3361__,
    new_new_n3362__, new_new_n3363__, new_new_n3364__, new_new_n3365__,
    new_new_n3366__, new_new_n3367__, new_new_n3368__, new_new_n3369__,
    new_new_n3370__, new_new_n3371__, new_new_n3372__, new_new_n3373__,
    new_new_n3374__, new_new_n3375__, new_new_n3376__, new_new_n3377__,
    new_new_n3378__, new_new_n3379__, new_new_n3380__, new_new_n3381__,
    new_new_n3382__, new_new_n3383__, new_new_n3384__, new_new_n3385__,
    new_new_n3386__, new_new_n3387__, new_new_n3388__, new_new_n3389__,
    new_new_n3390__, new_new_n3391__, new_new_n3392__, new_new_n3393__,
    new_new_n3394__, new_new_n3395__, new_new_n3396__, new_new_n3397__,
    new_new_n3398__, new_new_n3399__, new_new_n3400__, new_new_n3401__,
    new_new_n3402__, new_new_n3403__, new_new_n3404__, new_new_n3405__,
    new_new_n3406__, new_new_n3407__, new_new_n3408__, new_new_n3409__,
    new_new_n3410__, new_new_n3411__, new_new_n3412__, new_new_n3413__,
    new_new_n3414__, new_new_n3415__, new_new_n3416__, new_new_n3417__,
    new_new_n3418__, new_new_n3419__, new_new_n3420__, new_new_n3421__,
    new_new_n3422__, new_new_n3423__, new_new_n3424__, new_new_n3425__,
    new_new_n3426__, new_new_n3427__, new_new_n3428__, new_new_n3429__,
    new_new_n3430__, new_new_n3431__, new_new_n3432__, new_new_n3433__,
    new_new_n3434__, new_new_n3435__, new_new_n3436__, new_new_n3437__,
    new_new_n3438__, new_new_n3439__, new_new_n3440__, new_new_n3441__,
    new_new_n3442__, new_new_n3443__, new_new_n3444__, new_new_n3445__,
    new_new_n3446__, new_new_n3447__, new_new_n3448__, new_new_n3449__,
    new_new_n3450__, new_new_n3451__, new_new_n3452__, new_new_n3453__,
    new_new_n3454__, new_new_n3455__, new_new_n3456__, new_new_n3457__,
    new_new_n3458__, new_new_n3459__, new_new_n3460__, new_new_n3461__,
    new_new_n3462__, new_new_n3463__, new_new_n3464__, new_new_n3465__,
    new_new_n3466__, new_new_n3467__, new_new_n3468__, new_new_n3469__,
    new_new_n3470__, new_new_n3471__, new_new_n3472__, new_new_n3473__,
    new_new_n3474__, new_new_n3475__, new_new_n3476__, new_new_n3477__,
    new_new_n3478__, new_new_n3479__, new_new_n3480__, new_new_n3481__,
    new_new_n3482__, new_new_n3483__, new_new_n3484__, new_new_n3485__,
    new_new_n3486__, new_new_n3487__, new_new_n3488__, new_new_n3489__,
    new_new_n3490__, new_new_n3491__, new_new_n3492__, new_new_n3493__,
    new_new_n3494__, new_new_n3495__, new_new_n3496__, new_new_n3497__,
    new_new_n3498__, new_new_n3499__, new_new_n3500__, new_new_n3501__,
    new_new_n3502__, new_new_n3503__, new_new_n3504__, new_new_n3505__,
    new_new_n3506__, new_new_n3507__, new_new_n3508__, new_new_n3509__,
    new_new_n3510__, new_new_n3511__, new_new_n3512__, new_new_n3513__,
    new_new_n3514__, new_new_n3515__, new_new_n3516__, new_new_n3517__,
    new_new_n3518__, new_new_n3519__, new_new_n3520__, new_new_n3521__,
    new_new_n3522__, new_new_n3523__, new_new_n3524__, new_new_n3525__,
    new_new_n3526__, new_new_n3527__, new_new_n3528__, new_new_n3529__,
    new_new_n3530__, new_new_n3531__, new_new_n3532__, new_new_n3533__,
    new_new_n3534__, new_new_n3535__, new_new_n3536__, new_new_n3537__,
    new_new_n3538__, new_new_n3539__, new_new_n3540__, new_new_n3541__,
    new_new_n3542__, new_new_n3543__, new_new_n3544__, new_new_n3545__,
    new_new_n3546__, new_new_n3547__, new_new_n3548__, new_new_n3549__,
    new_new_n3550__, new_new_n3551__, new_new_n3552__, new_new_n3553__,
    new_new_n3554__, new_new_n3555__, new_new_n3556__, new_new_n3557__,
    new_new_n3558__, new_new_n3559__, new_new_n3560__, new_new_n3561__,
    new_new_n3562__, new_new_n3563__, new_new_n3564__, new_new_n3565__,
    new_new_n3566__, new_new_n3567__, new_new_n3568__, new_new_n3569__,
    new_new_n3570__, new_new_n3571__, new_new_n3572__, new_new_n3573__,
    new_new_n3574__, new_new_n3575__, new_new_n3576__, new_new_n3577__,
    new_new_n3578__, new_new_n3579__, new_new_n3580__, new_new_n3581__,
    new_new_n3582__, new_new_n3583__, new_new_n3584__, new_new_n3585__,
    new_new_n3586__, new_new_n3587__, new_new_n3588__, new_new_n3589__,
    new_new_n3590__, new_new_n3591__, new_new_n3592__, new_new_n3593__,
    new_new_n3594__, new_new_n3595__, new_new_n3596__, new_new_n3597__,
    new_new_n3598__, new_new_n3599__, new_new_n3600__, new_new_n3601__,
    new_new_n3602__, new_new_n3603__, new_new_n3605__, new_new_n3606__,
    new_new_n3607__, new_new_n3608__, new_new_n3609__, new_new_n3610__,
    new_new_n3611__, new_new_n3612__, new_new_n3613__, new_new_n3614__,
    new_new_n3615__, new_new_n3616__, new_new_n3617__, new_new_n3618__,
    new_new_n3619__, new_new_n3620__, new_new_n3621__, new_new_n3622__,
    new_new_n3623__, new_new_n3624__, new_new_n3625__, new_new_n3626__,
    new_new_n3627__, new_new_n3628__, new_new_n3629__, new_new_n3630__,
    new_new_n3631__, new_new_n3632__, new_new_n3633__, new_new_n3634__,
    new_new_n3635__, new_new_n3636__, new_new_n3637__, new_new_n3638__,
    new_new_n3639__, new_new_n3640__, new_new_n3641__, new_new_n3642__,
    new_new_n3643__, new_new_n3644__, new_new_n3645__, new_new_n3646__,
    new_new_n3647__, new_new_n3648__, new_new_n3649__, new_new_n3650__,
    new_new_n3651__, new_new_n3652__, new_new_n3653__, new_new_n3654__,
    new_new_n3655__, new_new_n3656__, new_new_n3657__, new_new_n3658__,
    new_new_n3659__, new_new_n3660__, new_new_n3661__, new_new_n3662__,
    new_new_n3663__, new_new_n3664__, new_new_n3665__, new_new_n3666__,
    new_new_n3667__, new_new_n3668__, new_new_n3669__, new_new_n3670__,
    new_new_n3671__, new_new_n3672__, new_new_n3673__, new_new_n3674__,
    new_new_n3675__, new_new_n3676__, new_new_n3677__, new_new_n3678__,
    new_new_n3679__, new_new_n3680__, new_new_n3681__, new_new_n3682__,
    new_new_n3683__, new_new_n3684__, new_new_n3685__, new_new_n3686__,
    new_new_n3687__, new_new_n3688__, new_new_n3689__, new_new_n3690__,
    new_new_n3691__, new_new_n3692__, new_new_n3693__, new_new_n3694__,
    new_new_n3695__, new_new_n3696__, new_new_n3697__, new_new_n3698__,
    new_new_n3699__, new_new_n3700__, new_new_n3701__, new_new_n3702__,
    new_new_n3703__, new_new_n3704__, new_new_n3705__, new_new_n3706__,
    new_new_n3707__, new_new_n3708__, new_new_n3709__, new_new_n3710__,
    new_new_n3711__, new_new_n3712__, new_new_n3713__, new_new_n3714__,
    new_new_n3715__, new_new_n3716__, new_new_n3717__, new_new_n3718__,
    new_new_n3719__, new_new_n3720__, new_new_n3721__, new_new_n3722__,
    new_new_n3723__, new_new_n3724__, new_new_n3725__, new_new_n3726__,
    new_new_n3727__, new_new_n3728__, new_new_n3729__, new_new_n3730__,
    new_new_n3731__, new_new_n3732__, new_new_n3733__, new_new_n3734__,
    new_new_n3735__, new_new_n3736__, new_new_n3737__, new_new_n3738__,
    new_new_n3739__, new_new_n3740__, new_new_n3741__, new_new_n3742__,
    new_new_n3743__, new_new_n3744__, new_new_n3745__, new_new_n3746__,
    new_new_n3747__, new_new_n3748__, new_new_n3749__, new_new_n3750__,
    new_new_n3751__, new_new_n3752__, new_new_n3753__, new_new_n3754__,
    new_new_n3755__, new_new_n3756__, new_new_n3757__, new_new_n3758__,
    new_new_n3759__, new_new_n3760__, new_new_n3761__, new_new_n3762__,
    new_new_n3763__, new_new_n3764__, new_new_n3765__, new_new_n3766__,
    new_new_n3767__, new_new_n3768__, new_new_n3769__, new_new_n3770__,
    new_new_n3771__, new_new_n3772__, new_new_n3773__, new_new_n3774__,
    new_new_n3775__, new_new_n3776__, new_new_n3777__, new_new_n3778__,
    new_new_n3779__, new_new_n3780__, new_new_n3781__, new_new_n3782__,
    new_new_n3783__, new_new_n3784__, new_new_n3785__, new_new_n3786__,
    new_new_n3787__, new_new_n3788__, new_new_n3789__, new_new_n3790__,
    new_new_n3791__, new_new_n3792__, new_new_n3793__, new_new_n3794__,
    new_new_n3795__, new_new_n3796__, new_new_n3797__, new_new_n3798__,
    new_new_n3799__, new_new_n3800__, new_new_n3801__, new_new_n3802__,
    new_new_n3803__, new_new_n3804__, new_new_n3805__, new_new_n3806__,
    new_new_n3807__, new_new_n3808__, new_new_n3809__, new_new_n3810__,
    new_new_n3811__, new_new_n3812__, new_new_n3813__, new_new_n3814__,
    new_new_n3815__, new_new_n3816__, new_new_n3817__, new_new_n3818__,
    new_new_n3819__, new_new_n3820__, new_new_n3821__, new_new_n3822__,
    new_new_n3823__, new_new_n3824__, new_new_n3825__, new_new_n3826__,
    new_new_n3827__, new_new_n3828__, new_new_n3829__, new_new_n3830__,
    new_new_n3831__, new_new_n3832__, new_new_n3833__, new_new_n3834__,
    new_new_n3835__, new_new_n3836__, new_new_n3837__, new_new_n3838__,
    new_new_n3839__, new_new_n3840__, new_new_n3841__, new_new_n3842__,
    new_new_n3843__, new_new_n3844__, new_new_n3845__, new_new_n3846__,
    new_new_n3847__, new_new_n3848__, new_new_n3849__, new_new_n3850__,
    new_new_n3851__, new_new_n3852__, new_new_n3853__, new_new_n3854__,
    new_new_n3855__, new_new_n3856__, new_new_n3857__, new_new_n3858__,
    new_new_n3859__, new_new_n3860__, new_new_n3861__, new_new_n3862__,
    new_new_n3863__, new_new_n3864__, new_new_n3865__, new_new_n3866__,
    new_new_n3867__, new_new_n3868__, new_new_n3869__, new_new_n3870__,
    new_new_n3871__, new_new_n3872__, new_new_n3873__, new_new_n3874__,
    new_new_n3875__, new_new_n3876__, new_new_n3877__, new_new_n3878__,
    new_new_n3879__, new_new_n3880__, new_new_n3881__, new_new_n3882__,
    new_new_n3884__, new_new_n3885__, new_new_n3886__, new_new_n3887__,
    new_new_n3888__, new_new_n3889__, new_new_n3890__, new_new_n3891__,
    new_new_n3892__, new_new_n3893__, new_new_n3894__, new_new_n3895__,
    new_new_n3896__, new_new_n3897__, new_new_n3898__, new_new_n3899__,
    new_new_n3900__, new_new_n3901__, new_new_n3902__, new_new_n3903__,
    new_new_n3904__, new_new_n3905__, new_new_n3906__, new_new_n3907__,
    new_new_n3908__, new_new_n3909__, new_new_n3910__, new_new_n3911__,
    new_new_n3912__, new_new_n3913__, new_new_n3914__, new_new_n3915__,
    new_new_n3916__, new_new_n3917__, new_new_n3918__, new_new_n3919__,
    new_new_n3920__, new_new_n3921__, new_new_n3922__, new_new_n3923__,
    new_new_n3924__, new_new_n3925__, new_new_n3926__, new_new_n3927__,
    new_new_n3928__, new_new_n3929__, new_new_n3930__, new_new_n3931__,
    new_new_n3932__, new_new_n3933__, new_new_n3934__, new_new_n3935__,
    new_new_n3936__, new_new_n3937__, new_new_n3938__, new_new_n3939__,
    new_new_n3940__, new_new_n3941__, new_new_n3942__, new_new_n3943__,
    new_new_n3944__, new_new_n3945__, new_new_n3946__, new_new_n3947__,
    new_new_n3948__, new_new_n3949__, new_new_n3950__, new_new_n3951__,
    new_new_n3952__, new_new_n3953__, new_new_n3954__, new_new_n3955__,
    new_new_n3956__, new_new_n3957__, new_new_n3958__, new_new_n3959__,
    new_new_n3960__, new_new_n3961__, new_new_n3962__, new_new_n3963__,
    new_new_n3964__, new_new_n3965__, new_new_n3966__, new_new_n3967__,
    new_new_n3968__, new_new_n3969__, new_new_n3970__, new_new_n3971__,
    new_new_n3972__, new_new_n3973__, new_new_n3974__, new_new_n3975__,
    new_new_n3976__, new_new_n3977__, new_new_n3978__, new_new_n3979__,
    new_new_n3980__, new_new_n3981__, new_new_n3982__, new_new_n3983__,
    new_new_n3984__, new_new_n3985__, new_new_n3986__, new_new_n3987__,
    new_new_n3988__, new_new_n3989__, new_new_n3990__, new_new_n3991__,
    new_new_n3992__, new_new_n3993__, new_new_n3994__, new_new_n3995__,
    new_new_n3996__, new_new_n3997__, new_new_n3998__, new_new_n3999__,
    new_new_n4000__, new_new_n4001__, new_new_n4002__, new_new_n4003__,
    new_new_n4004__, new_new_n4005__, new_new_n4006__, new_new_n4007__,
    new_new_n4008__, new_new_n4009__, new_new_n4010__, new_new_n4011__,
    new_new_n4012__, new_new_n4013__, new_new_n4014__, new_new_n4015__,
    new_new_n4016__, new_new_n4017__, new_new_n4018__, new_new_n4019__,
    new_new_n4020__, new_new_n4021__, new_new_n4022__, new_new_n4023__,
    new_new_n4024__, new_new_n4025__, new_new_n4026__, new_new_n4027__,
    new_new_n4028__, new_new_n4029__, new_new_n4030__, new_new_n4031__,
    new_new_n4032__, new_new_n4033__, new_new_n4034__, new_new_n4035__,
    new_new_n4036__, new_new_n4037__, new_new_n4038__, new_new_n4039__,
    new_new_n4040__, new_new_n4041__, new_new_n4042__, new_new_n4043__,
    new_new_n4044__, new_new_n4045__, new_new_n4046__, new_new_n4047__,
    new_new_n4048__, new_new_n4049__, new_new_n4050__, new_new_n4051__,
    new_new_n4052__, new_new_n4053__, new_new_n4054__, new_new_n4055__,
    new_new_n4056__, new_new_n4057__, new_new_n4058__, new_new_n4059__,
    new_new_n4060__, new_new_n4061__, new_new_n4062__, new_new_n4063__,
    new_new_n4064__, new_new_n4065__, new_new_n4066__, new_new_n4067__,
    new_new_n4068__, new_new_n4069__, new_new_n4070__, new_new_n4071__,
    new_new_n4072__, new_new_n4073__, new_new_n4074__, new_new_n4075__,
    new_new_n4076__, new_new_n4077__, new_new_n4078__, new_new_n4079__,
    new_new_n4080__, new_new_n4081__, new_new_n4082__, new_new_n4083__,
    new_new_n4084__, new_new_n4085__, new_new_n4086__, new_new_n4087__,
    new_new_n4088__, new_new_n4089__, new_new_n4090__, new_new_n4091__,
    new_new_n4092__, new_new_n4093__, new_new_n4094__, new_new_n4095__,
    new_new_n4096__, new_new_n4097__, new_new_n4098__, new_new_n4099__,
    new_new_n4100__, new_new_n4101__, new_new_n4102__, new_new_n4103__,
    new_new_n4104__, new_new_n4105__, new_new_n4106__, new_new_n4107__,
    new_new_n4108__, new_new_n4109__, new_new_n4110__, new_new_n4111__,
    new_new_n4112__, new_new_n4113__, new_new_n4114__, new_new_n4115__,
    new_new_n4116__, new_new_n4117__, new_new_n4118__, new_new_n4119__,
    new_new_n4120__, new_new_n4121__, new_new_n4122__, new_new_n4123__,
    new_new_n4124__, new_new_n4125__, new_new_n4126__, new_new_n4127__,
    new_new_n4128__, new_new_n4129__, new_new_n4130__, new_new_n4131__,
    new_new_n4132__, new_new_n4133__, new_new_n4134__, new_new_n4135__,
    new_new_n4136__, new_new_n4137__, new_new_n4138__, new_new_n4139__,
    new_new_n4140__, new_new_n4141__, new_new_n4142__, new_new_n4143__,
    new_new_n4144__, new_new_n4145__, new_new_n4146__, new_new_n4147__,
    new_new_n4148__, new_new_n4149__, new_new_n4150__, new_new_n4151__,
    new_new_n4152__, new_new_n4153__, new_new_n4154__, new_new_n4155__,
    new_new_n4156__, new_new_n4157__, new_new_n4158__, new_new_n4159__,
    new_new_n4160__, new_new_n4161__, new_new_n4162__, new_new_n4163__,
    new_new_n4164__, new_new_n4165__, new_new_n4166__, new_new_n4167__,
    new_new_n4168__, new_new_n4169__, new_new_n4170__, new_new_n4171__,
    new_new_n4172__, new_new_n4173__, new_new_n4175__, new_new_n4176__,
    new_new_n4177__, new_new_n4178__, new_new_n4179__, new_new_n4180__,
    new_new_n4181__, new_new_n4182__, new_new_n4183__, new_new_n4184__,
    new_new_n4185__, new_new_n4186__, new_new_n4187__, new_new_n4188__,
    new_new_n4189__, new_new_n4190__, new_new_n4191__, new_new_n4192__,
    new_new_n4193__, new_new_n4194__, new_new_n4195__, new_new_n4196__,
    new_new_n4197__, new_new_n4198__, new_new_n4199__, new_new_n4200__,
    new_new_n4201__, new_new_n4202__, new_new_n4203__, new_new_n4204__,
    new_new_n4205__, new_new_n4206__, new_new_n4207__, new_new_n4208__,
    new_new_n4209__, new_new_n4210__, new_new_n4211__, new_new_n4212__,
    new_new_n4213__, new_new_n4214__, new_new_n4215__, new_new_n4216__,
    new_new_n4217__, new_new_n4218__, new_new_n4219__, new_new_n4220__,
    new_new_n4221__, new_new_n4222__, new_new_n4223__, new_new_n4224__,
    new_new_n4225__, new_new_n4226__, new_new_n4227__, new_new_n4228__,
    new_new_n4229__, new_new_n4230__, new_new_n4231__, new_new_n4232__,
    new_new_n4233__, new_new_n4234__, new_new_n4235__, new_new_n4236__,
    new_new_n4237__, new_new_n4238__, new_new_n4239__, new_new_n4240__,
    new_new_n4241__, new_new_n4242__, new_new_n4243__, new_new_n4244__,
    new_new_n4245__, new_new_n4246__, new_new_n4247__, new_new_n4248__,
    new_new_n4249__, new_new_n4250__, new_new_n4251__, new_new_n4252__,
    new_new_n4253__, new_new_n4254__, new_new_n4255__, new_new_n4256__,
    new_new_n4257__, new_new_n4258__, new_new_n4259__, new_new_n4260__,
    new_new_n4261__, new_new_n4262__, new_new_n4263__, new_new_n4264__,
    new_new_n4265__, new_new_n4266__, new_new_n4267__, new_new_n4268__,
    new_new_n4269__, new_new_n4270__, new_new_n4271__, new_new_n4272__,
    new_new_n4273__, new_new_n4274__, new_new_n4275__, new_new_n4276__,
    new_new_n4277__, new_new_n4278__, new_new_n4279__, new_new_n4280__,
    new_new_n4281__, new_new_n4282__, new_new_n4283__, new_new_n4284__,
    new_new_n4285__, new_new_n4286__, new_new_n4287__, new_new_n4288__,
    new_new_n4289__, new_new_n4290__, new_new_n4291__, new_new_n4292__,
    new_new_n4293__, new_new_n4294__, new_new_n4295__, new_new_n4296__,
    new_new_n4297__, new_new_n4298__, new_new_n4299__, new_new_n4300__,
    new_new_n4301__, new_new_n4302__, new_new_n4303__, new_new_n4304__,
    new_new_n4305__, new_new_n4306__, new_new_n4307__, new_new_n4308__,
    new_new_n4309__, new_new_n4310__, new_new_n4311__, new_new_n4312__,
    new_new_n4313__, new_new_n4314__, new_new_n4315__, new_new_n4316__,
    new_new_n4317__, new_new_n4318__, new_new_n4319__, new_new_n4320__,
    new_new_n4321__, new_new_n4322__, new_new_n4323__, new_new_n4324__,
    new_new_n4325__, new_new_n4326__, new_new_n4327__, new_new_n4328__,
    new_new_n4329__, new_new_n4330__, new_new_n4331__, new_new_n4332__,
    new_new_n4333__, new_new_n4334__, new_new_n4335__, new_new_n4336__,
    new_new_n4337__, new_new_n4338__, new_new_n4339__, new_new_n4340__,
    new_new_n4341__, new_new_n4342__, new_new_n4343__, new_new_n4344__,
    new_new_n4345__, new_new_n4346__, new_new_n4347__, new_new_n4348__,
    new_new_n4349__, new_new_n4350__, new_new_n4351__, new_new_n4352__,
    new_new_n4353__, new_new_n4354__, new_new_n4355__, new_new_n4356__,
    new_new_n4357__, new_new_n4358__, new_new_n4359__, new_new_n4360__,
    new_new_n4361__, new_new_n4362__, new_new_n4363__, new_new_n4364__,
    new_new_n4365__, new_new_n4366__, new_new_n4367__, new_new_n4368__,
    new_new_n4369__, new_new_n4370__, new_new_n4371__, new_new_n4372__,
    new_new_n4373__, new_new_n4374__, new_new_n4375__, new_new_n4376__,
    new_new_n4377__, new_new_n4378__, new_new_n4379__, new_new_n4380__,
    new_new_n4381__, new_new_n4382__, new_new_n4383__, new_new_n4384__,
    new_new_n4385__, new_new_n4386__, new_new_n4387__, new_new_n4388__,
    new_new_n4389__, new_new_n4390__, new_new_n4391__, new_new_n4392__,
    new_new_n4393__, new_new_n4394__, new_new_n4395__, new_new_n4396__,
    new_new_n4397__, new_new_n4398__, new_new_n4399__, new_new_n4400__,
    new_new_n4401__, new_new_n4402__, new_new_n4403__, new_new_n4404__,
    new_new_n4405__, new_new_n4406__, new_new_n4407__, new_new_n4408__,
    new_new_n4409__, new_new_n4410__, new_new_n4411__, new_new_n4412__,
    new_new_n4413__, new_new_n4414__, new_new_n4415__, new_new_n4416__,
    new_new_n4417__, new_new_n4418__, new_new_n4419__, new_new_n4420__,
    new_new_n4421__, new_new_n4422__, new_new_n4423__, new_new_n4424__,
    new_new_n4425__, new_new_n4426__, new_new_n4427__, new_new_n4428__,
    new_new_n4429__, new_new_n4430__, new_new_n4431__, new_new_n4432__,
    new_new_n4433__, new_new_n4434__, new_new_n4435__, new_new_n4436__,
    new_new_n4437__, new_new_n4438__, new_new_n4439__, new_new_n4440__,
    new_new_n4441__, new_new_n4442__, new_new_n4443__, new_new_n4444__,
    new_new_n4445__, new_new_n4446__, new_new_n4447__, new_new_n4448__,
    new_new_n4449__, new_new_n4450__, new_new_n4451__, new_new_n4452__,
    new_new_n4453__, new_new_n4454__, new_new_n4455__, new_new_n4456__,
    new_new_n4457__, new_new_n4458__, new_new_n4459__, new_new_n4460__,
    new_new_n4461__, new_new_n4462__, new_new_n4463__, new_new_n4464__,
    new_new_n4465__, new_new_n4466__, new_new_n4467__, new_new_n4468__,
    new_new_n4469__, new_new_n4470__, new_new_n4471__, new_new_n4473__,
    new_new_n4474__, new_new_n4475__, new_new_n4476__, new_new_n4477__,
    new_new_n4478__, new_new_n4479__, new_new_n4480__, new_new_n4481__,
    new_new_n4482__, new_new_n4483__, new_new_n4484__, new_new_n4485__,
    new_new_n4486__, new_new_n4487__, new_new_n4488__, new_new_n4489__,
    new_new_n4490__, new_new_n4491__, new_new_n4492__, new_new_n4493__,
    new_new_n4494__, new_new_n4495__, new_new_n4496__, new_new_n4497__,
    new_new_n4498__, new_new_n4499__, new_new_n4500__, new_new_n4501__,
    new_new_n4502__, new_new_n4503__, new_new_n4504__, new_new_n4505__,
    new_new_n4506__, new_new_n4507__, new_new_n4508__, new_new_n4509__,
    new_new_n4510__, new_new_n4511__, new_new_n4512__, new_new_n4513__,
    new_new_n4514__, new_new_n4515__, new_new_n4516__, new_new_n4517__,
    new_new_n4518__, new_new_n4519__, new_new_n4520__, new_new_n4521__,
    new_new_n4522__, new_new_n4523__, new_new_n4524__, new_new_n4525__,
    new_new_n4526__, new_new_n4527__, new_new_n4528__, new_new_n4529__,
    new_new_n4530__, new_new_n4531__, new_new_n4532__, new_new_n4533__,
    new_new_n4534__, new_new_n4535__, new_new_n4536__, new_new_n4537__,
    new_new_n4538__, new_new_n4539__, new_new_n4540__, new_new_n4541__,
    new_new_n4542__, new_new_n4543__, new_new_n4544__, new_new_n4545__,
    new_new_n4546__, new_new_n4547__, new_new_n4548__, new_new_n4549__,
    new_new_n4550__, new_new_n4551__, new_new_n4552__, new_new_n4553__,
    new_new_n4554__, new_new_n4555__, new_new_n4556__, new_new_n4557__,
    new_new_n4558__, new_new_n4559__, new_new_n4560__, new_new_n4561__,
    new_new_n4562__, new_new_n4563__, new_new_n4564__, new_new_n4565__,
    new_new_n4566__, new_new_n4567__, new_new_n4568__, new_new_n4569__,
    new_new_n4570__, new_new_n4571__, new_new_n4572__, new_new_n4573__,
    new_new_n4574__, new_new_n4575__, new_new_n4576__, new_new_n4577__,
    new_new_n4578__, new_new_n4579__, new_new_n4580__, new_new_n4581__,
    new_new_n4582__, new_new_n4583__, new_new_n4584__, new_new_n4585__,
    new_new_n4586__, new_new_n4587__, new_new_n4588__, new_new_n4589__,
    new_new_n4590__, new_new_n4591__, new_new_n4592__, new_new_n4593__,
    new_new_n4594__, new_new_n4595__, new_new_n4596__, new_new_n4597__,
    new_new_n4598__, new_new_n4599__, new_new_n4600__, new_new_n4601__,
    new_new_n4602__, new_new_n4603__, new_new_n4604__, new_new_n4605__,
    new_new_n4606__, new_new_n4607__, new_new_n4608__, new_new_n4609__,
    new_new_n4610__, new_new_n4611__, new_new_n4612__, new_new_n4613__,
    new_new_n4614__, new_new_n4615__, new_new_n4616__, new_new_n4617__,
    new_new_n4618__, new_new_n4619__, new_new_n4620__, new_new_n4621__,
    new_new_n4622__, new_new_n4623__, new_new_n4624__, new_new_n4625__,
    new_new_n4626__, new_new_n4627__, new_new_n4628__, new_new_n4629__,
    new_new_n4630__, new_new_n4631__, new_new_n4632__, new_new_n4633__,
    new_new_n4634__, new_new_n4635__, new_new_n4636__, new_new_n4637__,
    new_new_n4638__, new_new_n4639__, new_new_n4640__, new_new_n4641__,
    new_new_n4642__, new_new_n4643__, new_new_n4644__, new_new_n4645__,
    new_new_n4646__, new_new_n4647__, new_new_n4648__, new_new_n4649__,
    new_new_n4650__, new_new_n4651__, new_new_n4652__, new_new_n4653__,
    new_new_n4654__, new_new_n4655__, new_new_n4656__, new_new_n4657__,
    new_new_n4658__, new_new_n4659__, new_new_n4660__, new_new_n4661__,
    new_new_n4662__, new_new_n4663__, new_new_n4664__, new_new_n4665__,
    new_new_n4666__, new_new_n4667__, new_new_n4668__, new_new_n4669__,
    new_new_n4670__, new_new_n4671__, new_new_n4672__, new_new_n4673__,
    new_new_n4674__, new_new_n4675__, new_new_n4676__, new_new_n4677__,
    new_new_n4678__, new_new_n4679__, new_new_n4680__, new_new_n4681__,
    new_new_n4682__, new_new_n4683__, new_new_n4684__, new_new_n4685__,
    new_new_n4686__, new_new_n4687__, new_new_n4688__, new_new_n4689__,
    new_new_n4690__, new_new_n4691__, new_new_n4692__, new_new_n4693__,
    new_new_n4694__, new_new_n4695__, new_new_n4696__, new_new_n4697__,
    new_new_n4698__, new_new_n4699__, new_new_n4700__, new_new_n4701__,
    new_new_n4702__, new_new_n4703__, new_new_n4704__, new_new_n4705__,
    new_new_n4706__, new_new_n4707__, new_new_n4708__, new_new_n4709__,
    new_new_n4710__, new_new_n4711__, new_new_n4712__, new_new_n4713__,
    new_new_n4714__, new_new_n4715__, new_new_n4716__, new_new_n4717__,
    new_new_n4718__, new_new_n4719__, new_new_n4720__, new_new_n4721__,
    new_new_n4722__, new_new_n4723__, new_new_n4724__, new_new_n4725__,
    new_new_n4726__, new_new_n4727__, new_new_n4728__, new_new_n4729__,
    new_new_n4730__, new_new_n4731__, new_new_n4732__, new_new_n4733__,
    new_new_n4734__, new_new_n4735__, new_new_n4736__, new_new_n4737__,
    new_new_n4738__, new_new_n4739__, new_new_n4740__, new_new_n4741__,
    new_new_n4742__, new_new_n4743__, new_new_n4744__, new_new_n4745__,
    new_new_n4746__, new_new_n4747__, new_new_n4748__, new_new_n4749__,
    new_new_n4750__, new_new_n4751__, new_new_n4752__, new_new_n4753__,
    new_new_n4754__, new_new_n4755__, new_new_n4756__, new_new_n4757__,
    new_new_n4758__, new_new_n4759__, new_new_n4760__, new_new_n4761__,
    new_new_n4762__, new_new_n4763__, new_new_n4764__, new_new_n4765__,
    new_new_n4766__, new_new_n4767__, new_new_n4768__, new_new_n4769__,
    new_new_n4770__, new_new_n4771__, new_new_n4772__, new_new_n4773__,
    new_new_n4775__, new_new_n4776__, new_new_n4777__, new_new_n4778__,
    new_new_n4779__, new_new_n4780__, new_new_n4781__, new_new_n4782__,
    new_new_n4783__, new_new_n4784__, new_new_n4785__, new_new_n4786__,
    new_new_n4787__, new_new_n4788__, new_new_n4789__, new_new_n4790__,
    new_new_n4791__, new_new_n4792__, new_new_n4793__, new_new_n4794__,
    new_new_n4795__, new_new_n4796__, new_new_n4797__, new_new_n4798__,
    new_new_n4799__, new_new_n4800__, new_new_n4801__, new_new_n4802__,
    new_new_n4803__, new_new_n4804__, new_new_n4805__, new_new_n4806__,
    new_new_n4807__, new_new_n4808__, new_new_n4809__, new_new_n4810__,
    new_new_n4811__, new_new_n4812__, new_new_n4813__, new_new_n4814__,
    new_new_n4815__, new_new_n4816__, new_new_n4817__, new_new_n4818__,
    new_new_n4819__, new_new_n4820__, new_new_n4821__, new_new_n4822__,
    new_new_n4823__, new_new_n4824__, new_new_n4825__, new_new_n4826__,
    new_new_n4827__, new_new_n4828__, new_new_n4829__, new_new_n4830__,
    new_new_n4831__, new_new_n4832__, new_new_n4833__, new_new_n4834__,
    new_new_n4835__, new_new_n4836__, new_new_n4837__, new_new_n4838__,
    new_new_n4839__, new_new_n4840__, new_new_n4841__, new_new_n4842__,
    new_new_n4843__, new_new_n4844__, new_new_n4845__, new_new_n4846__,
    new_new_n4847__, new_new_n4848__, new_new_n4849__, new_new_n4850__,
    new_new_n4851__, new_new_n4852__, new_new_n4853__, new_new_n4854__,
    new_new_n4855__, new_new_n4856__, new_new_n4857__, new_new_n4858__,
    new_new_n4859__, new_new_n4860__, new_new_n4861__, new_new_n4862__,
    new_new_n4863__, new_new_n4864__, new_new_n4865__, new_new_n4866__,
    new_new_n4867__, new_new_n4868__, new_new_n4869__, new_new_n4870__,
    new_new_n4871__, new_new_n4872__, new_new_n4873__, new_new_n4874__,
    new_new_n4875__, new_new_n4876__, new_new_n4877__, new_new_n4878__,
    new_new_n4879__, new_new_n4880__, new_new_n4881__, new_new_n4882__,
    new_new_n4883__, new_new_n4884__, new_new_n4885__, new_new_n4886__,
    new_new_n4887__, new_new_n4888__, new_new_n4889__, new_new_n4890__,
    new_new_n4891__, new_new_n4892__, new_new_n4893__, new_new_n4894__,
    new_new_n4895__, new_new_n4896__, new_new_n4897__, new_new_n4898__,
    new_new_n4899__, new_new_n4900__, new_new_n4901__, new_new_n4902__,
    new_new_n4903__, new_new_n4904__, new_new_n4905__, new_new_n4906__,
    new_new_n4907__, new_new_n4908__, new_new_n4909__, new_new_n4910__,
    new_new_n4911__, new_new_n4912__, new_new_n4913__, new_new_n4914__,
    new_new_n4915__, new_new_n4916__, new_new_n4917__, new_new_n4918__,
    new_new_n4919__, new_new_n4920__, new_new_n4921__, new_new_n4922__,
    new_new_n4923__, new_new_n4924__, new_new_n4925__, new_new_n4926__,
    new_new_n4927__, new_new_n4928__, new_new_n4929__, new_new_n4930__,
    new_new_n4931__, new_new_n4932__, new_new_n4933__, new_new_n4934__,
    new_new_n4935__, new_new_n4936__, new_new_n4937__, new_new_n4938__,
    new_new_n4939__, new_new_n4940__, new_new_n4941__, new_new_n4942__,
    new_new_n4943__, new_new_n4944__, new_new_n4945__, new_new_n4946__,
    new_new_n4947__, new_new_n4948__, new_new_n4949__, new_new_n4950__,
    new_new_n4951__, new_new_n4952__, new_new_n4953__, new_new_n4954__,
    new_new_n4955__, new_new_n4956__, new_new_n4957__, new_new_n4958__,
    new_new_n4959__, new_new_n4960__, new_new_n4961__, new_new_n4962__,
    new_new_n4963__, new_new_n4964__, new_new_n4965__, new_new_n4966__,
    new_new_n4967__, new_new_n4968__, new_new_n4969__, new_new_n4970__,
    new_new_n4971__, new_new_n4972__, new_new_n4973__, new_new_n4974__,
    new_new_n4975__, new_new_n4976__, new_new_n4977__, new_new_n4978__,
    new_new_n4979__, new_new_n4980__, new_new_n4981__, new_new_n4982__,
    new_new_n4983__, new_new_n4984__, new_new_n4985__, new_new_n4986__,
    new_new_n4987__, new_new_n4988__, new_new_n4989__, new_new_n4990__,
    new_new_n4991__, new_new_n4992__, new_new_n4993__, new_new_n4994__,
    new_new_n4995__, new_new_n4996__, new_new_n4997__, new_new_n4998__,
    new_new_n4999__, new_new_n5000__, new_new_n5001__, new_new_n5002__,
    new_new_n5003__, new_new_n5004__, new_new_n5005__, new_new_n5006__,
    new_new_n5007__, new_new_n5008__, new_new_n5009__, new_new_n5010__,
    new_new_n5011__, new_new_n5012__, new_new_n5013__, new_new_n5014__,
    new_new_n5015__, new_new_n5016__, new_new_n5017__, new_new_n5018__,
    new_new_n5019__, new_new_n5020__, new_new_n5021__, new_new_n5022__,
    new_new_n5023__, new_new_n5024__, new_new_n5025__, new_new_n5026__,
    new_new_n5027__, new_new_n5028__, new_new_n5029__, new_new_n5030__,
    new_new_n5031__, new_new_n5032__, new_new_n5033__, new_new_n5034__,
    new_new_n5035__, new_new_n5036__, new_new_n5037__, new_new_n5038__,
    new_new_n5039__, new_new_n5040__, new_new_n5041__, new_new_n5042__,
    new_new_n5043__, new_new_n5044__, new_new_n5045__, new_new_n5046__,
    new_new_n5047__, new_new_n5048__, new_new_n5049__, new_new_n5050__,
    new_new_n5051__, new_new_n5052__, new_new_n5053__, new_new_n5054__,
    new_new_n5055__, new_new_n5056__, new_new_n5057__, new_new_n5058__,
    new_new_n5059__, new_new_n5060__, new_new_n5061__, new_new_n5062__,
    new_new_n5063__, new_new_n5064__, new_new_n5065__, new_new_n5066__,
    new_new_n5067__, new_new_n5068__, new_new_n5069__, new_new_n5070__,
    new_new_n5071__, new_new_n5072__, new_new_n5073__, new_new_n5074__,
    new_new_n5075__, new_new_n5076__, new_new_n5077__, new_new_n5078__,
    new_new_n5079__, new_new_n5080__, new_new_n5081__, new_new_n5082__,
    new_new_n5083__, new_new_n5084__, new_new_n5085__, new_new_n5086__,
    new_new_n5087__, new_new_n5088__, new_new_n5089__, new_new_n5090__,
    new_new_n5091__, new_new_n5092__, new_new_n5093__, new_new_n5094__,
    new_new_n5095__, new_new_n5096__, new_new_n5097__, new_new_n5099__,
    new_new_n5100__, new_new_n5101__, new_new_n5102__, new_new_n5103__,
    new_new_n5104__, new_new_n5105__, new_new_n5106__, new_new_n5107__,
    new_new_n5108__, new_new_n5109__, new_new_n5110__, new_new_n5111__,
    new_new_n5112__, new_new_n5113__, new_new_n5114__, new_new_n5115__,
    new_new_n5116__, new_new_n5117__, new_new_n5118__, new_new_n5119__,
    new_new_n5120__, new_new_n5121__, new_new_n5122__, new_new_n5123__,
    new_new_n5124__, new_new_n5125__, new_new_n5126__, new_new_n5127__,
    new_new_n5128__, new_new_n5129__, new_new_n5130__, new_new_n5131__,
    new_new_n5132__, new_new_n5133__, new_new_n5134__, new_new_n5135__,
    new_new_n5136__, new_new_n5137__, new_new_n5138__, new_new_n5139__,
    new_new_n5140__, new_new_n5141__, new_new_n5142__, new_new_n5143__,
    new_new_n5144__, new_new_n5145__, new_new_n5146__, new_new_n5147__,
    new_new_n5148__, new_new_n5149__, new_new_n5150__, new_new_n5151__,
    new_new_n5152__, new_new_n5153__, new_new_n5154__, new_new_n5155__,
    new_new_n5156__, new_new_n5157__, new_new_n5158__, new_new_n5159__,
    new_new_n5160__, new_new_n5161__, new_new_n5162__, new_new_n5163__,
    new_new_n5164__, new_new_n5165__, new_new_n5166__, new_new_n5167__,
    new_new_n5168__, new_new_n5169__, new_new_n5170__, new_new_n5171__,
    new_new_n5172__, new_new_n5173__, new_new_n5174__, new_new_n5175__,
    new_new_n5176__, new_new_n5177__, new_new_n5178__, new_new_n5179__,
    new_new_n5180__, new_new_n5181__, new_new_n5182__, new_new_n5183__,
    new_new_n5184__, new_new_n5185__, new_new_n5186__, new_new_n5187__,
    new_new_n5188__, new_new_n5189__, new_new_n5190__, new_new_n5191__,
    new_new_n5192__, new_new_n5193__, new_new_n5194__, new_new_n5195__,
    new_new_n5196__, new_new_n5197__, new_new_n5198__, new_new_n5199__,
    new_new_n5200__, new_new_n5201__, new_new_n5202__, new_new_n5203__,
    new_new_n5204__, new_new_n5205__, new_new_n5206__, new_new_n5207__,
    new_new_n5208__, new_new_n5209__, new_new_n5210__, new_new_n5211__,
    new_new_n5212__, new_new_n5213__, new_new_n5214__, new_new_n5215__,
    new_new_n5216__, new_new_n5217__, new_new_n5218__, new_new_n5219__,
    new_new_n5220__, new_new_n5221__, new_new_n5222__, new_new_n5223__,
    new_new_n5224__, new_new_n5225__, new_new_n5226__, new_new_n5227__,
    new_new_n5228__, new_new_n5229__, new_new_n5230__, new_new_n5231__,
    new_new_n5232__, new_new_n5233__, new_new_n5234__, new_new_n5235__,
    new_new_n5236__, new_new_n5237__, new_new_n5238__, new_new_n5239__,
    new_new_n5240__, new_new_n5241__, new_new_n5242__, new_new_n5243__,
    new_new_n5244__, new_new_n5245__, new_new_n5246__, new_new_n5247__,
    new_new_n5248__, new_new_n5249__, new_new_n5250__, new_new_n5251__,
    new_new_n5252__, new_new_n5253__, new_new_n5254__, new_new_n5255__,
    new_new_n5256__, new_new_n5257__, new_new_n5258__, new_new_n5259__,
    new_new_n5260__, new_new_n5261__, new_new_n5262__, new_new_n5263__,
    new_new_n5264__, new_new_n5265__, new_new_n5266__, new_new_n5267__,
    new_new_n5268__, new_new_n5269__, new_new_n5270__, new_new_n5271__,
    new_new_n5272__, new_new_n5273__, new_new_n5274__, new_new_n5275__,
    new_new_n5276__, new_new_n5277__, new_new_n5278__, new_new_n5279__,
    new_new_n5280__, new_new_n5281__, new_new_n5282__, new_new_n5283__,
    new_new_n5284__, new_new_n5285__, new_new_n5286__, new_new_n5287__,
    new_new_n5288__, new_new_n5289__, new_new_n5290__, new_new_n5291__,
    new_new_n5292__, new_new_n5293__, new_new_n5294__, new_new_n5295__,
    new_new_n5296__, new_new_n5297__, new_new_n5298__, new_new_n5299__,
    new_new_n5300__, new_new_n5301__, new_new_n5302__, new_new_n5303__,
    new_new_n5304__, new_new_n5305__, new_new_n5306__, new_new_n5307__,
    new_new_n5308__, new_new_n5309__, new_new_n5310__, new_new_n5311__,
    new_new_n5312__, new_new_n5313__, new_new_n5314__, new_new_n5315__,
    new_new_n5316__, new_new_n5317__, new_new_n5318__, new_new_n5319__,
    new_new_n5320__, new_new_n5321__, new_new_n5322__, new_new_n5323__,
    new_new_n5324__, new_new_n5325__, new_new_n5326__, new_new_n5327__,
    new_new_n5328__, new_new_n5329__, new_new_n5330__, new_new_n5331__,
    new_new_n5332__, new_new_n5333__, new_new_n5334__, new_new_n5335__,
    new_new_n5336__, new_new_n5337__, new_new_n5338__, new_new_n5339__,
    new_new_n5340__, new_new_n5341__, new_new_n5342__, new_new_n5343__,
    new_new_n5344__, new_new_n5345__, new_new_n5346__, new_new_n5347__,
    new_new_n5348__, new_new_n5349__, new_new_n5350__, new_new_n5351__,
    new_new_n5352__, new_new_n5353__, new_new_n5354__, new_new_n5355__,
    new_new_n5356__, new_new_n5357__, new_new_n5358__, new_new_n5359__,
    new_new_n5360__, new_new_n5361__, new_new_n5362__, new_new_n5363__,
    new_new_n5364__, new_new_n5365__, new_new_n5366__, new_new_n5367__,
    new_new_n5368__, new_new_n5369__, new_new_n5370__, new_new_n5371__,
    new_new_n5372__, new_new_n5373__, new_new_n5374__, new_new_n5375__,
    new_new_n5376__, new_new_n5377__, new_new_n5378__, new_new_n5379__,
    new_new_n5380__, new_new_n5381__, new_new_n5382__, new_new_n5383__,
    new_new_n5384__, new_new_n5385__, new_new_n5386__, new_new_n5387__,
    new_new_n5388__, new_new_n5389__, new_new_n5390__, new_new_n5391__,
    new_new_n5392__, new_new_n5393__, new_new_n5394__, new_new_n5395__,
    new_new_n5396__, new_new_n5397__, new_new_n5398__, new_new_n5399__,
    new_new_n5400__, new_new_n5401__, new_new_n5402__, new_new_n5403__,
    new_new_n5404__, new_new_n5405__, new_new_n5406__, new_new_n5407__,
    new_new_n5408__, new_new_n5409__, new_new_n5410__, new_new_n5411__,
    new_new_n5412__, new_new_n5413__, new_new_n5414__, new_new_n5415__,
    new_new_n5416__, new_new_n5417__, new_new_n5418__, new_new_n5419__,
    new_new_n5420__, new_new_n5421__, new_new_n5422__, new_new_n5423__,
    new_new_n5424__, new_new_n5425__, new_new_n5426__, new_new_n5427__,
    new_new_n5428__, new_new_n5429__, new_new_n5430__, new_new_n5431__,
    new_new_n5432__, new_new_n5433__, new_new_n5434__, new_new_n5435__,
    new_new_n5436__, new_new_n5437__, new_new_n5439__, new_new_n5440__,
    new_new_n5441__, new_new_n5442__, new_new_n5443__, new_new_n5444__,
    new_new_n5445__, new_new_n5446__, new_new_n5447__, new_new_n5448__,
    new_new_n5449__, new_new_n5450__, new_new_n5451__, new_new_n5452__,
    new_new_n5453__, new_new_n5454__, new_new_n5455__, new_new_n5456__,
    new_new_n5457__, new_new_n5458__, new_new_n5459__, new_new_n5460__,
    new_new_n5461__, new_new_n5462__, new_new_n5463__, new_new_n5464__,
    new_new_n5465__, new_new_n5466__, new_new_n5467__, new_new_n5468__,
    new_new_n5469__, new_new_n5470__, new_new_n5471__, new_new_n5472__,
    new_new_n5473__, new_new_n5474__, new_new_n5475__, new_new_n5476__,
    new_new_n5477__, new_new_n5478__, new_new_n5479__, new_new_n5480__,
    new_new_n5481__, new_new_n5482__, new_new_n5483__, new_new_n5484__,
    new_new_n5485__, new_new_n5486__, new_new_n5487__, new_new_n5488__,
    new_new_n5489__, new_new_n5490__, new_new_n5491__, new_new_n5492__,
    new_new_n5493__, new_new_n5494__, new_new_n5495__, new_new_n5496__,
    new_new_n5497__, new_new_n5498__, new_new_n5499__, new_new_n5500__,
    new_new_n5501__, new_new_n5502__, new_new_n5503__, new_new_n5504__,
    new_new_n5505__, new_new_n5506__, new_new_n5507__, new_new_n5508__,
    new_new_n5509__, new_new_n5510__, new_new_n5511__, new_new_n5512__,
    new_new_n5513__, new_new_n5514__, new_new_n5515__, new_new_n5516__,
    new_new_n5517__, new_new_n5518__, new_new_n5519__, new_new_n5520__,
    new_new_n5521__, new_new_n5522__, new_new_n5523__, new_new_n5524__,
    new_new_n5525__, new_new_n5526__, new_new_n5527__, new_new_n5528__,
    new_new_n5529__, new_new_n5530__, new_new_n5531__, new_new_n5532__,
    new_new_n5533__, new_new_n5534__, new_new_n5535__, new_new_n5536__,
    new_new_n5537__, new_new_n5538__, new_new_n5539__, new_new_n5540__,
    new_new_n5541__, new_new_n5542__, new_new_n5543__, new_new_n5544__,
    new_new_n5545__, new_new_n5546__, new_new_n5547__, new_new_n5548__,
    new_new_n5549__, new_new_n5550__, new_new_n5551__, new_new_n5552__,
    new_new_n5553__, new_new_n5554__, new_new_n5555__, new_new_n5556__,
    new_new_n5557__, new_new_n5558__, new_new_n5559__, new_new_n5560__,
    new_new_n5561__, new_new_n5562__, new_new_n5563__, new_new_n5564__,
    new_new_n5565__, new_new_n5566__, new_new_n5567__, new_new_n5568__,
    new_new_n5569__, new_new_n5570__, new_new_n5571__, new_new_n5572__,
    new_new_n5573__, new_new_n5574__, new_new_n5575__, new_new_n5576__,
    new_new_n5577__, new_new_n5578__, new_new_n5579__, new_new_n5580__,
    new_new_n5581__, new_new_n5582__, new_new_n5583__, new_new_n5584__,
    new_new_n5585__, new_new_n5586__, new_new_n5587__, new_new_n5588__,
    new_new_n5589__, new_new_n5590__, new_new_n5591__, new_new_n5592__,
    new_new_n5593__, new_new_n5594__, new_new_n5595__, new_new_n5596__,
    new_new_n5597__, new_new_n5598__, new_new_n5599__, new_new_n5600__,
    new_new_n5601__, new_new_n5602__, new_new_n5603__, new_new_n5604__,
    new_new_n5605__, new_new_n5606__, new_new_n5607__, new_new_n5608__,
    new_new_n5609__, new_new_n5610__, new_new_n5611__, new_new_n5612__,
    new_new_n5613__, new_new_n5614__, new_new_n5615__, new_new_n5616__,
    new_new_n5617__, new_new_n5618__, new_new_n5619__, new_new_n5620__,
    new_new_n5621__, new_new_n5622__, new_new_n5623__, new_new_n5624__,
    new_new_n5625__, new_new_n5626__, new_new_n5627__, new_new_n5628__,
    new_new_n5629__, new_new_n5630__, new_new_n5631__, new_new_n5632__,
    new_new_n5633__, new_new_n5634__, new_new_n5635__, new_new_n5636__,
    new_new_n5637__, new_new_n5638__, new_new_n5639__, new_new_n5640__,
    new_new_n5641__, new_new_n5642__, new_new_n5643__, new_new_n5644__,
    new_new_n5645__, new_new_n5646__, new_new_n5647__, new_new_n5648__,
    new_new_n5649__, new_new_n5650__, new_new_n5651__, new_new_n5652__,
    new_new_n5653__, new_new_n5654__, new_new_n5655__, new_new_n5656__,
    new_new_n5657__, new_new_n5658__, new_new_n5659__, new_new_n5660__,
    new_new_n5661__, new_new_n5662__, new_new_n5663__, new_new_n5664__,
    new_new_n5665__, new_new_n5666__, new_new_n5667__, new_new_n5668__,
    new_new_n5669__, new_new_n5670__, new_new_n5671__, new_new_n5672__,
    new_new_n5673__, new_new_n5674__, new_new_n5675__, new_new_n5676__,
    new_new_n5677__, new_new_n5678__, new_new_n5679__, new_new_n5680__,
    new_new_n5681__, new_new_n5682__, new_new_n5683__, new_new_n5684__,
    new_new_n5685__, new_new_n5686__, new_new_n5687__, new_new_n5688__,
    new_new_n5689__, new_new_n5690__, new_new_n5691__, new_new_n5692__,
    new_new_n5693__, new_new_n5694__, new_new_n5695__, new_new_n5696__,
    new_new_n5697__, new_new_n5698__, new_new_n5699__, new_new_n5700__,
    new_new_n5701__, new_new_n5702__, new_new_n5703__, new_new_n5704__,
    new_new_n5705__, new_new_n5706__, new_new_n5707__, new_new_n5708__,
    new_new_n5709__, new_new_n5710__, new_new_n5711__, new_new_n5712__,
    new_new_n5713__, new_new_n5714__, new_new_n5715__, new_new_n5716__,
    new_new_n5717__, new_new_n5718__, new_new_n5719__, new_new_n5720__,
    new_new_n5721__, new_new_n5722__, new_new_n5723__, new_new_n5724__,
    new_new_n5725__, new_new_n5726__, new_new_n5727__, new_new_n5728__,
    new_new_n5729__, new_new_n5730__, new_new_n5731__, new_new_n5732__,
    new_new_n5733__, new_new_n5734__, new_new_n5735__, new_new_n5736__,
    new_new_n5737__, new_new_n5738__, new_new_n5739__, new_new_n5740__,
    new_new_n5741__, new_new_n5742__, new_new_n5743__, new_new_n5744__,
    new_new_n5745__, new_new_n5746__, new_new_n5747__, new_new_n5748__,
    new_new_n5749__, new_new_n5750__, new_new_n5751__, new_new_n5752__,
    new_new_n5753__, new_new_n5754__, new_new_n5755__, new_new_n5756__,
    new_new_n5757__, new_new_n5758__, new_new_n5759__, new_new_n5760__,
    new_new_n5761__, new_new_n5762__, new_new_n5763__, new_new_n5764__,
    new_new_n5765__, new_new_n5766__, new_new_n5767__, new_new_n5768__,
    new_new_n5769__, new_new_n5771__, new_new_n5772__, new_new_n5773__,
    new_new_n5774__, new_new_n5775__, new_new_n5776__, new_new_n5777__,
    new_new_n5778__, new_new_n5779__, new_new_n5780__, new_new_n5781__,
    new_new_n5782__, new_new_n5783__, new_new_n5784__, new_new_n5785__,
    new_new_n5786__, new_new_n5787__, new_new_n5788__, new_new_n5789__,
    new_new_n5790__, new_new_n5791__, new_new_n5792__, new_new_n5793__,
    new_new_n5794__, new_new_n5795__, new_new_n5796__, new_new_n5797__,
    new_new_n5798__, new_new_n5799__, new_new_n5800__, new_new_n5801__,
    new_new_n5802__, new_new_n5803__, new_new_n5804__, new_new_n5805__,
    new_new_n5806__, new_new_n5807__, new_new_n5808__, new_new_n5809__,
    new_new_n5810__, new_new_n5811__, new_new_n5812__, new_new_n5813__,
    new_new_n5814__, new_new_n5815__, new_new_n5816__, new_new_n5817__,
    new_new_n5818__, new_new_n5819__, new_new_n5820__, new_new_n5821__,
    new_new_n5822__, new_new_n5823__, new_new_n5824__, new_new_n5825__,
    new_new_n5826__, new_new_n5827__, new_new_n5828__, new_new_n5829__,
    new_new_n5830__, new_new_n5831__, new_new_n5832__, new_new_n5833__,
    new_new_n5834__, new_new_n5835__, new_new_n5836__, new_new_n5837__,
    new_new_n5838__, new_new_n5839__, new_new_n5840__, new_new_n5841__,
    new_new_n5842__, new_new_n5843__, new_new_n5844__, new_new_n5845__,
    new_new_n5846__, new_new_n5847__, new_new_n5848__, new_new_n5849__,
    new_new_n5850__, new_new_n5851__, new_new_n5852__, new_new_n5853__,
    new_new_n5854__, new_new_n5855__, new_new_n5856__, new_new_n5857__,
    new_new_n5858__, new_new_n5859__, new_new_n5860__, new_new_n5861__,
    new_new_n5862__, new_new_n5863__, new_new_n5864__, new_new_n5865__,
    new_new_n5866__, new_new_n5867__, new_new_n5868__, new_new_n5869__,
    new_new_n5870__, new_new_n5871__, new_new_n5872__, new_new_n5873__,
    new_new_n5874__, new_new_n5875__, new_new_n5876__, new_new_n5877__,
    new_new_n5878__, new_new_n5879__, new_new_n5880__, new_new_n5881__,
    new_new_n5882__, new_new_n5883__, new_new_n5884__, new_new_n5885__,
    new_new_n5886__, new_new_n5887__, new_new_n5888__, new_new_n5889__,
    new_new_n5890__, new_new_n5891__, new_new_n5892__, new_new_n5893__,
    new_new_n5894__, new_new_n5895__, new_new_n5896__, new_new_n5897__,
    new_new_n5898__, new_new_n5899__, new_new_n5900__, new_new_n5901__,
    new_new_n5902__, new_new_n5903__, new_new_n5904__, new_new_n5905__,
    new_new_n5906__, new_new_n5907__, new_new_n5908__, new_new_n5909__,
    new_new_n5910__, new_new_n5911__, new_new_n5912__, new_new_n5913__,
    new_new_n5914__, new_new_n5915__, new_new_n5916__, new_new_n5917__,
    new_new_n5918__, new_new_n5919__, new_new_n5920__, new_new_n5921__,
    new_new_n5922__, new_new_n5923__, new_new_n5924__, new_new_n5925__,
    new_new_n5926__, new_new_n5927__, new_new_n5928__, new_new_n5929__,
    new_new_n5930__, new_new_n5931__, new_new_n5932__, new_new_n5933__,
    new_new_n5934__, new_new_n5935__, new_new_n5936__, new_new_n5937__,
    new_new_n5938__, new_new_n5939__, new_new_n5940__, new_new_n5941__,
    new_new_n5942__, new_new_n5943__, new_new_n5944__, new_new_n5945__,
    new_new_n5946__, new_new_n5947__, new_new_n5948__, new_new_n5949__,
    new_new_n5950__, new_new_n5951__, new_new_n5952__, new_new_n5953__,
    new_new_n5954__, new_new_n5955__, new_new_n5956__, new_new_n5957__,
    new_new_n5958__, new_new_n5959__, new_new_n5960__, new_new_n5961__,
    new_new_n5962__, new_new_n5963__, new_new_n5964__, new_new_n5965__,
    new_new_n5966__, new_new_n5967__, new_new_n5968__, new_new_n5969__,
    new_new_n5970__, new_new_n5971__, new_new_n5972__, new_new_n5973__,
    new_new_n5974__, new_new_n5975__, new_new_n5976__, new_new_n5977__,
    new_new_n5978__, new_new_n5979__, new_new_n5980__, new_new_n5981__,
    new_new_n5982__, new_new_n5983__, new_new_n5984__, new_new_n5985__,
    new_new_n5986__, new_new_n5987__, new_new_n5988__, new_new_n5989__,
    new_new_n5990__, new_new_n5991__, new_new_n5992__, new_new_n5993__,
    new_new_n5994__, new_new_n5995__, new_new_n5996__, new_new_n5997__,
    new_new_n5998__, new_new_n5999__, new_new_n6000__, new_new_n6001__,
    new_new_n6002__, new_new_n6003__, new_new_n6004__, new_new_n6005__,
    new_new_n6006__, new_new_n6007__, new_new_n6008__, new_new_n6009__,
    new_new_n6010__, new_new_n6011__, new_new_n6012__, new_new_n6013__,
    new_new_n6014__, new_new_n6015__, new_new_n6016__, new_new_n6017__,
    new_new_n6018__, new_new_n6019__, new_new_n6020__, new_new_n6021__,
    new_new_n6022__, new_new_n6023__, new_new_n6024__, new_new_n6025__,
    new_new_n6026__, new_new_n6027__, new_new_n6028__, new_new_n6029__,
    new_new_n6030__, new_new_n6031__, new_new_n6032__, new_new_n6033__,
    new_new_n6034__, new_new_n6035__, new_new_n6036__, new_new_n6037__,
    new_new_n6038__, new_new_n6039__, new_new_n6040__, new_new_n6041__,
    new_new_n6042__, new_new_n6043__, new_new_n6044__, new_new_n6045__,
    new_new_n6046__, new_new_n6047__, new_new_n6048__, new_new_n6049__,
    new_new_n6050__, new_new_n6051__, new_new_n6052__, new_new_n6053__,
    new_new_n6054__, new_new_n6055__, new_new_n6056__, new_new_n6057__,
    new_new_n6058__, new_new_n6059__, new_new_n6060__, new_new_n6061__,
    new_new_n6062__, new_new_n6063__, new_new_n6064__, new_new_n6065__,
    new_new_n6066__, new_new_n6067__, new_new_n6068__, new_new_n6069__,
    new_new_n6070__, new_new_n6071__, new_new_n6072__, new_new_n6073__,
    new_new_n6074__, new_new_n6075__, new_new_n6076__, new_new_n6077__,
    new_new_n6078__, new_new_n6079__, new_new_n6080__, new_new_n6081__,
    new_new_n6082__, new_new_n6083__, new_new_n6084__, new_new_n6085__,
    new_new_n6086__, new_new_n6087__, new_new_n6088__, new_new_n6089__,
    new_new_n6090__, new_new_n6091__, new_new_n6092__, new_new_n6093__,
    new_new_n6094__, new_new_n6095__, new_new_n6096__, new_new_n6097__,
    new_new_n6098__, new_new_n6099__, new_new_n6100__, new_new_n6101__,
    new_new_n6102__, new_new_n6103__, new_new_n6104__, new_new_n6105__,
    new_new_n6106__, new_new_n6107__, new_new_n6108__, new_new_n6109__,
    new_new_n6110__, new_new_n6111__, new_new_n6112__, new_new_n6113__,
    new_new_n6114__, new_new_n6115__, new_new_n6116__, new_new_n6117__,
    new_new_n6118__, new_new_n6119__, new_new_n6120__, new_new_n6121__,
    new_new_n6122__, new_new_n6123__, new_new_n6124__, new_new_n6125__,
    new_new_n6126__, new_new_n6127__, new_new_n6128__, new_new_n6129__,
    new_new_n6130__, new_new_n6131__, new_new_n6132__, new_new_n6133__,
    new_new_n6134__, new_new_n6135__, new_new_n6137__, new_new_n6138__,
    new_new_n6139__, new_new_n6140__, new_new_n6141__, new_new_n6142__,
    new_new_n6143__, new_new_n6144__, new_new_n6145__, new_new_n6146__,
    new_new_n6147__, new_new_n6148__, new_new_n6149__, new_new_n6150__,
    new_new_n6151__, new_new_n6152__, new_new_n6153__, new_new_n6154__,
    new_new_n6155__, new_new_n6156__, new_new_n6157__, new_new_n6158__,
    new_new_n6159__, new_new_n6160__, new_new_n6161__, new_new_n6162__,
    new_new_n6163__, new_new_n6164__, new_new_n6165__, new_new_n6166__,
    new_new_n6167__, new_new_n6168__, new_new_n6169__, new_new_n6170__,
    new_new_n6171__, new_new_n6172__, new_new_n6173__, new_new_n6174__,
    new_new_n6175__, new_new_n6176__, new_new_n6177__, new_new_n6178__,
    new_new_n6179__, new_new_n6180__, new_new_n6181__, new_new_n6182__,
    new_new_n6183__, new_new_n6184__, new_new_n6185__, new_new_n6186__,
    new_new_n6187__, new_new_n6188__, new_new_n6189__, new_new_n6190__,
    new_new_n6191__, new_new_n6192__, new_new_n6193__, new_new_n6194__,
    new_new_n6195__, new_new_n6196__, new_new_n6197__, new_new_n6198__,
    new_new_n6199__, new_new_n6200__, new_new_n6201__, new_new_n6202__,
    new_new_n6203__, new_new_n6204__, new_new_n6205__, new_new_n6206__,
    new_new_n6207__, new_new_n6208__, new_new_n6209__, new_new_n6210__,
    new_new_n6211__, new_new_n6212__, new_new_n6213__, new_new_n6214__,
    new_new_n6215__, new_new_n6216__, new_new_n6217__, new_new_n6218__,
    new_new_n6219__, new_new_n6220__, new_new_n6221__, new_new_n6222__,
    new_new_n6223__, new_new_n6224__, new_new_n6225__, new_new_n6226__,
    new_new_n6227__, new_new_n6228__, new_new_n6229__, new_new_n6230__,
    new_new_n6231__, new_new_n6232__, new_new_n6233__, new_new_n6234__,
    new_new_n6235__, new_new_n6236__, new_new_n6237__, new_new_n6238__,
    new_new_n6239__, new_new_n6240__, new_new_n6241__, new_new_n6242__,
    new_new_n6243__, new_new_n6244__, new_new_n6245__, new_new_n6246__,
    new_new_n6247__, new_new_n6248__, new_new_n6249__, new_new_n6250__,
    new_new_n6251__, new_new_n6252__, new_new_n6253__, new_new_n6254__,
    new_new_n6255__, new_new_n6256__, new_new_n6257__, new_new_n6258__,
    new_new_n6259__, new_new_n6260__, new_new_n6261__, new_new_n6262__,
    new_new_n6263__, new_new_n6264__, new_new_n6265__, new_new_n6266__,
    new_new_n6267__, new_new_n6268__, new_new_n6269__, new_new_n6270__,
    new_new_n6271__, new_new_n6272__, new_new_n6273__, new_new_n6274__,
    new_new_n6275__, new_new_n6276__, new_new_n6277__, new_new_n6278__,
    new_new_n6279__, new_new_n6280__, new_new_n6281__, new_new_n6282__,
    new_new_n6283__, new_new_n6284__, new_new_n6285__, new_new_n6286__,
    new_new_n6287__, new_new_n6288__, new_new_n6289__, new_new_n6290__,
    new_new_n6291__, new_new_n6292__, new_new_n6293__, new_new_n6294__,
    new_new_n6295__, new_new_n6296__, new_new_n6297__, new_new_n6298__,
    new_new_n6299__, new_new_n6300__, new_new_n6301__, new_new_n6302__,
    new_new_n6303__, new_new_n6304__, new_new_n6305__, new_new_n6306__,
    new_new_n6307__, new_new_n6308__, new_new_n6309__, new_new_n6310__,
    new_new_n6311__, new_new_n6312__, new_new_n6313__, new_new_n6314__,
    new_new_n6315__, new_new_n6316__, new_new_n6317__, new_new_n6318__,
    new_new_n6319__, new_new_n6320__, new_new_n6321__, new_new_n6322__,
    new_new_n6323__, new_new_n6324__, new_new_n6325__, new_new_n6326__,
    new_new_n6327__, new_new_n6328__, new_new_n6329__, new_new_n6330__,
    new_new_n6331__, new_new_n6332__, new_new_n6333__, new_new_n6334__,
    new_new_n6335__, new_new_n6336__, new_new_n6337__, new_new_n6338__,
    new_new_n6339__, new_new_n6340__, new_new_n6341__, new_new_n6342__,
    new_new_n6343__, new_new_n6344__, new_new_n6345__, new_new_n6346__,
    new_new_n6347__, new_new_n6348__, new_new_n6349__, new_new_n6350__,
    new_new_n6351__, new_new_n6352__, new_new_n6353__, new_new_n6354__,
    new_new_n6355__, new_new_n6356__, new_new_n6357__, new_new_n6358__,
    new_new_n6359__, new_new_n6360__, new_new_n6361__, new_new_n6362__,
    new_new_n6363__, new_new_n6364__, new_new_n6365__, new_new_n6366__,
    new_new_n6367__, new_new_n6368__, new_new_n6369__, new_new_n6370__,
    new_new_n6371__, new_new_n6372__, new_new_n6373__, new_new_n6374__,
    new_new_n6375__, new_new_n6376__, new_new_n6377__, new_new_n6378__,
    new_new_n6379__, new_new_n6380__, new_new_n6381__, new_new_n6382__,
    new_new_n6383__, new_new_n6384__, new_new_n6385__, new_new_n6386__,
    new_new_n6387__, new_new_n6388__, new_new_n6389__, new_new_n6390__,
    new_new_n6391__, new_new_n6392__, new_new_n6393__, new_new_n6394__,
    new_new_n6395__, new_new_n6396__, new_new_n6397__, new_new_n6398__,
    new_new_n6399__, new_new_n6400__, new_new_n6401__, new_new_n6402__,
    new_new_n6403__, new_new_n6404__, new_new_n6405__, new_new_n6406__,
    new_new_n6407__, new_new_n6408__, new_new_n6409__, new_new_n6410__,
    new_new_n6411__, new_new_n6412__, new_new_n6413__, new_new_n6414__,
    new_new_n6415__, new_new_n6416__, new_new_n6417__, new_new_n6418__,
    new_new_n6419__, new_new_n6420__, new_new_n6421__, new_new_n6422__,
    new_new_n6423__, new_new_n6424__, new_new_n6425__, new_new_n6426__,
    new_new_n6427__, new_new_n6428__, new_new_n6429__, new_new_n6430__,
    new_new_n6431__, new_new_n6432__, new_new_n6433__, new_new_n6434__,
    new_new_n6435__, new_new_n6436__, new_new_n6437__, new_new_n6438__,
    new_new_n6439__, new_new_n6440__, new_new_n6441__, new_new_n6442__,
    new_new_n6443__, new_new_n6444__, new_new_n6445__, new_new_n6446__,
    new_new_n6447__, new_new_n6448__, new_new_n6449__, new_new_n6450__,
    new_new_n6451__, new_new_n6452__, new_new_n6453__, new_new_n6454__,
    new_new_n6455__, new_new_n6456__, new_new_n6457__, new_new_n6458__,
    new_new_n6459__, new_new_n6460__, new_new_n6461__, new_new_n6462__,
    new_new_n6463__, new_new_n6464__, new_new_n6465__, new_new_n6466__,
    new_new_n6467__, new_new_n6468__, new_new_n6469__, new_new_n6470__,
    new_new_n6471__, new_new_n6472__, new_new_n6473__, new_new_n6474__,
    new_new_n6475__, new_new_n6476__, new_new_n6477__, new_new_n6478__,
    new_new_n6479__, new_new_n6480__, new_new_n6481__, new_new_n6482__,
    new_new_n6483__, new_new_n6484__, new_new_n6485__, new_new_n6486__,
    new_new_n6487__, new_new_n6488__, new_new_n6489__, new_new_n6490__,
    new_new_n6491__, new_new_n6492__, new_new_n6494__, new_new_n6495__,
    new_new_n6496__, new_new_n6497__, new_new_n6498__, new_new_n6499__,
    new_new_n6500__, new_new_n6501__, new_new_n6502__, new_new_n6503__,
    new_new_n6504__, new_new_n6505__, new_new_n6506__, new_new_n6507__,
    new_new_n6508__, new_new_n6509__, new_new_n6510__, new_new_n6511__,
    new_new_n6512__, new_new_n6513__, new_new_n6514__, new_new_n6515__,
    new_new_n6516__, new_new_n6517__, new_new_n6518__, new_new_n6519__,
    new_new_n6520__, new_new_n6521__, new_new_n6522__, new_new_n6523__,
    new_new_n6524__, new_new_n6525__, new_new_n6526__, new_new_n6527__,
    new_new_n6528__, new_new_n6529__, new_new_n6530__, new_new_n6531__,
    new_new_n6532__, new_new_n6533__, new_new_n6534__, new_new_n6535__,
    new_new_n6536__, new_new_n6537__, new_new_n6538__, new_new_n6539__,
    new_new_n6540__, new_new_n6541__, new_new_n6542__, new_new_n6543__,
    new_new_n6544__, new_new_n6545__, new_new_n6546__, new_new_n6547__,
    new_new_n6548__, new_new_n6549__, new_new_n6550__, new_new_n6551__,
    new_new_n6552__, new_new_n6553__, new_new_n6554__, new_new_n6555__,
    new_new_n6556__, new_new_n6557__, new_new_n6558__, new_new_n6559__,
    new_new_n6560__, new_new_n6561__, new_new_n6562__, new_new_n6563__,
    new_new_n6564__, new_new_n6565__, new_new_n6566__, new_new_n6567__,
    new_new_n6568__, new_new_n6569__, new_new_n6570__, new_new_n6571__,
    new_new_n6572__, new_new_n6573__, new_new_n6574__, new_new_n6575__,
    new_new_n6576__, new_new_n6577__, new_new_n6578__, new_new_n6579__,
    new_new_n6580__, new_new_n6581__, new_new_n6582__, new_new_n6583__,
    new_new_n6584__, new_new_n6585__, new_new_n6586__, new_new_n6587__,
    new_new_n6588__, new_new_n6589__, new_new_n6590__, new_new_n6591__,
    new_new_n6592__, new_new_n6593__, new_new_n6594__, new_new_n6595__,
    new_new_n6596__, new_new_n6597__, new_new_n6598__, new_new_n6599__,
    new_new_n6600__, new_new_n6601__, new_new_n6602__, new_new_n6603__,
    new_new_n6604__, new_new_n6605__, new_new_n6606__, new_new_n6607__,
    new_new_n6608__, new_new_n6609__, new_new_n6610__, new_new_n6611__,
    new_new_n6612__, new_new_n6613__, new_new_n6614__, new_new_n6615__,
    new_new_n6616__, new_new_n6617__, new_new_n6618__, new_new_n6619__,
    new_new_n6620__, new_new_n6621__, new_new_n6622__, new_new_n6623__,
    new_new_n6624__, new_new_n6625__, new_new_n6626__, new_new_n6627__,
    new_new_n6628__, new_new_n6629__, new_new_n6630__, new_new_n6631__,
    new_new_n6632__, new_new_n6633__, new_new_n6634__, new_new_n6635__,
    new_new_n6636__, new_new_n6637__, new_new_n6638__, new_new_n6639__,
    new_new_n6640__, new_new_n6641__, new_new_n6642__, new_new_n6643__,
    new_new_n6644__, new_new_n6645__, new_new_n6646__, new_new_n6647__,
    new_new_n6648__, new_new_n6649__, new_new_n6650__, new_new_n6651__,
    new_new_n6652__, new_new_n6653__, new_new_n6654__, new_new_n6655__,
    new_new_n6656__, new_new_n6657__, new_new_n6658__, new_new_n6659__,
    new_new_n6660__, new_new_n6661__, new_new_n6662__, new_new_n6663__,
    new_new_n6664__, new_new_n6665__, new_new_n6666__, new_new_n6667__,
    new_new_n6668__, new_new_n6669__, new_new_n6670__, new_new_n6671__,
    new_new_n6672__, new_new_n6673__, new_new_n6674__, new_new_n6675__,
    new_new_n6676__, new_new_n6677__, new_new_n6678__, new_new_n6679__,
    new_new_n6680__, new_new_n6681__, new_new_n6682__, new_new_n6683__,
    new_new_n6684__, new_new_n6685__, new_new_n6686__, new_new_n6687__,
    new_new_n6688__, new_new_n6689__, new_new_n6690__, new_new_n6691__,
    new_new_n6692__, new_new_n6693__, new_new_n6694__, new_new_n6695__,
    new_new_n6696__, new_new_n6697__, new_new_n6698__, new_new_n6699__,
    new_new_n6700__, new_new_n6701__, new_new_n6702__, new_new_n6703__,
    new_new_n6704__, new_new_n6705__, new_new_n6706__, new_new_n6707__,
    new_new_n6708__, new_new_n6709__, new_new_n6710__, new_new_n6711__,
    new_new_n6712__, new_new_n6713__, new_new_n6714__, new_new_n6715__,
    new_new_n6716__, new_new_n6717__, new_new_n6718__, new_new_n6719__,
    new_new_n6720__, new_new_n6721__, new_new_n6722__, new_new_n6723__,
    new_new_n6724__, new_new_n6725__, new_new_n6726__, new_new_n6727__,
    new_new_n6728__, new_new_n6729__, new_new_n6730__, new_new_n6731__,
    new_new_n6732__, new_new_n6733__, new_new_n6734__, new_new_n6735__,
    new_new_n6736__, new_new_n6737__, new_new_n6738__, new_new_n6739__,
    new_new_n6740__, new_new_n6741__, new_new_n6742__, new_new_n6743__,
    new_new_n6744__, new_new_n6745__, new_new_n6746__, new_new_n6747__,
    new_new_n6748__, new_new_n6749__, new_new_n6750__, new_new_n6751__,
    new_new_n6752__, new_new_n6753__, new_new_n6754__, new_new_n6755__,
    new_new_n6756__, new_new_n6757__, new_new_n6758__, new_new_n6759__,
    new_new_n6760__, new_new_n6761__, new_new_n6762__, new_new_n6763__,
    new_new_n6764__, new_new_n6765__, new_new_n6766__, new_new_n6767__,
    new_new_n6768__, new_new_n6769__, new_new_n6770__, new_new_n6771__,
    new_new_n6772__, new_new_n6773__, new_new_n6774__, new_new_n6775__,
    new_new_n6776__, new_new_n6777__, new_new_n6778__, new_new_n6779__,
    new_new_n6780__, new_new_n6781__, new_new_n6782__, new_new_n6783__,
    new_new_n6784__, new_new_n6785__, new_new_n6786__, new_new_n6787__,
    new_new_n6788__, new_new_n6789__, new_new_n6790__, new_new_n6791__,
    new_new_n6792__, new_new_n6793__, new_new_n6794__, new_new_n6795__,
    new_new_n6796__, new_new_n6797__, new_new_n6798__, new_new_n6799__,
    new_new_n6800__, new_new_n6801__, new_new_n6802__, new_new_n6803__,
    new_new_n6804__, new_new_n6805__, new_new_n6806__, new_new_n6807__,
    new_new_n6808__, new_new_n6809__, new_new_n6810__, new_new_n6811__,
    new_new_n6812__, new_new_n6813__, new_new_n6814__, new_new_n6815__,
    new_new_n6816__, new_new_n6817__, new_new_n6818__, new_new_n6819__,
    new_new_n6820__, new_new_n6821__, new_new_n6822__, new_new_n6823__,
    new_new_n6824__, new_new_n6825__, new_new_n6826__, new_new_n6827__,
    new_new_n6828__, new_new_n6829__, new_new_n6830__, new_new_n6831__,
    new_new_n6832__, new_new_n6833__, new_new_n6834__, new_new_n6835__,
    new_new_n6836__, new_new_n6837__, new_new_n6838__, new_new_n6839__,
    new_new_n6840__, new_new_n6841__, new_new_n6842__, new_new_n6843__,
    new_new_n6844__, new_new_n6845__, new_new_n6846__, new_new_n6847__,
    new_new_n6848__, new_new_n6849__, new_new_n6850__, new_new_n6851__,
    new_new_n6852__, new_new_n6853__, new_new_n6854__, new_new_n6855__,
    new_new_n6856__, new_new_n6857__, new_new_n6858__, new_new_n6859__,
    new_new_n6860__, new_new_n6861__, new_new_n6862__, new_new_n6863__,
    new_new_n6864__, new_new_n6865__, new_new_n6866__, new_new_n6867__,
    new_new_n6869__, new_new_n6870__, new_new_n6871__, new_new_n6872__,
    new_new_n6873__, new_new_n6874__, new_new_n6875__, new_new_n6876__,
    new_new_n6877__, new_new_n6878__, new_new_n6879__, new_new_n6880__,
    new_new_n6881__, new_new_n6882__, new_new_n6883__, new_new_n6884__,
    new_new_n6885__, new_new_n6886__, new_new_n6887__, new_new_n6888__,
    new_new_n6889__, new_new_n6890__, new_new_n6891__, new_new_n6892__,
    new_new_n6893__, new_new_n6894__, new_new_n6895__, new_new_n6896__,
    new_new_n6897__, new_new_n6898__, new_new_n6899__, new_new_n6900__,
    new_new_n6901__, new_new_n6902__, new_new_n6903__, new_new_n6904__,
    new_new_n6905__, new_new_n6906__, new_new_n6907__, new_new_n6908__,
    new_new_n6909__, new_new_n6910__, new_new_n6911__, new_new_n6912__,
    new_new_n6913__, new_new_n6914__, new_new_n6915__, new_new_n6916__,
    new_new_n6917__, new_new_n6918__, new_new_n6919__, new_new_n6920__,
    new_new_n6921__, new_new_n6922__, new_new_n6923__, new_new_n6924__,
    new_new_n6925__, new_new_n6926__, new_new_n6927__, new_new_n6928__,
    new_new_n6929__, new_new_n6930__, new_new_n6931__, new_new_n6932__,
    new_new_n6933__, new_new_n6934__, new_new_n6935__, new_new_n6936__,
    new_new_n6937__, new_new_n6938__, new_new_n6939__, new_new_n6940__,
    new_new_n6941__, new_new_n6942__, new_new_n6943__, new_new_n6944__,
    new_new_n6945__, new_new_n6946__, new_new_n6947__, new_new_n6948__,
    new_new_n6949__, new_new_n6950__, new_new_n6951__, new_new_n6952__,
    new_new_n6953__, new_new_n6954__, new_new_n6955__, new_new_n6956__,
    new_new_n6957__, new_new_n6958__, new_new_n6959__, new_new_n6960__,
    new_new_n6961__, new_new_n6962__, new_new_n6963__, new_new_n6964__,
    new_new_n6965__, new_new_n6966__, new_new_n6967__, new_new_n6968__,
    new_new_n6969__, new_new_n6970__, new_new_n6971__, new_new_n6972__,
    new_new_n6973__, new_new_n6974__, new_new_n6975__, new_new_n6976__,
    new_new_n6977__, new_new_n6978__, new_new_n6979__, new_new_n6980__,
    new_new_n6981__, new_new_n6982__, new_new_n6983__, new_new_n6984__,
    new_new_n6985__, new_new_n6986__, new_new_n6987__, new_new_n6988__,
    new_new_n6989__, new_new_n6990__, new_new_n6991__, new_new_n6992__,
    new_new_n6993__, new_new_n6994__, new_new_n6995__, new_new_n6996__,
    new_new_n6997__, new_new_n6998__, new_new_n6999__, new_new_n7000__,
    new_new_n7001__, new_new_n7002__, new_new_n7003__, new_new_n7004__,
    new_new_n7005__, new_new_n7006__, new_new_n7007__, new_new_n7008__,
    new_new_n7009__, new_new_n7010__, new_new_n7011__, new_new_n7012__,
    new_new_n7013__, new_new_n7014__, new_new_n7015__, new_new_n7016__,
    new_new_n7017__, new_new_n7018__, new_new_n7019__, new_new_n7020__,
    new_new_n7021__, new_new_n7022__, new_new_n7023__, new_new_n7024__,
    new_new_n7025__, new_new_n7026__, new_new_n7027__, new_new_n7028__,
    new_new_n7029__, new_new_n7030__, new_new_n7031__, new_new_n7032__,
    new_new_n7033__, new_new_n7034__, new_new_n7035__, new_new_n7036__,
    new_new_n7037__, new_new_n7038__, new_new_n7039__, new_new_n7040__,
    new_new_n7041__, new_new_n7042__, new_new_n7043__, new_new_n7044__,
    new_new_n7045__, new_new_n7046__, new_new_n7047__, new_new_n7048__,
    new_new_n7049__, new_new_n7050__, new_new_n7051__, new_new_n7052__,
    new_new_n7053__, new_new_n7054__, new_new_n7055__, new_new_n7056__,
    new_new_n7057__, new_new_n7058__, new_new_n7059__, new_new_n7060__,
    new_new_n7061__, new_new_n7062__, new_new_n7063__, new_new_n7064__,
    new_new_n7065__, new_new_n7066__, new_new_n7067__, new_new_n7068__,
    new_new_n7069__, new_new_n7070__, new_new_n7071__, new_new_n7072__,
    new_new_n7073__, new_new_n7074__, new_new_n7075__, new_new_n7076__,
    new_new_n7077__, new_new_n7078__, new_new_n7079__, new_new_n7080__,
    new_new_n7081__, new_new_n7082__, new_new_n7083__, new_new_n7084__,
    new_new_n7085__, new_new_n7086__, new_new_n7087__, new_new_n7088__,
    new_new_n7089__, new_new_n7090__, new_new_n7091__, new_new_n7092__,
    new_new_n7093__, new_new_n7094__, new_new_n7095__, new_new_n7096__,
    new_new_n7097__, new_new_n7098__, new_new_n7099__, new_new_n7100__,
    new_new_n7101__, new_new_n7102__, new_new_n7103__, new_new_n7104__,
    new_new_n7105__, new_new_n7106__, new_new_n7107__, new_new_n7108__,
    new_new_n7109__, new_new_n7110__, new_new_n7111__, new_new_n7112__,
    new_new_n7113__, new_new_n7114__, new_new_n7115__, new_new_n7116__,
    new_new_n7117__, new_new_n7118__, new_new_n7119__, new_new_n7120__,
    new_new_n7121__, new_new_n7122__, new_new_n7123__, new_new_n7124__,
    new_new_n7125__, new_new_n7126__, new_new_n7127__, new_new_n7128__,
    new_new_n7129__, new_new_n7130__, new_new_n7131__, new_new_n7132__,
    new_new_n7133__, new_new_n7134__, new_new_n7135__, new_new_n7136__,
    new_new_n7137__, new_new_n7138__, new_new_n7139__, new_new_n7140__,
    new_new_n7141__, new_new_n7142__, new_new_n7143__, new_new_n7144__,
    new_new_n7145__, new_new_n7146__, new_new_n7147__, new_new_n7148__,
    new_new_n7149__, new_new_n7150__, new_new_n7151__, new_new_n7152__,
    new_new_n7153__, new_new_n7154__, new_new_n7155__, new_new_n7156__,
    new_new_n7157__, new_new_n7158__, new_new_n7159__, new_new_n7160__,
    new_new_n7161__, new_new_n7162__, new_new_n7163__, new_new_n7164__,
    new_new_n7165__, new_new_n7166__, new_new_n7167__, new_new_n7168__,
    new_new_n7169__, new_new_n7170__, new_new_n7171__, new_new_n7172__,
    new_new_n7173__, new_new_n7174__, new_new_n7175__, new_new_n7176__,
    new_new_n7177__, new_new_n7178__, new_new_n7179__, new_new_n7180__,
    new_new_n7181__, new_new_n7182__, new_new_n7183__, new_new_n7184__,
    new_new_n7185__, new_new_n7186__, new_new_n7187__, new_new_n7188__,
    new_new_n7189__, new_new_n7190__, new_new_n7191__, new_new_n7192__,
    new_new_n7193__, new_new_n7194__, new_new_n7195__, new_new_n7196__,
    new_new_n7197__, new_new_n7198__, new_new_n7199__, new_new_n7200__,
    new_new_n7201__, new_new_n7202__, new_new_n7203__, new_new_n7204__,
    new_new_n7205__, new_new_n7206__, new_new_n7207__, new_new_n7208__,
    new_new_n7209__, new_new_n7210__, new_new_n7211__, new_new_n7212__,
    new_new_n7213__, new_new_n7214__, new_new_n7215__, new_new_n7216__,
    new_new_n7217__, new_new_n7218__, new_new_n7219__, new_new_n7220__,
    new_new_n7221__, new_new_n7222__, new_new_n7223__, new_new_n7224__,
    new_new_n7225__, new_new_n7226__, new_new_n7227__, new_new_n7228__,
    new_new_n7229__, new_new_n7230__, new_new_n7231__, new_new_n7232__,
    new_new_n7233__, new_new_n7234__, new_new_n7235__, new_new_n7236__,
    new_new_n7237__, new_new_n7238__, new_new_n7239__, new_new_n7240__,
    new_new_n7241__, new_new_n7242__, new_new_n7243__, new_new_n7244__,
    new_new_n7245__, new_new_n7246__, new_new_n7247__, new_new_n7248__,
    new_new_n7249__, new_new_n7250__, new_new_n7251__, new_new_n7252__,
    new_new_n7253__, new_new_n7254__, new_new_n7256__, new_new_n7257__,
    new_new_n7258__, new_new_n7259__, new_new_n7260__, new_new_n7261__,
    new_new_n7262__, new_new_n7263__, new_new_n7264__, new_new_n7265__,
    new_new_n7266__, new_new_n7267__, new_new_n7268__, new_new_n7269__,
    new_new_n7270__, new_new_n7271__, new_new_n7272__, new_new_n7273__,
    new_new_n7274__, new_new_n7275__, new_new_n7276__, new_new_n7277__,
    new_new_n7278__, new_new_n7279__, new_new_n7280__, new_new_n7281__,
    new_new_n7282__, new_new_n7283__, new_new_n7284__, new_new_n7285__,
    new_new_n7286__, new_new_n7287__, new_new_n7288__, new_new_n7289__,
    new_new_n7290__, new_new_n7291__, new_new_n7292__, new_new_n7293__,
    new_new_n7294__, new_new_n7295__, new_new_n7296__, new_new_n7297__,
    new_new_n7298__, new_new_n7299__, new_new_n7300__, new_new_n7301__,
    new_new_n7302__, new_new_n7303__, new_new_n7304__, new_new_n7305__,
    new_new_n7306__, new_new_n7307__, new_new_n7308__, new_new_n7309__,
    new_new_n7310__, new_new_n7311__, new_new_n7312__, new_new_n7313__,
    new_new_n7314__, new_new_n7315__, new_new_n7316__, new_new_n7317__,
    new_new_n7318__, new_new_n7319__, new_new_n7320__, new_new_n7321__,
    new_new_n7322__, new_new_n7323__, new_new_n7324__, new_new_n7325__,
    new_new_n7326__, new_new_n7327__, new_new_n7328__, new_new_n7329__,
    new_new_n7330__, new_new_n7331__, new_new_n7332__, new_new_n7333__,
    new_new_n7334__, new_new_n7335__, new_new_n7336__, new_new_n7337__,
    new_new_n7338__, new_new_n7339__, new_new_n7340__, new_new_n7341__,
    new_new_n7342__, new_new_n7343__, new_new_n7344__, new_new_n7345__,
    new_new_n7346__, new_new_n7347__, new_new_n7348__, new_new_n7349__,
    new_new_n7350__, new_new_n7351__, new_new_n7352__, new_new_n7353__,
    new_new_n7354__, new_new_n7355__, new_new_n7356__, new_new_n7357__,
    new_new_n7358__, new_new_n7359__, new_new_n7360__, new_new_n7361__,
    new_new_n7362__, new_new_n7363__, new_new_n7364__, new_new_n7365__,
    new_new_n7366__, new_new_n7367__, new_new_n7368__, new_new_n7369__,
    new_new_n7370__, new_new_n7371__, new_new_n7372__, new_new_n7373__,
    new_new_n7374__, new_new_n7375__, new_new_n7376__, new_new_n7377__,
    new_new_n7378__, new_new_n7379__, new_new_n7380__, new_new_n7381__,
    new_new_n7382__, new_new_n7383__, new_new_n7384__, new_new_n7385__,
    new_new_n7386__, new_new_n7387__, new_new_n7388__, new_new_n7389__,
    new_new_n7390__, new_new_n7391__, new_new_n7392__, new_new_n7393__,
    new_new_n7394__, new_new_n7395__, new_new_n7396__, new_new_n7397__,
    new_new_n7398__, new_new_n7399__, new_new_n7400__, new_new_n7401__,
    new_new_n7402__, new_new_n7403__, new_new_n7404__, new_new_n7405__,
    new_new_n7406__, new_new_n7407__, new_new_n7408__, new_new_n7409__,
    new_new_n7410__, new_new_n7411__, new_new_n7412__, new_new_n7413__,
    new_new_n7414__, new_new_n7415__, new_new_n7416__, new_new_n7417__,
    new_new_n7418__, new_new_n7419__, new_new_n7420__, new_new_n7421__,
    new_new_n7422__, new_new_n7423__, new_new_n7424__, new_new_n7425__,
    new_new_n7426__, new_new_n7427__, new_new_n7428__, new_new_n7429__,
    new_new_n7430__, new_new_n7431__, new_new_n7432__, new_new_n7433__,
    new_new_n7434__, new_new_n7435__, new_new_n7436__, new_new_n7437__,
    new_new_n7438__, new_new_n7439__, new_new_n7440__, new_new_n7441__,
    new_new_n7442__, new_new_n7443__, new_new_n7444__, new_new_n7445__,
    new_new_n7446__, new_new_n7447__, new_new_n7448__, new_new_n7449__,
    new_new_n7450__, new_new_n7451__, new_new_n7452__, new_new_n7453__,
    new_new_n7454__, new_new_n7455__, new_new_n7456__, new_new_n7457__,
    new_new_n7458__, new_new_n7459__, new_new_n7460__, new_new_n7461__,
    new_new_n7462__, new_new_n7463__, new_new_n7464__, new_new_n7465__,
    new_new_n7466__, new_new_n7467__, new_new_n7468__, new_new_n7469__,
    new_new_n7470__, new_new_n7471__, new_new_n7472__, new_new_n7473__,
    new_new_n7474__, new_new_n7475__, new_new_n7476__, new_new_n7477__,
    new_new_n7478__, new_new_n7479__, new_new_n7480__, new_new_n7481__,
    new_new_n7482__, new_new_n7483__, new_new_n7484__, new_new_n7485__,
    new_new_n7486__, new_new_n7487__, new_new_n7488__, new_new_n7489__,
    new_new_n7490__, new_new_n7491__, new_new_n7492__, new_new_n7493__,
    new_new_n7494__, new_new_n7495__, new_new_n7496__, new_new_n7497__,
    new_new_n7498__, new_new_n7499__, new_new_n7500__, new_new_n7501__,
    new_new_n7502__, new_new_n7503__, new_new_n7504__, new_new_n7505__,
    new_new_n7506__, new_new_n7507__, new_new_n7508__, new_new_n7509__,
    new_new_n7510__, new_new_n7511__, new_new_n7512__, new_new_n7513__,
    new_new_n7514__, new_new_n7515__, new_new_n7516__, new_new_n7517__,
    new_new_n7518__, new_new_n7519__, new_new_n7520__, new_new_n7521__,
    new_new_n7522__, new_new_n7523__, new_new_n7524__, new_new_n7525__,
    new_new_n7526__, new_new_n7527__, new_new_n7528__, new_new_n7529__,
    new_new_n7530__, new_new_n7531__, new_new_n7532__, new_new_n7533__,
    new_new_n7534__, new_new_n7535__, new_new_n7536__, new_new_n7537__,
    new_new_n7538__, new_new_n7539__, new_new_n7540__, new_new_n7541__,
    new_new_n7542__, new_new_n7543__, new_new_n7544__, new_new_n7545__,
    new_new_n7546__, new_new_n7547__, new_new_n7548__, new_new_n7549__,
    new_new_n7550__, new_new_n7551__, new_new_n7552__, new_new_n7553__,
    new_new_n7554__, new_new_n7555__, new_new_n7556__, new_new_n7557__,
    new_new_n7558__, new_new_n7559__, new_new_n7560__, new_new_n7561__,
    new_new_n7562__, new_new_n7563__, new_new_n7564__, new_new_n7565__,
    new_new_n7566__, new_new_n7567__, new_new_n7568__, new_new_n7569__,
    new_new_n7570__, new_new_n7571__, new_new_n7572__, new_new_n7573__,
    new_new_n7574__, new_new_n7575__, new_new_n7576__, new_new_n7577__,
    new_new_n7578__, new_new_n7579__, new_new_n7580__, new_new_n7581__,
    new_new_n7582__, new_new_n7583__, new_new_n7584__, new_new_n7585__,
    new_new_n7586__, new_new_n7587__, new_new_n7588__, new_new_n7589__,
    new_new_n7590__, new_new_n7591__, new_new_n7592__, new_new_n7593__,
    new_new_n7594__, new_new_n7595__, new_new_n7596__, new_new_n7597__,
    new_new_n7598__, new_new_n7599__, new_new_n7600__, new_new_n7601__,
    new_new_n7602__, new_new_n7603__, new_new_n7604__, new_new_n7605__,
    new_new_n7606__, new_new_n7607__, new_new_n7608__, new_new_n7609__,
    new_new_n7610__, new_new_n7611__, new_new_n7612__, new_new_n7613__,
    new_new_n7614__, new_new_n7615__, new_new_n7616__, new_new_n7617__,
    new_new_n7618__, new_new_n7619__, new_new_n7620__, new_new_n7621__,
    new_new_n7622__, new_new_n7623__, new_new_n7624__, new_new_n7625__,
    new_new_n7626__, new_new_n7627__, new_new_n7628__, new_new_n7629__,
    new_new_n7630__, new_new_n7631__, new_new_n7632__, new_new_n7633__,
    new_new_n7634__, new_new_n7635__, new_new_n7636__, new_new_n7637__,
    new_new_n7638__, new_new_n7639__, new_new_n7640__, new_new_n7641__,
    new_new_n7642__, new_new_n7643__, new_new_n7644__, new_new_n7645__,
    new_new_n7646__, new_new_n7647__, new_new_n7648__, new_new_n7649__,
    new_new_n7650__, new_new_n7651__, new_new_n7652__, new_new_n7653__,
    new_new_n7654__, new_new_n7655__, new_new_n7657__, new_new_n7658__,
    new_new_n7659__, new_new_n7660__, new_new_n7661__, new_new_n7662__,
    new_new_n7663__, new_new_n7664__, new_new_n7665__, new_new_n7666__,
    new_new_n7667__, new_new_n7668__, new_new_n7669__, new_new_n7670__,
    new_new_n7671__, new_new_n7672__, new_new_n7673__, new_new_n7674__,
    new_new_n7675__, new_new_n7676__, new_new_n7677__, new_new_n7678__,
    new_new_n7679__, new_new_n7680__, new_new_n7681__, new_new_n7682__,
    new_new_n7683__, new_new_n7684__, new_new_n7685__, new_new_n7686__,
    new_new_n7687__, new_new_n7688__, new_new_n7689__, new_new_n7690__,
    new_new_n7691__, new_new_n7692__, new_new_n7693__, new_new_n7694__,
    new_new_n7695__, new_new_n7696__, new_new_n7697__, new_new_n7698__,
    new_new_n7699__, new_new_n7700__, new_new_n7701__, new_new_n7702__,
    new_new_n7703__, new_new_n7704__, new_new_n7705__, new_new_n7706__,
    new_new_n7707__, new_new_n7708__, new_new_n7709__, new_new_n7710__,
    new_new_n7711__, new_new_n7712__, new_new_n7713__, new_new_n7714__,
    new_new_n7715__, new_new_n7716__, new_new_n7717__, new_new_n7718__,
    new_new_n7719__, new_new_n7720__, new_new_n7721__, new_new_n7722__,
    new_new_n7723__, new_new_n7724__, new_new_n7725__, new_new_n7726__,
    new_new_n7727__, new_new_n7728__, new_new_n7729__, new_new_n7730__,
    new_new_n7731__, new_new_n7732__, new_new_n7733__, new_new_n7734__,
    new_new_n7735__, new_new_n7736__, new_new_n7737__, new_new_n7738__,
    new_new_n7739__, new_new_n7740__, new_new_n7741__, new_new_n7742__,
    new_new_n7743__, new_new_n7744__, new_new_n7745__, new_new_n7746__,
    new_new_n7747__, new_new_n7748__, new_new_n7749__, new_new_n7750__,
    new_new_n7751__, new_new_n7752__, new_new_n7753__, new_new_n7754__,
    new_new_n7755__, new_new_n7756__, new_new_n7757__, new_new_n7758__,
    new_new_n7759__, new_new_n7760__, new_new_n7761__, new_new_n7762__,
    new_new_n7763__, new_new_n7764__, new_new_n7765__, new_new_n7766__,
    new_new_n7767__, new_new_n7768__, new_new_n7769__, new_new_n7770__,
    new_new_n7771__, new_new_n7772__, new_new_n7773__, new_new_n7774__,
    new_new_n7775__, new_new_n7776__, new_new_n7777__, new_new_n7778__,
    new_new_n7779__, new_new_n7780__, new_new_n7781__, new_new_n7782__,
    new_new_n7783__, new_new_n7784__, new_new_n7785__, new_new_n7786__,
    new_new_n7787__, new_new_n7788__, new_new_n7789__, new_new_n7790__,
    new_new_n7791__, new_new_n7792__, new_new_n7793__, new_new_n7794__,
    new_new_n7795__, new_new_n7796__, new_new_n7797__, new_new_n7798__,
    new_new_n7799__, new_new_n7800__, new_new_n7801__, new_new_n7802__,
    new_new_n7803__, new_new_n7804__, new_new_n7805__, new_new_n7806__,
    new_new_n7807__, new_new_n7808__, new_new_n7809__, new_new_n7810__,
    new_new_n7811__, new_new_n7812__, new_new_n7813__, new_new_n7814__,
    new_new_n7815__, new_new_n7816__, new_new_n7817__, new_new_n7818__,
    new_new_n7819__, new_new_n7820__, new_new_n7821__, new_new_n7822__,
    new_new_n7823__, new_new_n7824__, new_new_n7825__, new_new_n7826__,
    new_new_n7827__, new_new_n7828__, new_new_n7829__, new_new_n7830__,
    new_new_n7831__, new_new_n7832__, new_new_n7833__, new_new_n7834__,
    new_new_n7835__, new_new_n7836__, new_new_n7837__, new_new_n7838__,
    new_new_n7839__, new_new_n7840__, new_new_n7841__, new_new_n7842__,
    new_new_n7843__, new_new_n7844__, new_new_n7845__, new_new_n7846__,
    new_new_n7847__, new_new_n7848__, new_new_n7849__, new_new_n7850__,
    new_new_n7851__, new_new_n7852__, new_new_n7853__, new_new_n7854__,
    new_new_n7855__, new_new_n7856__, new_new_n7857__, new_new_n7858__,
    new_new_n7859__, new_new_n7860__, new_new_n7861__, new_new_n7862__,
    new_new_n7863__, new_new_n7864__, new_new_n7865__, new_new_n7866__,
    new_new_n7867__, new_new_n7868__, new_new_n7869__, new_new_n7870__,
    new_new_n7871__, new_new_n7872__, new_new_n7873__, new_new_n7874__,
    new_new_n7875__, new_new_n7876__, new_new_n7877__, new_new_n7878__,
    new_new_n7879__, new_new_n7880__, new_new_n7881__, new_new_n7882__,
    new_new_n7883__, new_new_n7884__, new_new_n7885__, new_new_n7886__,
    new_new_n7887__, new_new_n7888__, new_new_n7889__, new_new_n7890__,
    new_new_n7891__, new_new_n7892__, new_new_n7893__, new_new_n7894__,
    new_new_n7895__, new_new_n7896__, new_new_n7897__, new_new_n7898__,
    new_new_n7899__, new_new_n7900__, new_new_n7901__, new_new_n7902__,
    new_new_n7903__, new_new_n7904__, new_new_n7905__, new_new_n7906__,
    new_new_n7907__, new_new_n7908__, new_new_n7909__, new_new_n7910__,
    new_new_n7911__, new_new_n7912__, new_new_n7913__, new_new_n7914__,
    new_new_n7915__, new_new_n7916__, new_new_n7917__, new_new_n7918__,
    new_new_n7919__, new_new_n7920__, new_new_n7921__, new_new_n7922__,
    new_new_n7923__, new_new_n7924__, new_new_n7925__, new_new_n7926__,
    new_new_n7927__, new_new_n7928__, new_new_n7929__, new_new_n7930__,
    new_new_n7931__, new_new_n7932__, new_new_n7933__, new_new_n7934__,
    new_new_n7935__, new_new_n7936__, new_new_n7937__, new_new_n7938__,
    new_new_n7939__, new_new_n7940__, new_new_n7941__, new_new_n7942__,
    new_new_n7943__, new_new_n7944__, new_new_n7945__, new_new_n7946__,
    new_new_n7947__, new_new_n7948__, new_new_n7949__, new_new_n7950__,
    new_new_n7951__, new_new_n7952__, new_new_n7953__, new_new_n7954__,
    new_new_n7955__, new_new_n7956__, new_new_n7957__, new_new_n7958__,
    new_new_n7959__, new_new_n7960__, new_new_n7961__, new_new_n7962__,
    new_new_n7963__, new_new_n7964__, new_new_n7965__, new_new_n7966__,
    new_new_n7967__, new_new_n7968__, new_new_n7969__, new_new_n7970__,
    new_new_n7971__, new_new_n7972__, new_new_n7973__, new_new_n7974__,
    new_new_n7975__, new_new_n7976__, new_new_n7977__, new_new_n7978__,
    new_new_n7979__, new_new_n7980__, new_new_n7981__, new_new_n7982__,
    new_new_n7983__, new_new_n7984__, new_new_n7985__, new_new_n7986__,
    new_new_n7987__, new_new_n7988__, new_new_n7989__, new_new_n7990__,
    new_new_n7991__, new_new_n7992__, new_new_n7993__, new_new_n7994__,
    new_new_n7995__, new_new_n7996__, new_new_n7997__, new_new_n7998__,
    new_new_n7999__, new_new_n8000__, new_new_n8001__, new_new_n8002__,
    new_new_n8003__, new_new_n8004__, new_new_n8005__, new_new_n8006__,
    new_new_n8007__, new_new_n8008__, new_new_n8009__, new_new_n8010__,
    new_new_n8011__, new_new_n8012__, new_new_n8013__, new_new_n8014__,
    new_new_n8015__, new_new_n8016__, new_new_n8017__, new_new_n8018__,
    new_new_n8019__, new_new_n8020__, new_new_n8021__, new_new_n8022__,
    new_new_n8023__, new_new_n8024__, new_new_n8025__, new_new_n8026__,
    new_new_n8027__, new_new_n8028__, new_new_n8029__, new_new_n8030__,
    new_new_n8031__, new_new_n8032__, new_new_n8033__, new_new_n8034__,
    new_new_n8035__, new_new_n8036__, new_new_n8037__, new_new_n8038__,
    new_new_n8039__, new_new_n8040__, new_new_n8041__, new_new_n8042__,
    new_new_n8043__, new_new_n8044__, new_new_n8045__, new_new_n8046__,
    new_new_n8047__, new_new_n8048__, new_new_n8049__, new_new_n8050__,
    new_new_n8051__, new_new_n8052__, new_new_n8053__, new_new_n8054__,
    new_new_n8055__, new_new_n8056__, new_new_n8057__, new_new_n8058__,
    new_new_n8059__, new_new_n8060__, new_new_n8061__, new_new_n8063__,
    new_new_n8064__, new_new_n8065__, new_new_n8066__, new_new_n8067__,
    new_new_n8068__, new_new_n8069__, new_new_n8070__, new_new_n8071__,
    new_new_n8072__, new_new_n8073__, new_new_n8074__, new_new_n8075__,
    new_new_n8076__, new_new_n8077__, new_new_n8078__, new_new_n8079__,
    new_new_n8080__, new_new_n8081__, new_new_n8082__, new_new_n8083__,
    new_new_n8084__, new_new_n8085__, new_new_n8086__, new_new_n8087__,
    new_new_n8088__, new_new_n8089__, new_new_n8090__, new_new_n8091__,
    new_new_n8092__, new_new_n8093__, new_new_n8094__, new_new_n8095__,
    new_new_n8096__, new_new_n8097__, new_new_n8098__, new_new_n8099__,
    new_new_n8100__, new_new_n8101__, new_new_n8102__, new_new_n8103__,
    new_new_n8104__, new_new_n8105__, new_new_n8106__, new_new_n8107__,
    new_new_n8108__, new_new_n8109__, new_new_n8110__, new_new_n8111__,
    new_new_n8112__, new_new_n8113__, new_new_n8114__, new_new_n8115__,
    new_new_n8116__, new_new_n8117__, new_new_n8118__, new_new_n8119__,
    new_new_n8120__, new_new_n8121__, new_new_n8122__, new_new_n8123__,
    new_new_n8124__, new_new_n8125__, new_new_n8126__, new_new_n8127__,
    new_new_n8128__, new_new_n8129__, new_new_n8130__, new_new_n8131__,
    new_new_n8132__, new_new_n8133__, new_new_n8134__, new_new_n8135__,
    new_new_n8136__, new_new_n8137__, new_new_n8138__, new_new_n8139__,
    new_new_n8140__, new_new_n8141__, new_new_n8142__, new_new_n8143__,
    new_new_n8144__, new_new_n8145__, new_new_n8146__, new_new_n8147__,
    new_new_n8148__, new_new_n8149__, new_new_n8150__, new_new_n8151__,
    new_new_n8152__, new_new_n8153__, new_new_n8154__, new_new_n8155__,
    new_new_n8156__, new_new_n8157__, new_new_n8158__, new_new_n8159__,
    new_new_n8160__, new_new_n8161__, new_new_n8162__, new_new_n8163__,
    new_new_n8164__, new_new_n8165__, new_new_n8166__, new_new_n8167__,
    new_new_n8168__, new_new_n8169__, new_new_n8170__, new_new_n8171__,
    new_new_n8172__, new_new_n8173__, new_new_n8174__, new_new_n8175__,
    new_new_n8176__, new_new_n8177__, new_new_n8178__, new_new_n8179__,
    new_new_n8180__, new_new_n8181__, new_new_n8182__, new_new_n8183__,
    new_new_n8184__, new_new_n8185__, new_new_n8186__, new_new_n8187__,
    new_new_n8188__, new_new_n8189__, new_new_n8190__, new_new_n8191__,
    new_new_n8192__, new_new_n8193__, new_new_n8194__, new_new_n8195__,
    new_new_n8196__, new_new_n8197__, new_new_n8198__, new_new_n8199__,
    new_new_n8200__, new_new_n8201__, new_new_n8202__, new_new_n8203__,
    new_new_n8204__, new_new_n8205__, new_new_n8206__, new_new_n8207__,
    new_new_n8208__, new_new_n8209__, new_new_n8210__, new_new_n8211__,
    new_new_n8212__, new_new_n8213__, new_new_n8214__, new_new_n8215__,
    new_new_n8216__, new_new_n8217__, new_new_n8218__, new_new_n8219__,
    new_new_n8220__, new_new_n8221__, new_new_n8222__, new_new_n8223__,
    new_new_n8224__, new_new_n8225__, new_new_n8226__, new_new_n8227__,
    new_new_n8228__, new_new_n8229__, new_new_n8230__, new_new_n8231__,
    new_new_n8232__, new_new_n8233__, new_new_n8234__, new_new_n8235__,
    new_new_n8236__, new_new_n8237__, new_new_n8238__, new_new_n8239__,
    new_new_n8240__, new_new_n8241__, new_new_n8242__, new_new_n8243__,
    new_new_n8244__, new_new_n8245__, new_new_n8246__, new_new_n8247__,
    new_new_n8248__, new_new_n8249__, new_new_n8250__, new_new_n8251__,
    new_new_n8252__, new_new_n8253__, new_new_n8254__, new_new_n8255__,
    new_new_n8256__, new_new_n8257__, new_new_n8258__, new_new_n8259__,
    new_new_n8260__, new_new_n8261__, new_new_n8262__, new_new_n8263__,
    new_new_n8264__, new_new_n8265__, new_new_n8266__, new_new_n8267__,
    new_new_n8268__, new_new_n8269__, new_new_n8270__, new_new_n8271__,
    new_new_n8272__, new_new_n8273__, new_new_n8274__, new_new_n8275__,
    new_new_n8276__, new_new_n8277__, new_new_n8278__, new_new_n8279__,
    new_new_n8280__, new_new_n8281__, new_new_n8282__, new_new_n8283__,
    new_new_n8284__, new_new_n8285__, new_new_n8286__, new_new_n8287__,
    new_new_n8288__, new_new_n8289__, new_new_n8290__, new_new_n8291__,
    new_new_n8292__, new_new_n8293__, new_new_n8294__, new_new_n8295__,
    new_new_n8296__, new_new_n8297__, new_new_n8298__, new_new_n8299__,
    new_new_n8300__, new_new_n8301__, new_new_n8302__, new_new_n8303__,
    new_new_n8304__, new_new_n8305__, new_new_n8306__, new_new_n8307__,
    new_new_n8308__, new_new_n8309__, new_new_n8310__, new_new_n8311__,
    new_new_n8312__, new_new_n8313__, new_new_n8314__, new_new_n8315__,
    new_new_n8316__, new_new_n8317__, new_new_n8318__, new_new_n8319__,
    new_new_n8320__, new_new_n8321__, new_new_n8322__, new_new_n8323__,
    new_new_n8324__, new_new_n8325__, new_new_n8326__, new_new_n8327__,
    new_new_n8328__, new_new_n8329__, new_new_n8330__, new_new_n8331__,
    new_new_n8332__, new_new_n8333__, new_new_n8334__, new_new_n8335__,
    new_new_n8336__, new_new_n8337__, new_new_n8338__, new_new_n8339__,
    new_new_n8340__, new_new_n8341__, new_new_n8342__, new_new_n8343__,
    new_new_n8344__, new_new_n8345__, new_new_n8346__, new_new_n8347__,
    new_new_n8348__, new_new_n8349__, new_new_n8350__, new_new_n8351__,
    new_new_n8352__, new_new_n8353__, new_new_n8354__, new_new_n8355__,
    new_new_n8356__, new_new_n8357__, new_new_n8358__, new_new_n8359__,
    new_new_n8360__, new_new_n8361__, new_new_n8362__, new_new_n8363__,
    new_new_n8364__, new_new_n8365__, new_new_n8366__, new_new_n8367__,
    new_new_n8368__, new_new_n8369__, new_new_n8370__, new_new_n8371__,
    new_new_n8372__, new_new_n8373__, new_new_n8374__, new_new_n8375__,
    new_new_n8376__, new_new_n8377__, new_new_n8378__, new_new_n8379__,
    new_new_n8380__, new_new_n8381__, new_new_n8382__, new_new_n8383__,
    new_new_n8384__, new_new_n8385__, new_new_n8386__, new_new_n8387__,
    new_new_n8388__, new_new_n8389__, new_new_n8390__, new_new_n8391__,
    new_new_n8392__, new_new_n8393__, new_new_n8394__, new_new_n8395__,
    new_new_n8396__, new_new_n8397__, new_new_n8398__, new_new_n8399__,
    new_new_n8400__, new_new_n8401__, new_new_n8402__, new_new_n8403__,
    new_new_n8404__, new_new_n8405__, new_new_n8406__, new_new_n8407__,
    new_new_n8408__, new_new_n8409__, new_new_n8410__, new_new_n8411__,
    new_new_n8412__, new_new_n8413__, new_new_n8414__, new_new_n8415__,
    new_new_n8416__, new_new_n8417__, new_new_n8418__, new_new_n8419__,
    new_new_n8420__, new_new_n8421__, new_new_n8422__, new_new_n8423__,
    new_new_n8424__, new_new_n8425__, new_new_n8426__, new_new_n8427__,
    new_new_n8428__, new_new_n8429__, new_new_n8430__, new_new_n8431__,
    new_new_n8432__, new_new_n8433__, new_new_n8434__, new_new_n8435__,
    new_new_n8436__, new_new_n8437__, new_new_n8438__, new_new_n8439__,
    new_new_n8440__, new_new_n8441__, new_new_n8442__, new_new_n8443__,
    new_new_n8444__, new_new_n8445__, new_new_n8446__, new_new_n8447__,
    new_new_n8448__, new_new_n8449__, new_new_n8450__, new_new_n8451__,
    new_new_n8452__, new_new_n8453__, new_new_n8454__, new_new_n8455__,
    new_new_n8456__, new_new_n8457__, new_new_n8458__, new_new_n8459__,
    new_new_n8460__, new_new_n8461__, new_new_n8462__, new_new_n8463__,
    new_new_n8464__, new_new_n8465__, new_new_n8466__, new_new_n8467__,
    new_new_n8468__, new_new_n8469__, new_new_n8470__, new_new_n8471__,
    new_new_n8472__, new_new_n8473__, new_new_n8474__, new_new_n8475__,
    new_new_n8476__, new_new_n8477__, new_new_n8478__, new_new_n8479__,
    new_new_n8480__, new_new_n8481__, new_new_n8482__, new_new_n8483__,
    new_new_n8484__, new_new_n8485__, new_new_n8486__, new_new_n8487__,
    new_new_n8488__, new_new_n8489__, new_new_n8490__, new_new_n8491__,
    new_new_n8492__, new_new_n8493__, new_new_n8495__, new_new_n8496__,
    new_new_n8497__, new_new_n8498__, new_new_n8499__, new_new_n8500__,
    new_new_n8501__, new_new_n8502__, new_new_n8503__, new_new_n8504__,
    new_new_n8505__, new_new_n8506__, new_new_n8507__, new_new_n8508__,
    new_new_n8509__, new_new_n8510__, new_new_n8511__, new_new_n8512__,
    new_new_n8513__, new_new_n8514__, new_new_n8515__, new_new_n8516__,
    new_new_n8517__, new_new_n8518__, new_new_n8519__, new_new_n8520__,
    new_new_n8521__, new_new_n8522__, new_new_n8523__, new_new_n8524__,
    new_new_n8525__, new_new_n8526__, new_new_n8527__, new_new_n8528__,
    new_new_n8529__, new_new_n8530__, new_new_n8531__, new_new_n8532__,
    new_new_n8533__, new_new_n8534__, new_new_n8535__, new_new_n8536__,
    new_new_n8537__, new_new_n8538__, new_new_n8539__, new_new_n8540__,
    new_new_n8541__, new_new_n8542__, new_new_n8543__, new_new_n8544__,
    new_new_n8545__, new_new_n8546__, new_new_n8547__, new_new_n8548__,
    new_new_n8549__, new_new_n8550__, new_new_n8551__, new_new_n8552__,
    new_new_n8553__, new_new_n8554__, new_new_n8555__, new_new_n8556__,
    new_new_n8557__, new_new_n8558__, new_new_n8559__, new_new_n8560__,
    new_new_n8561__, new_new_n8562__, new_new_n8563__, new_new_n8564__,
    new_new_n8565__, new_new_n8566__, new_new_n8567__, new_new_n8568__,
    new_new_n8569__, new_new_n8570__, new_new_n8571__, new_new_n8572__,
    new_new_n8573__, new_new_n8574__, new_new_n8575__, new_new_n8576__,
    new_new_n8577__, new_new_n8578__, new_new_n8579__, new_new_n8580__,
    new_new_n8581__, new_new_n8582__, new_new_n8583__, new_new_n8584__,
    new_new_n8585__, new_new_n8586__, new_new_n8587__, new_new_n8588__,
    new_new_n8589__, new_new_n8590__, new_new_n8591__, new_new_n8592__,
    new_new_n8593__, new_new_n8594__, new_new_n8595__, new_new_n8596__,
    new_new_n8597__, new_new_n8598__, new_new_n8599__, new_new_n8600__,
    new_new_n8601__, new_new_n8602__, new_new_n8603__, new_new_n8604__,
    new_new_n8605__, new_new_n8606__, new_new_n8607__, new_new_n8608__,
    new_new_n8609__, new_new_n8610__, new_new_n8611__, new_new_n8612__,
    new_new_n8613__, new_new_n8614__, new_new_n8615__, new_new_n8616__,
    new_new_n8617__, new_new_n8618__, new_new_n8619__, new_new_n8620__,
    new_new_n8621__, new_new_n8622__, new_new_n8623__, new_new_n8624__,
    new_new_n8625__, new_new_n8626__, new_new_n8627__, new_new_n8628__,
    new_new_n8629__, new_new_n8630__, new_new_n8631__, new_new_n8632__,
    new_new_n8633__, new_new_n8634__, new_new_n8635__, new_new_n8636__,
    new_new_n8637__, new_new_n8638__, new_new_n8639__, new_new_n8640__,
    new_new_n8641__, new_new_n8642__, new_new_n8643__, new_new_n8644__,
    new_new_n8645__, new_new_n8646__, new_new_n8647__, new_new_n8648__,
    new_new_n8649__, new_new_n8650__, new_new_n8651__, new_new_n8652__,
    new_new_n8653__, new_new_n8654__, new_new_n8655__, new_new_n8656__,
    new_new_n8657__, new_new_n8658__, new_new_n8659__, new_new_n8660__,
    new_new_n8661__, new_new_n8662__, new_new_n8663__, new_new_n8664__,
    new_new_n8665__, new_new_n8666__, new_new_n8667__, new_new_n8668__,
    new_new_n8669__, new_new_n8670__, new_new_n8671__, new_new_n8672__,
    new_new_n8673__, new_new_n8674__, new_new_n8675__, new_new_n8676__,
    new_new_n8677__, new_new_n8678__, new_new_n8679__, new_new_n8680__,
    new_new_n8681__, new_new_n8682__, new_new_n8683__, new_new_n8684__,
    new_new_n8685__, new_new_n8686__, new_new_n8687__, new_new_n8688__,
    new_new_n8689__, new_new_n8690__, new_new_n8691__, new_new_n8692__,
    new_new_n8693__, new_new_n8694__, new_new_n8695__, new_new_n8696__,
    new_new_n8697__, new_new_n8698__, new_new_n8699__, new_new_n8700__,
    new_new_n8701__, new_new_n8702__, new_new_n8703__, new_new_n8704__,
    new_new_n8705__, new_new_n8706__, new_new_n8707__, new_new_n8708__,
    new_new_n8709__, new_new_n8710__, new_new_n8711__, new_new_n8712__,
    new_new_n8713__, new_new_n8714__, new_new_n8715__, new_new_n8716__,
    new_new_n8717__, new_new_n8718__, new_new_n8719__, new_new_n8720__,
    new_new_n8721__, new_new_n8722__, new_new_n8723__, new_new_n8724__,
    new_new_n8725__, new_new_n8726__, new_new_n8727__, new_new_n8728__,
    new_new_n8729__, new_new_n8730__, new_new_n8731__, new_new_n8732__,
    new_new_n8733__, new_new_n8734__, new_new_n8735__, new_new_n8736__,
    new_new_n8737__, new_new_n8738__, new_new_n8739__, new_new_n8740__,
    new_new_n8741__, new_new_n8742__, new_new_n8743__, new_new_n8744__,
    new_new_n8745__, new_new_n8746__, new_new_n8747__, new_new_n8748__,
    new_new_n8749__, new_new_n8750__, new_new_n8751__, new_new_n8752__,
    new_new_n8753__, new_new_n8754__, new_new_n8755__, new_new_n8756__,
    new_new_n8757__, new_new_n8758__, new_new_n8759__, new_new_n8760__,
    new_new_n8761__, new_new_n8762__, new_new_n8763__, new_new_n8764__,
    new_new_n8765__, new_new_n8766__, new_new_n8767__, new_new_n8768__,
    new_new_n8769__, new_new_n8770__, new_new_n8771__, new_new_n8772__,
    new_new_n8773__, new_new_n8774__, new_new_n8775__, new_new_n8776__,
    new_new_n8777__, new_new_n8778__, new_new_n8779__, new_new_n8780__,
    new_new_n8781__, new_new_n8782__, new_new_n8783__, new_new_n8784__,
    new_new_n8785__, new_new_n8786__, new_new_n8787__, new_new_n8788__,
    new_new_n8789__, new_new_n8790__, new_new_n8791__, new_new_n8792__,
    new_new_n8793__, new_new_n8794__, new_new_n8795__, new_new_n8796__,
    new_new_n8797__, new_new_n8798__, new_new_n8799__, new_new_n8800__,
    new_new_n8801__, new_new_n8802__, new_new_n8803__, new_new_n8804__,
    new_new_n8805__, new_new_n8806__, new_new_n8807__, new_new_n8808__,
    new_new_n8809__, new_new_n8810__, new_new_n8811__, new_new_n8812__,
    new_new_n8813__, new_new_n8814__, new_new_n8815__, new_new_n8816__,
    new_new_n8817__, new_new_n8818__, new_new_n8819__, new_new_n8820__,
    new_new_n8821__, new_new_n8822__, new_new_n8823__, new_new_n8824__,
    new_new_n8825__, new_new_n8826__, new_new_n8827__, new_new_n8828__,
    new_new_n8829__, new_new_n8830__, new_new_n8831__, new_new_n8832__,
    new_new_n8833__, new_new_n8834__, new_new_n8835__, new_new_n8836__,
    new_new_n8837__, new_new_n8838__, new_new_n8839__, new_new_n8840__,
    new_new_n8841__, new_new_n8842__, new_new_n8843__, new_new_n8844__,
    new_new_n8845__, new_new_n8846__, new_new_n8847__, new_new_n8848__,
    new_new_n8849__, new_new_n8850__, new_new_n8851__, new_new_n8852__,
    new_new_n8853__, new_new_n8854__, new_new_n8855__, new_new_n8856__,
    new_new_n8857__, new_new_n8858__, new_new_n8859__, new_new_n8860__,
    new_new_n8861__, new_new_n8862__, new_new_n8863__, new_new_n8864__,
    new_new_n8865__, new_new_n8866__, new_new_n8867__, new_new_n8868__,
    new_new_n8869__, new_new_n8870__, new_new_n8871__, new_new_n8872__,
    new_new_n8873__, new_new_n8874__, new_new_n8875__, new_new_n8876__,
    new_new_n8877__, new_new_n8878__, new_new_n8879__, new_new_n8880__,
    new_new_n8881__, new_new_n8882__, new_new_n8883__, new_new_n8884__,
    new_new_n8885__, new_new_n8886__, new_new_n8887__, new_new_n8888__,
    new_new_n8889__, new_new_n8890__, new_new_n8891__, new_new_n8892__,
    new_new_n8893__, new_new_n8894__, new_new_n8895__, new_new_n8896__,
    new_new_n8897__, new_new_n8898__, new_new_n8899__, new_new_n8900__,
    new_new_n8901__, new_new_n8902__, new_new_n8903__, new_new_n8904__,
    new_new_n8905__, new_new_n8906__, new_new_n8907__, new_new_n8908__,
    new_new_n8909__, new_new_n8910__, new_new_n8911__, new_new_n8912__,
    new_new_n8913__, new_new_n8914__, new_new_n8915__, new_new_n8916__,
    new_new_n8917__, new_new_n8918__, new_new_n8919__, new_new_n8920__,
    new_new_n8921__, new_new_n8922__, new_new_n8923__, new_new_n8924__,
    new_new_n8925__, new_new_n8926__, new_new_n8927__, new_new_n8929__,
    new_new_n8930__, new_new_n8931__, new_new_n8932__, new_new_n8933__,
    new_new_n8934__, new_new_n8935__, new_new_n8936__, new_new_n8937__,
    new_new_n8938__, new_new_n8939__, new_new_n8940__, new_new_n8941__,
    new_new_n8942__, new_new_n8943__, new_new_n8944__, new_new_n8945__,
    new_new_n8946__, new_new_n8947__, new_new_n8948__, new_new_n8949__,
    new_new_n8950__, new_new_n8951__, new_new_n8952__, new_new_n8953__,
    new_new_n8954__, new_new_n8955__, new_new_n8956__, new_new_n8957__,
    new_new_n8958__, new_new_n8959__, new_new_n8960__, new_new_n8961__,
    new_new_n8962__, new_new_n8963__, new_new_n8964__, new_new_n8965__,
    new_new_n8966__, new_new_n8967__, new_new_n8968__, new_new_n8969__,
    new_new_n8970__, new_new_n8971__, new_new_n8972__, new_new_n8973__,
    new_new_n8974__, new_new_n8975__, new_new_n8976__, new_new_n8977__,
    new_new_n8978__, new_new_n8979__, new_new_n8980__, new_new_n8981__,
    new_new_n8982__, new_new_n8983__, new_new_n8984__, new_new_n8985__,
    new_new_n8986__, new_new_n8987__, new_new_n8988__, new_new_n8989__,
    new_new_n8990__, new_new_n8991__, new_new_n8992__, new_new_n8993__,
    new_new_n8994__, new_new_n8995__, new_new_n8996__, new_new_n8997__,
    new_new_n8998__, new_new_n8999__, new_new_n9000__, new_new_n9001__,
    new_new_n9002__, new_new_n9003__, new_new_n9004__, new_new_n9005__,
    new_new_n9006__, new_new_n9007__, new_new_n9008__, new_new_n9009__,
    new_new_n9010__, new_new_n9011__, new_new_n9012__, new_new_n9013__,
    new_new_n9014__, new_new_n9015__, new_new_n9016__, new_new_n9017__,
    new_new_n9018__, new_new_n9019__, new_new_n9020__, new_new_n9021__,
    new_new_n9022__, new_new_n9023__, new_new_n9024__, new_new_n9025__,
    new_new_n9026__, new_new_n9027__, new_new_n9028__, new_new_n9029__,
    new_new_n9030__, new_new_n9031__, new_new_n9032__, new_new_n9033__,
    new_new_n9034__, new_new_n9035__, new_new_n9036__, new_new_n9037__,
    new_new_n9038__, new_new_n9039__, new_new_n9040__, new_new_n9041__,
    new_new_n9042__, new_new_n9043__, new_new_n9044__, new_new_n9045__,
    new_new_n9046__, new_new_n9047__, new_new_n9048__, new_new_n9049__,
    new_new_n9050__, new_new_n9051__, new_new_n9052__, new_new_n9053__,
    new_new_n9054__, new_new_n9055__, new_new_n9056__, new_new_n9057__,
    new_new_n9058__, new_new_n9059__, new_new_n9060__, new_new_n9061__,
    new_new_n9062__, new_new_n9063__, new_new_n9064__, new_new_n9065__,
    new_new_n9066__, new_new_n9067__, new_new_n9068__, new_new_n9069__,
    new_new_n9070__, new_new_n9071__, new_new_n9072__, new_new_n9073__,
    new_new_n9074__, new_new_n9075__, new_new_n9076__, new_new_n9077__,
    new_new_n9078__, new_new_n9079__, new_new_n9080__, new_new_n9081__,
    new_new_n9082__, new_new_n9083__, new_new_n9084__, new_new_n9085__,
    new_new_n9086__, new_new_n9087__, new_new_n9088__, new_new_n9089__,
    new_new_n9090__, new_new_n9091__, new_new_n9092__, new_new_n9093__,
    new_new_n9094__, new_new_n9095__, new_new_n9096__, new_new_n9097__,
    new_new_n9098__, new_new_n9099__, new_new_n9100__, new_new_n9101__,
    new_new_n9102__, new_new_n9103__, new_new_n9104__, new_new_n9105__,
    new_new_n9106__, new_new_n9107__, new_new_n9108__, new_new_n9109__,
    new_new_n9110__, new_new_n9111__, new_new_n9112__, new_new_n9113__,
    new_new_n9114__, new_new_n9115__, new_new_n9116__, new_new_n9117__,
    new_new_n9118__, new_new_n9119__, new_new_n9120__, new_new_n9121__,
    new_new_n9122__, new_new_n9123__, new_new_n9124__, new_new_n9125__,
    new_new_n9126__, new_new_n9127__, new_new_n9128__, new_new_n9129__,
    new_new_n9130__, new_new_n9131__, new_new_n9132__, new_new_n9133__,
    new_new_n9134__, new_new_n9135__, new_new_n9136__, new_new_n9137__,
    new_new_n9138__, new_new_n9139__, new_new_n9140__, new_new_n9141__,
    new_new_n9142__, new_new_n9143__, new_new_n9144__, new_new_n9145__,
    new_new_n9146__, new_new_n9147__, new_new_n9148__, new_new_n9149__,
    new_new_n9150__, new_new_n9151__, new_new_n9152__, new_new_n9153__,
    new_new_n9154__, new_new_n9155__, new_new_n9156__, new_new_n9157__,
    new_new_n9158__, new_new_n9159__, new_new_n9160__, new_new_n9161__,
    new_new_n9162__, new_new_n9163__, new_new_n9164__, new_new_n9165__,
    new_new_n9166__, new_new_n9167__, new_new_n9168__, new_new_n9169__,
    new_new_n9170__, new_new_n9171__, new_new_n9172__, new_new_n9173__,
    new_new_n9174__, new_new_n9175__, new_new_n9176__, new_new_n9177__,
    new_new_n9178__, new_new_n9179__, new_new_n9180__, new_new_n9181__,
    new_new_n9182__, new_new_n9183__, new_new_n9184__, new_new_n9185__,
    new_new_n9186__, new_new_n9187__, new_new_n9188__, new_new_n9189__,
    new_new_n9190__, new_new_n9191__, new_new_n9192__, new_new_n9193__,
    new_new_n9194__, new_new_n9195__, new_new_n9196__, new_new_n9197__,
    new_new_n9198__, new_new_n9199__, new_new_n9200__, new_new_n9201__,
    new_new_n9202__, new_new_n9203__, new_new_n9204__, new_new_n9205__,
    new_new_n9206__, new_new_n9207__, new_new_n9208__, new_new_n9209__,
    new_new_n9210__, new_new_n9211__, new_new_n9212__, new_new_n9213__,
    new_new_n9214__, new_new_n9215__, new_new_n9216__, new_new_n9217__,
    new_new_n9218__, new_new_n9219__, new_new_n9220__, new_new_n9221__,
    new_new_n9222__, new_new_n9223__, new_new_n9224__, new_new_n9225__,
    new_new_n9226__, new_new_n9227__, new_new_n9228__, new_new_n9229__,
    new_new_n9230__, new_new_n9231__, new_new_n9232__, new_new_n9233__,
    new_new_n9234__, new_new_n9235__, new_new_n9236__, new_new_n9237__,
    new_new_n9238__, new_new_n9239__, new_new_n9240__, new_new_n9241__,
    new_new_n9242__, new_new_n9243__, new_new_n9244__, new_new_n9245__,
    new_new_n9246__, new_new_n9247__, new_new_n9248__, new_new_n9249__,
    new_new_n9250__, new_new_n9251__, new_new_n9252__, new_new_n9253__,
    new_new_n9254__, new_new_n9255__, new_new_n9256__, new_new_n9257__,
    new_new_n9258__, new_new_n9259__, new_new_n9260__, new_new_n9261__,
    new_new_n9262__, new_new_n9263__, new_new_n9264__, new_new_n9265__,
    new_new_n9266__, new_new_n9267__, new_new_n9268__, new_new_n9269__,
    new_new_n9270__, new_new_n9271__, new_new_n9272__, new_new_n9273__,
    new_new_n9274__, new_new_n9275__, new_new_n9276__, new_new_n9277__,
    new_new_n9278__, new_new_n9279__, new_new_n9280__, new_new_n9281__,
    new_new_n9282__, new_new_n9283__, new_new_n9284__, new_new_n9285__,
    new_new_n9286__, new_new_n9287__, new_new_n9288__, new_new_n9289__,
    new_new_n9290__, new_new_n9291__, new_new_n9292__, new_new_n9293__,
    new_new_n9294__, new_new_n9295__, new_new_n9296__, new_new_n9297__,
    new_new_n9298__, new_new_n9299__, new_new_n9300__, new_new_n9301__,
    new_new_n9302__, new_new_n9303__, new_new_n9304__, new_new_n9305__,
    new_new_n9306__, new_new_n9307__, new_new_n9308__, new_new_n9309__,
    new_new_n9310__, new_new_n9311__, new_new_n9312__, new_new_n9313__,
    new_new_n9314__, new_new_n9315__, new_new_n9316__, new_new_n9317__,
    new_new_n9318__, new_new_n9319__, new_new_n9320__, new_new_n9321__,
    new_new_n9322__, new_new_n9323__, new_new_n9324__, new_new_n9325__,
    new_new_n9326__, new_new_n9327__, new_new_n9328__, new_new_n9329__,
    new_new_n9330__, new_new_n9331__, new_new_n9332__, new_new_n9333__,
    new_new_n9334__, new_new_n9335__, new_new_n9336__, new_new_n9337__,
    new_new_n9338__, new_new_n9339__, new_new_n9340__, new_new_n9341__,
    new_new_n9342__, new_new_n9343__, new_new_n9344__, new_new_n9345__,
    new_new_n9346__, new_new_n9347__, new_new_n9348__, new_new_n9349__,
    new_new_n9350__, new_new_n9351__, new_new_n9352__, new_new_n9353__,
    new_new_n9354__, new_new_n9355__, new_new_n9356__, new_new_n9357__,
    new_new_n9358__, new_new_n9360__, new_new_n9361__, new_new_n9362__,
    new_new_n9363__, new_new_n9364__, new_new_n9365__, new_new_n9366__,
    new_new_n9367__, new_new_n9368__, new_new_n9369__, new_new_n9370__,
    new_new_n9371__, new_new_n9372__, new_new_n9373__, new_new_n9374__,
    new_new_n9375__, new_new_n9376__, new_new_n9377__, new_new_n9378__,
    new_new_n9379__, new_new_n9380__, new_new_n9381__, new_new_n9382__,
    new_new_n9383__, new_new_n9384__, new_new_n9385__, new_new_n9386__,
    new_new_n9387__, new_new_n9388__, new_new_n9389__, new_new_n9390__,
    new_new_n9391__, new_new_n9392__, new_new_n9393__, new_new_n9394__,
    new_new_n9395__, new_new_n9396__, new_new_n9397__, new_new_n9398__,
    new_new_n9399__, new_new_n9400__, new_new_n9401__, new_new_n9402__,
    new_new_n9403__, new_new_n9404__, new_new_n9405__, new_new_n9406__,
    new_new_n9407__, new_new_n9408__, new_new_n9409__, new_new_n9410__,
    new_new_n9411__, new_new_n9412__, new_new_n9413__, new_new_n9414__,
    new_new_n9415__, new_new_n9416__, new_new_n9417__, new_new_n9418__,
    new_new_n9419__, new_new_n9420__, new_new_n9421__, new_new_n9422__,
    new_new_n9423__, new_new_n9424__, new_new_n9425__, new_new_n9426__,
    new_new_n9427__, new_new_n9428__, new_new_n9429__, new_new_n9430__,
    new_new_n9431__, new_new_n9432__, new_new_n9433__, new_new_n9434__,
    new_new_n9435__, new_new_n9436__, new_new_n9437__, new_new_n9438__,
    new_new_n9439__, new_new_n9440__, new_new_n9441__, new_new_n9442__,
    new_new_n9443__, new_new_n9444__, new_new_n9445__, new_new_n9446__,
    new_new_n9447__, new_new_n9448__, new_new_n9449__, new_new_n9450__,
    new_new_n9451__, new_new_n9452__, new_new_n9453__, new_new_n9454__,
    new_new_n9455__, new_new_n9456__, new_new_n9457__, new_new_n9458__,
    new_new_n9459__, new_new_n9460__, new_new_n9461__, new_new_n9462__,
    new_new_n9463__, new_new_n9464__, new_new_n9465__, new_new_n9466__,
    new_new_n9467__, new_new_n9468__, new_new_n9469__, new_new_n9470__,
    new_new_n9471__, new_new_n9472__, new_new_n9473__, new_new_n9474__,
    new_new_n9475__, new_new_n9476__, new_new_n9477__, new_new_n9478__,
    new_new_n9479__, new_new_n9480__, new_new_n9481__, new_new_n9482__,
    new_new_n9483__, new_new_n9484__, new_new_n9485__, new_new_n9486__,
    new_new_n9487__, new_new_n9488__, new_new_n9489__, new_new_n9490__,
    new_new_n9491__, new_new_n9492__, new_new_n9493__, new_new_n9494__,
    new_new_n9495__, new_new_n9496__, new_new_n9497__, new_new_n9498__,
    new_new_n9499__, new_new_n9500__, new_new_n9501__, new_new_n9502__,
    new_new_n9503__, new_new_n9504__, new_new_n9505__, new_new_n9506__,
    new_new_n9507__, new_new_n9508__, new_new_n9509__, new_new_n9510__,
    new_new_n9511__, new_new_n9512__, new_new_n9513__, new_new_n9514__,
    new_new_n9515__, new_new_n9516__, new_new_n9517__, new_new_n9518__,
    new_new_n9519__, new_new_n9520__, new_new_n9521__, new_new_n9522__,
    new_new_n9523__, new_new_n9524__, new_new_n9525__, new_new_n9526__,
    new_new_n9527__, new_new_n9528__, new_new_n9529__, new_new_n9530__,
    new_new_n9531__, new_new_n9532__, new_new_n9533__, new_new_n9534__,
    new_new_n9535__, new_new_n9536__, new_new_n9537__, new_new_n9538__,
    new_new_n9539__, new_new_n9540__, new_new_n9541__, new_new_n9542__,
    new_new_n9543__, new_new_n9544__, new_new_n9545__, new_new_n9546__,
    new_new_n9547__, new_new_n9548__, new_new_n9549__, new_new_n9550__,
    new_new_n9551__, new_new_n9552__, new_new_n9553__, new_new_n9554__,
    new_new_n9555__, new_new_n9556__, new_new_n9557__, new_new_n9558__,
    new_new_n9559__, new_new_n9560__, new_new_n9561__, new_new_n9562__,
    new_new_n9563__, new_new_n9564__, new_new_n9565__, new_new_n9566__,
    new_new_n9567__, new_new_n9568__, new_new_n9569__, new_new_n9570__,
    new_new_n9571__, new_new_n9572__, new_new_n9573__, new_new_n9574__,
    new_new_n9575__, new_new_n9576__, new_new_n9577__, new_new_n9578__,
    new_new_n9579__, new_new_n9580__, new_new_n9581__, new_new_n9582__,
    new_new_n9583__, new_new_n9584__, new_new_n9585__, new_new_n9586__,
    new_new_n9587__, new_new_n9588__, new_new_n9589__, new_new_n9590__,
    new_new_n9591__, new_new_n9592__, new_new_n9593__, new_new_n9594__,
    new_new_n9595__, new_new_n9596__, new_new_n9597__, new_new_n9598__,
    new_new_n9599__, new_new_n9600__, new_new_n9601__, new_new_n9602__,
    new_new_n9603__, new_new_n9604__, new_new_n9605__, new_new_n9606__,
    new_new_n9607__, new_new_n9608__, new_new_n9609__, new_new_n9610__,
    new_new_n9611__, new_new_n9612__, new_new_n9613__, new_new_n9614__,
    new_new_n9615__, new_new_n9616__, new_new_n9617__, new_new_n9618__,
    new_new_n9619__, new_new_n9620__, new_new_n9621__, new_new_n9622__,
    new_new_n9623__, new_new_n9624__, new_new_n9625__, new_new_n9626__,
    new_new_n9627__, new_new_n9628__, new_new_n9629__, new_new_n9630__,
    new_new_n9631__, new_new_n9632__, new_new_n9633__, new_new_n9634__,
    new_new_n9635__, new_new_n9636__, new_new_n9637__, new_new_n9638__,
    new_new_n9639__, new_new_n9640__, new_new_n9641__, new_new_n9642__,
    new_new_n9643__, new_new_n9644__, new_new_n9645__, new_new_n9646__,
    new_new_n9647__, new_new_n9648__, new_new_n9649__, new_new_n9650__,
    new_new_n9651__, new_new_n9652__, new_new_n9653__, new_new_n9654__,
    new_new_n9655__, new_new_n9656__, new_new_n9657__, new_new_n9658__,
    new_new_n9659__, new_new_n9660__, new_new_n9661__, new_new_n9662__,
    new_new_n9663__, new_new_n9664__, new_new_n9665__, new_new_n9666__,
    new_new_n9667__, new_new_n9668__, new_new_n9669__, new_new_n9670__,
    new_new_n9671__, new_new_n9672__, new_new_n9673__, new_new_n9674__,
    new_new_n9675__, new_new_n9676__, new_new_n9677__, new_new_n9678__,
    new_new_n9679__, new_new_n9680__, new_new_n9681__, new_new_n9682__,
    new_new_n9683__, new_new_n9684__, new_new_n9685__, new_new_n9686__,
    new_new_n9687__, new_new_n9688__, new_new_n9689__, new_new_n9690__,
    new_new_n9691__, new_new_n9692__, new_new_n9693__, new_new_n9694__,
    new_new_n9695__, new_new_n9696__, new_new_n9697__, new_new_n9698__,
    new_new_n9699__, new_new_n9700__, new_new_n9701__, new_new_n9702__,
    new_new_n9703__, new_new_n9704__, new_new_n9705__, new_new_n9706__,
    new_new_n9707__, new_new_n9708__, new_new_n9709__, new_new_n9710__,
    new_new_n9711__, new_new_n9712__, new_new_n9713__, new_new_n9714__,
    new_new_n9715__, new_new_n9716__, new_new_n9717__, new_new_n9718__,
    new_new_n9719__, new_new_n9720__, new_new_n9721__, new_new_n9722__,
    new_new_n9723__, new_new_n9724__, new_new_n9725__, new_new_n9726__,
    new_new_n9727__, new_new_n9728__, new_new_n9729__, new_new_n9730__,
    new_new_n9731__, new_new_n9732__, new_new_n9733__, new_new_n9734__,
    new_new_n9735__, new_new_n9736__, new_new_n9737__, new_new_n9738__,
    new_new_n9739__, new_new_n9740__, new_new_n9741__, new_new_n9742__,
    new_new_n9743__, new_new_n9744__, new_new_n9745__, new_new_n9746__,
    new_new_n9747__, new_new_n9748__, new_new_n9749__, new_new_n9750__,
    new_new_n9751__, new_new_n9752__, new_new_n9753__, new_new_n9754__,
    new_new_n9755__, new_new_n9756__, new_new_n9757__, new_new_n9758__,
    new_new_n9759__, new_new_n9760__, new_new_n9761__, new_new_n9762__,
    new_new_n9763__, new_new_n9764__, new_new_n9765__, new_new_n9766__,
    new_new_n9767__, new_new_n9768__, new_new_n9769__, new_new_n9770__,
    new_new_n9771__, new_new_n9772__, new_new_n9773__, new_new_n9774__,
    new_new_n9775__, new_new_n9776__, new_new_n9777__, new_new_n9778__,
    new_new_n9779__, new_new_n9780__, new_new_n9781__, new_new_n9782__,
    new_new_n9783__, new_new_n9784__, new_new_n9785__, new_new_n9786__,
    new_new_n9787__, new_new_n9788__, new_new_n9789__, new_new_n9790__,
    new_new_n9791__, new_new_n9792__, new_new_n9793__, new_new_n9794__,
    new_new_n9795__, new_new_n9796__, new_new_n9797__, new_new_n9798__,
    new_new_n9799__, new_new_n9800__, new_new_n9801__, new_new_n9802__,
    new_new_n9803__, new_new_n9804__, new_new_n9805__, new_new_n9806__,
    new_new_n9807__, new_new_n9808__, new_new_n9809__, new_new_n9810__,
    new_new_n9811__, new_new_n9812__, new_new_n9813__, new_new_n9815__,
    new_new_n9816__, new_new_n9817__, new_new_n9818__, new_new_n9819__,
    new_new_n9820__, new_new_n9821__, new_new_n9822__, new_new_n9823__,
    new_new_n9824__, new_new_n9825__, new_new_n9826__, new_new_n9827__,
    new_new_n9828__, new_new_n9829__, new_new_n9830__, new_new_n9831__,
    new_new_n9832__, new_new_n9833__, new_new_n9834__, new_new_n9835__,
    new_new_n9836__, new_new_n9837__, new_new_n9838__, new_new_n9839__,
    new_new_n9840__, new_new_n9841__, new_new_n9842__, new_new_n9843__,
    new_new_n9844__, new_new_n9845__, new_new_n9846__, new_new_n9847__,
    new_new_n9848__, new_new_n9849__, new_new_n9850__, new_new_n9851__,
    new_new_n9852__, new_new_n9853__, new_new_n9854__, new_new_n9855__,
    new_new_n9856__, new_new_n9857__, new_new_n9858__, new_new_n9859__,
    new_new_n9860__, new_new_n9861__, new_new_n9862__, new_new_n9863__,
    new_new_n9864__, new_new_n9865__, new_new_n9866__, new_new_n9867__,
    new_new_n9868__, new_new_n9869__, new_new_n9870__, new_new_n9871__,
    new_new_n9872__, new_new_n9873__, new_new_n9874__, new_new_n9875__,
    new_new_n9876__, new_new_n9877__, new_new_n9878__, new_new_n9879__,
    new_new_n9880__, new_new_n9881__, new_new_n9882__, new_new_n9883__,
    new_new_n9884__, new_new_n9885__, new_new_n9886__, new_new_n9887__,
    new_new_n9888__, new_new_n9889__, new_new_n9890__, new_new_n9891__,
    new_new_n9892__, new_new_n9893__, new_new_n9894__, new_new_n9895__,
    new_new_n9896__, new_new_n9897__, new_new_n9898__, new_new_n9899__,
    new_new_n9900__, new_new_n9901__, new_new_n9902__, new_new_n9903__,
    new_new_n9904__, new_new_n9905__, new_new_n9906__, new_new_n9907__,
    new_new_n9908__, new_new_n9909__, new_new_n9910__, new_new_n9911__,
    new_new_n9912__, new_new_n9913__, new_new_n9914__, new_new_n9915__,
    new_new_n9916__, new_new_n9917__, new_new_n9918__, new_new_n9919__,
    new_new_n9920__, new_new_n9921__, new_new_n9922__, new_new_n9923__,
    new_new_n9924__, new_new_n9925__, new_new_n9926__, new_new_n9927__,
    new_new_n9928__, new_new_n9929__, new_new_n9930__, new_new_n9931__,
    new_new_n9932__, new_new_n9933__, new_new_n9934__, new_new_n9935__,
    new_new_n9936__, new_new_n9937__, new_new_n9938__, new_new_n9939__,
    new_new_n9940__, new_new_n9941__, new_new_n9942__, new_new_n9943__,
    new_new_n9944__, new_new_n9945__, new_new_n9946__, new_new_n9947__,
    new_new_n9948__, new_new_n9949__, new_new_n9950__, new_new_n9951__,
    new_new_n9952__, new_new_n9953__, new_new_n9954__, new_new_n9955__,
    new_new_n9956__, new_new_n9957__, new_new_n9958__, new_new_n9959__,
    new_new_n9960__, new_new_n9961__, new_new_n9962__, new_new_n9963__,
    new_new_n9964__, new_new_n9965__, new_new_n9966__, new_new_n9967__,
    new_new_n9968__, new_new_n9969__, new_new_n9970__, new_new_n9971__,
    new_new_n9972__, new_new_n9973__, new_new_n9974__, new_new_n9975__,
    new_new_n9976__, new_new_n9977__, new_new_n9978__, new_new_n9979__,
    new_new_n9980__, new_new_n9981__, new_new_n9982__, new_new_n9983__,
    new_new_n9984__, new_new_n9985__, new_new_n9986__, new_new_n9987__,
    new_new_n9988__, new_new_n9989__, new_new_n9990__, new_new_n9991__,
    new_new_n9992__, new_new_n9993__, new_new_n9994__, new_new_n9995__,
    new_new_n9996__, new_new_n9997__, new_new_n9998__, new_new_n9999__,
    new_new_n10000__, new_new_n10001__, new_new_n10002__, new_new_n10003__,
    new_new_n10004__, new_new_n10005__, new_new_n10006__, new_new_n10007__,
    new_new_n10008__, new_new_n10009__, new_new_n10010__, new_new_n10011__,
    new_new_n10012__, new_new_n10013__, new_new_n10014__, new_new_n10015__,
    new_new_n10016__, new_new_n10017__, new_new_n10018__, new_new_n10019__,
    new_new_n10020__, new_new_n10021__, new_new_n10022__, new_new_n10023__,
    new_new_n10024__, new_new_n10025__, new_new_n10026__, new_new_n10027__,
    new_new_n10028__, new_new_n10029__, new_new_n10030__, new_new_n10031__,
    new_new_n10032__, new_new_n10033__, new_new_n10034__, new_new_n10035__,
    new_new_n10036__, new_new_n10037__, new_new_n10038__, new_new_n10039__,
    new_new_n10040__, new_new_n10041__, new_new_n10042__, new_new_n10043__,
    new_new_n10044__, new_new_n10045__, new_new_n10046__, new_new_n10047__,
    new_new_n10048__, new_new_n10049__, new_new_n10050__, new_new_n10051__,
    new_new_n10052__, new_new_n10053__, new_new_n10054__, new_new_n10055__,
    new_new_n10056__, new_new_n10057__, new_new_n10058__, new_new_n10059__,
    new_new_n10060__, new_new_n10061__, new_new_n10062__, new_new_n10063__,
    new_new_n10064__, new_new_n10065__, new_new_n10066__, new_new_n10067__,
    new_new_n10068__, new_new_n10069__, new_new_n10070__, new_new_n10071__,
    new_new_n10072__, new_new_n10073__, new_new_n10074__, new_new_n10075__,
    new_new_n10076__, new_new_n10077__, new_new_n10078__, new_new_n10079__,
    new_new_n10080__, new_new_n10081__, new_new_n10082__, new_new_n10083__,
    new_new_n10084__, new_new_n10085__, new_new_n10086__, new_new_n10087__,
    new_new_n10088__, new_new_n10089__, new_new_n10090__, new_new_n10091__,
    new_new_n10092__, new_new_n10093__, new_new_n10094__, new_new_n10095__,
    new_new_n10096__, new_new_n10097__, new_new_n10098__, new_new_n10099__,
    new_new_n10100__, new_new_n10101__, new_new_n10102__, new_new_n10103__,
    new_new_n10104__, new_new_n10105__, new_new_n10106__, new_new_n10107__,
    new_new_n10108__, new_new_n10109__, new_new_n10110__, new_new_n10111__,
    new_new_n10112__, new_new_n10113__, new_new_n10114__, new_new_n10115__,
    new_new_n10116__, new_new_n10117__, new_new_n10118__, new_new_n10119__,
    new_new_n10120__, new_new_n10121__, new_new_n10122__, new_new_n10123__,
    new_new_n10124__, new_new_n10125__, new_new_n10126__, new_new_n10127__,
    new_new_n10128__, new_new_n10129__, new_new_n10130__, new_new_n10131__,
    new_new_n10132__, new_new_n10133__, new_new_n10134__, new_new_n10135__,
    new_new_n10136__, new_new_n10137__, new_new_n10138__, new_new_n10139__,
    new_new_n10140__, new_new_n10141__, new_new_n10142__, new_new_n10143__,
    new_new_n10144__, new_new_n10145__, new_new_n10146__, new_new_n10147__,
    new_new_n10148__, new_new_n10149__, new_new_n10150__, new_new_n10151__,
    new_new_n10152__, new_new_n10153__, new_new_n10154__, new_new_n10155__,
    new_new_n10156__, new_new_n10157__, new_new_n10158__, new_new_n10159__,
    new_new_n10160__, new_new_n10161__, new_new_n10162__, new_new_n10163__,
    new_new_n10164__, new_new_n10165__, new_new_n10166__, new_new_n10167__,
    new_new_n10168__, new_new_n10169__, new_new_n10170__, new_new_n10171__,
    new_new_n10172__, new_new_n10173__, new_new_n10174__, new_new_n10175__,
    new_new_n10176__, new_new_n10177__, new_new_n10178__, new_new_n10179__,
    new_new_n10180__, new_new_n10181__, new_new_n10182__, new_new_n10183__,
    new_new_n10184__, new_new_n10185__, new_new_n10186__, new_new_n10187__,
    new_new_n10188__, new_new_n10189__, new_new_n10190__, new_new_n10191__,
    new_new_n10192__, new_new_n10193__, new_new_n10194__, new_new_n10195__,
    new_new_n10196__, new_new_n10197__, new_new_n10198__, new_new_n10199__,
    new_new_n10200__, new_new_n10201__, new_new_n10202__, new_new_n10203__,
    new_new_n10204__, new_new_n10205__, new_new_n10206__, new_new_n10207__,
    new_new_n10208__, new_new_n10209__, new_new_n10210__, new_new_n10211__,
    new_new_n10212__, new_new_n10213__, new_new_n10214__, new_new_n10215__,
    new_new_n10216__, new_new_n10217__, new_new_n10218__, new_new_n10219__,
    new_new_n10220__, new_new_n10221__, new_new_n10222__, new_new_n10223__,
    new_new_n10224__, new_new_n10225__, new_new_n10226__, new_new_n10227__,
    new_new_n10228__, new_new_n10229__, new_new_n10230__, new_new_n10231__,
    new_new_n10232__, new_new_n10233__, new_new_n10234__, new_new_n10235__,
    new_new_n10236__, new_new_n10237__, new_new_n10238__, new_new_n10239__,
    new_new_n10240__, new_new_n10241__, new_new_n10242__, new_new_n10243__,
    new_new_n10244__, new_new_n10245__, new_new_n10246__, new_new_n10247__,
    new_new_n10248__, new_new_n10249__, new_new_n10250__, new_new_n10251__,
    new_new_n10252__, new_new_n10253__, new_new_n10254__, new_new_n10255__,
    new_new_n10256__, new_new_n10257__, new_new_n10258__, new_new_n10259__,
    new_new_n10260__, new_new_n10261__, new_new_n10262__, new_new_n10263__,
    new_new_n10264__, new_new_n10265__, new_new_n10266__, new_new_n10267__,
    new_new_n10268__, new_new_n10269__, new_new_n10270__, new_new_n10271__,
    new_new_n10272__, new_new_n10273__, new_new_n10274__, new_new_n10275__,
    new_new_n10277__, new_new_n10278__, new_new_n10279__, new_new_n10280__,
    new_new_n10281__, new_new_n10282__, new_new_n10283__, new_new_n10284__,
    new_new_n10285__, new_new_n10286__, new_new_n10287__, new_new_n10288__,
    new_new_n10289__, new_new_n10290__, new_new_n10291__, new_new_n10292__,
    new_new_n10293__, new_new_n10294__, new_new_n10295__, new_new_n10296__,
    new_new_n10297__, new_new_n10298__, new_new_n10299__, new_new_n10300__,
    new_new_n10301__, new_new_n10302__, new_new_n10303__, new_new_n10304__,
    new_new_n10305__, new_new_n10306__, new_new_n10307__, new_new_n10308__,
    new_new_n10309__, new_new_n10310__, new_new_n10311__, new_new_n10312__,
    new_new_n10313__, new_new_n10314__, new_new_n10315__, new_new_n10316__,
    new_new_n10317__, new_new_n10318__, new_new_n10319__, new_new_n10320__,
    new_new_n10321__, new_new_n10322__, new_new_n10323__, new_new_n10324__,
    new_new_n10325__, new_new_n10326__, new_new_n10327__, new_new_n10328__,
    new_new_n10329__, new_new_n10330__, new_new_n10331__, new_new_n10332__,
    new_new_n10333__, new_new_n10334__, new_new_n10335__, new_new_n10336__,
    new_new_n10337__, new_new_n10338__, new_new_n10339__, new_new_n10340__,
    new_new_n10341__, new_new_n10342__, new_new_n10343__, new_new_n10344__,
    new_new_n10345__, new_new_n10346__, new_new_n10347__, new_new_n10348__,
    new_new_n10349__, new_new_n10350__, new_new_n10351__, new_new_n10352__,
    new_new_n10353__, new_new_n10354__, new_new_n10355__, new_new_n10356__,
    new_new_n10357__, new_new_n10358__, new_new_n10359__, new_new_n10360__,
    new_new_n10361__, new_new_n10362__, new_new_n10363__, new_new_n10364__,
    new_new_n10365__, new_new_n10366__, new_new_n10367__, new_new_n10368__,
    new_new_n10369__, new_new_n10370__, new_new_n10371__, new_new_n10372__,
    new_new_n10373__, new_new_n10374__, new_new_n10375__, new_new_n10376__,
    new_new_n10377__, new_new_n10378__, new_new_n10379__, new_new_n10380__,
    new_new_n10381__, new_new_n10382__, new_new_n10383__, new_new_n10384__,
    new_new_n10385__, new_new_n10386__, new_new_n10387__, new_new_n10388__,
    new_new_n10389__, new_new_n10390__, new_new_n10391__, new_new_n10392__,
    new_new_n10393__, new_new_n10394__, new_new_n10395__, new_new_n10396__,
    new_new_n10397__, new_new_n10398__, new_new_n10399__, new_new_n10400__,
    new_new_n10401__, new_new_n10402__, new_new_n10403__, new_new_n10404__,
    new_new_n10405__, new_new_n10406__, new_new_n10407__, new_new_n10408__,
    new_new_n10409__, new_new_n10410__, new_new_n10411__, new_new_n10412__,
    new_new_n10413__, new_new_n10414__, new_new_n10415__, new_new_n10416__,
    new_new_n10417__, new_new_n10418__, new_new_n10419__, new_new_n10420__,
    new_new_n10421__, new_new_n10422__, new_new_n10423__, new_new_n10424__,
    new_new_n10425__, new_new_n10426__, new_new_n10427__, new_new_n10428__,
    new_new_n10429__, new_new_n10430__, new_new_n10431__, new_new_n10432__,
    new_new_n10433__, new_new_n10434__, new_new_n10435__, new_new_n10436__,
    new_new_n10437__, new_new_n10438__, new_new_n10439__, new_new_n10440__,
    new_new_n10441__, new_new_n10442__, new_new_n10443__, new_new_n10444__,
    new_new_n10445__, new_new_n10446__, new_new_n10447__, new_new_n10448__,
    new_new_n10449__, new_new_n10450__, new_new_n10451__, new_new_n10452__,
    new_new_n10453__, new_new_n10454__, new_new_n10455__, new_new_n10456__,
    new_new_n10457__, new_new_n10458__, new_new_n10459__, new_new_n10460__,
    new_new_n10461__, new_new_n10462__, new_new_n10463__, new_new_n10464__,
    new_new_n10465__, new_new_n10466__, new_new_n10467__, new_new_n10468__,
    new_new_n10469__, new_new_n10470__, new_new_n10471__, new_new_n10472__,
    new_new_n10473__, new_new_n10474__, new_new_n10475__, new_new_n10476__,
    new_new_n10477__, new_new_n10478__, new_new_n10479__, new_new_n10480__,
    new_new_n10481__, new_new_n10482__, new_new_n10483__, new_new_n10484__,
    new_new_n10485__, new_new_n10486__, new_new_n10487__, new_new_n10488__,
    new_new_n10489__, new_new_n10490__, new_new_n10491__, new_new_n10492__,
    new_new_n10493__, new_new_n10494__, new_new_n10495__, new_new_n10496__,
    new_new_n10497__, new_new_n10498__, new_new_n10499__, new_new_n10500__,
    new_new_n10501__, new_new_n10502__, new_new_n10503__, new_new_n10504__,
    new_new_n10505__, new_new_n10506__, new_new_n10507__, new_new_n10508__,
    new_new_n10509__, new_new_n10510__, new_new_n10511__, new_new_n10512__,
    new_new_n10513__, new_new_n10514__, new_new_n10515__, new_new_n10516__,
    new_new_n10517__, new_new_n10518__, new_new_n10519__, new_new_n10520__,
    new_new_n10521__, new_new_n10522__, new_new_n10523__, new_new_n10524__,
    new_new_n10525__, new_new_n10526__, new_new_n10527__, new_new_n10528__,
    new_new_n10529__, new_new_n10530__, new_new_n10531__, new_new_n10532__,
    new_new_n10533__, new_new_n10534__, new_new_n10535__, new_new_n10536__,
    new_new_n10537__, new_new_n10538__, new_new_n10539__, new_new_n10540__,
    new_new_n10541__, new_new_n10542__, new_new_n10543__, new_new_n10544__,
    new_new_n10545__, new_new_n10546__, new_new_n10547__, new_new_n10548__,
    new_new_n10549__, new_new_n10550__, new_new_n10551__, new_new_n10552__,
    new_new_n10553__, new_new_n10554__, new_new_n10555__, new_new_n10556__,
    new_new_n10557__, new_new_n10558__, new_new_n10559__, new_new_n10560__,
    new_new_n10561__, new_new_n10562__, new_new_n10563__, new_new_n10564__,
    new_new_n10565__, new_new_n10566__, new_new_n10567__, new_new_n10568__,
    new_new_n10569__, new_new_n10570__, new_new_n10571__, new_new_n10572__,
    new_new_n10573__, new_new_n10574__, new_new_n10575__, new_new_n10576__,
    new_new_n10577__, new_new_n10578__, new_new_n10579__, new_new_n10580__,
    new_new_n10581__, new_new_n10582__, new_new_n10583__, new_new_n10584__,
    new_new_n10585__, new_new_n10586__, new_new_n10587__, new_new_n10588__,
    new_new_n10589__, new_new_n10590__, new_new_n10591__, new_new_n10592__,
    new_new_n10593__, new_new_n10594__, new_new_n10595__, new_new_n10596__,
    new_new_n10597__, new_new_n10598__, new_new_n10599__, new_new_n10600__,
    new_new_n10601__, new_new_n10602__, new_new_n10603__, new_new_n10604__,
    new_new_n10605__, new_new_n10606__, new_new_n10607__, new_new_n10608__,
    new_new_n10609__, new_new_n10610__, new_new_n10611__, new_new_n10612__,
    new_new_n10613__, new_new_n10614__, new_new_n10615__, new_new_n10616__,
    new_new_n10617__, new_new_n10618__, new_new_n10619__, new_new_n10620__,
    new_new_n10621__, new_new_n10622__, new_new_n10623__, new_new_n10624__,
    new_new_n10625__, new_new_n10626__, new_new_n10627__, new_new_n10628__,
    new_new_n10629__, new_new_n10630__, new_new_n10631__, new_new_n10632__,
    new_new_n10633__, new_new_n10634__, new_new_n10635__, new_new_n10636__,
    new_new_n10637__, new_new_n10638__, new_new_n10639__, new_new_n10640__,
    new_new_n10641__, new_new_n10642__, new_new_n10643__, new_new_n10644__,
    new_new_n10645__, new_new_n10646__, new_new_n10647__, new_new_n10648__,
    new_new_n10649__, new_new_n10650__, new_new_n10651__, new_new_n10652__,
    new_new_n10653__, new_new_n10654__, new_new_n10655__, new_new_n10656__,
    new_new_n10657__, new_new_n10658__, new_new_n10659__, new_new_n10660__,
    new_new_n10661__, new_new_n10662__, new_new_n10663__, new_new_n10664__,
    new_new_n10665__, new_new_n10666__, new_new_n10667__, new_new_n10668__,
    new_new_n10669__, new_new_n10670__, new_new_n10671__, new_new_n10672__,
    new_new_n10673__, new_new_n10674__, new_new_n10675__, new_new_n10676__,
    new_new_n10677__, new_new_n10678__, new_new_n10679__, new_new_n10680__,
    new_new_n10681__, new_new_n10682__, new_new_n10683__, new_new_n10684__,
    new_new_n10685__, new_new_n10686__, new_new_n10687__, new_new_n10688__,
    new_new_n10689__, new_new_n10690__, new_new_n10691__, new_new_n10692__,
    new_new_n10693__, new_new_n10694__, new_new_n10695__, new_new_n10696__,
    new_new_n10697__, new_new_n10698__, new_new_n10699__, new_new_n10700__,
    new_new_n10701__, new_new_n10702__, new_new_n10703__, new_new_n10704__,
    new_new_n10705__, new_new_n10706__, new_new_n10707__, new_new_n10708__,
    new_new_n10709__, new_new_n10710__, new_new_n10711__, new_new_n10712__,
    new_new_n10713__, new_new_n10714__, new_new_n10715__, new_new_n10716__,
    new_new_n10717__, new_new_n10718__, new_new_n10719__, new_new_n10720__,
    new_new_n10721__, new_new_n10722__, new_new_n10723__, new_new_n10724__,
    new_new_n10725__, new_new_n10726__, new_new_n10727__, new_new_n10728__,
    new_new_n10729__, new_new_n10730__, new_new_n10731__, new_new_n10732__,
    new_new_n10733__, new_new_n10734__, new_new_n10735__, new_new_n10736__,
    new_new_n10737__, new_new_n10738__, new_new_n10739__, new_new_n10740__,
    new_new_n10741__, new_new_n10742__, new_new_n10743__, new_new_n10744__,
    new_new_n10745__, new_new_n10746__, new_new_n10747__, new_new_n10748__,
    new_new_n10749__, new_new_n10750__, new_new_n10751__, new_new_n10752__,
    new_new_n10753__, new_new_n10754__, new_new_n10755__, new_new_n10756__,
    new_new_n10757__, new_new_n10758__, new_new_n10760__, new_new_n10761__,
    new_new_n10762__, new_new_n10763__, new_new_n10764__, new_new_n10765__,
    new_new_n10766__, new_new_n10767__, new_new_n10768__, new_new_n10769__,
    new_new_n10770__, new_new_n10771__, new_new_n10772__, new_new_n10773__,
    new_new_n10774__, new_new_n10775__, new_new_n10776__, new_new_n10777__,
    new_new_n10778__, new_new_n10779__, new_new_n10780__, new_new_n10781__,
    new_new_n10782__, new_new_n10783__, new_new_n10784__, new_new_n10785__,
    new_new_n10786__, new_new_n10787__, new_new_n10788__, new_new_n10789__,
    new_new_n10790__, new_new_n10791__, new_new_n10792__, new_new_n10793__,
    new_new_n10794__, new_new_n10795__, new_new_n10796__, new_new_n10797__,
    new_new_n10798__, new_new_n10799__, new_new_n10800__, new_new_n10801__,
    new_new_n10802__, new_new_n10803__, new_new_n10804__, new_new_n10805__,
    new_new_n10806__, new_new_n10807__, new_new_n10808__, new_new_n10809__,
    new_new_n10810__, new_new_n10811__, new_new_n10812__, new_new_n10813__,
    new_new_n10814__, new_new_n10815__, new_new_n10816__, new_new_n10817__,
    new_new_n10818__, new_new_n10819__, new_new_n10820__, new_new_n10821__,
    new_new_n10822__, new_new_n10823__, new_new_n10824__, new_new_n10825__,
    new_new_n10826__, new_new_n10827__, new_new_n10828__, new_new_n10829__,
    new_new_n10830__, new_new_n10831__, new_new_n10832__, new_new_n10833__,
    new_new_n10834__, new_new_n10835__, new_new_n10836__, new_new_n10837__,
    new_new_n10838__, new_new_n10839__, new_new_n10840__, new_new_n10841__,
    new_new_n10842__, new_new_n10843__, new_new_n10844__, new_new_n10845__,
    new_new_n10846__, new_new_n10847__, new_new_n10848__, new_new_n10849__,
    new_new_n10850__, new_new_n10851__, new_new_n10852__, new_new_n10853__,
    new_new_n10854__, new_new_n10855__, new_new_n10856__, new_new_n10857__,
    new_new_n10858__, new_new_n10859__, new_new_n10860__, new_new_n10861__,
    new_new_n10862__, new_new_n10863__, new_new_n10864__, new_new_n10865__,
    new_new_n10866__, new_new_n10867__, new_new_n10868__, new_new_n10869__,
    new_new_n10870__, new_new_n10871__, new_new_n10872__, new_new_n10873__,
    new_new_n10874__, new_new_n10875__, new_new_n10876__, new_new_n10877__,
    new_new_n10878__, new_new_n10879__, new_new_n10880__, new_new_n10881__,
    new_new_n10882__, new_new_n10883__, new_new_n10884__, new_new_n10885__,
    new_new_n10886__, new_new_n10887__, new_new_n10888__, new_new_n10889__,
    new_new_n10890__, new_new_n10891__, new_new_n10892__, new_new_n10893__,
    new_new_n10894__, new_new_n10895__, new_new_n10896__, new_new_n10897__,
    new_new_n10898__, new_new_n10899__, new_new_n10900__, new_new_n10901__,
    new_new_n10902__, new_new_n10903__, new_new_n10904__, new_new_n10905__,
    new_new_n10906__, new_new_n10907__, new_new_n10908__, new_new_n10909__,
    new_new_n10910__, new_new_n10911__, new_new_n10912__, new_new_n10913__,
    new_new_n10914__, new_new_n10915__, new_new_n10916__, new_new_n10917__,
    new_new_n10918__, new_new_n10919__, new_new_n10920__, new_new_n10921__,
    new_new_n10922__, new_new_n10923__, new_new_n10924__, new_new_n10925__,
    new_new_n10926__, new_new_n10927__, new_new_n10928__, new_new_n10929__,
    new_new_n10930__, new_new_n10931__, new_new_n10932__, new_new_n10933__,
    new_new_n10934__, new_new_n10935__, new_new_n10936__, new_new_n10937__,
    new_new_n10938__, new_new_n10939__, new_new_n10940__, new_new_n10941__,
    new_new_n10942__, new_new_n10943__, new_new_n10944__, new_new_n10945__,
    new_new_n10946__, new_new_n10947__, new_new_n10948__, new_new_n10949__,
    new_new_n10950__, new_new_n10951__, new_new_n10952__, new_new_n10953__,
    new_new_n10954__, new_new_n10955__, new_new_n10956__, new_new_n10957__,
    new_new_n10958__, new_new_n10959__, new_new_n10960__, new_new_n10961__,
    new_new_n10962__, new_new_n10963__, new_new_n10964__, new_new_n10965__,
    new_new_n10966__, new_new_n10967__, new_new_n10968__, new_new_n10969__,
    new_new_n10970__, new_new_n10971__, new_new_n10972__, new_new_n10973__,
    new_new_n10974__, new_new_n10975__, new_new_n10976__, new_new_n10977__,
    new_new_n10978__, new_new_n10979__, new_new_n10980__, new_new_n10981__,
    new_new_n10982__, new_new_n10983__, new_new_n10984__, new_new_n10985__,
    new_new_n10986__, new_new_n10987__, new_new_n10988__, new_new_n10989__,
    new_new_n10990__, new_new_n10991__, new_new_n10992__, new_new_n10993__,
    new_new_n10994__, new_new_n10995__, new_new_n10996__, new_new_n10997__,
    new_new_n10998__, new_new_n10999__, new_new_n11000__, new_new_n11001__,
    new_new_n11002__, new_new_n11003__, new_new_n11004__, new_new_n11005__,
    new_new_n11006__, new_new_n11007__, new_new_n11008__, new_new_n11009__,
    new_new_n11010__, new_new_n11011__, new_new_n11012__, new_new_n11013__,
    new_new_n11014__, new_new_n11015__, new_new_n11016__, new_new_n11017__,
    new_new_n11018__, new_new_n11019__, new_new_n11020__, new_new_n11021__,
    new_new_n11022__, new_new_n11023__, new_new_n11024__, new_new_n11025__,
    new_new_n11026__, new_new_n11027__, new_new_n11028__, new_new_n11029__,
    new_new_n11030__, new_new_n11031__, new_new_n11032__, new_new_n11033__,
    new_new_n11034__, new_new_n11035__, new_new_n11036__, new_new_n11037__,
    new_new_n11038__, new_new_n11039__, new_new_n11040__, new_new_n11041__,
    new_new_n11042__, new_new_n11043__, new_new_n11044__, new_new_n11045__,
    new_new_n11046__, new_new_n11047__, new_new_n11048__, new_new_n11049__,
    new_new_n11050__, new_new_n11051__, new_new_n11052__, new_new_n11053__,
    new_new_n11054__, new_new_n11055__, new_new_n11056__, new_new_n11057__,
    new_new_n11058__, new_new_n11059__, new_new_n11060__, new_new_n11061__,
    new_new_n11062__, new_new_n11063__, new_new_n11064__, new_new_n11065__,
    new_new_n11066__, new_new_n11067__, new_new_n11068__, new_new_n11069__,
    new_new_n11070__, new_new_n11071__, new_new_n11072__, new_new_n11073__,
    new_new_n11074__, new_new_n11075__, new_new_n11076__, new_new_n11077__,
    new_new_n11078__, new_new_n11079__, new_new_n11080__, new_new_n11081__,
    new_new_n11082__, new_new_n11083__, new_new_n11084__, new_new_n11085__,
    new_new_n11086__, new_new_n11087__, new_new_n11088__, new_new_n11089__,
    new_new_n11090__, new_new_n11091__, new_new_n11092__, new_new_n11093__,
    new_new_n11094__, new_new_n11095__, new_new_n11096__, new_new_n11097__,
    new_new_n11098__, new_new_n11099__, new_new_n11100__, new_new_n11101__,
    new_new_n11102__, new_new_n11103__, new_new_n11104__, new_new_n11105__,
    new_new_n11106__, new_new_n11107__, new_new_n11108__, new_new_n11109__,
    new_new_n11110__, new_new_n11111__, new_new_n11112__, new_new_n11113__,
    new_new_n11114__, new_new_n11115__, new_new_n11116__, new_new_n11117__,
    new_new_n11118__, new_new_n11119__, new_new_n11120__, new_new_n11121__,
    new_new_n11122__, new_new_n11123__, new_new_n11124__, new_new_n11125__,
    new_new_n11126__, new_new_n11127__, new_new_n11128__, new_new_n11129__,
    new_new_n11130__, new_new_n11131__, new_new_n11132__, new_new_n11133__,
    new_new_n11134__, new_new_n11135__, new_new_n11136__, new_new_n11137__,
    new_new_n11138__, new_new_n11139__, new_new_n11140__, new_new_n11141__,
    new_new_n11142__, new_new_n11143__, new_new_n11144__, new_new_n11145__,
    new_new_n11146__, new_new_n11147__, new_new_n11148__, new_new_n11149__,
    new_new_n11150__, new_new_n11151__, new_new_n11152__, new_new_n11153__,
    new_new_n11154__, new_new_n11155__, new_new_n11156__, new_new_n11157__,
    new_new_n11158__, new_new_n11159__, new_new_n11160__, new_new_n11161__,
    new_new_n11162__, new_new_n11163__, new_new_n11164__, new_new_n11165__,
    new_new_n11166__, new_new_n11167__, new_new_n11168__, new_new_n11169__,
    new_new_n11170__, new_new_n11171__, new_new_n11172__, new_new_n11173__,
    new_new_n11174__, new_new_n11175__, new_new_n11176__, new_new_n11177__,
    new_new_n11178__, new_new_n11179__, new_new_n11180__, new_new_n11181__,
    new_new_n11182__, new_new_n11183__, new_new_n11184__, new_new_n11185__,
    new_new_n11186__, new_new_n11187__, new_new_n11188__, new_new_n11189__,
    new_new_n11190__, new_new_n11191__, new_new_n11192__, new_new_n11193__,
    new_new_n11194__, new_new_n11195__, new_new_n11196__, new_new_n11197__,
    new_new_n11198__, new_new_n11199__, new_new_n11200__, new_new_n11201__,
    new_new_n11202__, new_new_n11203__, new_new_n11204__, new_new_n11205__,
    new_new_n11206__, new_new_n11207__, new_new_n11208__, new_new_n11209__,
    new_new_n11210__, new_new_n11211__, new_new_n11212__, new_new_n11213__,
    new_new_n11214__, new_new_n11215__, new_new_n11216__, new_new_n11217__,
    new_new_n11218__, new_new_n11219__, new_new_n11220__, new_new_n11221__,
    new_new_n11222__, new_new_n11223__, new_new_n11224__, new_new_n11225__,
    new_new_n11226__, new_new_n11227__, new_new_n11228__, new_new_n11229__,
    new_new_n11230__, new_new_n11231__, new_new_n11232__, new_new_n11233__,
    new_new_n11234__, new_new_n11235__, new_new_n11236__, new_new_n11237__,
    new_new_n11238__, new_new_n11239__, new_new_n11240__, new_new_n11241__,
    new_new_n11242__, new_new_n11243__, new_new_n11244__, new_new_n11245__,
    new_new_n11246__, new_new_n11247__, new_new_n11248__, new_new_n11249__,
    new_new_n11250__, new_new_n11251__, new_new_n11252__, new_new_n11253__,
    new_new_n11254__, new_new_n11255__, new_new_n11256__, new_new_n11257__,
    new_new_n11258__, new_new_n11259__, new_new_n11260__, new_new_n11261__,
    new_new_n11262__, new_new_n11263__, new_new_n11264__, new_new_n11265__,
    new_new_n11266__, new_new_n11267__, new_new_n11268__, new_new_n11269__,
    new_new_n11270__, new_new_n11271__, new_new_n11272__, new_new_n11273__,
    new_new_n11274__, new_new_n11275__, new_new_n11276__, new_new_n11277__,
    new_new_n11278__, new_new_n11279__, new_new_n11280__, new_new_n11281__,
    new_new_n11282__, new_new_n11283__, new_new_n11284__, new_new_n11285__,
    new_new_n11287__, new_new_n11288__, new_new_n11289__, new_new_n11290__,
    new_new_n11291__, new_new_n11292__, new_new_n11293__, new_new_n11294__,
    new_new_n11295__, new_new_n11296__, new_new_n11297__, new_new_n11298__,
    new_new_n11299__, new_new_n11300__, new_new_n11301__, new_new_n11302__,
    new_new_n11303__, new_new_n11304__, new_new_n11305__, new_new_n11306__,
    new_new_n11307__, new_new_n11308__, new_new_n11309__, new_new_n11310__,
    new_new_n11311__, new_new_n11312__, new_new_n11313__, new_new_n11314__,
    new_new_n11315__, new_new_n11316__, new_new_n11317__, new_new_n11318__,
    new_new_n11319__, new_new_n11320__, new_new_n11321__, new_new_n11322__,
    new_new_n11323__, new_new_n11324__, new_new_n11325__, new_new_n11326__,
    new_new_n11327__, new_new_n11328__, new_new_n11329__, new_new_n11330__,
    new_new_n11331__, new_new_n11332__, new_new_n11333__, new_new_n11334__,
    new_new_n11335__, new_new_n11336__, new_new_n11337__, new_new_n11338__,
    new_new_n11339__, new_new_n11340__, new_new_n11341__, new_new_n11342__,
    new_new_n11343__, new_new_n11344__, new_new_n11345__, new_new_n11346__,
    new_new_n11347__, new_new_n11348__, new_new_n11349__, new_new_n11350__,
    new_new_n11351__, new_new_n11352__, new_new_n11353__, new_new_n11354__,
    new_new_n11355__, new_new_n11356__, new_new_n11357__, new_new_n11358__,
    new_new_n11359__, new_new_n11360__, new_new_n11361__, new_new_n11362__,
    new_new_n11363__, new_new_n11364__, new_new_n11365__, new_new_n11366__,
    new_new_n11367__, new_new_n11368__, new_new_n11369__, new_new_n11370__,
    new_new_n11371__, new_new_n11372__, new_new_n11373__, new_new_n11374__,
    new_new_n11375__, new_new_n11376__, new_new_n11377__, new_new_n11378__,
    new_new_n11379__, new_new_n11380__, new_new_n11381__, new_new_n11382__,
    new_new_n11383__, new_new_n11384__, new_new_n11385__, new_new_n11386__,
    new_new_n11387__, new_new_n11388__, new_new_n11389__, new_new_n11390__,
    new_new_n11391__, new_new_n11392__, new_new_n11393__, new_new_n11394__,
    new_new_n11395__, new_new_n11396__, new_new_n11397__, new_new_n11398__,
    new_new_n11399__, new_new_n11400__, new_new_n11401__, new_new_n11402__,
    new_new_n11403__, new_new_n11404__, new_new_n11405__, new_new_n11406__,
    new_new_n11407__, new_new_n11408__, new_new_n11409__, new_new_n11410__,
    new_new_n11411__, new_new_n11412__, new_new_n11413__, new_new_n11414__,
    new_new_n11415__, new_new_n11416__, new_new_n11417__, new_new_n11418__,
    new_new_n11419__, new_new_n11420__, new_new_n11421__, new_new_n11422__,
    new_new_n11423__, new_new_n11424__, new_new_n11425__, new_new_n11426__,
    new_new_n11427__, new_new_n11428__, new_new_n11429__, new_new_n11430__,
    new_new_n11431__, new_new_n11432__, new_new_n11433__, new_new_n11434__,
    new_new_n11435__, new_new_n11436__, new_new_n11437__, new_new_n11438__,
    new_new_n11439__, new_new_n11440__, new_new_n11441__, new_new_n11442__,
    new_new_n11443__, new_new_n11444__, new_new_n11445__, new_new_n11446__,
    new_new_n11447__, new_new_n11448__, new_new_n11449__, new_new_n11450__,
    new_new_n11451__, new_new_n11452__, new_new_n11453__, new_new_n11454__,
    new_new_n11455__, new_new_n11456__, new_new_n11457__, new_new_n11458__,
    new_new_n11459__, new_new_n11460__, new_new_n11461__, new_new_n11462__,
    new_new_n11463__, new_new_n11464__, new_new_n11465__, new_new_n11466__,
    new_new_n11467__, new_new_n11468__, new_new_n11469__, new_new_n11470__,
    new_new_n11471__, new_new_n11472__, new_new_n11473__, new_new_n11474__,
    new_new_n11475__, new_new_n11476__, new_new_n11477__, new_new_n11478__,
    new_new_n11479__, new_new_n11480__, new_new_n11481__, new_new_n11482__,
    new_new_n11483__, new_new_n11484__, new_new_n11485__, new_new_n11486__,
    new_new_n11487__, new_new_n11488__, new_new_n11489__, new_new_n11490__,
    new_new_n11491__, new_new_n11492__, new_new_n11493__, new_new_n11494__,
    new_new_n11495__, new_new_n11496__, new_new_n11497__, new_new_n11498__,
    new_new_n11499__, new_new_n11500__, new_new_n11501__, new_new_n11502__,
    new_new_n11503__, new_new_n11504__, new_new_n11505__, new_new_n11506__,
    new_new_n11507__, new_new_n11508__, new_new_n11509__, new_new_n11510__,
    new_new_n11511__, new_new_n11512__, new_new_n11513__, new_new_n11514__,
    new_new_n11515__, new_new_n11516__, new_new_n11517__, new_new_n11518__,
    new_new_n11519__, new_new_n11520__, new_new_n11521__, new_new_n11522__,
    new_new_n11523__, new_new_n11524__, new_new_n11525__, new_new_n11526__,
    new_new_n11527__, new_new_n11528__, new_new_n11529__, new_new_n11530__,
    new_new_n11531__, new_new_n11532__, new_new_n11533__, new_new_n11534__,
    new_new_n11535__, new_new_n11536__, new_new_n11537__, new_new_n11538__,
    new_new_n11539__, new_new_n11540__, new_new_n11541__, new_new_n11542__,
    new_new_n11543__, new_new_n11544__, new_new_n11545__, new_new_n11546__,
    new_new_n11547__, new_new_n11548__, new_new_n11549__, new_new_n11550__,
    new_new_n11551__, new_new_n11552__, new_new_n11553__, new_new_n11554__,
    new_new_n11555__, new_new_n11556__, new_new_n11557__, new_new_n11558__,
    new_new_n11559__, new_new_n11560__, new_new_n11561__, new_new_n11562__,
    new_new_n11563__, new_new_n11564__, new_new_n11565__, new_new_n11566__,
    new_new_n11567__, new_new_n11568__, new_new_n11569__, new_new_n11570__,
    new_new_n11571__, new_new_n11572__, new_new_n11573__, new_new_n11574__,
    new_new_n11575__, new_new_n11576__, new_new_n11577__, new_new_n11578__,
    new_new_n11579__, new_new_n11580__, new_new_n11581__, new_new_n11582__,
    new_new_n11583__, new_new_n11584__, new_new_n11585__, new_new_n11586__,
    new_new_n11587__, new_new_n11588__, new_new_n11589__, new_new_n11590__,
    new_new_n11591__, new_new_n11592__, new_new_n11593__, new_new_n11594__,
    new_new_n11595__, new_new_n11596__, new_new_n11597__, new_new_n11598__,
    new_new_n11599__, new_new_n11600__, new_new_n11601__, new_new_n11602__,
    new_new_n11603__, new_new_n11604__, new_new_n11605__, new_new_n11606__,
    new_new_n11607__, new_new_n11608__, new_new_n11609__, new_new_n11610__,
    new_new_n11611__, new_new_n11612__, new_new_n11613__, new_new_n11614__,
    new_new_n11615__, new_new_n11616__, new_new_n11617__, new_new_n11618__,
    new_new_n11619__, new_new_n11620__, new_new_n11621__, new_new_n11622__,
    new_new_n11623__, new_new_n11624__, new_new_n11625__, new_new_n11626__,
    new_new_n11627__, new_new_n11628__, new_new_n11629__, new_new_n11630__,
    new_new_n11631__, new_new_n11632__, new_new_n11633__, new_new_n11634__,
    new_new_n11635__, new_new_n11636__, new_new_n11637__, new_new_n11638__,
    new_new_n11639__, new_new_n11640__, new_new_n11641__, new_new_n11642__,
    new_new_n11643__, new_new_n11644__, new_new_n11645__, new_new_n11646__,
    new_new_n11647__, new_new_n11648__, new_new_n11649__, new_new_n11650__,
    new_new_n11651__, new_new_n11652__, new_new_n11653__, new_new_n11654__,
    new_new_n11655__, new_new_n11656__, new_new_n11657__, new_new_n11658__,
    new_new_n11659__, new_new_n11660__, new_new_n11661__, new_new_n11662__,
    new_new_n11663__, new_new_n11664__, new_new_n11665__, new_new_n11666__,
    new_new_n11667__, new_new_n11668__, new_new_n11669__, new_new_n11670__,
    new_new_n11671__, new_new_n11672__, new_new_n11673__, new_new_n11674__,
    new_new_n11675__, new_new_n11676__, new_new_n11677__, new_new_n11678__,
    new_new_n11679__, new_new_n11680__, new_new_n11681__, new_new_n11682__,
    new_new_n11683__, new_new_n11684__, new_new_n11685__, new_new_n11686__,
    new_new_n11687__, new_new_n11688__, new_new_n11689__, new_new_n11690__,
    new_new_n11691__, new_new_n11692__, new_new_n11693__, new_new_n11694__,
    new_new_n11695__, new_new_n11696__, new_new_n11697__, new_new_n11698__,
    new_new_n11699__, new_new_n11700__, new_new_n11701__, new_new_n11702__,
    new_new_n11703__, new_new_n11704__, new_new_n11705__, new_new_n11706__,
    new_new_n11707__, new_new_n11708__, new_new_n11709__, new_new_n11710__,
    new_new_n11711__, new_new_n11712__, new_new_n11713__, new_new_n11714__,
    new_new_n11715__, new_new_n11716__, new_new_n11717__, new_new_n11718__,
    new_new_n11719__, new_new_n11720__, new_new_n11721__, new_new_n11722__,
    new_new_n11723__, new_new_n11724__, new_new_n11725__, new_new_n11726__,
    new_new_n11727__, new_new_n11728__, new_new_n11729__, new_new_n11730__,
    new_new_n11731__, new_new_n11732__, new_new_n11733__, new_new_n11734__,
    new_new_n11735__, new_new_n11736__, new_new_n11737__, new_new_n11738__,
    new_new_n11739__, new_new_n11740__, new_new_n11741__, new_new_n11742__,
    new_new_n11743__, new_new_n11744__, new_new_n11745__, new_new_n11746__,
    new_new_n11747__, new_new_n11748__, new_new_n11749__, new_new_n11750__,
    new_new_n11751__, new_new_n11752__, new_new_n11753__, new_new_n11754__,
    new_new_n11755__, new_new_n11756__, new_new_n11757__, new_new_n11758__,
    new_new_n11759__, new_new_n11760__, new_new_n11761__, new_new_n11762__,
    new_new_n11763__, new_new_n11764__, new_new_n11765__, new_new_n11766__,
    new_new_n11767__, new_new_n11768__, new_new_n11769__, new_new_n11770__,
    new_new_n11771__, new_new_n11772__, new_new_n11773__, new_new_n11774__,
    new_new_n11775__, new_new_n11776__, new_new_n11777__, new_new_n11778__,
    new_new_n11779__, new_new_n11780__, new_new_n11781__, new_new_n11782__,
    new_new_n11783__, new_new_n11784__, new_new_n11785__, new_new_n11786__,
    new_new_n11787__, new_new_n11788__, new_new_n11789__, new_new_n11791__,
    new_new_n11792__, new_new_n11793__, new_new_n11794__, new_new_n11795__,
    new_new_n11796__, new_new_n11797__, new_new_n11798__, new_new_n11799__,
    new_new_n11800__, new_new_n11801__, new_new_n11802__, new_new_n11803__,
    new_new_n11804__, new_new_n11805__, new_new_n11806__, new_new_n11807__,
    new_new_n11808__, new_new_n11809__, new_new_n11810__, new_new_n11811__,
    new_new_n11812__, new_new_n11813__, new_new_n11814__, new_new_n11815__,
    new_new_n11816__, new_new_n11817__, new_new_n11818__, new_new_n11819__,
    new_new_n11820__, new_new_n11821__, new_new_n11822__, new_new_n11823__,
    new_new_n11824__, new_new_n11825__, new_new_n11826__, new_new_n11827__,
    new_new_n11828__, new_new_n11829__, new_new_n11830__, new_new_n11831__,
    new_new_n11832__, new_new_n11833__, new_new_n11834__, new_new_n11835__,
    new_new_n11836__, new_new_n11837__, new_new_n11838__, new_new_n11839__,
    new_new_n11840__, new_new_n11841__, new_new_n11842__, new_new_n11843__,
    new_new_n11844__, new_new_n11845__, new_new_n11846__, new_new_n11847__,
    new_new_n11848__, new_new_n11849__, new_new_n11850__, new_new_n11851__,
    new_new_n11852__, new_new_n11853__, new_new_n11854__, new_new_n11855__,
    new_new_n11856__, new_new_n11857__, new_new_n11858__, new_new_n11859__,
    new_new_n11860__, new_new_n11861__, new_new_n11862__, new_new_n11863__,
    new_new_n11864__, new_new_n11865__, new_new_n11866__, new_new_n11867__,
    new_new_n11868__, new_new_n11869__, new_new_n11870__, new_new_n11871__,
    new_new_n11872__, new_new_n11873__, new_new_n11874__, new_new_n11875__,
    new_new_n11876__, new_new_n11877__, new_new_n11878__, new_new_n11879__,
    new_new_n11880__, new_new_n11881__, new_new_n11882__, new_new_n11883__,
    new_new_n11884__, new_new_n11885__, new_new_n11886__, new_new_n11887__,
    new_new_n11888__, new_new_n11889__, new_new_n11890__, new_new_n11891__,
    new_new_n11892__, new_new_n11893__, new_new_n11894__, new_new_n11895__,
    new_new_n11896__, new_new_n11897__, new_new_n11898__, new_new_n11899__,
    new_new_n11900__, new_new_n11901__, new_new_n11902__, new_new_n11903__,
    new_new_n11904__, new_new_n11905__, new_new_n11906__, new_new_n11907__,
    new_new_n11908__, new_new_n11909__, new_new_n11910__, new_new_n11911__,
    new_new_n11912__, new_new_n11913__, new_new_n11914__, new_new_n11915__,
    new_new_n11916__, new_new_n11917__, new_new_n11918__, new_new_n11919__,
    new_new_n11920__, new_new_n11921__, new_new_n11922__, new_new_n11923__,
    new_new_n11924__, new_new_n11925__, new_new_n11926__, new_new_n11927__,
    new_new_n11928__, new_new_n11929__, new_new_n11930__, new_new_n11931__,
    new_new_n11932__, new_new_n11933__, new_new_n11934__, new_new_n11935__,
    new_new_n11936__, new_new_n11937__, new_new_n11938__, new_new_n11939__,
    new_new_n11940__, new_new_n11941__, new_new_n11942__, new_new_n11943__,
    new_new_n11944__, new_new_n11945__, new_new_n11946__, new_new_n11947__,
    new_new_n11948__, new_new_n11949__, new_new_n11950__, new_new_n11951__,
    new_new_n11952__, new_new_n11953__, new_new_n11954__, new_new_n11955__,
    new_new_n11956__, new_new_n11957__, new_new_n11958__, new_new_n11959__,
    new_new_n11960__, new_new_n11961__, new_new_n11962__, new_new_n11963__,
    new_new_n11964__, new_new_n11965__, new_new_n11966__, new_new_n11967__,
    new_new_n11968__, new_new_n11969__, new_new_n11970__, new_new_n11971__,
    new_new_n11972__, new_new_n11973__, new_new_n11974__, new_new_n11975__,
    new_new_n11976__, new_new_n11977__, new_new_n11978__, new_new_n11979__,
    new_new_n11980__, new_new_n11981__, new_new_n11982__, new_new_n11983__,
    new_new_n11984__, new_new_n11985__, new_new_n11986__, new_new_n11987__,
    new_new_n11988__, new_new_n11989__, new_new_n11990__, new_new_n11991__,
    new_new_n11992__, new_new_n11993__, new_new_n11994__, new_new_n11995__,
    new_new_n11996__, new_new_n11997__, new_new_n11998__, new_new_n11999__,
    new_new_n12000__, new_new_n12001__, new_new_n12002__, new_new_n12003__,
    new_new_n12004__, new_new_n12005__, new_new_n12006__, new_new_n12007__,
    new_new_n12008__, new_new_n12009__, new_new_n12010__, new_new_n12011__,
    new_new_n12012__, new_new_n12013__, new_new_n12014__, new_new_n12015__,
    new_new_n12016__, new_new_n12017__, new_new_n12018__, new_new_n12019__,
    new_new_n12020__, new_new_n12021__, new_new_n12022__, new_new_n12023__,
    new_new_n12024__, new_new_n12025__, new_new_n12026__, new_new_n12027__,
    new_new_n12028__, new_new_n12029__, new_new_n12030__, new_new_n12031__,
    new_new_n12032__, new_new_n12033__, new_new_n12034__, new_new_n12035__,
    new_new_n12036__, new_new_n12037__, new_new_n12038__, new_new_n12039__,
    new_new_n12040__, new_new_n12041__, new_new_n12042__, new_new_n12043__,
    new_new_n12044__, new_new_n12045__, new_new_n12046__, new_new_n12047__,
    new_new_n12048__, new_new_n12049__, new_new_n12050__, new_new_n12051__,
    new_new_n12052__, new_new_n12053__, new_new_n12054__, new_new_n12055__,
    new_new_n12056__, new_new_n12057__, new_new_n12058__, new_new_n12059__,
    new_new_n12060__, new_new_n12061__, new_new_n12062__, new_new_n12063__,
    new_new_n12064__, new_new_n12065__, new_new_n12066__, new_new_n12067__,
    new_new_n12068__, new_new_n12069__, new_new_n12070__, new_new_n12071__,
    new_new_n12072__, new_new_n12073__, new_new_n12074__, new_new_n12075__,
    new_new_n12076__, new_new_n12077__, new_new_n12078__, new_new_n12079__,
    new_new_n12080__, new_new_n12081__, new_new_n12082__, new_new_n12083__,
    new_new_n12084__, new_new_n12085__, new_new_n12086__, new_new_n12087__,
    new_new_n12088__, new_new_n12089__, new_new_n12090__, new_new_n12091__,
    new_new_n12092__, new_new_n12093__, new_new_n12094__, new_new_n12095__,
    new_new_n12096__, new_new_n12097__, new_new_n12098__, new_new_n12099__,
    new_new_n12100__, new_new_n12101__, new_new_n12102__, new_new_n12103__,
    new_new_n12104__, new_new_n12105__, new_new_n12106__, new_new_n12107__,
    new_new_n12108__, new_new_n12109__, new_new_n12110__, new_new_n12111__,
    new_new_n12112__, new_new_n12113__, new_new_n12114__, new_new_n12115__,
    new_new_n12116__, new_new_n12117__, new_new_n12118__, new_new_n12119__,
    new_new_n12120__, new_new_n12121__, new_new_n12122__, new_new_n12123__,
    new_new_n12124__, new_new_n12125__, new_new_n12126__, new_new_n12127__,
    new_new_n12128__, new_new_n12129__, new_new_n12130__, new_new_n12131__,
    new_new_n12132__, new_new_n12133__, new_new_n12134__, new_new_n12135__,
    new_new_n12136__, new_new_n12137__, new_new_n12138__, new_new_n12139__,
    new_new_n12140__, new_new_n12141__, new_new_n12142__, new_new_n12143__,
    new_new_n12144__, new_new_n12145__, new_new_n12146__, new_new_n12147__,
    new_new_n12148__, new_new_n12149__, new_new_n12150__, new_new_n12151__,
    new_new_n12152__, new_new_n12153__, new_new_n12154__, new_new_n12155__,
    new_new_n12156__, new_new_n12157__, new_new_n12158__, new_new_n12159__,
    new_new_n12160__, new_new_n12161__, new_new_n12162__, new_new_n12163__,
    new_new_n12164__, new_new_n12165__, new_new_n12166__, new_new_n12167__,
    new_new_n12168__, new_new_n12169__, new_new_n12170__, new_new_n12171__,
    new_new_n12172__, new_new_n12173__, new_new_n12174__, new_new_n12175__,
    new_new_n12176__, new_new_n12177__, new_new_n12178__, new_new_n12179__,
    new_new_n12180__, new_new_n12181__, new_new_n12182__, new_new_n12183__,
    new_new_n12184__, new_new_n12185__, new_new_n12186__, new_new_n12187__,
    new_new_n12188__, new_new_n12189__, new_new_n12190__, new_new_n12191__,
    new_new_n12192__, new_new_n12193__, new_new_n12194__, new_new_n12195__,
    new_new_n12196__, new_new_n12197__, new_new_n12198__, new_new_n12199__,
    new_new_n12200__, new_new_n12201__, new_new_n12202__, new_new_n12203__,
    new_new_n12204__, new_new_n12205__, new_new_n12206__, new_new_n12207__,
    new_new_n12208__, new_new_n12209__, new_new_n12210__, new_new_n12211__,
    new_new_n12212__, new_new_n12213__, new_new_n12214__, new_new_n12215__,
    new_new_n12216__, new_new_n12217__, new_new_n12218__, new_new_n12219__,
    new_new_n12220__, new_new_n12221__, new_new_n12222__, new_new_n12223__,
    new_new_n12224__, new_new_n12225__, new_new_n12226__, new_new_n12227__,
    new_new_n12228__, new_new_n12229__, new_new_n12230__, new_new_n12231__,
    new_new_n12232__, new_new_n12233__, new_new_n12234__, new_new_n12235__,
    new_new_n12236__, new_new_n12237__, new_new_n12238__, new_new_n12239__,
    new_new_n12240__, new_new_n12241__, new_new_n12242__, new_new_n12243__,
    new_new_n12244__, new_new_n12245__, new_new_n12246__, new_new_n12247__,
    new_new_n12248__, new_new_n12249__, new_new_n12250__, new_new_n12251__,
    new_new_n12252__, new_new_n12253__, new_new_n12254__, new_new_n12255__,
    new_new_n12256__, new_new_n12257__, new_new_n12258__, new_new_n12259__,
    new_new_n12260__, new_new_n12261__, new_new_n12262__, new_new_n12263__,
    new_new_n12264__, new_new_n12265__, new_new_n12266__, new_new_n12267__,
    new_new_n12268__, new_new_n12269__, new_new_n12270__, new_new_n12271__,
    new_new_n12272__, new_new_n12273__, new_new_n12274__, new_new_n12275__,
    new_new_n12276__, new_new_n12277__, new_new_n12278__, new_new_n12279__,
    new_new_n12280__, new_new_n12281__, new_new_n12282__, new_new_n12283__,
    new_new_n12284__, new_new_n12285__, new_new_n12286__, new_new_n12287__,
    new_new_n12288__, new_new_n12289__, new_new_n12290__, new_new_n12291__,
    new_new_n12292__, new_new_n12293__, new_new_n12294__, new_new_n12295__,
    new_new_n12296__, new_new_n12297__, new_new_n12298__, new_new_n12299__,
    new_new_n12300__, new_new_n12301__, new_new_n12302__, new_new_n12303__,
    new_new_n12304__, new_new_n12305__, new_new_n12306__, new_new_n12307__,
    new_new_n12308__, new_new_n12309__, new_new_n12310__, new_new_n12311__,
    new_new_n12312__, new_new_n12313__, new_new_n12314__, new_new_n12315__,
    new_new_n12316__, new_new_n12317__, new_new_n12318__, new_new_n12319__,
    new_new_n12320__, new_new_n12321__, new_new_n12322__, new_new_n12323__,
    new_new_n12324__, new_new_n12325__, new_new_n12326__, new_new_n12327__,
    new_new_n12329__, new_new_n12330__, new_new_n12331__, new_new_n12332__,
    new_new_n12333__, new_new_n12334__, new_new_n12335__, new_new_n12336__,
    new_new_n12337__, new_new_n12338__, new_new_n12339__, new_new_n12340__,
    new_new_n12341__, new_new_n12342__, new_new_n12343__, new_new_n12344__,
    new_new_n12345__, new_new_n12346__, new_new_n12347__, new_new_n12348__,
    new_new_n12349__, new_new_n12350__, new_new_n12351__, new_new_n12352__,
    new_new_n12353__, new_new_n12354__, new_new_n12355__, new_new_n12356__,
    new_new_n12357__, new_new_n12358__, new_new_n12359__, new_new_n12360__,
    new_new_n12361__, new_new_n12362__, new_new_n12363__, new_new_n12364__,
    new_new_n12365__, new_new_n12366__, new_new_n12367__, new_new_n12368__,
    new_new_n12369__, new_new_n12370__, new_new_n12371__, new_new_n12372__,
    new_new_n12373__, new_new_n12374__, new_new_n12375__, new_new_n12376__,
    new_new_n12377__, new_new_n12378__, new_new_n12379__, new_new_n12380__,
    new_new_n12381__, new_new_n12382__, new_new_n12383__, new_new_n12384__,
    new_new_n12385__, new_new_n12386__, new_new_n12387__, new_new_n12388__,
    new_new_n12389__, new_new_n12390__, new_new_n12391__, new_new_n12392__,
    new_new_n12393__, new_new_n12394__, new_new_n12395__, new_new_n12396__,
    new_new_n12397__, new_new_n12398__, new_new_n12399__, new_new_n12400__,
    new_new_n12401__, new_new_n12402__, new_new_n12403__, new_new_n12404__,
    new_new_n12405__, new_new_n12406__, new_new_n12407__, new_new_n12408__,
    new_new_n12409__, new_new_n12410__, new_new_n12411__, new_new_n12412__,
    new_new_n12413__, new_new_n12414__, new_new_n12415__, new_new_n12416__,
    new_new_n12417__, new_new_n12418__, new_new_n12419__, new_new_n12420__,
    new_new_n12421__, new_new_n12422__, new_new_n12423__, new_new_n12424__,
    new_new_n12425__, new_new_n12426__, new_new_n12427__, new_new_n12428__,
    new_new_n12429__, new_new_n12430__, new_new_n12431__, new_new_n12432__,
    new_new_n12433__, new_new_n12434__, new_new_n12435__, new_new_n12436__,
    new_new_n12437__, new_new_n12438__, new_new_n12439__, new_new_n12440__,
    new_new_n12441__, new_new_n12442__, new_new_n12443__, new_new_n12444__,
    new_new_n12445__, new_new_n12446__, new_new_n12447__, new_new_n12448__,
    new_new_n12449__, new_new_n12450__, new_new_n12451__, new_new_n12452__,
    new_new_n12453__, new_new_n12454__, new_new_n12455__, new_new_n12456__,
    new_new_n12457__, new_new_n12458__, new_new_n12459__, new_new_n12460__,
    new_new_n12461__, new_new_n12462__, new_new_n12463__, new_new_n12464__,
    new_new_n12465__, new_new_n12466__, new_new_n12467__, new_new_n12468__,
    new_new_n12469__, new_new_n12470__, new_new_n12471__, new_new_n12472__,
    new_new_n12473__, new_new_n12474__, new_new_n12475__, new_new_n12476__,
    new_new_n12477__, new_new_n12478__, new_new_n12479__, new_new_n12480__,
    new_new_n12481__, new_new_n12482__, new_new_n12483__, new_new_n12484__,
    new_new_n12485__, new_new_n12486__, new_new_n12487__, new_new_n12488__,
    new_new_n12489__, new_new_n12490__, new_new_n12491__, new_new_n12492__,
    new_new_n12493__, new_new_n12494__, new_new_n12495__, new_new_n12496__,
    new_new_n12497__, new_new_n12498__, new_new_n12499__, new_new_n12500__,
    new_new_n12501__, new_new_n12502__, new_new_n12503__, new_new_n12504__,
    new_new_n12505__, new_new_n12506__, new_new_n12507__, new_new_n12508__,
    new_new_n12509__, new_new_n12510__, new_new_n12511__, new_new_n12512__,
    new_new_n12513__, new_new_n12514__, new_new_n12515__, new_new_n12516__,
    new_new_n12517__, new_new_n12518__, new_new_n12519__, new_new_n12520__,
    new_new_n12521__, new_new_n12522__, new_new_n12523__, new_new_n12524__,
    new_new_n12525__, new_new_n12526__, new_new_n12527__, new_new_n12528__,
    new_new_n12529__, new_new_n12530__, new_new_n12531__, new_new_n12532__,
    new_new_n12533__, new_new_n12534__, new_new_n12535__, new_new_n12536__,
    new_new_n12537__, new_new_n12538__, new_new_n12539__, new_new_n12540__,
    new_new_n12541__, new_new_n12542__, new_new_n12543__, new_new_n12544__,
    new_new_n12545__, new_new_n12546__, new_new_n12547__, new_new_n12548__,
    new_new_n12549__, new_new_n12550__, new_new_n12551__, new_new_n12552__,
    new_new_n12553__, new_new_n12554__, new_new_n12555__, new_new_n12556__,
    new_new_n12557__, new_new_n12558__, new_new_n12559__, new_new_n12560__,
    new_new_n12561__, new_new_n12562__, new_new_n12563__, new_new_n12564__,
    new_new_n12565__, new_new_n12566__, new_new_n12567__, new_new_n12568__,
    new_new_n12569__, new_new_n12570__, new_new_n12571__, new_new_n12572__,
    new_new_n12573__, new_new_n12574__, new_new_n12575__, new_new_n12576__,
    new_new_n12577__, new_new_n12578__, new_new_n12579__, new_new_n12580__,
    new_new_n12581__, new_new_n12582__, new_new_n12583__, new_new_n12584__,
    new_new_n12585__, new_new_n12586__, new_new_n12587__, new_new_n12588__,
    new_new_n12589__, new_new_n12590__, new_new_n12591__, new_new_n12592__,
    new_new_n12593__, new_new_n12594__, new_new_n12595__, new_new_n12596__,
    new_new_n12597__, new_new_n12598__, new_new_n12599__, new_new_n12600__,
    new_new_n12601__, new_new_n12602__, new_new_n12603__, new_new_n12604__,
    new_new_n12605__, new_new_n12606__, new_new_n12607__, new_new_n12608__,
    new_new_n12609__, new_new_n12610__, new_new_n12611__, new_new_n12612__,
    new_new_n12613__, new_new_n12614__, new_new_n12615__, new_new_n12616__,
    new_new_n12617__, new_new_n12618__, new_new_n12619__, new_new_n12620__,
    new_new_n12621__, new_new_n12622__, new_new_n12623__, new_new_n12624__,
    new_new_n12625__, new_new_n12626__, new_new_n12627__, new_new_n12628__,
    new_new_n12629__, new_new_n12630__, new_new_n12631__, new_new_n12632__,
    new_new_n12633__, new_new_n12634__, new_new_n12635__, new_new_n12636__,
    new_new_n12637__, new_new_n12638__, new_new_n12639__, new_new_n12640__,
    new_new_n12641__, new_new_n12642__, new_new_n12643__, new_new_n12644__,
    new_new_n12645__, new_new_n12646__, new_new_n12647__, new_new_n12648__,
    new_new_n12649__, new_new_n12650__, new_new_n12651__, new_new_n12652__,
    new_new_n12653__, new_new_n12654__, new_new_n12655__, new_new_n12656__,
    new_new_n12657__, new_new_n12658__, new_new_n12659__, new_new_n12660__,
    new_new_n12661__, new_new_n12662__, new_new_n12663__, new_new_n12664__,
    new_new_n12665__, new_new_n12666__, new_new_n12667__, new_new_n12668__,
    new_new_n12669__, new_new_n12670__, new_new_n12671__, new_new_n12672__,
    new_new_n12673__, new_new_n12674__, new_new_n12675__, new_new_n12676__,
    new_new_n12677__, new_new_n12678__, new_new_n12679__, new_new_n12680__,
    new_new_n12681__, new_new_n12682__, new_new_n12683__, new_new_n12684__,
    new_new_n12685__, new_new_n12686__, new_new_n12687__, new_new_n12688__,
    new_new_n12689__, new_new_n12690__, new_new_n12691__, new_new_n12692__,
    new_new_n12693__, new_new_n12694__, new_new_n12695__, new_new_n12696__,
    new_new_n12697__, new_new_n12698__, new_new_n12699__, new_new_n12700__,
    new_new_n12701__, new_new_n12702__, new_new_n12703__, new_new_n12704__,
    new_new_n12705__, new_new_n12706__, new_new_n12707__, new_new_n12708__,
    new_new_n12709__, new_new_n12710__, new_new_n12711__, new_new_n12712__,
    new_new_n12713__, new_new_n12714__, new_new_n12715__, new_new_n12716__,
    new_new_n12717__, new_new_n12718__, new_new_n12719__, new_new_n12720__,
    new_new_n12721__, new_new_n12722__, new_new_n12723__, new_new_n12724__,
    new_new_n12725__, new_new_n12726__, new_new_n12727__, new_new_n12728__,
    new_new_n12729__, new_new_n12730__, new_new_n12731__, new_new_n12732__,
    new_new_n12733__, new_new_n12734__, new_new_n12735__, new_new_n12736__,
    new_new_n12737__, new_new_n12738__, new_new_n12739__, new_new_n12740__,
    new_new_n12741__, new_new_n12742__, new_new_n12743__, new_new_n12744__,
    new_new_n12745__, new_new_n12746__, new_new_n12747__, new_new_n12748__,
    new_new_n12749__, new_new_n12750__, new_new_n12751__, new_new_n12752__,
    new_new_n12753__, new_new_n12754__, new_new_n12755__, new_new_n12756__,
    new_new_n12757__, new_new_n12758__, new_new_n12759__, new_new_n12760__,
    new_new_n12761__, new_new_n12762__, new_new_n12763__, new_new_n12764__,
    new_new_n12765__, new_new_n12766__, new_new_n12767__, new_new_n12768__,
    new_new_n12769__, new_new_n12770__, new_new_n12771__, new_new_n12772__,
    new_new_n12773__, new_new_n12774__, new_new_n12775__, new_new_n12776__,
    new_new_n12777__, new_new_n12778__, new_new_n12779__, new_new_n12780__,
    new_new_n12781__, new_new_n12782__, new_new_n12783__, new_new_n12784__,
    new_new_n12785__, new_new_n12786__, new_new_n12787__, new_new_n12788__,
    new_new_n12789__, new_new_n12790__, new_new_n12791__, new_new_n12792__,
    new_new_n12793__, new_new_n12794__, new_new_n12795__, new_new_n12796__,
    new_new_n12797__, new_new_n12798__, new_new_n12799__, new_new_n12800__,
    new_new_n12801__, new_new_n12802__, new_new_n12803__, new_new_n12804__,
    new_new_n12805__, new_new_n12806__, new_new_n12807__, new_new_n12808__,
    new_new_n12809__, new_new_n12810__, new_new_n12811__, new_new_n12812__,
    new_new_n12813__, new_new_n12814__, new_new_n12815__, new_new_n12816__,
    new_new_n12817__, new_new_n12818__, new_new_n12819__, new_new_n12820__,
    new_new_n12821__, new_new_n12822__, new_new_n12823__, new_new_n12824__,
    new_new_n12825__, new_new_n12826__, new_new_n12827__, new_new_n12828__,
    new_new_n12829__, new_new_n12830__, new_new_n12831__, new_new_n12832__,
    new_new_n12833__, new_new_n12834__, new_new_n12835__, new_new_n12836__,
    new_new_n12837__, new_new_n12838__, new_new_n12839__, new_new_n12840__,
    new_new_n12841__, new_new_n12842__, new_new_n12843__, new_new_n12844__,
    new_new_n12845__, new_new_n12846__, new_new_n12847__, new_new_n12848__,
    new_new_n12849__, new_new_n12850__, new_new_n12852__, new_new_n12853__,
    new_new_n12854__, new_new_n12855__, new_new_n12856__, new_new_n12857__,
    new_new_n12858__, new_new_n12859__, new_new_n12860__, new_new_n12861__,
    new_new_n12862__, new_new_n12863__, new_new_n12864__, new_new_n12865__,
    new_new_n12866__, new_new_n12867__, new_new_n12868__, new_new_n12869__,
    new_new_n12870__, new_new_n12871__, new_new_n12872__, new_new_n12873__,
    new_new_n12874__, new_new_n12875__, new_new_n12876__, new_new_n12877__,
    new_new_n12878__, new_new_n12879__, new_new_n12880__, new_new_n12881__,
    new_new_n12882__, new_new_n12883__, new_new_n12884__, new_new_n12885__,
    new_new_n12886__, new_new_n12887__, new_new_n12888__, new_new_n12889__,
    new_new_n12890__, new_new_n12891__, new_new_n12892__, new_new_n12893__,
    new_new_n12894__, new_new_n12895__, new_new_n12896__, new_new_n12897__,
    new_new_n12898__, new_new_n12899__, new_new_n12900__, new_new_n12901__,
    new_new_n12902__, new_new_n12903__, new_new_n12904__, new_new_n12905__,
    new_new_n12906__, new_new_n12907__, new_new_n12908__, new_new_n12909__,
    new_new_n12910__, new_new_n12911__, new_new_n12912__, new_new_n12913__,
    new_new_n12914__, new_new_n12915__, new_new_n12916__, new_new_n12917__,
    new_new_n12918__, new_new_n12919__, new_new_n12920__, new_new_n12921__,
    new_new_n12922__, new_new_n12923__, new_new_n12924__, new_new_n12925__,
    new_new_n12926__, new_new_n12927__, new_new_n12928__, new_new_n12929__,
    new_new_n12930__, new_new_n12931__, new_new_n12932__, new_new_n12933__,
    new_new_n12934__, new_new_n12935__, new_new_n12936__, new_new_n12937__,
    new_new_n12938__, new_new_n12939__, new_new_n12940__, new_new_n12941__,
    new_new_n12942__, new_new_n12943__, new_new_n12944__, new_new_n12945__,
    new_new_n12946__, new_new_n12947__, new_new_n12948__, new_new_n12949__,
    new_new_n12950__, new_new_n12951__, new_new_n12952__, new_new_n12953__,
    new_new_n12954__, new_new_n12955__, new_new_n12956__, new_new_n12957__,
    new_new_n12958__, new_new_n12959__, new_new_n12960__, new_new_n12961__,
    new_new_n12962__, new_new_n12963__, new_new_n12964__, new_new_n12965__,
    new_new_n12966__, new_new_n12967__, new_new_n12968__, new_new_n12969__,
    new_new_n12970__, new_new_n12971__, new_new_n12972__, new_new_n12973__,
    new_new_n12974__, new_new_n12975__, new_new_n12976__, new_new_n12977__,
    new_new_n12978__, new_new_n12979__, new_new_n12980__, new_new_n12981__,
    new_new_n12982__, new_new_n12983__, new_new_n12984__, new_new_n12985__,
    new_new_n12986__, new_new_n12987__, new_new_n12988__, new_new_n12989__,
    new_new_n12990__, new_new_n12991__, new_new_n12992__, new_new_n12993__,
    new_new_n12994__, new_new_n12995__, new_new_n12996__, new_new_n12997__,
    new_new_n12998__, new_new_n12999__, new_new_n13000__, new_new_n13001__,
    new_new_n13002__, new_new_n13003__, new_new_n13004__, new_new_n13005__,
    new_new_n13006__, new_new_n13007__, new_new_n13008__, new_new_n13009__,
    new_new_n13010__, new_new_n13011__, new_new_n13012__, new_new_n13013__,
    new_new_n13014__, new_new_n13015__, new_new_n13016__, new_new_n13017__,
    new_new_n13018__, new_new_n13019__, new_new_n13020__, new_new_n13021__,
    new_new_n13022__, new_new_n13023__, new_new_n13024__, new_new_n13025__,
    new_new_n13026__, new_new_n13027__, new_new_n13028__, new_new_n13029__,
    new_new_n13030__, new_new_n13031__, new_new_n13032__, new_new_n13033__,
    new_new_n13034__, new_new_n13035__, new_new_n13036__, new_new_n13037__,
    new_new_n13038__, new_new_n13039__, new_new_n13040__, new_new_n13041__,
    new_new_n13042__, new_new_n13043__, new_new_n13044__, new_new_n13045__,
    new_new_n13046__, new_new_n13047__, new_new_n13048__, new_new_n13049__,
    new_new_n13050__, new_new_n13051__, new_new_n13052__, new_new_n13053__,
    new_new_n13054__, new_new_n13055__, new_new_n13056__, new_new_n13057__,
    new_new_n13058__, new_new_n13059__, new_new_n13060__, new_new_n13061__,
    new_new_n13062__, new_new_n13063__, new_new_n13064__, new_new_n13065__,
    new_new_n13066__, new_new_n13067__, new_new_n13068__, new_new_n13069__,
    new_new_n13070__, new_new_n13071__, new_new_n13072__, new_new_n13073__,
    new_new_n13074__, new_new_n13075__, new_new_n13076__, new_new_n13077__,
    new_new_n13078__, new_new_n13079__, new_new_n13080__, new_new_n13081__,
    new_new_n13082__, new_new_n13083__, new_new_n13084__, new_new_n13085__,
    new_new_n13086__, new_new_n13087__, new_new_n13088__, new_new_n13089__,
    new_new_n13090__, new_new_n13091__, new_new_n13092__, new_new_n13093__,
    new_new_n13094__, new_new_n13095__, new_new_n13096__, new_new_n13097__,
    new_new_n13098__, new_new_n13099__, new_new_n13100__, new_new_n13101__,
    new_new_n13102__, new_new_n13103__, new_new_n13104__, new_new_n13105__,
    new_new_n13106__, new_new_n13107__, new_new_n13108__, new_new_n13109__,
    new_new_n13110__, new_new_n13111__, new_new_n13112__, new_new_n13113__,
    new_new_n13114__, new_new_n13115__, new_new_n13116__, new_new_n13117__,
    new_new_n13118__, new_new_n13119__, new_new_n13120__, new_new_n13121__,
    new_new_n13122__, new_new_n13123__, new_new_n13124__, new_new_n13125__,
    new_new_n13126__, new_new_n13127__, new_new_n13128__, new_new_n13129__,
    new_new_n13130__, new_new_n13131__, new_new_n13132__, new_new_n13133__,
    new_new_n13134__, new_new_n13135__, new_new_n13136__, new_new_n13137__,
    new_new_n13138__, new_new_n13139__, new_new_n13140__, new_new_n13141__,
    new_new_n13142__, new_new_n13143__, new_new_n13144__, new_new_n13145__,
    new_new_n13146__, new_new_n13147__, new_new_n13148__, new_new_n13149__,
    new_new_n13150__, new_new_n13151__, new_new_n13152__, new_new_n13153__,
    new_new_n13154__, new_new_n13155__, new_new_n13156__, new_new_n13157__,
    new_new_n13158__, new_new_n13159__, new_new_n13160__, new_new_n13161__,
    new_new_n13162__, new_new_n13163__, new_new_n13164__, new_new_n13165__,
    new_new_n13166__, new_new_n13167__, new_new_n13168__, new_new_n13169__,
    new_new_n13170__, new_new_n13171__, new_new_n13172__, new_new_n13173__,
    new_new_n13174__, new_new_n13175__, new_new_n13176__, new_new_n13177__,
    new_new_n13178__, new_new_n13179__, new_new_n13180__, new_new_n13181__,
    new_new_n13182__, new_new_n13183__, new_new_n13184__, new_new_n13185__,
    new_new_n13186__, new_new_n13187__, new_new_n13188__, new_new_n13189__,
    new_new_n13190__, new_new_n13191__, new_new_n13192__, new_new_n13193__,
    new_new_n13194__, new_new_n13195__, new_new_n13196__, new_new_n13197__,
    new_new_n13198__, new_new_n13199__, new_new_n13200__, new_new_n13201__,
    new_new_n13202__, new_new_n13203__, new_new_n13204__, new_new_n13205__,
    new_new_n13206__, new_new_n13207__, new_new_n13208__, new_new_n13209__,
    new_new_n13210__, new_new_n13211__, new_new_n13212__, new_new_n13213__,
    new_new_n13214__, new_new_n13215__, new_new_n13216__, new_new_n13217__,
    new_new_n13218__, new_new_n13219__, new_new_n13220__, new_new_n13221__,
    new_new_n13222__, new_new_n13223__, new_new_n13224__, new_new_n13225__,
    new_new_n13226__, new_new_n13227__, new_new_n13228__, new_new_n13229__,
    new_new_n13230__, new_new_n13231__, new_new_n13232__, new_new_n13233__,
    new_new_n13234__, new_new_n13235__, new_new_n13236__, new_new_n13237__,
    new_new_n13238__, new_new_n13239__, new_new_n13240__, new_new_n13241__,
    new_new_n13242__, new_new_n13243__, new_new_n13244__, new_new_n13245__,
    new_new_n13246__, new_new_n13247__, new_new_n13248__, new_new_n13249__,
    new_new_n13250__, new_new_n13251__, new_new_n13252__, new_new_n13253__,
    new_new_n13254__, new_new_n13255__, new_new_n13256__, new_new_n13257__,
    new_new_n13258__, new_new_n13259__, new_new_n13260__, new_new_n13261__,
    new_new_n13262__, new_new_n13263__, new_new_n13264__, new_new_n13265__,
    new_new_n13266__, new_new_n13267__, new_new_n13268__, new_new_n13269__,
    new_new_n13270__, new_new_n13271__, new_new_n13272__, new_new_n13273__,
    new_new_n13274__, new_new_n13275__, new_new_n13276__, new_new_n13277__,
    new_new_n13278__, new_new_n13279__, new_new_n13280__, new_new_n13281__,
    new_new_n13282__, new_new_n13283__, new_new_n13284__, new_new_n13285__,
    new_new_n13286__, new_new_n13287__, new_new_n13288__, new_new_n13289__,
    new_new_n13290__, new_new_n13291__, new_new_n13292__, new_new_n13293__,
    new_new_n13294__, new_new_n13295__, new_new_n13296__, new_new_n13297__,
    new_new_n13298__, new_new_n13299__, new_new_n13300__, new_new_n13301__,
    new_new_n13302__, new_new_n13303__, new_new_n13304__, new_new_n13305__,
    new_new_n13306__, new_new_n13307__, new_new_n13308__, new_new_n13309__,
    new_new_n13310__, new_new_n13311__, new_new_n13312__, new_new_n13313__,
    new_new_n13314__, new_new_n13315__, new_new_n13316__, new_new_n13317__,
    new_new_n13318__, new_new_n13319__, new_new_n13320__, new_new_n13321__,
    new_new_n13322__, new_new_n13323__, new_new_n13324__, new_new_n13325__,
    new_new_n13326__, new_new_n13327__, new_new_n13328__, new_new_n13329__,
    new_new_n13330__, new_new_n13331__, new_new_n13332__, new_new_n13333__,
    new_new_n13334__, new_new_n13335__, new_new_n13336__, new_new_n13337__,
    new_new_n13338__, new_new_n13339__, new_new_n13340__, new_new_n13341__,
    new_new_n13342__, new_new_n13343__, new_new_n13344__, new_new_n13345__,
    new_new_n13346__, new_new_n13347__, new_new_n13348__, new_new_n13349__,
    new_new_n13350__, new_new_n13351__, new_new_n13352__, new_new_n13353__,
    new_new_n13354__, new_new_n13355__, new_new_n13356__, new_new_n13357__,
    new_new_n13358__, new_new_n13359__, new_new_n13360__, new_new_n13361__,
    new_new_n13362__, new_new_n13363__, new_new_n13364__, new_new_n13365__,
    new_new_n13366__, new_new_n13367__, new_new_n13368__, new_new_n13369__,
    new_new_n13370__, new_new_n13371__, new_new_n13372__, new_new_n13373__,
    new_new_n13374__, new_new_n13375__, new_new_n13376__, new_new_n13377__,
    new_new_n13378__, new_new_n13379__, new_new_n13380__, new_new_n13381__,
    new_new_n13382__, new_new_n13383__, new_new_n13384__, new_new_n13386__,
    new_new_n13387__, new_new_n13388__, new_new_n13389__, new_new_n13390__,
    new_new_n13391__, new_new_n13392__, new_new_n13393__, new_new_n13394__,
    new_new_n13395__, new_new_n13396__, new_new_n13397__, new_new_n13398__,
    new_new_n13399__, new_new_n13400__, new_new_n13401__, new_new_n13402__,
    new_new_n13403__, new_new_n13404__, new_new_n13405__, new_new_n13406__,
    new_new_n13407__, new_new_n13408__, new_new_n13409__, new_new_n13410__,
    new_new_n13411__, new_new_n13412__, new_new_n13413__, new_new_n13414__,
    new_new_n13415__, new_new_n13416__, new_new_n13417__, new_new_n13418__,
    new_new_n13419__, new_new_n13420__, new_new_n13421__, new_new_n13422__,
    new_new_n13423__, new_new_n13424__, new_new_n13425__, new_new_n13426__,
    new_new_n13427__, new_new_n13428__, new_new_n13429__, new_new_n13430__,
    new_new_n13431__, new_new_n13432__, new_new_n13433__, new_new_n13434__,
    new_new_n13435__, new_new_n13436__, new_new_n13437__, new_new_n13438__,
    new_new_n13439__, new_new_n13440__, new_new_n13441__, new_new_n13442__,
    new_new_n13443__, new_new_n13444__, new_new_n13445__, new_new_n13446__,
    new_new_n13447__, new_new_n13448__, new_new_n13449__, new_new_n13450__,
    new_new_n13451__, new_new_n13452__, new_new_n13453__, new_new_n13454__,
    new_new_n13455__, new_new_n13456__, new_new_n13457__, new_new_n13458__,
    new_new_n13459__, new_new_n13460__, new_new_n13461__, new_new_n13462__,
    new_new_n13463__, new_new_n13464__, new_new_n13465__, new_new_n13466__,
    new_new_n13467__, new_new_n13468__, new_new_n13469__, new_new_n13470__,
    new_new_n13471__, new_new_n13472__, new_new_n13473__, new_new_n13474__,
    new_new_n13475__, new_new_n13476__, new_new_n13477__, new_new_n13478__,
    new_new_n13479__, new_new_n13480__, new_new_n13481__, new_new_n13482__,
    new_new_n13483__, new_new_n13484__, new_new_n13485__, new_new_n13486__,
    new_new_n13487__, new_new_n13488__, new_new_n13489__, new_new_n13490__,
    new_new_n13491__, new_new_n13492__, new_new_n13493__, new_new_n13494__,
    new_new_n13495__, new_new_n13496__, new_new_n13497__, new_new_n13498__,
    new_new_n13499__, new_new_n13500__, new_new_n13501__, new_new_n13502__,
    new_new_n13503__, new_new_n13504__, new_new_n13505__, new_new_n13506__,
    new_new_n13507__, new_new_n13508__, new_new_n13509__, new_new_n13510__,
    new_new_n13511__, new_new_n13512__, new_new_n13513__, new_new_n13514__,
    new_new_n13515__, new_new_n13516__, new_new_n13517__, new_new_n13518__,
    new_new_n13519__, new_new_n13520__, new_new_n13521__, new_new_n13522__,
    new_new_n13523__, new_new_n13524__, new_new_n13525__, new_new_n13526__,
    new_new_n13527__, new_new_n13528__, new_new_n13529__, new_new_n13530__,
    new_new_n13531__, new_new_n13532__, new_new_n13533__, new_new_n13534__,
    new_new_n13535__, new_new_n13536__, new_new_n13537__, new_new_n13538__,
    new_new_n13539__, new_new_n13540__, new_new_n13541__, new_new_n13542__,
    new_new_n13543__, new_new_n13544__, new_new_n13545__, new_new_n13546__,
    new_new_n13547__, new_new_n13548__, new_new_n13549__, new_new_n13550__,
    new_new_n13551__, new_new_n13552__, new_new_n13553__, new_new_n13554__,
    new_new_n13555__, new_new_n13556__, new_new_n13557__, new_new_n13558__,
    new_new_n13559__, new_new_n13560__, new_new_n13561__, new_new_n13562__,
    new_new_n13563__, new_new_n13564__, new_new_n13565__, new_new_n13566__,
    new_new_n13567__, new_new_n13568__, new_new_n13569__, new_new_n13570__,
    new_new_n13571__, new_new_n13572__, new_new_n13573__, new_new_n13574__,
    new_new_n13575__, new_new_n13576__, new_new_n13577__, new_new_n13578__,
    new_new_n13579__, new_new_n13580__, new_new_n13581__, new_new_n13582__,
    new_new_n13583__, new_new_n13584__, new_new_n13585__, new_new_n13586__,
    new_new_n13587__, new_new_n13588__, new_new_n13589__, new_new_n13590__,
    new_new_n13591__, new_new_n13592__, new_new_n13593__, new_new_n13594__,
    new_new_n13595__, new_new_n13596__, new_new_n13597__, new_new_n13598__,
    new_new_n13599__, new_new_n13600__, new_new_n13601__, new_new_n13602__,
    new_new_n13603__, new_new_n13604__, new_new_n13605__, new_new_n13606__,
    new_new_n13607__, new_new_n13608__, new_new_n13609__, new_new_n13610__,
    new_new_n13611__, new_new_n13612__, new_new_n13613__, new_new_n13614__,
    new_new_n13615__, new_new_n13616__, new_new_n13617__, new_new_n13618__,
    new_new_n13619__, new_new_n13620__, new_new_n13621__, new_new_n13622__,
    new_new_n13623__, new_new_n13624__, new_new_n13625__, new_new_n13626__,
    new_new_n13627__, new_new_n13628__, new_new_n13629__, new_new_n13630__,
    new_new_n13631__, new_new_n13632__, new_new_n13633__, new_new_n13634__,
    new_new_n13635__, new_new_n13636__, new_new_n13637__, new_new_n13638__,
    new_new_n13639__, new_new_n13640__, new_new_n13641__, new_new_n13642__,
    new_new_n13643__, new_new_n13644__, new_new_n13645__, new_new_n13646__,
    new_new_n13647__, new_new_n13648__, new_new_n13649__, new_new_n13650__,
    new_new_n13651__, new_new_n13652__, new_new_n13653__, new_new_n13654__,
    new_new_n13655__, new_new_n13656__, new_new_n13657__, new_new_n13658__,
    new_new_n13659__, new_new_n13660__, new_new_n13661__, new_new_n13662__,
    new_new_n13663__, new_new_n13664__, new_new_n13665__, new_new_n13666__,
    new_new_n13667__, new_new_n13668__, new_new_n13669__, new_new_n13670__,
    new_new_n13671__, new_new_n13672__, new_new_n13673__, new_new_n13674__,
    new_new_n13675__, new_new_n13676__, new_new_n13677__, new_new_n13678__,
    new_new_n13679__, new_new_n13680__, new_new_n13681__, new_new_n13682__,
    new_new_n13683__, new_new_n13684__, new_new_n13685__, new_new_n13686__,
    new_new_n13687__, new_new_n13688__, new_new_n13689__, new_new_n13690__,
    new_new_n13691__, new_new_n13692__, new_new_n13693__, new_new_n13694__,
    new_new_n13695__, new_new_n13696__, new_new_n13697__, new_new_n13698__,
    new_new_n13699__, new_new_n13700__, new_new_n13701__, new_new_n13702__,
    new_new_n13703__, new_new_n13704__, new_new_n13705__, new_new_n13706__,
    new_new_n13707__, new_new_n13708__, new_new_n13709__, new_new_n13710__,
    new_new_n13711__, new_new_n13712__, new_new_n13713__, new_new_n13714__,
    new_new_n13715__, new_new_n13716__, new_new_n13717__, new_new_n13718__,
    new_new_n13719__, new_new_n13720__, new_new_n13721__, new_new_n13722__,
    new_new_n13723__, new_new_n13724__, new_new_n13725__, new_new_n13726__,
    new_new_n13727__, new_new_n13728__, new_new_n13729__, new_new_n13730__,
    new_new_n13731__, new_new_n13732__, new_new_n13733__, new_new_n13734__,
    new_new_n13735__, new_new_n13736__, new_new_n13737__, new_new_n13738__,
    new_new_n13739__, new_new_n13740__, new_new_n13741__, new_new_n13742__,
    new_new_n13743__, new_new_n13744__, new_new_n13745__, new_new_n13746__,
    new_new_n13747__, new_new_n13748__, new_new_n13749__, new_new_n13750__,
    new_new_n13751__, new_new_n13752__, new_new_n13753__, new_new_n13754__,
    new_new_n13755__, new_new_n13756__, new_new_n13757__, new_new_n13758__,
    new_new_n13759__, new_new_n13760__, new_new_n13761__, new_new_n13762__,
    new_new_n13763__, new_new_n13764__, new_new_n13765__, new_new_n13766__,
    new_new_n13767__, new_new_n13768__, new_new_n13769__, new_new_n13770__,
    new_new_n13771__, new_new_n13772__, new_new_n13773__, new_new_n13774__,
    new_new_n13775__, new_new_n13776__, new_new_n13777__, new_new_n13778__,
    new_new_n13779__, new_new_n13780__, new_new_n13781__, new_new_n13782__,
    new_new_n13783__, new_new_n13784__, new_new_n13785__, new_new_n13786__,
    new_new_n13787__, new_new_n13788__, new_new_n13789__, new_new_n13790__,
    new_new_n13791__, new_new_n13792__, new_new_n13793__, new_new_n13794__,
    new_new_n13795__, new_new_n13796__, new_new_n13797__, new_new_n13798__,
    new_new_n13799__, new_new_n13800__, new_new_n13801__, new_new_n13802__,
    new_new_n13803__, new_new_n13804__, new_new_n13805__, new_new_n13806__,
    new_new_n13807__, new_new_n13808__, new_new_n13809__, new_new_n13810__,
    new_new_n13811__, new_new_n13812__, new_new_n13813__, new_new_n13814__,
    new_new_n13815__, new_new_n13816__, new_new_n13817__, new_new_n13818__,
    new_new_n13819__, new_new_n13820__, new_new_n13821__, new_new_n13822__,
    new_new_n13823__, new_new_n13824__, new_new_n13825__, new_new_n13826__,
    new_new_n13827__, new_new_n13828__, new_new_n13829__, new_new_n13830__,
    new_new_n13831__, new_new_n13832__, new_new_n13833__, new_new_n13834__,
    new_new_n13835__, new_new_n13836__, new_new_n13837__, new_new_n13838__,
    new_new_n13839__, new_new_n13840__, new_new_n13841__, new_new_n13842__,
    new_new_n13843__, new_new_n13844__, new_new_n13845__, new_new_n13846__,
    new_new_n13847__, new_new_n13848__, new_new_n13849__, new_new_n13850__,
    new_new_n13851__, new_new_n13852__, new_new_n13853__, new_new_n13854__,
    new_new_n13855__, new_new_n13856__, new_new_n13857__, new_new_n13858__,
    new_new_n13859__, new_new_n13860__, new_new_n13861__, new_new_n13862__,
    new_new_n13863__, new_new_n13864__, new_new_n13865__, new_new_n13866__,
    new_new_n13867__, new_new_n13868__, new_new_n13869__, new_new_n13870__,
    new_new_n13871__, new_new_n13872__, new_new_n13873__, new_new_n13874__,
    new_new_n13875__, new_new_n13876__, new_new_n13877__, new_new_n13878__,
    new_new_n13879__, new_new_n13880__, new_new_n13881__, new_new_n13882__,
    new_new_n13883__, new_new_n13884__, new_new_n13885__, new_new_n13886__,
    new_new_n13887__, new_new_n13888__, new_new_n13889__, new_new_n13890__,
    new_new_n13891__, new_new_n13892__, new_new_n13893__, new_new_n13894__,
    new_new_n13895__, new_new_n13896__, new_new_n13897__, new_new_n13898__,
    new_new_n13899__, new_new_n13900__, new_new_n13901__, new_new_n13902__,
    new_new_n13903__, new_new_n13904__, new_new_n13905__, new_new_n13906__,
    new_new_n13907__, new_new_n13908__, new_new_n13909__, new_new_n13910__,
    new_new_n13911__, new_new_n13912__, new_new_n13913__, new_new_n13914__,
    new_new_n13915__, new_new_n13916__, new_new_n13917__, new_new_n13918__,
    new_new_n13919__, new_new_n13920__, new_new_n13921__, new_new_n13922__,
    new_new_n13923__, new_new_n13924__, new_new_n13925__, new_new_n13926__,
    new_new_n13927__, new_new_n13928__, new_new_n13929__, new_new_n13930__,
    new_new_n13931__, new_new_n13932__, new_new_n13933__, new_new_n13934__,
    new_new_n13935__, new_new_n13936__, new_new_n13937__, new_new_n13938__,
    new_new_n13939__, new_new_n13940__, new_new_n13941__, new_new_n13942__,
    new_new_n13943__, new_new_n13944__, new_new_n13946__, new_new_n13947__,
    new_new_n13948__, new_new_n13949__, new_new_n13950__, new_new_n13951__,
    new_new_n13952__, new_new_n13953__, new_new_n13954__, new_new_n13955__,
    new_new_n13956__, new_new_n13957__, new_new_n13958__, new_new_n13959__,
    new_new_n13960__, new_new_n13961__, new_new_n13962__, new_new_n13963__,
    new_new_n13964__, new_new_n13965__, new_new_n13966__, new_new_n13967__,
    new_new_n13968__, new_new_n13969__, new_new_n13970__, new_new_n13971__,
    new_new_n13972__, new_new_n13973__, new_new_n13974__, new_new_n13975__,
    new_new_n13976__, new_new_n13977__, new_new_n13978__, new_new_n13979__,
    new_new_n13980__, new_new_n13981__, new_new_n13982__, new_new_n13983__,
    new_new_n13984__, new_new_n13985__, new_new_n13986__, new_new_n13987__,
    new_new_n13988__, new_new_n13989__, new_new_n13990__, new_new_n13991__,
    new_new_n13992__, new_new_n13993__, new_new_n13994__, new_new_n13995__,
    new_new_n13996__, new_new_n13997__, new_new_n13998__, new_new_n13999__,
    new_new_n14000__, new_new_n14001__, new_new_n14002__, new_new_n14003__,
    new_new_n14004__, new_new_n14005__, new_new_n14006__, new_new_n14007__,
    new_new_n14008__, new_new_n14009__, new_new_n14010__, new_new_n14011__,
    new_new_n14012__, new_new_n14013__, new_new_n14014__, new_new_n14015__,
    new_new_n14016__, new_new_n14017__, new_new_n14018__, new_new_n14019__,
    new_new_n14020__, new_new_n14021__, new_new_n14022__, new_new_n14023__,
    new_new_n14024__, new_new_n14025__, new_new_n14026__, new_new_n14027__,
    new_new_n14028__, new_new_n14029__, new_new_n14030__, new_new_n14031__,
    new_new_n14032__, new_new_n14033__, new_new_n14034__, new_new_n14035__,
    new_new_n14036__, new_new_n14037__, new_new_n14038__, new_new_n14039__,
    new_new_n14040__, new_new_n14041__, new_new_n14042__, new_new_n14043__,
    new_new_n14044__, new_new_n14045__, new_new_n14046__, new_new_n14047__,
    new_new_n14048__, new_new_n14049__, new_new_n14050__, new_new_n14051__,
    new_new_n14052__, new_new_n14053__, new_new_n14054__, new_new_n14055__,
    new_new_n14056__, new_new_n14057__, new_new_n14058__, new_new_n14059__,
    new_new_n14060__, new_new_n14061__, new_new_n14062__, new_new_n14063__,
    new_new_n14064__, new_new_n14065__, new_new_n14066__, new_new_n14067__,
    new_new_n14068__, new_new_n14069__, new_new_n14070__, new_new_n14071__,
    new_new_n14072__, new_new_n14073__, new_new_n14074__, new_new_n14075__,
    new_new_n14076__, new_new_n14077__, new_new_n14078__, new_new_n14079__,
    new_new_n14080__, new_new_n14081__, new_new_n14082__, new_new_n14083__,
    new_new_n14084__, new_new_n14085__, new_new_n14086__, new_new_n14087__,
    new_new_n14088__, new_new_n14089__, new_new_n14090__, new_new_n14091__,
    new_new_n14092__, new_new_n14093__, new_new_n14094__, new_new_n14095__,
    new_new_n14096__, new_new_n14097__, new_new_n14098__, new_new_n14099__,
    new_new_n14100__, new_new_n14101__, new_new_n14102__, new_new_n14103__,
    new_new_n14104__, new_new_n14105__, new_new_n14106__, new_new_n14107__,
    new_new_n14108__, new_new_n14109__, new_new_n14110__, new_new_n14111__,
    new_new_n14112__, new_new_n14113__, new_new_n14114__, new_new_n14115__,
    new_new_n14116__, new_new_n14117__, new_new_n14118__, new_new_n14119__,
    new_new_n14120__, new_new_n14121__, new_new_n14122__, new_new_n14123__,
    new_new_n14124__, new_new_n14125__, new_new_n14126__, new_new_n14127__,
    new_new_n14128__, new_new_n14129__, new_new_n14130__, new_new_n14131__,
    new_new_n14132__, new_new_n14133__, new_new_n14134__, new_new_n14135__,
    new_new_n14136__, new_new_n14137__, new_new_n14138__, new_new_n14139__,
    new_new_n14140__, new_new_n14141__, new_new_n14142__, new_new_n14143__,
    new_new_n14144__, new_new_n14145__, new_new_n14146__, new_new_n14147__,
    new_new_n14148__, new_new_n14149__, new_new_n14150__, new_new_n14151__,
    new_new_n14152__, new_new_n14153__, new_new_n14154__, new_new_n14155__,
    new_new_n14156__, new_new_n14157__, new_new_n14158__, new_new_n14159__,
    new_new_n14160__, new_new_n14161__, new_new_n14162__, new_new_n14163__,
    new_new_n14164__, new_new_n14165__, new_new_n14166__, new_new_n14167__,
    new_new_n14168__, new_new_n14169__, new_new_n14170__, new_new_n14171__,
    new_new_n14172__, new_new_n14173__, new_new_n14174__, new_new_n14175__,
    new_new_n14176__, new_new_n14177__, new_new_n14178__, new_new_n14179__,
    new_new_n14180__, new_new_n14181__, new_new_n14182__, new_new_n14183__,
    new_new_n14184__, new_new_n14185__, new_new_n14186__, new_new_n14187__,
    new_new_n14188__, new_new_n14189__, new_new_n14190__, new_new_n14191__,
    new_new_n14192__, new_new_n14193__, new_new_n14194__, new_new_n14195__,
    new_new_n14196__, new_new_n14197__, new_new_n14198__, new_new_n14199__,
    new_new_n14200__, new_new_n14201__, new_new_n14202__, new_new_n14203__,
    new_new_n14204__, new_new_n14205__, new_new_n14206__, new_new_n14207__,
    new_new_n14208__, new_new_n14209__, new_new_n14210__, new_new_n14211__,
    new_new_n14212__, new_new_n14213__, new_new_n14214__, new_new_n14215__,
    new_new_n14216__, new_new_n14217__, new_new_n14218__, new_new_n14219__,
    new_new_n14220__, new_new_n14221__, new_new_n14222__, new_new_n14223__,
    new_new_n14224__, new_new_n14225__, new_new_n14226__, new_new_n14227__,
    new_new_n14228__, new_new_n14229__, new_new_n14230__, new_new_n14231__,
    new_new_n14232__, new_new_n14233__, new_new_n14234__, new_new_n14235__,
    new_new_n14236__, new_new_n14237__, new_new_n14238__, new_new_n14239__,
    new_new_n14240__, new_new_n14241__, new_new_n14242__, new_new_n14243__,
    new_new_n14244__, new_new_n14245__, new_new_n14246__, new_new_n14247__,
    new_new_n14248__, new_new_n14249__, new_new_n14250__, new_new_n14251__,
    new_new_n14252__, new_new_n14253__, new_new_n14254__, new_new_n14255__,
    new_new_n14256__, new_new_n14257__, new_new_n14258__, new_new_n14259__,
    new_new_n14260__, new_new_n14261__, new_new_n14262__, new_new_n14263__,
    new_new_n14264__, new_new_n14265__, new_new_n14266__, new_new_n14267__,
    new_new_n14268__, new_new_n14269__, new_new_n14270__, new_new_n14271__,
    new_new_n14272__, new_new_n14273__, new_new_n14274__, new_new_n14275__,
    new_new_n14276__, new_new_n14277__, new_new_n14278__, new_new_n14279__,
    new_new_n14280__, new_new_n14281__, new_new_n14282__, new_new_n14283__,
    new_new_n14284__, new_new_n14285__, new_new_n14286__, new_new_n14287__,
    new_new_n14288__, new_new_n14289__, new_new_n14290__, new_new_n14291__,
    new_new_n14292__, new_new_n14293__, new_new_n14294__, new_new_n14295__,
    new_new_n14296__, new_new_n14297__, new_new_n14298__, new_new_n14299__,
    new_new_n14300__, new_new_n14301__, new_new_n14302__, new_new_n14303__,
    new_new_n14304__, new_new_n14305__, new_new_n14306__, new_new_n14307__,
    new_new_n14308__, new_new_n14309__, new_new_n14310__, new_new_n14311__,
    new_new_n14312__, new_new_n14313__, new_new_n14314__, new_new_n14315__,
    new_new_n14316__, new_new_n14317__, new_new_n14318__, new_new_n14319__,
    new_new_n14320__, new_new_n14321__, new_new_n14322__, new_new_n14323__,
    new_new_n14324__, new_new_n14325__, new_new_n14326__, new_new_n14327__,
    new_new_n14328__, new_new_n14329__, new_new_n14330__, new_new_n14331__,
    new_new_n14332__, new_new_n14333__, new_new_n14334__, new_new_n14335__,
    new_new_n14336__, new_new_n14337__, new_new_n14338__, new_new_n14339__,
    new_new_n14340__, new_new_n14341__, new_new_n14342__, new_new_n14343__,
    new_new_n14344__, new_new_n14345__, new_new_n14346__, new_new_n14347__,
    new_new_n14348__, new_new_n14349__, new_new_n14350__, new_new_n14351__,
    new_new_n14352__, new_new_n14353__, new_new_n14354__, new_new_n14355__,
    new_new_n14356__, new_new_n14357__, new_new_n14358__, new_new_n14359__,
    new_new_n14360__, new_new_n14361__, new_new_n14362__, new_new_n14363__,
    new_new_n14364__, new_new_n14365__, new_new_n14366__, new_new_n14367__,
    new_new_n14368__, new_new_n14369__, new_new_n14370__, new_new_n14371__,
    new_new_n14372__, new_new_n14373__, new_new_n14374__, new_new_n14375__,
    new_new_n14376__, new_new_n14377__, new_new_n14378__, new_new_n14379__,
    new_new_n14380__, new_new_n14381__, new_new_n14382__, new_new_n14383__,
    new_new_n14384__, new_new_n14385__, new_new_n14386__, new_new_n14387__,
    new_new_n14388__, new_new_n14389__, new_new_n14390__, new_new_n14391__,
    new_new_n14392__, new_new_n14393__, new_new_n14394__, new_new_n14395__,
    new_new_n14396__, new_new_n14397__, new_new_n14398__, new_new_n14399__,
    new_new_n14400__, new_new_n14401__, new_new_n14402__, new_new_n14403__,
    new_new_n14404__, new_new_n14405__, new_new_n14406__, new_new_n14407__,
    new_new_n14408__, new_new_n14409__, new_new_n14410__, new_new_n14411__,
    new_new_n14412__, new_new_n14413__, new_new_n14414__, new_new_n14415__,
    new_new_n14416__, new_new_n14417__, new_new_n14418__, new_new_n14419__,
    new_new_n14420__, new_new_n14421__, new_new_n14422__, new_new_n14423__,
    new_new_n14424__, new_new_n14425__, new_new_n14426__, new_new_n14427__,
    new_new_n14428__, new_new_n14429__, new_new_n14430__, new_new_n14431__,
    new_new_n14432__, new_new_n14433__, new_new_n14434__, new_new_n14435__,
    new_new_n14436__, new_new_n14437__, new_new_n14438__, new_new_n14439__,
    new_new_n14440__, new_new_n14441__, new_new_n14442__, new_new_n14443__,
    new_new_n14444__, new_new_n14445__, new_new_n14446__, new_new_n14447__,
    new_new_n14448__, new_new_n14449__, new_new_n14450__, new_new_n14451__,
    new_new_n14452__, new_new_n14453__, new_new_n14454__, new_new_n14455__,
    new_new_n14456__, new_new_n14457__, new_new_n14458__, new_new_n14459__,
    new_new_n14460__, new_new_n14461__, new_new_n14462__, new_new_n14463__,
    new_new_n14464__, new_new_n14465__, new_new_n14466__, new_new_n14467__,
    new_new_n14468__, new_new_n14469__, new_new_n14470__, new_new_n14471__,
    new_new_n14472__, new_new_n14473__, new_new_n14474__, new_new_n14475__,
    new_new_n14476__, new_new_n14477__, new_new_n14478__, new_new_n14479__,
    new_new_n14480__, new_new_n14481__, new_new_n14482__, new_new_n14483__,
    new_new_n14484__, new_new_n14485__, new_new_n14486__, new_new_n14487__,
    new_new_n14488__, new_new_n14489__, new_new_n14490__, new_new_n14491__,
    new_new_n14492__, new_new_n14493__, new_new_n14494__, new_new_n14495__,
    new_new_n14496__, new_new_n14498__, new_new_n14499__, new_new_n14500__,
    new_new_n14501__, new_new_n14502__, new_new_n14503__, new_new_n14504__,
    new_new_n14505__, new_new_n14506__, new_new_n14507__, new_new_n14508__,
    new_new_n14509__, new_new_n14510__, new_new_n14511__, new_new_n14512__,
    new_new_n14513__, new_new_n14514__, new_new_n14515__, new_new_n14516__,
    new_new_n14517__, new_new_n14518__, new_new_n14519__, new_new_n14520__,
    new_new_n14521__, new_new_n14522__, new_new_n14523__, new_new_n14524__,
    new_new_n14525__, new_new_n14526__, new_new_n14527__, new_new_n14528__,
    new_new_n14529__, new_new_n14530__, new_new_n14531__, new_new_n14532__,
    new_new_n14533__, new_new_n14534__, new_new_n14535__, new_new_n14536__,
    new_new_n14537__, new_new_n14538__, new_new_n14539__, new_new_n14540__,
    new_new_n14541__, new_new_n14542__, new_new_n14543__, new_new_n14544__,
    new_new_n14545__, new_new_n14546__, new_new_n14547__, new_new_n14548__,
    new_new_n14549__, new_new_n14550__, new_new_n14551__, new_new_n14552__,
    new_new_n14553__, new_new_n14554__, new_new_n14555__, new_new_n14556__,
    new_new_n14557__, new_new_n14558__, new_new_n14559__, new_new_n14560__,
    new_new_n14561__, new_new_n14562__, new_new_n14563__, new_new_n14564__,
    new_new_n14565__, new_new_n14566__, new_new_n14567__, new_new_n14568__,
    new_new_n14569__, new_new_n14570__, new_new_n14571__, new_new_n14572__,
    new_new_n14573__, new_new_n14574__, new_new_n14575__, new_new_n14576__,
    new_new_n14577__, new_new_n14578__, new_new_n14579__, new_new_n14580__,
    new_new_n14581__, new_new_n14582__, new_new_n14583__, new_new_n14584__,
    new_new_n14585__, new_new_n14586__, new_new_n14587__, new_new_n14588__,
    new_new_n14589__, new_new_n14590__, new_new_n14591__, new_new_n14592__,
    new_new_n14593__, new_new_n14594__, new_new_n14595__, new_new_n14596__,
    new_new_n14597__, new_new_n14598__, new_new_n14599__, new_new_n14600__,
    new_new_n14601__, new_new_n14602__, new_new_n14603__, new_new_n14604__,
    new_new_n14605__, new_new_n14606__, new_new_n14607__, new_new_n14608__,
    new_new_n14609__, new_new_n14610__, new_new_n14611__, new_new_n14612__,
    new_new_n14613__, new_new_n14614__, new_new_n14615__, new_new_n14616__,
    new_new_n14617__, new_new_n14618__, new_new_n14619__, new_new_n14620__,
    new_new_n14621__, new_new_n14622__, new_new_n14623__, new_new_n14624__,
    new_new_n14625__, new_new_n14626__, new_new_n14627__, new_new_n14628__,
    new_new_n14629__, new_new_n14630__, new_new_n14631__, new_new_n14632__,
    new_new_n14633__, new_new_n14634__, new_new_n14635__, new_new_n14636__,
    new_new_n14637__, new_new_n14638__, new_new_n14639__, new_new_n14640__,
    new_new_n14641__, new_new_n14642__, new_new_n14643__, new_new_n14644__,
    new_new_n14645__, new_new_n14646__, new_new_n14647__, new_new_n14648__,
    new_new_n14649__, new_new_n14650__, new_new_n14651__, new_new_n14652__,
    new_new_n14653__, new_new_n14654__, new_new_n14655__, new_new_n14656__,
    new_new_n14657__, new_new_n14658__, new_new_n14659__, new_new_n14660__,
    new_new_n14661__, new_new_n14662__, new_new_n14663__, new_new_n14664__,
    new_new_n14665__, new_new_n14666__, new_new_n14667__, new_new_n14668__,
    new_new_n14669__, new_new_n14670__, new_new_n14671__, new_new_n14672__,
    new_new_n14673__, new_new_n14674__, new_new_n14675__, new_new_n14676__,
    new_new_n14677__, new_new_n14678__, new_new_n14679__, new_new_n14680__,
    new_new_n14681__, new_new_n14682__, new_new_n14683__, new_new_n14684__,
    new_new_n14685__, new_new_n14686__, new_new_n14687__, new_new_n14688__,
    new_new_n14689__, new_new_n14690__, new_new_n14691__, new_new_n14692__,
    new_new_n14693__, new_new_n14694__, new_new_n14695__, new_new_n14696__,
    new_new_n14697__, new_new_n14698__, new_new_n14699__, new_new_n14700__,
    new_new_n14701__, new_new_n14702__, new_new_n14703__, new_new_n14704__,
    new_new_n14705__, new_new_n14706__, new_new_n14707__, new_new_n14708__,
    new_new_n14709__, new_new_n14710__, new_new_n14711__, new_new_n14712__,
    new_new_n14713__, new_new_n14714__, new_new_n14715__, new_new_n14716__,
    new_new_n14717__, new_new_n14718__, new_new_n14719__, new_new_n14720__,
    new_new_n14721__, new_new_n14722__, new_new_n14723__, new_new_n14724__,
    new_new_n14725__, new_new_n14726__, new_new_n14727__, new_new_n14728__,
    new_new_n14729__, new_new_n14730__, new_new_n14731__, new_new_n14732__,
    new_new_n14733__, new_new_n14734__, new_new_n14735__, new_new_n14736__,
    new_new_n14737__, new_new_n14738__, new_new_n14739__, new_new_n14740__,
    new_new_n14741__, new_new_n14742__, new_new_n14743__, new_new_n14744__,
    new_new_n14745__, new_new_n14746__, new_new_n14747__, new_new_n14748__,
    new_new_n14749__, new_new_n14750__, new_new_n14751__, new_new_n14752__,
    new_new_n14753__, new_new_n14754__, new_new_n14755__, new_new_n14756__,
    new_new_n14757__, new_new_n14758__, new_new_n14759__, new_new_n14760__,
    new_new_n14761__, new_new_n14762__, new_new_n14763__, new_new_n14764__,
    new_new_n14765__, new_new_n14766__, new_new_n14767__, new_new_n14768__,
    new_new_n14769__, new_new_n14770__, new_new_n14771__, new_new_n14772__,
    new_new_n14773__, new_new_n14774__, new_new_n14775__, new_new_n14776__,
    new_new_n14777__, new_new_n14778__, new_new_n14779__, new_new_n14780__,
    new_new_n14781__, new_new_n14782__, new_new_n14783__, new_new_n14784__,
    new_new_n14785__, new_new_n14786__, new_new_n14787__, new_new_n14788__,
    new_new_n14789__, new_new_n14790__, new_new_n14791__, new_new_n14792__,
    new_new_n14793__, new_new_n14794__, new_new_n14795__, new_new_n14796__,
    new_new_n14797__, new_new_n14798__, new_new_n14799__, new_new_n14800__,
    new_new_n14801__, new_new_n14802__, new_new_n14803__, new_new_n14804__,
    new_new_n14805__, new_new_n14806__, new_new_n14807__, new_new_n14808__,
    new_new_n14809__, new_new_n14810__, new_new_n14811__, new_new_n14812__,
    new_new_n14813__, new_new_n14814__, new_new_n14815__, new_new_n14816__,
    new_new_n14817__, new_new_n14818__, new_new_n14819__, new_new_n14820__,
    new_new_n14821__, new_new_n14822__, new_new_n14823__, new_new_n14824__,
    new_new_n14825__, new_new_n14826__, new_new_n14827__, new_new_n14828__,
    new_new_n14829__, new_new_n14830__, new_new_n14831__, new_new_n14832__,
    new_new_n14833__, new_new_n14834__, new_new_n14835__, new_new_n14836__,
    new_new_n14837__, new_new_n14838__, new_new_n14839__, new_new_n14840__,
    new_new_n14841__, new_new_n14842__, new_new_n14843__, new_new_n14844__,
    new_new_n14845__, new_new_n14846__, new_new_n14847__, new_new_n14848__,
    new_new_n14849__, new_new_n14850__, new_new_n14851__, new_new_n14852__,
    new_new_n14853__, new_new_n14854__, new_new_n14855__, new_new_n14856__,
    new_new_n14857__, new_new_n14858__, new_new_n14859__, new_new_n14860__,
    new_new_n14861__, new_new_n14862__, new_new_n14863__, new_new_n14864__,
    new_new_n14865__, new_new_n14866__, new_new_n14867__, new_new_n14868__,
    new_new_n14869__, new_new_n14870__, new_new_n14871__, new_new_n14872__,
    new_new_n14873__, new_new_n14874__, new_new_n14875__, new_new_n14876__,
    new_new_n14877__, new_new_n14878__, new_new_n14879__, new_new_n14880__,
    new_new_n14881__, new_new_n14882__, new_new_n14883__, new_new_n14884__,
    new_new_n14885__, new_new_n14886__, new_new_n14887__, new_new_n14888__,
    new_new_n14889__, new_new_n14890__, new_new_n14891__, new_new_n14892__,
    new_new_n14893__, new_new_n14894__, new_new_n14895__, new_new_n14896__,
    new_new_n14897__, new_new_n14898__, new_new_n14899__, new_new_n14900__,
    new_new_n14901__, new_new_n14902__, new_new_n14903__, new_new_n14904__,
    new_new_n14905__, new_new_n14906__, new_new_n14907__, new_new_n14908__,
    new_new_n14909__, new_new_n14910__, new_new_n14911__, new_new_n14912__,
    new_new_n14913__, new_new_n14914__, new_new_n14915__, new_new_n14916__,
    new_new_n14917__, new_new_n14918__, new_new_n14919__, new_new_n14920__,
    new_new_n14921__, new_new_n14922__, new_new_n14923__, new_new_n14924__,
    new_new_n14925__, new_new_n14926__, new_new_n14927__, new_new_n14928__,
    new_new_n14929__, new_new_n14930__, new_new_n14931__, new_new_n14932__,
    new_new_n14933__, new_new_n14934__, new_new_n14935__, new_new_n14936__,
    new_new_n14937__, new_new_n14938__, new_new_n14939__, new_new_n14940__,
    new_new_n14941__, new_new_n14942__, new_new_n14943__, new_new_n14944__,
    new_new_n14945__, new_new_n14946__, new_new_n14947__, new_new_n14948__,
    new_new_n14949__, new_new_n14950__, new_new_n14951__, new_new_n14952__,
    new_new_n14953__, new_new_n14954__, new_new_n14955__, new_new_n14956__,
    new_new_n14957__, new_new_n14958__, new_new_n14959__, new_new_n14960__,
    new_new_n14961__, new_new_n14962__, new_new_n14963__, new_new_n14964__,
    new_new_n14965__, new_new_n14966__, new_new_n14967__, new_new_n14968__,
    new_new_n14969__, new_new_n14970__, new_new_n14971__, new_new_n14972__,
    new_new_n14973__, new_new_n14974__, new_new_n14975__, new_new_n14976__,
    new_new_n14977__, new_new_n14978__, new_new_n14979__, new_new_n14980__,
    new_new_n14981__, new_new_n14982__, new_new_n14983__, new_new_n14984__,
    new_new_n14985__, new_new_n14986__, new_new_n14987__, new_new_n14988__,
    new_new_n14989__, new_new_n14990__, new_new_n14991__, new_new_n14992__,
    new_new_n14993__, new_new_n14994__, new_new_n14995__, new_new_n14996__,
    new_new_n14997__, new_new_n14998__, new_new_n14999__, new_new_n15000__,
    new_new_n15001__, new_new_n15002__, new_new_n15003__, new_new_n15004__,
    new_new_n15005__, new_new_n15006__, new_new_n15007__, new_new_n15008__,
    new_new_n15009__, new_new_n15010__, new_new_n15011__, new_new_n15012__,
    new_new_n15013__, new_new_n15014__, new_new_n15015__, new_new_n15016__,
    new_new_n15017__, new_new_n15018__, new_new_n15019__, new_new_n15020__,
    new_new_n15021__, new_new_n15022__, new_new_n15023__, new_new_n15024__,
    new_new_n15025__, new_new_n15026__, new_new_n15027__, new_new_n15028__,
    new_new_n15029__, new_new_n15030__, new_new_n15031__, new_new_n15032__,
    new_new_n15033__, new_new_n15034__, new_new_n15035__, new_new_n15036__,
    new_new_n15037__, new_new_n15038__, new_new_n15039__, new_new_n15040__,
    new_new_n15041__, new_new_n15042__, new_new_n15043__, new_new_n15044__,
    new_new_n15045__, new_new_n15046__, new_new_n15047__, new_new_n15048__,
    new_new_n15049__, new_new_n15050__, new_new_n15051__, new_new_n15052__,
    new_new_n15053__, new_new_n15054__, new_new_n15055__, new_new_n15056__,
    new_new_n15057__, new_new_n15058__, new_new_n15059__, new_new_n15060__,
    new_new_n15061__, new_new_n15062__, new_new_n15063__, new_new_n15064__,
    new_new_n15065__, new_new_n15066__, new_new_n15067__, new_new_n15068__,
    new_new_n15069__, new_new_n15070__, new_new_n15071__, new_new_n15072__,
    new_new_n15073__, new_new_n15074__, new_new_n15075__, new_new_n15076__,
    new_new_n15077__, new_new_n15078__, new_new_n15080__, new_new_n15081__,
    new_new_n15082__, new_new_n15083__, new_new_n15084__, new_new_n15085__,
    new_new_n15086__, new_new_n15087__, new_new_n15088__, new_new_n15089__,
    new_new_n15090__, new_new_n15091__, new_new_n15092__, new_new_n15093__,
    new_new_n15094__, new_new_n15095__, new_new_n15096__, new_new_n15097__,
    new_new_n15098__, new_new_n15099__, new_new_n15100__, new_new_n15101__,
    new_new_n15102__, new_new_n15103__, new_new_n15104__, new_new_n15105__,
    new_new_n15106__, new_new_n15107__, new_new_n15108__, new_new_n15109__,
    new_new_n15110__, new_new_n15111__, new_new_n15112__, new_new_n15113__,
    new_new_n15114__, new_new_n15115__, new_new_n15116__, new_new_n15117__,
    new_new_n15118__, new_new_n15119__, new_new_n15120__, new_new_n15121__,
    new_new_n15122__, new_new_n15123__, new_new_n15124__, new_new_n15125__,
    new_new_n15126__, new_new_n15127__, new_new_n15128__, new_new_n15129__,
    new_new_n15130__, new_new_n15131__, new_new_n15132__, new_new_n15133__,
    new_new_n15134__, new_new_n15135__, new_new_n15136__, new_new_n15137__,
    new_new_n15138__, new_new_n15139__, new_new_n15140__, new_new_n15141__,
    new_new_n15142__, new_new_n15143__, new_new_n15144__, new_new_n15145__,
    new_new_n15146__, new_new_n15147__, new_new_n15148__, new_new_n15149__,
    new_new_n15150__, new_new_n15151__, new_new_n15152__, new_new_n15153__,
    new_new_n15154__, new_new_n15155__, new_new_n15156__, new_new_n15157__,
    new_new_n15158__, new_new_n15159__, new_new_n15160__, new_new_n15161__,
    new_new_n15162__, new_new_n15163__, new_new_n15164__, new_new_n15165__,
    new_new_n15166__, new_new_n15167__, new_new_n15168__, new_new_n15169__,
    new_new_n15170__, new_new_n15171__, new_new_n15172__, new_new_n15173__,
    new_new_n15174__, new_new_n15175__, new_new_n15176__, new_new_n15177__,
    new_new_n15178__, new_new_n15179__, new_new_n15180__, new_new_n15181__,
    new_new_n15182__, new_new_n15183__, new_new_n15184__, new_new_n15185__,
    new_new_n15186__, new_new_n15187__, new_new_n15188__, new_new_n15189__,
    new_new_n15190__, new_new_n15191__, new_new_n15192__, new_new_n15193__,
    new_new_n15194__, new_new_n15195__, new_new_n15196__, new_new_n15197__,
    new_new_n15198__, new_new_n15199__, new_new_n15200__, new_new_n15201__,
    new_new_n15202__, new_new_n15203__, new_new_n15204__, new_new_n15205__,
    new_new_n15206__, new_new_n15207__, new_new_n15208__, new_new_n15209__,
    new_new_n15210__, new_new_n15211__, new_new_n15212__, new_new_n15213__,
    new_new_n15214__, new_new_n15215__, new_new_n15216__, new_new_n15217__,
    new_new_n15218__, new_new_n15219__, new_new_n15220__, new_new_n15221__,
    new_new_n15222__, new_new_n15223__, new_new_n15224__, new_new_n15225__,
    new_new_n15226__, new_new_n15227__, new_new_n15228__, new_new_n15229__,
    new_new_n15230__, new_new_n15231__, new_new_n15232__, new_new_n15233__,
    new_new_n15234__, new_new_n15235__, new_new_n15236__, new_new_n15237__,
    new_new_n15238__, new_new_n15239__, new_new_n15240__, new_new_n15241__,
    new_new_n15242__, new_new_n15243__, new_new_n15244__, new_new_n15245__,
    new_new_n15246__, new_new_n15247__, new_new_n15248__, new_new_n15249__,
    new_new_n15250__, new_new_n15251__, new_new_n15252__, new_new_n15253__,
    new_new_n15254__, new_new_n15255__, new_new_n15256__, new_new_n15257__,
    new_new_n15258__, new_new_n15259__, new_new_n15260__, new_new_n15261__,
    new_new_n15262__, new_new_n15263__, new_new_n15264__, new_new_n15265__,
    new_new_n15266__, new_new_n15267__, new_new_n15268__, new_new_n15269__,
    new_new_n15270__, new_new_n15271__, new_new_n15272__, new_new_n15273__,
    new_new_n15274__, new_new_n15275__, new_new_n15276__, new_new_n15277__,
    new_new_n15278__, new_new_n15279__, new_new_n15280__, new_new_n15281__,
    new_new_n15282__, new_new_n15283__, new_new_n15284__, new_new_n15285__,
    new_new_n15286__, new_new_n15287__, new_new_n15288__, new_new_n15289__,
    new_new_n15290__, new_new_n15291__, new_new_n15292__, new_new_n15293__,
    new_new_n15294__, new_new_n15295__, new_new_n15296__, new_new_n15297__,
    new_new_n15298__, new_new_n15299__, new_new_n15300__, new_new_n15301__,
    new_new_n15302__, new_new_n15303__, new_new_n15304__, new_new_n15305__,
    new_new_n15306__, new_new_n15307__, new_new_n15308__, new_new_n15309__,
    new_new_n15310__, new_new_n15311__, new_new_n15312__, new_new_n15313__,
    new_new_n15314__, new_new_n15315__, new_new_n15316__, new_new_n15317__,
    new_new_n15318__, new_new_n15319__, new_new_n15320__, new_new_n15321__,
    new_new_n15322__, new_new_n15323__, new_new_n15324__, new_new_n15325__,
    new_new_n15326__, new_new_n15327__, new_new_n15328__, new_new_n15329__,
    new_new_n15330__, new_new_n15331__, new_new_n15332__, new_new_n15333__,
    new_new_n15334__, new_new_n15335__, new_new_n15336__, new_new_n15337__,
    new_new_n15338__, new_new_n15339__, new_new_n15340__, new_new_n15341__,
    new_new_n15342__, new_new_n15343__, new_new_n15344__, new_new_n15345__,
    new_new_n15346__, new_new_n15347__, new_new_n15348__, new_new_n15349__,
    new_new_n15350__, new_new_n15351__, new_new_n15352__, new_new_n15353__,
    new_new_n15354__, new_new_n15355__, new_new_n15356__, new_new_n15357__,
    new_new_n15358__, new_new_n15359__, new_new_n15360__, new_new_n15361__,
    new_new_n15362__, new_new_n15363__, new_new_n15364__, new_new_n15365__,
    new_new_n15366__, new_new_n15367__, new_new_n15368__, new_new_n15369__,
    new_new_n15370__, new_new_n15371__, new_new_n15372__, new_new_n15373__,
    new_new_n15374__, new_new_n15375__, new_new_n15376__, new_new_n15377__,
    new_new_n15378__, new_new_n15379__, new_new_n15380__, new_new_n15381__,
    new_new_n15382__, new_new_n15383__, new_new_n15384__, new_new_n15385__,
    new_new_n15386__, new_new_n15387__, new_new_n15388__, new_new_n15389__,
    new_new_n15390__, new_new_n15391__, new_new_n15392__, new_new_n15393__,
    new_new_n15394__, new_new_n15395__, new_new_n15396__, new_new_n15397__,
    new_new_n15398__, new_new_n15399__, new_new_n15400__, new_new_n15401__,
    new_new_n15402__, new_new_n15403__, new_new_n15404__, new_new_n15405__,
    new_new_n15406__, new_new_n15407__, new_new_n15408__, new_new_n15409__,
    new_new_n15410__, new_new_n15411__, new_new_n15412__, new_new_n15413__,
    new_new_n15414__, new_new_n15415__, new_new_n15416__, new_new_n15417__,
    new_new_n15418__, new_new_n15419__, new_new_n15420__, new_new_n15421__,
    new_new_n15422__, new_new_n15423__, new_new_n15424__, new_new_n15425__,
    new_new_n15426__, new_new_n15427__, new_new_n15428__, new_new_n15429__,
    new_new_n15430__, new_new_n15431__, new_new_n15432__, new_new_n15433__,
    new_new_n15434__, new_new_n15435__, new_new_n15436__, new_new_n15437__,
    new_new_n15438__, new_new_n15439__, new_new_n15440__, new_new_n15441__,
    new_new_n15442__, new_new_n15443__, new_new_n15444__, new_new_n15445__,
    new_new_n15446__, new_new_n15447__, new_new_n15448__, new_new_n15449__,
    new_new_n15450__, new_new_n15451__, new_new_n15452__, new_new_n15453__,
    new_new_n15454__, new_new_n15455__, new_new_n15456__, new_new_n15457__,
    new_new_n15458__, new_new_n15459__, new_new_n15460__, new_new_n15461__,
    new_new_n15462__, new_new_n15463__, new_new_n15464__, new_new_n15465__,
    new_new_n15466__, new_new_n15467__, new_new_n15468__, new_new_n15469__,
    new_new_n15470__, new_new_n15471__, new_new_n15472__, new_new_n15473__,
    new_new_n15474__, new_new_n15475__, new_new_n15476__, new_new_n15477__,
    new_new_n15478__, new_new_n15479__, new_new_n15480__, new_new_n15481__,
    new_new_n15482__, new_new_n15483__, new_new_n15484__, new_new_n15485__,
    new_new_n15486__, new_new_n15487__, new_new_n15488__, new_new_n15489__,
    new_new_n15490__, new_new_n15491__, new_new_n15492__, new_new_n15493__,
    new_new_n15494__, new_new_n15495__, new_new_n15496__, new_new_n15497__,
    new_new_n15498__, new_new_n15499__, new_new_n15500__, new_new_n15501__,
    new_new_n15502__, new_new_n15503__, new_new_n15504__, new_new_n15505__,
    new_new_n15506__, new_new_n15507__, new_new_n15508__, new_new_n15509__,
    new_new_n15510__, new_new_n15511__, new_new_n15512__, new_new_n15513__,
    new_new_n15514__, new_new_n15515__, new_new_n15516__, new_new_n15517__,
    new_new_n15518__, new_new_n15519__, new_new_n15520__, new_new_n15521__,
    new_new_n15522__, new_new_n15523__, new_new_n15524__, new_new_n15525__,
    new_new_n15526__, new_new_n15527__, new_new_n15528__, new_new_n15529__,
    new_new_n15530__, new_new_n15531__, new_new_n15532__, new_new_n15533__,
    new_new_n15534__, new_new_n15535__, new_new_n15536__, new_new_n15537__,
    new_new_n15538__, new_new_n15539__, new_new_n15540__, new_new_n15541__,
    new_new_n15542__, new_new_n15543__, new_new_n15544__, new_new_n15545__,
    new_new_n15546__, new_new_n15547__, new_new_n15548__, new_new_n15549__,
    new_new_n15550__, new_new_n15551__, new_new_n15552__, new_new_n15553__,
    new_new_n15554__, new_new_n15555__, new_new_n15556__, new_new_n15557__,
    new_new_n15558__, new_new_n15559__, new_new_n15560__, new_new_n15561__,
    new_new_n15562__, new_new_n15563__, new_new_n15564__, new_new_n15565__,
    new_new_n15566__, new_new_n15567__, new_new_n15568__, new_new_n15569__,
    new_new_n15570__, new_new_n15571__, new_new_n15572__, new_new_n15573__,
    new_new_n15574__, new_new_n15575__, new_new_n15576__, new_new_n15577__,
    new_new_n15578__, new_new_n15579__, new_new_n15580__, new_new_n15581__,
    new_new_n15582__, new_new_n15583__, new_new_n15584__, new_new_n15585__,
    new_new_n15586__, new_new_n15587__, new_new_n15588__, new_new_n15589__,
    new_new_n15590__, new_new_n15591__, new_new_n15592__, new_new_n15593__,
    new_new_n15594__, new_new_n15595__, new_new_n15596__, new_new_n15597__,
    new_new_n15598__, new_new_n15599__, new_new_n15600__, new_new_n15601__,
    new_new_n15602__, new_new_n15603__, new_new_n15604__, new_new_n15605__,
    new_new_n15606__, new_new_n15607__, new_new_n15608__, new_new_n15609__,
    new_new_n15610__, new_new_n15611__, new_new_n15612__, new_new_n15613__,
    new_new_n15614__, new_new_n15615__, new_new_n15616__, new_new_n15617__,
    new_new_n15618__, new_new_n15619__, new_new_n15620__, new_new_n15621__,
    new_new_n15622__, new_new_n15623__, new_new_n15624__, new_new_n15625__,
    new_new_n15626__, new_new_n15627__, new_new_n15628__, new_new_n15629__,
    new_new_n15630__, new_new_n15631__, new_new_n15632__, new_new_n15633__,
    new_new_n15634__, new_new_n15635__, new_new_n15636__, new_new_n15637__,
    new_new_n15638__, new_new_n15639__, new_new_n15640__, new_new_n15641__,
    new_new_n15642__, new_new_n15643__, new_new_n15644__, new_new_n15645__,
    new_new_n15647__, new_new_n15648__, new_new_n15649__, new_new_n15650__,
    new_new_n15651__, new_new_n15652__, new_new_n15653__, new_new_n15654__,
    new_new_n15655__, new_new_n15656__, new_new_n15657__, new_new_n15658__,
    new_new_n15659__, new_new_n15660__, new_new_n15661__, new_new_n15662__,
    new_new_n15663__, new_new_n15664__, new_new_n15665__, new_new_n15666__,
    new_new_n15667__, new_new_n15668__, new_new_n15669__, new_new_n15670__,
    new_new_n15671__, new_new_n15672__, new_new_n15673__, new_new_n15674__,
    new_new_n15675__, new_new_n15676__, new_new_n15677__, new_new_n15678__,
    new_new_n15679__, new_new_n15680__, new_new_n15681__, new_new_n15682__,
    new_new_n15683__, new_new_n15684__, new_new_n15685__, new_new_n15686__,
    new_new_n15687__, new_new_n15688__, new_new_n15689__, new_new_n15690__,
    new_new_n15691__, new_new_n15692__, new_new_n15693__, new_new_n15694__,
    new_new_n15695__, new_new_n15696__, new_new_n15697__, new_new_n15698__,
    new_new_n15699__, new_new_n15700__, new_new_n15701__, new_new_n15702__,
    new_new_n15703__, new_new_n15704__, new_new_n15705__, new_new_n15706__,
    new_new_n15707__, new_new_n15708__, new_new_n15709__, new_new_n15710__,
    new_new_n15711__, new_new_n15712__, new_new_n15713__, new_new_n15714__,
    new_new_n15715__, new_new_n15716__, new_new_n15717__, new_new_n15718__,
    new_new_n15719__, new_new_n15720__, new_new_n15721__, new_new_n15722__,
    new_new_n15723__, new_new_n15724__, new_new_n15725__, new_new_n15726__,
    new_new_n15727__, new_new_n15728__, new_new_n15729__, new_new_n15730__,
    new_new_n15731__, new_new_n15732__, new_new_n15733__, new_new_n15734__,
    new_new_n15735__, new_new_n15736__, new_new_n15737__, new_new_n15738__,
    new_new_n15739__, new_new_n15740__, new_new_n15741__, new_new_n15742__,
    new_new_n15743__, new_new_n15744__, new_new_n15745__, new_new_n15746__,
    new_new_n15747__, new_new_n15748__, new_new_n15749__, new_new_n15750__,
    new_new_n15751__, new_new_n15752__, new_new_n15753__, new_new_n15754__,
    new_new_n15755__, new_new_n15756__, new_new_n15757__, new_new_n15758__,
    new_new_n15759__, new_new_n15760__, new_new_n15761__, new_new_n15762__,
    new_new_n15763__, new_new_n15764__, new_new_n15765__, new_new_n15766__,
    new_new_n15767__, new_new_n15768__, new_new_n15769__, new_new_n15770__,
    new_new_n15771__, new_new_n15772__, new_new_n15773__, new_new_n15774__,
    new_new_n15775__, new_new_n15776__, new_new_n15777__, new_new_n15778__,
    new_new_n15779__, new_new_n15780__, new_new_n15781__, new_new_n15782__,
    new_new_n15783__, new_new_n15784__, new_new_n15785__, new_new_n15786__,
    new_new_n15787__, new_new_n15788__, new_new_n15789__, new_new_n15790__,
    new_new_n15791__, new_new_n15792__, new_new_n15793__, new_new_n15794__,
    new_new_n15795__, new_new_n15796__, new_new_n15797__, new_new_n15798__,
    new_new_n15799__, new_new_n15800__, new_new_n15801__, new_new_n15802__,
    new_new_n15803__, new_new_n15804__, new_new_n15805__, new_new_n15806__,
    new_new_n15807__, new_new_n15808__, new_new_n15809__, new_new_n15810__,
    new_new_n15811__, new_new_n15812__, new_new_n15813__, new_new_n15814__,
    new_new_n15815__, new_new_n15816__, new_new_n15817__, new_new_n15818__,
    new_new_n15819__, new_new_n15820__, new_new_n15821__, new_new_n15822__,
    new_new_n15823__, new_new_n15824__, new_new_n15825__, new_new_n15826__,
    new_new_n15827__, new_new_n15828__, new_new_n15829__, new_new_n15830__,
    new_new_n15831__, new_new_n15832__, new_new_n15833__, new_new_n15834__,
    new_new_n15835__, new_new_n15836__, new_new_n15837__, new_new_n15838__,
    new_new_n15839__, new_new_n15840__, new_new_n15841__, new_new_n15842__,
    new_new_n15843__, new_new_n15844__, new_new_n15845__, new_new_n15846__,
    new_new_n15847__, new_new_n15848__, new_new_n15849__, new_new_n15850__,
    new_new_n15851__, new_new_n15852__, new_new_n15853__, new_new_n15854__,
    new_new_n15855__, new_new_n15856__, new_new_n15857__, new_new_n15858__,
    new_new_n15859__, new_new_n15860__, new_new_n15861__, new_new_n15862__,
    new_new_n15863__, new_new_n15864__, new_new_n15865__, new_new_n15866__,
    new_new_n15867__, new_new_n15868__, new_new_n15869__, new_new_n15870__,
    new_new_n15871__, new_new_n15872__, new_new_n15873__, new_new_n15874__,
    new_new_n15875__, new_new_n15876__, new_new_n15877__, new_new_n15878__,
    new_new_n15879__, new_new_n15880__, new_new_n15881__, new_new_n15882__,
    new_new_n15883__, new_new_n15884__, new_new_n15885__, new_new_n15886__,
    new_new_n15887__, new_new_n15888__, new_new_n15889__, new_new_n15890__,
    new_new_n15891__, new_new_n15892__, new_new_n15893__, new_new_n15894__,
    new_new_n15895__, new_new_n15896__, new_new_n15897__, new_new_n15898__,
    new_new_n15899__, new_new_n15900__, new_new_n15901__, new_new_n15902__,
    new_new_n15903__, new_new_n15904__, new_new_n15905__, new_new_n15906__,
    new_new_n15907__, new_new_n15908__, new_new_n15909__, new_new_n15910__,
    new_new_n15911__, new_new_n15912__, new_new_n15913__, new_new_n15914__,
    new_new_n15915__, new_new_n15916__, new_new_n15917__, new_new_n15918__,
    new_new_n15919__, new_new_n15920__, new_new_n15921__, new_new_n15922__,
    new_new_n15923__, new_new_n15924__, new_new_n15925__, new_new_n15926__,
    new_new_n15927__, new_new_n15928__, new_new_n15929__, new_new_n15930__,
    new_new_n15931__, new_new_n15932__, new_new_n15933__, new_new_n15934__,
    new_new_n15935__, new_new_n15936__, new_new_n15937__, new_new_n15938__,
    new_new_n15939__, new_new_n15940__, new_new_n15941__, new_new_n15942__,
    new_new_n15943__, new_new_n15944__, new_new_n15945__, new_new_n15946__,
    new_new_n15947__, new_new_n15948__, new_new_n15949__, new_new_n15950__,
    new_new_n15951__, new_new_n15952__, new_new_n15953__, new_new_n15954__,
    new_new_n15955__, new_new_n15956__, new_new_n15957__, new_new_n15958__,
    new_new_n15959__, new_new_n15960__, new_new_n15961__, new_new_n15962__,
    new_new_n15963__, new_new_n15964__, new_new_n15965__, new_new_n15966__,
    new_new_n15967__, new_new_n15968__, new_new_n15969__, new_new_n15970__,
    new_new_n15971__, new_new_n15972__, new_new_n15973__, new_new_n15974__,
    new_new_n15975__, new_new_n15976__, new_new_n15977__, new_new_n15978__,
    new_new_n15979__, new_new_n15980__, new_new_n15981__, new_new_n15982__,
    new_new_n15983__, new_new_n15984__, new_new_n15985__, new_new_n15986__,
    new_new_n15987__, new_new_n15988__, new_new_n15989__, new_new_n15990__,
    new_new_n15991__, new_new_n15992__, new_new_n15993__, new_new_n15994__,
    new_new_n15995__, new_new_n15996__, new_new_n15997__, new_new_n15998__,
    new_new_n15999__, new_new_n16000__, new_new_n16001__, new_new_n16002__,
    new_new_n16003__, new_new_n16004__, new_new_n16005__, new_new_n16006__,
    new_new_n16007__, new_new_n16008__, new_new_n16009__, new_new_n16010__,
    new_new_n16011__, new_new_n16012__, new_new_n16013__, new_new_n16014__,
    new_new_n16015__, new_new_n16016__, new_new_n16017__, new_new_n16018__,
    new_new_n16019__, new_new_n16020__, new_new_n16021__, new_new_n16022__,
    new_new_n16023__, new_new_n16024__, new_new_n16025__, new_new_n16026__,
    new_new_n16027__, new_new_n16028__, new_new_n16029__, new_new_n16030__,
    new_new_n16031__, new_new_n16032__, new_new_n16033__, new_new_n16034__,
    new_new_n16035__, new_new_n16036__, new_new_n16037__, new_new_n16038__,
    new_new_n16039__, new_new_n16040__, new_new_n16041__, new_new_n16042__,
    new_new_n16043__, new_new_n16044__, new_new_n16045__, new_new_n16046__,
    new_new_n16047__, new_new_n16048__, new_new_n16049__, new_new_n16050__,
    new_new_n16051__, new_new_n16052__, new_new_n16053__, new_new_n16054__,
    new_new_n16055__, new_new_n16056__, new_new_n16057__, new_new_n16058__,
    new_new_n16059__, new_new_n16060__, new_new_n16061__, new_new_n16062__,
    new_new_n16063__, new_new_n16064__, new_new_n16065__, new_new_n16066__,
    new_new_n16067__, new_new_n16068__, new_new_n16069__, new_new_n16070__,
    new_new_n16071__, new_new_n16072__, new_new_n16073__, new_new_n16074__,
    new_new_n16075__, new_new_n16076__, new_new_n16077__, new_new_n16078__,
    new_new_n16079__, new_new_n16080__, new_new_n16081__, new_new_n16082__,
    new_new_n16083__, new_new_n16084__, new_new_n16085__, new_new_n16086__,
    new_new_n16087__, new_new_n16088__, new_new_n16089__, new_new_n16090__,
    new_new_n16091__, new_new_n16092__, new_new_n16093__, new_new_n16094__,
    new_new_n16095__, new_new_n16096__, new_new_n16097__, new_new_n16098__,
    new_new_n16099__, new_new_n16100__, new_new_n16101__, new_new_n16102__,
    new_new_n16103__, new_new_n16104__, new_new_n16105__, new_new_n16106__,
    new_new_n16107__, new_new_n16108__, new_new_n16109__, new_new_n16110__,
    new_new_n16111__, new_new_n16112__, new_new_n16113__, new_new_n16114__,
    new_new_n16115__, new_new_n16116__, new_new_n16117__, new_new_n16118__,
    new_new_n16119__, new_new_n16120__, new_new_n16121__, new_new_n16122__,
    new_new_n16123__, new_new_n16124__, new_new_n16125__, new_new_n16126__,
    new_new_n16127__, new_new_n16128__, new_new_n16129__, new_new_n16130__,
    new_new_n16131__, new_new_n16132__, new_new_n16133__, new_new_n16134__,
    new_new_n16135__, new_new_n16136__, new_new_n16137__, new_new_n16138__,
    new_new_n16139__, new_new_n16140__, new_new_n16141__, new_new_n16142__,
    new_new_n16143__, new_new_n16144__, new_new_n16145__, new_new_n16146__,
    new_new_n16147__, new_new_n16148__, new_new_n16149__, new_new_n16150__,
    new_new_n16151__, new_new_n16152__, new_new_n16153__, new_new_n16154__,
    new_new_n16155__, new_new_n16156__, new_new_n16157__, new_new_n16158__,
    new_new_n16159__, new_new_n16160__, new_new_n16161__, new_new_n16162__,
    new_new_n16163__, new_new_n16164__, new_new_n16165__, new_new_n16166__,
    new_new_n16167__, new_new_n16168__, new_new_n16169__, new_new_n16170__,
    new_new_n16171__, new_new_n16172__, new_new_n16173__, new_new_n16174__,
    new_new_n16175__, new_new_n16176__, new_new_n16177__, new_new_n16178__,
    new_new_n16179__, new_new_n16180__, new_new_n16181__, new_new_n16182__,
    new_new_n16183__, new_new_n16184__, new_new_n16185__, new_new_n16186__,
    new_new_n16187__, new_new_n16188__, new_new_n16189__, new_new_n16190__,
    new_new_n16191__, new_new_n16192__, new_new_n16193__, new_new_n16194__,
    new_new_n16195__, new_new_n16196__, new_new_n16197__, new_new_n16198__,
    new_new_n16199__, new_new_n16200__, new_new_n16201__, new_new_n16202__,
    new_new_n16203__, new_new_n16204__, new_new_n16205__, new_new_n16206__,
    new_new_n16207__, new_new_n16208__, new_new_n16209__, new_new_n16210__,
    new_new_n16211__, new_new_n16212__, new_new_n16213__, new_new_n16214__,
    new_new_n16215__, new_new_n16216__, new_new_n16217__, new_new_n16218__,
    new_new_n16219__, new_new_n16220__, new_new_n16221__, new_new_n16222__,
    new_new_n16223__, new_new_n16224__, new_new_n16225__, new_new_n16226__,
    new_new_n16227__, new_new_n16228__, new_new_n16229__, new_new_n16230__,
    new_new_n16231__, new_new_n16232__, new_new_n16233__, new_new_n16234__,
    new_new_n16236__, new_new_n16237__, new_new_n16238__, new_new_n16239__,
    new_new_n16240__, new_new_n16241__, new_new_n16242__, new_new_n16243__,
    new_new_n16244__, new_new_n16245__, new_new_n16246__, new_new_n16247__,
    new_new_n16248__, new_new_n16249__, new_new_n16250__, new_new_n16251__,
    new_new_n16252__, new_new_n16253__, new_new_n16254__, new_new_n16255__,
    new_new_n16256__, new_new_n16257__, new_new_n16258__, new_new_n16259__,
    new_new_n16260__, new_new_n16261__, new_new_n16262__, new_new_n16263__,
    new_new_n16264__, new_new_n16265__, new_new_n16266__, new_new_n16267__,
    new_new_n16268__, new_new_n16269__, new_new_n16270__, new_new_n16271__,
    new_new_n16272__, new_new_n16273__, new_new_n16274__, new_new_n16275__,
    new_new_n16276__, new_new_n16277__, new_new_n16278__, new_new_n16279__,
    new_new_n16280__, new_new_n16281__, new_new_n16282__, new_new_n16283__,
    new_new_n16284__, new_new_n16285__, new_new_n16286__, new_new_n16287__,
    new_new_n16288__, new_new_n16289__, new_new_n16290__, new_new_n16291__,
    new_new_n16292__, new_new_n16293__, new_new_n16294__, new_new_n16295__,
    new_new_n16296__, new_new_n16297__, new_new_n16298__, new_new_n16299__,
    new_new_n16300__, new_new_n16301__, new_new_n16302__, new_new_n16303__,
    new_new_n16304__, new_new_n16305__, new_new_n16306__, new_new_n16307__,
    new_new_n16308__, new_new_n16309__, new_new_n16310__, new_new_n16311__,
    new_new_n16312__, new_new_n16313__, new_new_n16314__, new_new_n16315__,
    new_new_n16316__, new_new_n16317__, new_new_n16318__, new_new_n16319__,
    new_new_n16320__, new_new_n16321__, new_new_n16322__, new_new_n16323__,
    new_new_n16324__, new_new_n16325__, new_new_n16326__, new_new_n16327__,
    new_new_n16328__, new_new_n16329__, new_new_n16330__, new_new_n16331__,
    new_new_n16332__, new_new_n16333__, new_new_n16334__, new_new_n16335__,
    new_new_n16336__, new_new_n16337__, new_new_n16338__, new_new_n16339__,
    new_new_n16340__, new_new_n16341__, new_new_n16342__, new_new_n16343__,
    new_new_n16344__, new_new_n16345__, new_new_n16346__, new_new_n16347__,
    new_new_n16348__, new_new_n16349__, new_new_n16350__, new_new_n16351__,
    new_new_n16352__, new_new_n16353__, new_new_n16354__, new_new_n16355__,
    new_new_n16356__, new_new_n16357__, new_new_n16358__, new_new_n16359__,
    new_new_n16360__, new_new_n16361__, new_new_n16362__, new_new_n16363__,
    new_new_n16364__, new_new_n16365__, new_new_n16366__, new_new_n16367__,
    new_new_n16368__, new_new_n16369__, new_new_n16370__, new_new_n16371__,
    new_new_n16372__, new_new_n16373__, new_new_n16374__, new_new_n16375__,
    new_new_n16376__, new_new_n16377__, new_new_n16378__, new_new_n16379__,
    new_new_n16380__, new_new_n16381__, new_new_n16382__, new_new_n16383__,
    new_new_n16384__, new_new_n16385__, new_new_n16386__, new_new_n16387__,
    new_new_n16388__, new_new_n16389__, new_new_n16390__, new_new_n16391__,
    new_new_n16392__, new_new_n16393__, new_new_n16394__, new_new_n16395__,
    new_new_n16396__, new_new_n16397__, new_new_n16398__, new_new_n16399__,
    new_new_n16400__, new_new_n16401__, new_new_n16402__, new_new_n16403__,
    new_new_n16404__, new_new_n16405__, new_new_n16406__, new_new_n16407__,
    new_new_n16408__, new_new_n16409__, new_new_n16410__, new_new_n16411__,
    new_new_n16412__, new_new_n16413__, new_new_n16414__, new_new_n16415__,
    new_new_n16416__, new_new_n16417__, new_new_n16418__, new_new_n16419__,
    new_new_n16420__, new_new_n16421__, new_new_n16422__, new_new_n16423__,
    new_new_n16424__, new_new_n16425__, new_new_n16426__, new_new_n16427__,
    new_new_n16428__, new_new_n16429__, new_new_n16430__, new_new_n16431__,
    new_new_n16432__, new_new_n16433__, new_new_n16434__, new_new_n16435__,
    new_new_n16436__, new_new_n16437__, new_new_n16438__, new_new_n16439__,
    new_new_n16440__, new_new_n16441__, new_new_n16442__, new_new_n16443__,
    new_new_n16444__, new_new_n16445__, new_new_n16446__, new_new_n16447__,
    new_new_n16448__, new_new_n16449__, new_new_n16450__, new_new_n16451__,
    new_new_n16452__, new_new_n16453__, new_new_n16454__, new_new_n16455__,
    new_new_n16456__, new_new_n16457__, new_new_n16458__, new_new_n16459__,
    new_new_n16460__, new_new_n16461__, new_new_n16462__, new_new_n16463__,
    new_new_n16464__, new_new_n16465__, new_new_n16466__, new_new_n16467__,
    new_new_n16468__, new_new_n16469__, new_new_n16470__, new_new_n16471__,
    new_new_n16472__, new_new_n16473__, new_new_n16474__, new_new_n16475__,
    new_new_n16476__, new_new_n16477__, new_new_n16478__, new_new_n16479__,
    new_new_n16480__, new_new_n16481__, new_new_n16482__, new_new_n16483__,
    new_new_n16484__, new_new_n16485__, new_new_n16486__, new_new_n16487__,
    new_new_n16488__, new_new_n16489__, new_new_n16490__, new_new_n16491__,
    new_new_n16492__, new_new_n16493__, new_new_n16494__, new_new_n16495__,
    new_new_n16496__, new_new_n16497__, new_new_n16498__, new_new_n16499__,
    new_new_n16500__, new_new_n16501__, new_new_n16502__, new_new_n16503__,
    new_new_n16504__, new_new_n16505__, new_new_n16506__, new_new_n16507__,
    new_new_n16508__, new_new_n16509__, new_new_n16510__, new_new_n16511__,
    new_new_n16512__, new_new_n16513__, new_new_n16514__, new_new_n16515__,
    new_new_n16516__, new_new_n16517__, new_new_n16518__, new_new_n16519__,
    new_new_n16520__, new_new_n16521__, new_new_n16522__, new_new_n16523__,
    new_new_n16524__, new_new_n16525__, new_new_n16526__, new_new_n16527__,
    new_new_n16528__, new_new_n16529__, new_new_n16530__, new_new_n16531__,
    new_new_n16532__, new_new_n16533__, new_new_n16534__, new_new_n16535__,
    new_new_n16536__, new_new_n16537__, new_new_n16538__, new_new_n16539__,
    new_new_n16540__, new_new_n16541__, new_new_n16542__, new_new_n16543__,
    new_new_n16544__, new_new_n16545__, new_new_n16546__, new_new_n16547__,
    new_new_n16548__, new_new_n16549__, new_new_n16550__, new_new_n16551__,
    new_new_n16552__, new_new_n16553__, new_new_n16554__, new_new_n16555__,
    new_new_n16556__, new_new_n16557__, new_new_n16558__, new_new_n16559__,
    new_new_n16560__, new_new_n16561__, new_new_n16562__, new_new_n16563__,
    new_new_n16564__, new_new_n16565__, new_new_n16566__, new_new_n16567__,
    new_new_n16568__, new_new_n16569__, new_new_n16570__, new_new_n16571__,
    new_new_n16572__, new_new_n16573__, new_new_n16574__, new_new_n16575__,
    new_new_n16576__, new_new_n16577__, new_new_n16578__, new_new_n16579__,
    new_new_n16580__, new_new_n16581__, new_new_n16582__, new_new_n16583__,
    new_new_n16584__, new_new_n16585__, new_new_n16586__, new_new_n16587__,
    new_new_n16588__, new_new_n16589__, new_new_n16590__, new_new_n16591__,
    new_new_n16592__, new_new_n16593__, new_new_n16594__, new_new_n16595__,
    new_new_n16596__, new_new_n16597__, new_new_n16598__, new_new_n16599__,
    new_new_n16600__, new_new_n16601__, new_new_n16602__, new_new_n16603__,
    new_new_n16604__, new_new_n16605__, new_new_n16606__, new_new_n16607__,
    new_new_n16608__, new_new_n16609__, new_new_n16610__, new_new_n16611__,
    new_new_n16612__, new_new_n16613__, new_new_n16614__, new_new_n16615__,
    new_new_n16616__, new_new_n16617__, new_new_n16618__, new_new_n16619__,
    new_new_n16620__, new_new_n16621__, new_new_n16622__, new_new_n16623__,
    new_new_n16624__, new_new_n16625__, new_new_n16626__, new_new_n16627__,
    new_new_n16628__, new_new_n16629__, new_new_n16630__, new_new_n16631__,
    new_new_n16632__, new_new_n16633__, new_new_n16634__, new_new_n16635__,
    new_new_n16636__, new_new_n16637__, new_new_n16638__, new_new_n16639__,
    new_new_n16640__, new_new_n16641__, new_new_n16642__, new_new_n16643__,
    new_new_n16644__, new_new_n16645__, new_new_n16646__, new_new_n16647__,
    new_new_n16648__, new_new_n16649__, new_new_n16650__, new_new_n16651__,
    new_new_n16652__, new_new_n16653__, new_new_n16654__, new_new_n16655__,
    new_new_n16656__, new_new_n16657__, new_new_n16658__, new_new_n16659__,
    new_new_n16660__, new_new_n16661__, new_new_n16662__, new_new_n16663__,
    new_new_n16664__, new_new_n16665__, new_new_n16666__, new_new_n16667__,
    new_new_n16668__, new_new_n16669__, new_new_n16670__, new_new_n16671__,
    new_new_n16672__, new_new_n16673__, new_new_n16674__, new_new_n16675__,
    new_new_n16676__, new_new_n16677__, new_new_n16678__, new_new_n16679__,
    new_new_n16680__, new_new_n16681__, new_new_n16682__, new_new_n16683__,
    new_new_n16684__, new_new_n16685__, new_new_n16686__, new_new_n16687__,
    new_new_n16688__, new_new_n16689__, new_new_n16690__, new_new_n16691__,
    new_new_n16692__, new_new_n16693__, new_new_n16694__, new_new_n16695__,
    new_new_n16696__, new_new_n16697__, new_new_n16698__, new_new_n16699__,
    new_new_n16700__, new_new_n16701__, new_new_n16702__, new_new_n16703__,
    new_new_n16704__, new_new_n16705__, new_new_n16706__, new_new_n16707__,
    new_new_n16708__, new_new_n16709__, new_new_n16710__, new_new_n16711__,
    new_new_n16712__, new_new_n16713__, new_new_n16714__, new_new_n16715__,
    new_new_n16716__, new_new_n16717__, new_new_n16718__, new_new_n16719__,
    new_new_n16720__, new_new_n16721__, new_new_n16722__, new_new_n16723__,
    new_new_n16724__, new_new_n16725__, new_new_n16726__, new_new_n16727__,
    new_new_n16728__, new_new_n16729__, new_new_n16730__, new_new_n16731__,
    new_new_n16732__, new_new_n16733__, new_new_n16734__, new_new_n16735__,
    new_new_n16736__, new_new_n16737__, new_new_n16738__, new_new_n16739__,
    new_new_n16740__, new_new_n16741__, new_new_n16742__, new_new_n16743__,
    new_new_n16744__, new_new_n16745__, new_new_n16746__, new_new_n16747__,
    new_new_n16748__, new_new_n16749__, new_new_n16750__, new_new_n16751__,
    new_new_n16752__, new_new_n16753__, new_new_n16754__, new_new_n16755__,
    new_new_n16756__, new_new_n16757__, new_new_n16758__, new_new_n16759__,
    new_new_n16760__, new_new_n16761__, new_new_n16762__, new_new_n16763__,
    new_new_n16764__, new_new_n16765__, new_new_n16766__, new_new_n16767__,
    new_new_n16768__, new_new_n16769__, new_new_n16770__, new_new_n16771__,
    new_new_n16772__, new_new_n16773__, new_new_n16774__, new_new_n16775__,
    new_new_n16776__, new_new_n16777__, new_new_n16778__, new_new_n16779__,
    new_new_n16780__, new_new_n16781__, new_new_n16782__, new_new_n16783__,
    new_new_n16784__, new_new_n16785__, new_new_n16786__, new_new_n16787__,
    new_new_n16788__, new_new_n16789__, new_new_n16790__, new_new_n16791__,
    new_new_n16792__, new_new_n16793__, new_new_n16794__, new_new_n16795__,
    new_new_n16796__, new_new_n16797__, new_new_n16798__, new_new_n16799__,
    new_new_n16800__, new_new_n16801__, new_new_n16802__, new_new_n16803__,
    new_new_n16804__, new_new_n16805__, new_new_n16806__, new_new_n16807__,
    new_new_n16808__, new_new_n16809__, new_new_n16810__, new_new_n16811__,
    new_new_n16812__, new_new_n16813__, new_new_n16814__, new_new_n16815__,
    new_new_n16816__, new_new_n16817__, new_new_n16818__, new_new_n16819__,
    new_new_n16820__, new_new_n16821__, new_new_n16822__, new_new_n16823__,
    new_new_n16824__, new_new_n16825__, new_new_n16826__, new_new_n16827__,
    new_new_n16828__, new_new_n16829__, new_new_n16830__, new_new_n16831__,
    new_new_n16832__, new_new_n16834__, new_new_n16835__, new_new_n16836__,
    new_new_n16837__, new_new_n16838__, new_new_n16839__, new_new_n16840__,
    new_new_n16841__, new_new_n16842__, new_new_n16843__, new_new_n16844__,
    new_new_n16845__, new_new_n16846__, new_new_n16847__, new_new_n16848__,
    new_new_n16849__, new_new_n16850__, new_new_n16851__, new_new_n16852__,
    new_new_n16853__, new_new_n16854__, new_new_n16855__, new_new_n16856__,
    new_new_n16857__, new_new_n16858__, new_new_n16859__, new_new_n16860__,
    new_new_n16861__, new_new_n16862__, new_new_n16863__, new_new_n16864__,
    new_new_n16865__, new_new_n16866__, new_new_n16867__, new_new_n16868__,
    new_new_n16869__, new_new_n16870__, new_new_n16871__, new_new_n16872__,
    new_new_n16873__, new_new_n16874__, new_new_n16875__, new_new_n16876__,
    new_new_n16877__, new_new_n16878__, new_new_n16879__, new_new_n16880__,
    new_new_n16881__, new_new_n16882__, new_new_n16883__, new_new_n16884__,
    new_new_n16885__, new_new_n16886__, new_new_n16887__, new_new_n16888__,
    new_new_n16889__, new_new_n16890__, new_new_n16891__, new_new_n16892__,
    new_new_n16893__, new_new_n16894__, new_new_n16895__, new_new_n16896__,
    new_new_n16897__, new_new_n16898__, new_new_n16899__, new_new_n16900__,
    new_new_n16901__, new_new_n16902__, new_new_n16903__, new_new_n16904__,
    new_new_n16905__, new_new_n16906__, new_new_n16907__, new_new_n16908__,
    new_new_n16909__, new_new_n16910__, new_new_n16911__, new_new_n16912__,
    new_new_n16913__, new_new_n16914__, new_new_n16915__, new_new_n16916__,
    new_new_n16917__, new_new_n16918__, new_new_n16919__, new_new_n16920__,
    new_new_n16921__, new_new_n16922__, new_new_n16923__, new_new_n16924__,
    new_new_n16925__, new_new_n16926__, new_new_n16927__, new_new_n16928__,
    new_new_n16929__, new_new_n16930__, new_new_n16931__, new_new_n16932__,
    new_new_n16933__, new_new_n16934__, new_new_n16935__, new_new_n16936__,
    new_new_n16937__, new_new_n16938__, new_new_n16939__, new_new_n16940__,
    new_new_n16941__, new_new_n16942__, new_new_n16943__, new_new_n16944__,
    new_new_n16945__, new_new_n16946__, new_new_n16947__, new_new_n16948__,
    new_new_n16949__, new_new_n16950__, new_new_n16951__, new_new_n16952__,
    new_new_n16953__, new_new_n16954__, new_new_n16955__, new_new_n16956__,
    new_new_n16957__, new_new_n16958__, new_new_n16959__, new_new_n16960__,
    new_new_n16961__, new_new_n16962__, new_new_n16963__, new_new_n16964__,
    new_new_n16965__, new_new_n16966__, new_new_n16967__, new_new_n16968__,
    new_new_n16969__, new_new_n16970__, new_new_n16971__, new_new_n16972__,
    new_new_n16973__, new_new_n16974__, new_new_n16975__, new_new_n16976__,
    new_new_n16977__, new_new_n16978__, new_new_n16979__, new_new_n16980__,
    new_new_n16981__, new_new_n16982__, new_new_n16983__, new_new_n16984__,
    new_new_n16985__, new_new_n16986__, new_new_n16987__, new_new_n16988__,
    new_new_n16989__, new_new_n16990__, new_new_n16991__, new_new_n16992__,
    new_new_n16993__, new_new_n16994__, new_new_n16995__, new_new_n16996__,
    new_new_n16997__, new_new_n16998__, new_new_n16999__, new_new_n17000__,
    new_new_n17001__, new_new_n17002__, new_new_n17003__, new_new_n17004__,
    new_new_n17005__, new_new_n17006__, new_new_n17007__, new_new_n17008__,
    new_new_n17009__, new_new_n17010__, new_new_n17011__, new_new_n17012__,
    new_new_n17013__, new_new_n17014__, new_new_n17015__, new_new_n17016__,
    new_new_n17017__, new_new_n17018__, new_new_n17019__, new_new_n17020__,
    new_new_n17021__, new_new_n17022__, new_new_n17023__, new_new_n17024__,
    new_new_n17025__, new_new_n17026__, new_new_n17027__, new_new_n17028__,
    new_new_n17029__, new_new_n17030__, new_new_n17031__, new_new_n17032__,
    new_new_n17033__, new_new_n17034__, new_new_n17035__, new_new_n17036__,
    new_new_n17037__, new_new_n17038__, new_new_n17039__, new_new_n17040__,
    new_new_n17041__, new_new_n17042__, new_new_n17043__, new_new_n17044__,
    new_new_n17045__, new_new_n17046__, new_new_n17047__, new_new_n17048__,
    new_new_n17049__, new_new_n17050__, new_new_n17051__, new_new_n17052__,
    new_new_n17053__, new_new_n17054__, new_new_n17055__, new_new_n17056__,
    new_new_n17057__, new_new_n17058__, new_new_n17059__, new_new_n17060__,
    new_new_n17061__, new_new_n17062__, new_new_n17063__, new_new_n17064__,
    new_new_n17065__, new_new_n17066__, new_new_n17067__, new_new_n17068__,
    new_new_n17069__, new_new_n17070__, new_new_n17071__, new_new_n17072__,
    new_new_n17073__, new_new_n17074__, new_new_n17075__, new_new_n17076__,
    new_new_n17077__, new_new_n17078__, new_new_n17079__, new_new_n17080__,
    new_new_n17081__, new_new_n17082__, new_new_n17083__, new_new_n17084__,
    new_new_n17085__, new_new_n17086__, new_new_n17087__, new_new_n17088__,
    new_new_n17089__, new_new_n17090__, new_new_n17091__, new_new_n17092__,
    new_new_n17093__, new_new_n17094__, new_new_n17095__, new_new_n17096__,
    new_new_n17097__, new_new_n17098__, new_new_n17099__, new_new_n17100__,
    new_new_n17101__, new_new_n17102__, new_new_n17103__, new_new_n17104__,
    new_new_n17105__, new_new_n17106__, new_new_n17107__, new_new_n17108__,
    new_new_n17109__, new_new_n17110__, new_new_n17111__, new_new_n17112__,
    new_new_n17113__, new_new_n17114__, new_new_n17115__, new_new_n17116__,
    new_new_n17117__, new_new_n17118__, new_new_n17119__, new_new_n17120__,
    new_new_n17121__, new_new_n17122__, new_new_n17123__, new_new_n17124__,
    new_new_n17125__, new_new_n17126__, new_new_n17127__, new_new_n17128__,
    new_new_n17129__, new_new_n17130__, new_new_n17131__, new_new_n17132__,
    new_new_n17133__, new_new_n17134__, new_new_n17135__, new_new_n17136__,
    new_new_n17137__, new_new_n17138__, new_new_n17139__, new_new_n17140__,
    new_new_n17141__, new_new_n17142__, new_new_n17143__, new_new_n17144__,
    new_new_n17145__, new_new_n17146__, new_new_n17147__, new_new_n17148__,
    new_new_n17149__, new_new_n17150__, new_new_n17151__, new_new_n17152__,
    new_new_n17153__, new_new_n17154__, new_new_n17155__, new_new_n17156__,
    new_new_n17157__, new_new_n17158__, new_new_n17159__, new_new_n17160__,
    new_new_n17161__, new_new_n17162__, new_new_n17163__, new_new_n17164__,
    new_new_n17165__, new_new_n17166__, new_new_n17167__, new_new_n17168__,
    new_new_n17169__, new_new_n17170__, new_new_n17171__, new_new_n17172__,
    new_new_n17173__, new_new_n17174__, new_new_n17175__, new_new_n17176__,
    new_new_n17177__, new_new_n17178__, new_new_n17179__, new_new_n17180__,
    new_new_n17181__, new_new_n17182__, new_new_n17183__, new_new_n17184__,
    new_new_n17185__, new_new_n17186__, new_new_n17187__, new_new_n17188__,
    new_new_n17189__, new_new_n17190__, new_new_n17191__, new_new_n17192__,
    new_new_n17193__, new_new_n17194__, new_new_n17195__, new_new_n17196__,
    new_new_n17197__, new_new_n17198__, new_new_n17199__, new_new_n17200__,
    new_new_n17201__, new_new_n17202__, new_new_n17203__, new_new_n17204__,
    new_new_n17205__, new_new_n17206__, new_new_n17207__, new_new_n17208__,
    new_new_n17209__, new_new_n17210__, new_new_n17211__, new_new_n17212__,
    new_new_n17213__, new_new_n17214__, new_new_n17215__, new_new_n17216__,
    new_new_n17217__, new_new_n17218__, new_new_n17219__, new_new_n17220__,
    new_new_n17221__, new_new_n17222__, new_new_n17223__, new_new_n17224__,
    new_new_n17225__, new_new_n17226__, new_new_n17227__, new_new_n17228__,
    new_new_n17229__, new_new_n17230__, new_new_n17231__, new_new_n17232__,
    new_new_n17233__, new_new_n17234__, new_new_n17235__, new_new_n17236__,
    new_new_n17237__, new_new_n17238__, new_new_n17239__, new_new_n17240__,
    new_new_n17241__, new_new_n17242__, new_new_n17243__, new_new_n17244__,
    new_new_n17245__, new_new_n17246__, new_new_n17247__, new_new_n17248__,
    new_new_n17249__, new_new_n17250__, new_new_n17251__, new_new_n17252__,
    new_new_n17253__, new_new_n17254__, new_new_n17255__, new_new_n17256__,
    new_new_n17257__, new_new_n17258__, new_new_n17259__, new_new_n17260__,
    new_new_n17261__, new_new_n17262__, new_new_n17263__, new_new_n17264__,
    new_new_n17265__, new_new_n17266__, new_new_n17267__, new_new_n17268__,
    new_new_n17269__, new_new_n17270__, new_new_n17271__, new_new_n17272__,
    new_new_n17273__, new_new_n17274__, new_new_n17275__, new_new_n17276__,
    new_new_n17277__, new_new_n17278__, new_new_n17279__, new_new_n17280__,
    new_new_n17281__, new_new_n17282__, new_new_n17283__, new_new_n17284__,
    new_new_n17285__, new_new_n17286__, new_new_n17287__, new_new_n17288__,
    new_new_n17289__, new_new_n17290__, new_new_n17291__, new_new_n17292__,
    new_new_n17293__, new_new_n17294__, new_new_n17295__, new_new_n17296__,
    new_new_n17297__, new_new_n17298__, new_new_n17299__, new_new_n17300__,
    new_new_n17301__, new_new_n17302__, new_new_n17303__, new_new_n17304__,
    new_new_n17305__, new_new_n17306__, new_new_n17307__, new_new_n17308__,
    new_new_n17309__, new_new_n17310__, new_new_n17311__, new_new_n17312__,
    new_new_n17313__, new_new_n17314__, new_new_n17315__, new_new_n17316__,
    new_new_n17317__, new_new_n17318__, new_new_n17319__, new_new_n17320__,
    new_new_n17321__, new_new_n17322__, new_new_n17323__, new_new_n17324__,
    new_new_n17325__, new_new_n17326__, new_new_n17327__, new_new_n17328__,
    new_new_n17329__, new_new_n17330__, new_new_n17331__, new_new_n17332__,
    new_new_n17333__, new_new_n17334__, new_new_n17335__, new_new_n17336__,
    new_new_n17337__, new_new_n17338__, new_new_n17339__, new_new_n17340__,
    new_new_n17341__, new_new_n17342__, new_new_n17343__, new_new_n17344__,
    new_new_n17345__, new_new_n17346__, new_new_n17347__, new_new_n17348__,
    new_new_n17349__, new_new_n17350__, new_new_n17351__, new_new_n17352__,
    new_new_n17353__, new_new_n17354__, new_new_n17355__, new_new_n17356__,
    new_new_n17357__, new_new_n17358__, new_new_n17359__, new_new_n17360__,
    new_new_n17361__, new_new_n17362__, new_new_n17363__, new_new_n17364__,
    new_new_n17365__, new_new_n17366__, new_new_n17367__, new_new_n17368__,
    new_new_n17369__, new_new_n17370__, new_new_n17371__, new_new_n17372__,
    new_new_n17373__, new_new_n17374__, new_new_n17375__, new_new_n17376__,
    new_new_n17377__, new_new_n17378__, new_new_n17379__, new_new_n17380__,
    new_new_n17381__, new_new_n17382__, new_new_n17383__, new_new_n17384__,
    new_new_n17385__, new_new_n17386__, new_new_n17387__, new_new_n17388__,
    new_new_n17389__, new_new_n17390__, new_new_n17391__, new_new_n17392__,
    new_new_n17393__, new_new_n17394__, new_new_n17395__, new_new_n17396__,
    new_new_n17397__, new_new_n17398__, new_new_n17399__, new_new_n17400__,
    new_new_n17401__, new_new_n17402__, new_new_n17403__, new_new_n17404__,
    new_new_n17405__, new_new_n17406__, new_new_n17407__, new_new_n17408__,
    new_new_n17409__, new_new_n17410__, new_new_n17411__, new_new_n17412__,
    new_new_n17413__, new_new_n17414__, new_new_n17415__, new_new_n17416__,
    new_new_n17417__, new_new_n17418__, new_new_n17419__, new_new_n17420__,
    new_new_n17421__, new_new_n17422__, new_new_n17423__, new_new_n17424__,
    new_new_n17425__, new_new_n17426__, new_new_n17427__, new_new_n17428__,
    new_new_n17429__, new_new_n17430__, new_new_n17431__, new_new_n17432__,
    new_new_n17433__, new_new_n17434__, new_new_n17435__, new_new_n17436__,
    new_new_n17437__, new_new_n17438__, new_new_n17439__, new_new_n17440__,
    new_new_n17441__, new_new_n17442__, new_new_n17443__, new_new_n17444__,
    new_new_n17445__, new_new_n17446__, new_new_n17447__, new_new_n17448__,
    new_new_n17449__, new_new_n17450__, new_new_n17451__, new_new_n17452__,
    new_new_n17453__, new_new_n17454__, new_new_n17455__, new_new_n17456__,
    new_new_n17457__, new_new_n17458__, new_new_n17459__, new_new_n17461__,
    new_new_n17462__, new_new_n17463__, new_new_n17464__, new_new_n17465__,
    new_new_n17466__, new_new_n17467__, new_new_n17468__, new_new_n17469__,
    new_new_n17470__, new_new_n17471__, new_new_n17472__, new_new_n17473__,
    new_new_n17474__, new_new_n17475__, new_new_n17476__, new_new_n17477__,
    new_new_n17478__, new_new_n17479__, new_new_n17480__, new_new_n17481__,
    new_new_n17482__, new_new_n17483__, new_new_n17484__, new_new_n17485__,
    new_new_n17486__, new_new_n17487__, new_new_n17488__, new_new_n17489__,
    new_new_n17490__, new_new_n17491__, new_new_n17492__, new_new_n17493__,
    new_new_n17494__, new_new_n17495__, new_new_n17496__, new_new_n17497__,
    new_new_n17498__, new_new_n17499__, new_new_n17500__, new_new_n17501__,
    new_new_n17502__, new_new_n17503__, new_new_n17504__, new_new_n17505__,
    new_new_n17506__, new_new_n17507__, new_new_n17508__, new_new_n17509__,
    new_new_n17510__, new_new_n17511__, new_new_n17512__, new_new_n17513__,
    new_new_n17514__, new_new_n17515__, new_new_n17516__, new_new_n17517__,
    new_new_n17518__, new_new_n17519__, new_new_n17520__, new_new_n17521__,
    new_new_n17522__, new_new_n17523__, new_new_n17524__, new_new_n17525__,
    new_new_n17526__, new_new_n17527__, new_new_n17528__, new_new_n17529__,
    new_new_n17530__, new_new_n17531__, new_new_n17532__, new_new_n17533__,
    new_new_n17534__, new_new_n17535__, new_new_n17536__, new_new_n17537__,
    new_new_n17538__, new_new_n17539__, new_new_n17540__, new_new_n17541__,
    new_new_n17542__, new_new_n17543__, new_new_n17544__, new_new_n17545__,
    new_new_n17546__, new_new_n17547__, new_new_n17548__, new_new_n17549__,
    new_new_n17550__, new_new_n17551__, new_new_n17552__, new_new_n17553__,
    new_new_n17554__, new_new_n17555__, new_new_n17556__, new_new_n17557__,
    new_new_n17558__, new_new_n17559__, new_new_n17560__, new_new_n17561__,
    new_new_n17562__, new_new_n17563__, new_new_n17564__, new_new_n17565__,
    new_new_n17566__, new_new_n17567__, new_new_n17568__, new_new_n17569__,
    new_new_n17570__, new_new_n17571__, new_new_n17572__, new_new_n17573__,
    new_new_n17574__, new_new_n17575__, new_new_n17576__, new_new_n17577__,
    new_new_n17578__, new_new_n17579__, new_new_n17580__, new_new_n17581__,
    new_new_n17582__, new_new_n17583__, new_new_n17584__, new_new_n17585__,
    new_new_n17586__, new_new_n17587__, new_new_n17588__, new_new_n17589__,
    new_new_n17590__, new_new_n17591__, new_new_n17592__, new_new_n17593__,
    new_new_n17594__, new_new_n17595__, new_new_n17596__, new_new_n17597__,
    new_new_n17598__, new_new_n17599__, new_new_n17600__, new_new_n17601__,
    new_new_n17602__, new_new_n17603__, new_new_n17604__, new_new_n17605__,
    new_new_n17606__, new_new_n17607__, new_new_n17608__, new_new_n17609__,
    new_new_n17610__, new_new_n17611__, new_new_n17612__, new_new_n17613__,
    new_new_n17614__, new_new_n17615__, new_new_n17616__, new_new_n17617__,
    new_new_n17618__, new_new_n17619__, new_new_n17620__, new_new_n17621__,
    new_new_n17622__, new_new_n17623__, new_new_n17624__, new_new_n17625__,
    new_new_n17626__, new_new_n17627__, new_new_n17628__, new_new_n17629__,
    new_new_n17630__, new_new_n17631__, new_new_n17632__, new_new_n17633__,
    new_new_n17634__, new_new_n17635__, new_new_n17636__, new_new_n17637__,
    new_new_n17638__, new_new_n17639__, new_new_n17640__, new_new_n17641__,
    new_new_n17642__, new_new_n17643__, new_new_n17644__, new_new_n17645__,
    new_new_n17646__, new_new_n17647__, new_new_n17648__, new_new_n17649__,
    new_new_n17650__, new_new_n17651__, new_new_n17652__, new_new_n17653__,
    new_new_n17654__, new_new_n17655__, new_new_n17656__, new_new_n17657__,
    new_new_n17658__, new_new_n17659__, new_new_n17660__, new_new_n17661__,
    new_new_n17662__, new_new_n17663__, new_new_n17664__, new_new_n17665__,
    new_new_n17666__, new_new_n17667__, new_new_n17668__, new_new_n17669__,
    new_new_n17670__, new_new_n17671__, new_new_n17672__, new_new_n17673__,
    new_new_n17674__, new_new_n17675__, new_new_n17676__, new_new_n17677__,
    new_new_n17678__, new_new_n17679__, new_new_n17680__, new_new_n17681__,
    new_new_n17682__, new_new_n17683__, new_new_n17684__, new_new_n17685__,
    new_new_n17686__, new_new_n17687__, new_new_n17688__, new_new_n17689__,
    new_new_n17690__, new_new_n17691__, new_new_n17692__, new_new_n17693__,
    new_new_n17694__, new_new_n17695__, new_new_n17696__, new_new_n17697__,
    new_new_n17698__, new_new_n17699__, new_new_n17700__, new_new_n17701__,
    new_new_n17702__, new_new_n17703__, new_new_n17704__, new_new_n17705__,
    new_new_n17706__, new_new_n17707__, new_new_n17708__, new_new_n17709__,
    new_new_n17710__, new_new_n17711__, new_new_n17712__, new_new_n17713__,
    new_new_n17714__, new_new_n17715__, new_new_n17716__, new_new_n17717__,
    new_new_n17718__, new_new_n17719__, new_new_n17720__, new_new_n17721__,
    new_new_n17722__, new_new_n17723__, new_new_n17724__, new_new_n17725__,
    new_new_n17726__, new_new_n17727__, new_new_n17728__, new_new_n17729__,
    new_new_n17730__, new_new_n17731__, new_new_n17732__, new_new_n17733__,
    new_new_n17734__, new_new_n17735__, new_new_n17736__, new_new_n17737__,
    new_new_n17738__, new_new_n17739__, new_new_n17740__, new_new_n17741__,
    new_new_n17742__, new_new_n17743__, new_new_n17744__, new_new_n17745__,
    new_new_n17746__, new_new_n17747__, new_new_n17748__, new_new_n17749__,
    new_new_n17750__, new_new_n17751__, new_new_n17752__, new_new_n17753__,
    new_new_n17754__, new_new_n17755__, new_new_n17756__, new_new_n17757__,
    new_new_n17758__, new_new_n17759__, new_new_n17760__, new_new_n17761__,
    new_new_n17762__, new_new_n17763__, new_new_n17764__, new_new_n17765__,
    new_new_n17766__, new_new_n17767__, new_new_n17768__, new_new_n17769__,
    new_new_n17770__, new_new_n17771__, new_new_n17772__, new_new_n17773__,
    new_new_n17774__, new_new_n17775__, new_new_n17776__, new_new_n17777__,
    new_new_n17778__, new_new_n17779__, new_new_n17780__, new_new_n17781__,
    new_new_n17782__, new_new_n17783__, new_new_n17784__, new_new_n17785__,
    new_new_n17786__, new_new_n17787__, new_new_n17788__, new_new_n17789__,
    new_new_n17790__, new_new_n17791__, new_new_n17792__, new_new_n17793__,
    new_new_n17794__, new_new_n17795__, new_new_n17796__, new_new_n17797__,
    new_new_n17798__, new_new_n17799__, new_new_n17800__, new_new_n17801__,
    new_new_n17802__, new_new_n17803__, new_new_n17804__, new_new_n17805__,
    new_new_n17806__, new_new_n17807__, new_new_n17808__, new_new_n17809__,
    new_new_n17810__, new_new_n17811__, new_new_n17812__, new_new_n17813__,
    new_new_n17814__, new_new_n17815__, new_new_n17816__, new_new_n17817__,
    new_new_n17818__, new_new_n17819__, new_new_n17820__, new_new_n17821__,
    new_new_n17822__, new_new_n17823__, new_new_n17824__, new_new_n17825__,
    new_new_n17826__, new_new_n17827__, new_new_n17828__, new_new_n17829__,
    new_new_n17830__, new_new_n17831__, new_new_n17832__, new_new_n17833__,
    new_new_n17834__, new_new_n17835__, new_new_n17836__, new_new_n17837__,
    new_new_n17838__, new_new_n17839__, new_new_n17840__, new_new_n17841__,
    new_new_n17842__, new_new_n17843__, new_new_n17844__, new_new_n17845__,
    new_new_n17846__, new_new_n17847__, new_new_n17848__, new_new_n17849__,
    new_new_n17850__, new_new_n17851__, new_new_n17852__, new_new_n17853__,
    new_new_n17854__, new_new_n17855__, new_new_n17856__, new_new_n17857__,
    new_new_n17858__, new_new_n17859__, new_new_n17860__, new_new_n17861__,
    new_new_n17862__, new_new_n17863__, new_new_n17864__, new_new_n17865__,
    new_new_n17866__, new_new_n17867__, new_new_n17868__, new_new_n17869__,
    new_new_n17870__, new_new_n17871__, new_new_n17872__, new_new_n17873__,
    new_new_n17874__, new_new_n17875__, new_new_n17876__, new_new_n17877__,
    new_new_n17878__, new_new_n17879__, new_new_n17880__, new_new_n17881__,
    new_new_n17882__, new_new_n17883__, new_new_n17884__, new_new_n17885__,
    new_new_n17886__, new_new_n17887__, new_new_n17888__, new_new_n17889__,
    new_new_n17890__, new_new_n17891__, new_new_n17892__, new_new_n17893__,
    new_new_n17894__, new_new_n17895__, new_new_n17896__, new_new_n17897__,
    new_new_n17898__, new_new_n17899__, new_new_n17900__, new_new_n17901__,
    new_new_n17902__, new_new_n17903__, new_new_n17904__, new_new_n17905__,
    new_new_n17906__, new_new_n17907__, new_new_n17908__, new_new_n17909__,
    new_new_n17910__, new_new_n17911__, new_new_n17912__, new_new_n17913__,
    new_new_n17914__, new_new_n17915__, new_new_n17916__, new_new_n17917__,
    new_new_n17918__, new_new_n17919__, new_new_n17920__, new_new_n17921__,
    new_new_n17922__, new_new_n17923__, new_new_n17924__, new_new_n17925__,
    new_new_n17926__, new_new_n17927__, new_new_n17928__, new_new_n17929__,
    new_new_n17930__, new_new_n17931__, new_new_n17932__, new_new_n17933__,
    new_new_n17934__, new_new_n17935__, new_new_n17936__, new_new_n17937__,
    new_new_n17938__, new_new_n17939__, new_new_n17940__, new_new_n17941__,
    new_new_n17942__, new_new_n17943__, new_new_n17944__, new_new_n17945__,
    new_new_n17946__, new_new_n17947__, new_new_n17948__, new_new_n17949__,
    new_new_n17950__, new_new_n17951__, new_new_n17952__, new_new_n17953__,
    new_new_n17954__, new_new_n17955__, new_new_n17956__, new_new_n17957__,
    new_new_n17958__, new_new_n17959__, new_new_n17960__, new_new_n17961__,
    new_new_n17962__, new_new_n17963__, new_new_n17964__, new_new_n17965__,
    new_new_n17966__, new_new_n17967__, new_new_n17968__, new_new_n17969__,
    new_new_n17970__, new_new_n17971__, new_new_n17972__, new_new_n17973__,
    new_new_n17974__, new_new_n17975__, new_new_n17976__, new_new_n17977__,
    new_new_n17978__, new_new_n17979__, new_new_n17980__, new_new_n17981__,
    new_new_n17982__, new_new_n17983__, new_new_n17984__, new_new_n17985__,
    new_new_n17986__, new_new_n17987__, new_new_n17988__, new_new_n17989__,
    new_new_n17990__, new_new_n17991__, new_new_n17992__, new_new_n17993__,
    new_new_n17994__, new_new_n17995__, new_new_n17996__, new_new_n17997__,
    new_new_n17998__, new_new_n17999__, new_new_n18000__, new_new_n18001__,
    new_new_n18002__, new_new_n18003__, new_new_n18004__, new_new_n18005__,
    new_new_n18006__, new_new_n18007__, new_new_n18008__, new_new_n18009__,
    new_new_n18010__, new_new_n18011__, new_new_n18012__, new_new_n18013__,
    new_new_n18014__, new_new_n18015__, new_new_n18016__, new_new_n18017__,
    new_new_n18018__, new_new_n18019__, new_new_n18020__, new_new_n18021__,
    new_new_n18022__, new_new_n18023__, new_new_n18024__, new_new_n18025__,
    new_new_n18026__, new_new_n18027__, new_new_n18028__, new_new_n18029__,
    new_new_n18030__, new_new_n18031__, new_new_n18032__, new_new_n18033__,
    new_new_n18034__, new_new_n18035__, new_new_n18036__, new_new_n18037__,
    new_new_n18038__, new_new_n18039__, new_new_n18040__, new_new_n18041__,
    new_new_n18042__, new_new_n18043__, new_new_n18044__, new_new_n18045__,
    new_new_n18046__, new_new_n18047__, new_new_n18048__, new_new_n18049__,
    new_new_n18050__, new_new_n18051__, new_new_n18052__, new_new_n18053__,
    new_new_n18054__, new_new_n18055__, new_new_n18056__, new_new_n18057__,
    new_new_n18058__, new_new_n18059__, new_new_n18060__, new_new_n18061__,
    new_new_n18062__, new_new_n18063__, new_new_n18064__, new_new_n18065__,
    new_new_n18066__, new_new_n18067__, new_new_n18068__, new_new_n18069__,
    new_new_n18070__, new_new_n18071__, new_new_n18072__, new_new_n18073__,
    new_new_n18074__, new_new_n18075__, new_new_n18076__, new_new_n18077__,
    new_new_n18078__, new_new_n18079__, new_new_n18080__, new_new_n18081__,
    new_new_n18082__, new_new_n18083__, new_new_n18084__, new_new_n18085__,
    new_new_n18086__, new_new_n18087__, new_new_n18089__, new_new_n18090__,
    new_new_n18091__, new_new_n18092__, new_new_n18093__, new_new_n18094__,
    new_new_n18095__, new_new_n18096__, new_new_n18097__, new_new_n18098__,
    new_new_n18099__, new_new_n18100__, new_new_n18101__, new_new_n18102__,
    new_new_n18103__, new_new_n18104__, new_new_n18105__, new_new_n18106__,
    new_new_n18107__, new_new_n18108__, new_new_n18109__, new_new_n18110__,
    new_new_n18111__, new_new_n18112__, new_new_n18113__, new_new_n18114__,
    new_new_n18115__, new_new_n18116__, new_new_n18117__, new_new_n18118__,
    new_new_n18119__, new_new_n18120__, new_new_n18121__, new_new_n18122__,
    new_new_n18123__, new_new_n18124__, new_new_n18125__, new_new_n18126__,
    new_new_n18127__, new_new_n18128__, new_new_n18129__, new_new_n18130__,
    new_new_n18131__, new_new_n18132__, new_new_n18133__, new_new_n18134__,
    new_new_n18135__, new_new_n18136__, new_new_n18137__, new_new_n18138__,
    new_new_n18139__, new_new_n18140__, new_new_n18141__, new_new_n18142__,
    new_new_n18143__, new_new_n18144__, new_new_n18145__, new_new_n18146__,
    new_new_n18147__, new_new_n18148__, new_new_n18149__, new_new_n18150__,
    new_new_n18151__, new_new_n18152__, new_new_n18153__, new_new_n18154__,
    new_new_n18155__, new_new_n18156__, new_new_n18157__, new_new_n18158__,
    new_new_n18159__, new_new_n18160__, new_new_n18161__, new_new_n18162__,
    new_new_n18163__, new_new_n18164__, new_new_n18165__, new_new_n18166__,
    new_new_n18167__, new_new_n18168__, new_new_n18169__, new_new_n18170__,
    new_new_n18171__, new_new_n18172__, new_new_n18173__, new_new_n18174__,
    new_new_n18175__, new_new_n18176__, new_new_n18177__, new_new_n18178__,
    new_new_n18179__, new_new_n18180__, new_new_n18181__, new_new_n18182__,
    new_new_n18183__, new_new_n18184__, new_new_n18185__, new_new_n18186__,
    new_new_n18187__, new_new_n18188__, new_new_n18189__, new_new_n18190__,
    new_new_n18191__, new_new_n18192__, new_new_n18193__, new_new_n18194__,
    new_new_n18195__, new_new_n18196__, new_new_n18197__, new_new_n18198__,
    new_new_n18199__, new_new_n18200__, new_new_n18201__, new_new_n18202__,
    new_new_n18203__, new_new_n18204__, new_new_n18205__, new_new_n18206__,
    new_new_n18207__, new_new_n18208__, new_new_n18209__, new_new_n18210__,
    new_new_n18211__, new_new_n18212__, new_new_n18213__, new_new_n18214__,
    new_new_n18215__, new_new_n18216__, new_new_n18217__, new_new_n18218__,
    new_new_n18219__, new_new_n18220__, new_new_n18221__, new_new_n18222__,
    new_new_n18223__, new_new_n18224__, new_new_n18225__, new_new_n18226__,
    new_new_n18227__, new_new_n18228__, new_new_n18229__, new_new_n18230__,
    new_new_n18231__, new_new_n18232__, new_new_n18233__, new_new_n18234__,
    new_new_n18235__, new_new_n18236__, new_new_n18237__, new_new_n18238__,
    new_new_n18239__, new_new_n18240__, new_new_n18241__, new_new_n18242__,
    new_new_n18243__, new_new_n18244__, new_new_n18245__, new_new_n18246__,
    new_new_n18247__, new_new_n18248__, new_new_n18249__, new_new_n18250__,
    new_new_n18251__, new_new_n18252__, new_new_n18253__, new_new_n18254__,
    new_new_n18255__, new_new_n18256__, new_new_n18257__, new_new_n18258__,
    new_new_n18259__, new_new_n18260__, new_new_n18261__, new_new_n18262__,
    new_new_n18263__, new_new_n18264__, new_new_n18265__, new_new_n18266__,
    new_new_n18267__, new_new_n18268__, new_new_n18269__, new_new_n18270__,
    new_new_n18271__, new_new_n18272__, new_new_n18273__, new_new_n18274__,
    new_new_n18275__, new_new_n18276__, new_new_n18277__, new_new_n18278__,
    new_new_n18279__, new_new_n18280__, new_new_n18281__, new_new_n18282__,
    new_new_n18283__, new_new_n18284__, new_new_n18285__, new_new_n18286__,
    new_new_n18287__, new_new_n18288__, new_new_n18289__, new_new_n18290__,
    new_new_n18291__, new_new_n18292__, new_new_n18293__, new_new_n18294__,
    new_new_n18295__, new_new_n18296__, new_new_n18297__, new_new_n18298__,
    new_new_n18299__, new_new_n18300__, new_new_n18301__, new_new_n18302__,
    new_new_n18303__, new_new_n18304__, new_new_n18305__, new_new_n18306__,
    new_new_n18307__, new_new_n18308__, new_new_n18309__, new_new_n18310__,
    new_new_n18311__, new_new_n18312__, new_new_n18313__, new_new_n18314__,
    new_new_n18315__, new_new_n18316__, new_new_n18317__, new_new_n18318__,
    new_new_n18319__, new_new_n18320__, new_new_n18321__, new_new_n18322__,
    new_new_n18323__, new_new_n18324__, new_new_n18325__, new_new_n18326__,
    new_new_n18327__, new_new_n18328__, new_new_n18329__, new_new_n18330__,
    new_new_n18331__, new_new_n18332__, new_new_n18333__, new_new_n18334__,
    new_new_n18335__, new_new_n18336__, new_new_n18337__, new_new_n18338__,
    new_new_n18339__, new_new_n18340__, new_new_n18341__, new_new_n18342__,
    new_new_n18343__, new_new_n18344__, new_new_n18345__, new_new_n18346__,
    new_new_n18347__, new_new_n18348__, new_new_n18349__, new_new_n18350__,
    new_new_n18351__, new_new_n18352__, new_new_n18353__, new_new_n18354__,
    new_new_n18355__, new_new_n18356__, new_new_n18357__, new_new_n18358__,
    new_new_n18359__, new_new_n18360__, new_new_n18361__, new_new_n18362__,
    new_new_n18363__, new_new_n18364__, new_new_n18365__, new_new_n18366__,
    new_new_n18367__, new_new_n18368__, new_new_n18369__, new_new_n18370__,
    new_new_n18371__, new_new_n18372__, new_new_n18373__, new_new_n18374__,
    new_new_n18375__, new_new_n18376__, new_new_n18377__, new_new_n18378__,
    new_new_n18379__, new_new_n18380__, new_new_n18381__, new_new_n18382__,
    new_new_n18383__, new_new_n18384__, new_new_n18385__, new_new_n18386__,
    new_new_n18387__, new_new_n18388__, new_new_n18389__, new_new_n18390__,
    new_new_n18391__, new_new_n18392__, new_new_n18393__, new_new_n18394__,
    new_new_n18395__, new_new_n18396__, new_new_n18397__, new_new_n18398__,
    new_new_n18399__, new_new_n18400__, new_new_n18401__, new_new_n18402__,
    new_new_n18403__, new_new_n18404__, new_new_n18405__, new_new_n18406__,
    new_new_n18407__, new_new_n18408__, new_new_n18409__, new_new_n18410__,
    new_new_n18411__, new_new_n18412__, new_new_n18413__, new_new_n18414__,
    new_new_n18415__, new_new_n18416__, new_new_n18417__, new_new_n18418__,
    new_new_n18419__, new_new_n18420__, new_new_n18421__, new_new_n18422__,
    new_new_n18423__, new_new_n18424__, new_new_n18425__, new_new_n18426__,
    new_new_n18427__, new_new_n18428__, new_new_n18429__, new_new_n18430__,
    new_new_n18431__, new_new_n18432__, new_new_n18433__, new_new_n18434__,
    new_new_n18435__, new_new_n18436__, new_new_n18437__, new_new_n18438__,
    new_new_n18439__, new_new_n18440__, new_new_n18441__, new_new_n18442__,
    new_new_n18443__, new_new_n18444__, new_new_n18445__, new_new_n18446__,
    new_new_n18447__, new_new_n18448__, new_new_n18449__, new_new_n18450__,
    new_new_n18451__, new_new_n18452__, new_new_n18453__, new_new_n18454__,
    new_new_n18455__, new_new_n18456__, new_new_n18457__, new_new_n18458__,
    new_new_n18459__, new_new_n18460__, new_new_n18461__, new_new_n18462__,
    new_new_n18463__, new_new_n18464__, new_new_n18465__, new_new_n18466__,
    new_new_n18467__, new_new_n18468__, new_new_n18469__, new_new_n18470__,
    new_new_n18471__, new_new_n18472__, new_new_n18473__, new_new_n18474__,
    new_new_n18475__, new_new_n18476__, new_new_n18477__, new_new_n18478__,
    new_new_n18479__, new_new_n18480__, new_new_n18481__, new_new_n18482__,
    new_new_n18483__, new_new_n18484__, new_new_n18485__, new_new_n18486__,
    new_new_n18487__, new_new_n18488__, new_new_n18489__, new_new_n18490__,
    new_new_n18491__, new_new_n18492__, new_new_n18493__, new_new_n18494__,
    new_new_n18495__, new_new_n18496__, new_new_n18497__, new_new_n18498__,
    new_new_n18499__, new_new_n18500__, new_new_n18501__, new_new_n18502__,
    new_new_n18503__, new_new_n18504__, new_new_n18505__, new_new_n18506__,
    new_new_n18507__, new_new_n18508__, new_new_n18509__, new_new_n18510__,
    new_new_n18511__, new_new_n18512__, new_new_n18513__, new_new_n18514__,
    new_new_n18515__, new_new_n18516__, new_new_n18517__, new_new_n18518__,
    new_new_n18519__, new_new_n18520__, new_new_n18521__, new_new_n18522__,
    new_new_n18523__, new_new_n18524__, new_new_n18525__, new_new_n18526__,
    new_new_n18527__, new_new_n18528__, new_new_n18529__, new_new_n18530__,
    new_new_n18531__, new_new_n18532__, new_new_n18533__, new_new_n18534__,
    new_new_n18535__, new_new_n18536__, new_new_n18537__, new_new_n18538__,
    new_new_n18539__, new_new_n18540__, new_new_n18541__, new_new_n18542__,
    new_new_n18543__, new_new_n18544__, new_new_n18545__, new_new_n18546__,
    new_new_n18547__, new_new_n18548__, new_new_n18549__, new_new_n18550__,
    new_new_n18551__, new_new_n18552__, new_new_n18553__, new_new_n18554__,
    new_new_n18555__, new_new_n18556__, new_new_n18557__, new_new_n18558__,
    new_new_n18559__, new_new_n18560__, new_new_n18561__, new_new_n18562__,
    new_new_n18563__, new_new_n18564__, new_new_n18565__, new_new_n18566__,
    new_new_n18567__, new_new_n18568__, new_new_n18569__, new_new_n18570__,
    new_new_n18571__, new_new_n18572__, new_new_n18573__, new_new_n18574__,
    new_new_n18575__, new_new_n18576__, new_new_n18577__, new_new_n18578__,
    new_new_n18579__, new_new_n18580__, new_new_n18581__, new_new_n18582__,
    new_new_n18583__, new_new_n18584__, new_new_n18585__, new_new_n18586__,
    new_new_n18587__, new_new_n18588__, new_new_n18589__, new_new_n18590__,
    new_new_n18591__, new_new_n18592__, new_new_n18593__, new_new_n18594__,
    new_new_n18595__, new_new_n18596__, new_new_n18597__, new_new_n18598__,
    new_new_n18599__, new_new_n18600__, new_new_n18601__, new_new_n18602__,
    new_new_n18603__, new_new_n18604__, new_new_n18605__, new_new_n18606__,
    new_new_n18607__, new_new_n18608__, new_new_n18609__, new_new_n18610__,
    new_new_n18611__, new_new_n18612__, new_new_n18613__, new_new_n18614__,
    new_new_n18615__, new_new_n18616__, new_new_n18617__, new_new_n18618__,
    new_new_n18619__, new_new_n18620__, new_new_n18621__, new_new_n18622__,
    new_new_n18623__, new_new_n18624__, new_new_n18625__, new_new_n18626__,
    new_new_n18627__, new_new_n18628__, new_new_n18629__, new_new_n18630__,
    new_new_n18631__, new_new_n18632__, new_new_n18633__, new_new_n18634__,
    new_new_n18635__, new_new_n18636__, new_new_n18637__, new_new_n18638__,
    new_new_n18639__, new_new_n18640__, new_new_n18641__, new_new_n18642__,
    new_new_n18643__, new_new_n18644__, new_new_n18645__, new_new_n18646__,
    new_new_n18647__, new_new_n18648__, new_new_n18649__, new_new_n18650__,
    new_new_n18651__, new_new_n18652__, new_new_n18653__, new_new_n18654__,
    new_new_n18655__, new_new_n18656__, new_new_n18657__, new_new_n18658__,
    new_new_n18659__, new_new_n18660__, new_new_n18661__, new_new_n18662__,
    new_new_n18663__, new_new_n18664__, new_new_n18665__, new_new_n18666__,
    new_new_n18667__, new_new_n18668__, new_new_n18669__, new_new_n18670__,
    new_new_n18671__, new_new_n18672__, new_new_n18673__, new_new_n18674__,
    new_new_n18675__, new_new_n18676__, new_new_n18677__, new_new_n18678__,
    new_new_n18679__, new_new_n18680__, new_new_n18681__, new_new_n18682__,
    new_new_n18683__, new_new_n18684__, new_new_n18685__, new_new_n18686__,
    new_new_n18687__, new_new_n18688__, new_new_n18689__, new_new_n18690__,
    new_new_n18691__, new_new_n18692__, new_new_n18693__, new_new_n18694__,
    new_new_n18695__, new_new_n18696__, new_new_n18697__, new_new_n18698__,
    new_new_n18699__, new_new_n18700__, new_new_n18701__, new_new_n18702__,
    new_new_n18703__, new_new_n18704__, new_new_n18705__, new_new_n18706__,
    new_new_n18707__, new_new_n18708__, new_new_n18709__, new_new_n18710__,
    new_new_n18711__, new_new_n18712__, new_new_n18713__, new_new_n18714__,
    new_new_n18715__, new_new_n18716__, new_new_n18717__, new_new_n18718__,
    new_new_n18719__, new_new_n18720__, new_new_n18721__, new_new_n18722__,
    new_new_n18723__, new_new_n18724__, new_new_n18726__, new_new_n18727__,
    new_new_n18728__, new_new_n18729__, new_new_n18730__, new_new_n18731__,
    new_new_n18732__, new_new_n18733__, new_new_n18734__, new_new_n18735__,
    new_new_n18736__, new_new_n18737__, new_new_n18738__, new_new_n18739__,
    new_new_n18740__, new_new_n18741__, new_new_n18742__, new_new_n18743__,
    new_new_n18744__, new_new_n18745__, new_new_n18746__, new_new_n18747__,
    new_new_n18748__, new_new_n18749__, new_new_n18750__, new_new_n18751__,
    new_new_n18752__, new_new_n18753__, new_new_n18754__, new_new_n18755__,
    new_new_n18756__, new_new_n18757__, new_new_n18758__, new_new_n18759__,
    new_new_n18760__, new_new_n18761__, new_new_n18762__, new_new_n18763__,
    new_new_n18764__, new_new_n18765__, new_new_n18766__, new_new_n18767__,
    new_new_n18768__, new_new_n18769__, new_new_n18770__, new_new_n18771__,
    new_new_n18772__, new_new_n18773__, new_new_n18774__, new_new_n18775__,
    new_new_n18776__, new_new_n18777__, new_new_n18778__, new_new_n18779__,
    new_new_n18780__, new_new_n18781__, new_new_n18782__, new_new_n18783__,
    new_new_n18784__, new_new_n18785__, new_new_n18786__, new_new_n18787__,
    new_new_n18788__, new_new_n18789__, new_new_n18790__, new_new_n18791__,
    new_new_n18792__, new_new_n18793__, new_new_n18794__, new_new_n18795__,
    new_new_n18796__, new_new_n18797__, new_new_n18798__, new_new_n18799__,
    new_new_n18800__, new_new_n18801__, new_new_n18802__, new_new_n18803__,
    new_new_n18804__, new_new_n18805__, new_new_n18806__, new_new_n18807__,
    new_new_n18808__, new_new_n18809__, new_new_n18810__, new_new_n18811__,
    new_new_n18812__, new_new_n18813__, new_new_n18814__, new_new_n18815__,
    new_new_n18816__, new_new_n18817__, new_new_n18818__, new_new_n18819__,
    new_new_n18820__, new_new_n18821__, new_new_n18822__, new_new_n18823__,
    new_new_n18824__, new_new_n18825__, new_new_n18826__, new_new_n18827__,
    new_new_n18828__, new_new_n18829__, new_new_n18830__, new_new_n18831__,
    new_new_n18832__, new_new_n18833__, new_new_n18834__, new_new_n18835__,
    new_new_n18836__, new_new_n18837__, new_new_n18838__, new_new_n18839__,
    new_new_n18840__, new_new_n18841__, new_new_n18842__, new_new_n18843__,
    new_new_n18844__, new_new_n18845__, new_new_n18846__, new_new_n18847__,
    new_new_n18848__, new_new_n18849__, new_new_n18850__, new_new_n18851__,
    new_new_n18852__, new_new_n18853__, new_new_n18854__, new_new_n18855__,
    new_new_n18856__, new_new_n18857__, new_new_n18858__, new_new_n18859__,
    new_new_n18860__, new_new_n18861__, new_new_n18862__, new_new_n18863__,
    new_new_n18864__, new_new_n18865__, new_new_n18866__, new_new_n18867__,
    new_new_n18868__, new_new_n18869__, new_new_n18870__, new_new_n18871__,
    new_new_n18872__, new_new_n18873__, new_new_n18874__, new_new_n18875__,
    new_new_n18876__, new_new_n18877__, new_new_n18878__, new_new_n18879__,
    new_new_n18880__, new_new_n18881__, new_new_n18882__, new_new_n18883__,
    new_new_n18884__, new_new_n18885__, new_new_n18886__, new_new_n18887__,
    new_new_n18888__, new_new_n18889__, new_new_n18890__, new_new_n18891__,
    new_new_n18892__, new_new_n18893__, new_new_n18894__, new_new_n18895__,
    new_new_n18896__, new_new_n18897__, new_new_n18898__, new_new_n18899__,
    new_new_n18900__, new_new_n18901__, new_new_n18902__, new_new_n18903__,
    new_new_n18904__, new_new_n18905__, new_new_n18906__, new_new_n18907__,
    new_new_n18908__, new_new_n18909__, new_new_n18910__, new_new_n18911__,
    new_new_n18912__, new_new_n18913__, new_new_n18914__, new_new_n18915__,
    new_new_n18916__, new_new_n18917__, new_new_n18918__, new_new_n18919__,
    new_new_n18920__, new_new_n18921__, new_new_n18922__, new_new_n18923__,
    new_new_n18924__, new_new_n18925__, new_new_n18926__, new_new_n18927__,
    new_new_n18928__, new_new_n18929__, new_new_n18930__, new_new_n18931__,
    new_new_n18932__, new_new_n18933__, new_new_n18934__, new_new_n18935__,
    new_new_n18936__, new_new_n18937__, new_new_n18938__, new_new_n18939__,
    new_new_n18940__, new_new_n18941__, new_new_n18942__, new_new_n18943__,
    new_new_n18944__, new_new_n18945__, new_new_n18946__, new_new_n18947__,
    new_new_n18948__, new_new_n18949__, new_new_n18950__, new_new_n18951__,
    new_new_n18952__, new_new_n18953__, new_new_n18954__, new_new_n18955__,
    new_new_n18956__, new_new_n18957__, new_new_n18958__, new_new_n18959__,
    new_new_n18960__, new_new_n18961__, new_new_n18962__, new_new_n18963__,
    new_new_n18964__, new_new_n18965__, new_new_n18966__, new_new_n18967__,
    new_new_n18968__, new_new_n18969__, new_new_n18970__, new_new_n18971__,
    new_new_n18972__, new_new_n18973__, new_new_n18974__, new_new_n18975__,
    new_new_n18976__, new_new_n18977__, new_new_n18978__, new_new_n18979__,
    new_new_n18980__, new_new_n18981__, new_new_n18982__, new_new_n18983__,
    new_new_n18984__, new_new_n18985__, new_new_n18986__, new_new_n18987__,
    new_new_n18988__, new_new_n18989__, new_new_n18990__, new_new_n18991__,
    new_new_n18992__, new_new_n18993__, new_new_n18994__, new_new_n18995__,
    new_new_n18996__, new_new_n18997__, new_new_n18998__, new_new_n18999__,
    new_new_n19000__, new_new_n19001__, new_new_n19002__, new_new_n19003__,
    new_new_n19004__, new_new_n19005__, new_new_n19006__, new_new_n19007__,
    new_new_n19008__, new_new_n19009__, new_new_n19010__, new_new_n19011__,
    new_new_n19012__, new_new_n19013__, new_new_n19014__, new_new_n19015__,
    new_new_n19016__, new_new_n19017__, new_new_n19018__, new_new_n19019__,
    new_new_n19020__, new_new_n19021__, new_new_n19022__, new_new_n19023__,
    new_new_n19024__, new_new_n19025__, new_new_n19026__, new_new_n19027__,
    new_new_n19028__, new_new_n19029__, new_new_n19030__, new_new_n19031__,
    new_new_n19032__, new_new_n19033__, new_new_n19034__, new_new_n19035__,
    new_new_n19036__, new_new_n19037__, new_new_n19038__, new_new_n19039__,
    new_new_n19040__, new_new_n19041__, new_new_n19042__, new_new_n19043__,
    new_new_n19044__, new_new_n19045__, new_new_n19046__, new_new_n19047__,
    new_new_n19048__, new_new_n19049__, new_new_n19050__, new_new_n19051__,
    new_new_n19052__, new_new_n19053__, new_new_n19054__, new_new_n19055__,
    new_new_n19056__, new_new_n19057__, new_new_n19058__, new_new_n19059__,
    new_new_n19060__, new_new_n19061__, new_new_n19062__, new_new_n19063__,
    new_new_n19064__, new_new_n19065__, new_new_n19066__, new_new_n19067__,
    new_new_n19068__, new_new_n19069__, new_new_n19070__, new_new_n19071__,
    new_new_n19072__, new_new_n19073__, new_new_n19074__, new_new_n19075__,
    new_new_n19076__, new_new_n19077__, new_new_n19078__, new_new_n19079__,
    new_new_n19080__, new_new_n19081__, new_new_n19082__, new_new_n19083__,
    new_new_n19084__, new_new_n19085__, new_new_n19086__, new_new_n19087__,
    new_new_n19088__, new_new_n19089__, new_new_n19090__, new_new_n19091__,
    new_new_n19092__, new_new_n19093__, new_new_n19094__, new_new_n19095__,
    new_new_n19096__, new_new_n19097__, new_new_n19098__, new_new_n19099__,
    new_new_n19100__, new_new_n19101__, new_new_n19102__, new_new_n19103__,
    new_new_n19104__, new_new_n19105__, new_new_n19106__, new_new_n19107__,
    new_new_n19108__, new_new_n19109__, new_new_n19110__, new_new_n19111__,
    new_new_n19112__, new_new_n19113__, new_new_n19114__, new_new_n19115__,
    new_new_n19116__, new_new_n19117__, new_new_n19118__, new_new_n19119__,
    new_new_n19120__, new_new_n19121__, new_new_n19122__, new_new_n19123__,
    new_new_n19124__, new_new_n19125__, new_new_n19126__, new_new_n19127__,
    new_new_n19128__, new_new_n19129__, new_new_n19130__, new_new_n19131__,
    new_new_n19132__, new_new_n19133__, new_new_n19134__, new_new_n19135__,
    new_new_n19136__, new_new_n19137__, new_new_n19138__, new_new_n19139__,
    new_new_n19140__, new_new_n19141__, new_new_n19142__, new_new_n19143__,
    new_new_n19144__, new_new_n19145__, new_new_n19146__, new_new_n19147__,
    new_new_n19148__, new_new_n19149__, new_new_n19150__, new_new_n19151__,
    new_new_n19152__, new_new_n19153__, new_new_n19154__, new_new_n19155__,
    new_new_n19156__, new_new_n19157__, new_new_n19158__, new_new_n19159__,
    new_new_n19160__, new_new_n19161__, new_new_n19162__, new_new_n19163__,
    new_new_n19164__, new_new_n19165__, new_new_n19166__, new_new_n19167__,
    new_new_n19168__, new_new_n19169__, new_new_n19170__, new_new_n19171__,
    new_new_n19172__, new_new_n19173__, new_new_n19174__, new_new_n19175__,
    new_new_n19176__, new_new_n19177__, new_new_n19178__, new_new_n19179__,
    new_new_n19180__, new_new_n19181__, new_new_n19182__, new_new_n19183__,
    new_new_n19184__, new_new_n19185__, new_new_n19186__, new_new_n19187__,
    new_new_n19188__, new_new_n19189__, new_new_n19190__, new_new_n19191__,
    new_new_n19192__, new_new_n19193__, new_new_n19194__, new_new_n19195__,
    new_new_n19196__, new_new_n19197__, new_new_n19198__, new_new_n19199__,
    new_new_n19200__, new_new_n19201__, new_new_n19202__, new_new_n19203__,
    new_new_n19204__, new_new_n19205__, new_new_n19206__, new_new_n19207__,
    new_new_n19208__, new_new_n19209__, new_new_n19210__, new_new_n19211__,
    new_new_n19212__, new_new_n19213__, new_new_n19214__, new_new_n19215__,
    new_new_n19216__, new_new_n19217__, new_new_n19218__, new_new_n19219__,
    new_new_n19220__, new_new_n19221__, new_new_n19222__, new_new_n19223__,
    new_new_n19224__, new_new_n19225__, new_new_n19226__, new_new_n19227__,
    new_new_n19228__, new_new_n19229__, new_new_n19230__, new_new_n19231__,
    new_new_n19232__, new_new_n19233__, new_new_n19234__, new_new_n19235__,
    new_new_n19236__, new_new_n19237__, new_new_n19238__, new_new_n19239__,
    new_new_n19240__, new_new_n19241__, new_new_n19242__, new_new_n19243__,
    new_new_n19244__, new_new_n19245__, new_new_n19246__, new_new_n19247__,
    new_new_n19248__, new_new_n19249__, new_new_n19250__, new_new_n19251__,
    new_new_n19252__, new_new_n19253__, new_new_n19254__, new_new_n19255__,
    new_new_n19256__, new_new_n19257__, new_new_n19258__, new_new_n19259__,
    new_new_n19260__, new_new_n19261__, new_new_n19262__, new_new_n19263__,
    new_new_n19264__, new_new_n19265__, new_new_n19266__, new_new_n19267__,
    new_new_n19268__, new_new_n19269__, new_new_n19270__, new_new_n19271__,
    new_new_n19272__, new_new_n19273__, new_new_n19274__, new_new_n19275__,
    new_new_n19276__, new_new_n19277__, new_new_n19278__, new_new_n19279__,
    new_new_n19280__, new_new_n19281__, new_new_n19282__, new_new_n19283__,
    new_new_n19284__, new_new_n19285__, new_new_n19286__, new_new_n19287__,
    new_new_n19288__, new_new_n19289__, new_new_n19290__, new_new_n19291__,
    new_new_n19292__, new_new_n19293__, new_new_n19294__, new_new_n19295__,
    new_new_n19296__, new_new_n19297__, new_new_n19298__, new_new_n19299__,
    new_new_n19300__, new_new_n19301__, new_new_n19302__, new_new_n19303__,
    new_new_n19304__, new_new_n19305__, new_new_n19306__, new_new_n19307__,
    new_new_n19308__, new_new_n19309__, new_new_n19310__, new_new_n19311__,
    new_new_n19312__, new_new_n19313__, new_new_n19314__, new_new_n19315__,
    new_new_n19316__, new_new_n19317__, new_new_n19318__, new_new_n19319__,
    new_new_n19320__, new_new_n19321__, new_new_n19322__, new_new_n19323__,
    new_new_n19324__, new_new_n19325__, new_new_n19326__, new_new_n19327__,
    new_new_n19328__, new_new_n19329__, new_new_n19330__, new_new_n19331__,
    new_new_n19332__, new_new_n19333__, new_new_n19334__, new_new_n19335__,
    new_new_n19336__, new_new_n19337__, new_new_n19338__, new_new_n19339__,
    new_new_n19340__, new_new_n19341__, new_new_n19342__, new_new_n19343__,
    new_new_n19344__, new_new_n19345__, new_new_n19346__, new_new_n19347__,
    new_new_n19348__, new_new_n19349__, new_new_n19350__, new_new_n19351__,
    new_new_n19352__, new_new_n19353__, new_new_n19354__, new_new_n19355__,
    new_new_n19356__, new_new_n19357__, new_new_n19358__, new_new_n19359__,
    new_new_n19360__, new_new_n19361__, new_new_n19362__, new_new_n19363__,
    new_new_n19364__, new_new_n19366__, new_new_n19367__, new_new_n19368__,
    new_new_n19369__, new_new_n19370__, new_new_n19371__, new_new_n19372__,
    new_new_n19373__, new_new_n19374__, new_new_n19375__, new_new_n19376__,
    new_new_n19377__, new_new_n19378__, new_new_n19379__, new_new_n19380__,
    new_new_n19381__, new_new_n19382__, new_new_n19383__, new_new_n19384__,
    new_new_n19385__, new_new_n19386__, new_new_n19387__, new_new_n19388__,
    new_new_n19389__, new_new_n19390__, new_new_n19391__, new_new_n19392__,
    new_new_n19393__, new_new_n19394__, new_new_n19395__, new_new_n19396__,
    new_new_n19397__, new_new_n19398__, new_new_n19399__, new_new_n19400__,
    new_new_n19401__, new_new_n19402__, new_new_n19403__, new_new_n19404__,
    new_new_n19405__, new_new_n19406__, new_new_n19407__, new_new_n19408__,
    new_new_n19409__, new_new_n19410__, new_new_n19411__, new_new_n19412__,
    new_new_n19413__, new_new_n19414__, new_new_n19415__, new_new_n19416__,
    new_new_n19417__, new_new_n19418__, new_new_n19419__, new_new_n19420__,
    new_new_n19421__, new_new_n19422__, new_new_n19423__, new_new_n19424__,
    new_new_n19425__, new_new_n19426__, new_new_n19427__, new_new_n19428__,
    new_new_n19429__, new_new_n19430__, new_new_n19431__, new_new_n19432__,
    new_new_n19433__, new_new_n19434__, new_new_n19435__, new_new_n19436__,
    new_new_n19437__, new_new_n19438__, new_new_n19439__, new_new_n19440__,
    new_new_n19441__, new_new_n19442__, new_new_n19443__, new_new_n19444__,
    new_new_n19445__, new_new_n19446__, new_new_n19447__, new_new_n19448__,
    new_new_n19449__, new_new_n19450__, new_new_n19451__, new_new_n19452__,
    new_new_n19453__, new_new_n19454__, new_new_n19455__, new_new_n19456__,
    new_new_n19457__, new_new_n19458__, new_new_n19459__, new_new_n19460__,
    new_new_n19461__, new_new_n19462__, new_new_n19463__, new_new_n19464__,
    new_new_n19465__, new_new_n19466__, new_new_n19467__, new_new_n19468__,
    new_new_n19469__, new_new_n19470__, new_new_n19471__, new_new_n19472__,
    new_new_n19473__, new_new_n19474__, new_new_n19475__, new_new_n19476__,
    new_new_n19477__, new_new_n19478__, new_new_n19479__, new_new_n19480__,
    new_new_n19481__, new_new_n19482__, new_new_n19483__, new_new_n19484__,
    new_new_n19485__, new_new_n19486__, new_new_n19487__, new_new_n19488__,
    new_new_n19489__, new_new_n19490__, new_new_n19491__, new_new_n19492__,
    new_new_n19493__, new_new_n19494__, new_new_n19495__, new_new_n19496__,
    new_new_n19497__, new_new_n19498__, new_new_n19499__, new_new_n19500__,
    new_new_n19501__, new_new_n19502__, new_new_n19503__, new_new_n19504__,
    new_new_n19505__, new_new_n19506__, new_new_n19507__, new_new_n19508__,
    new_new_n19509__, new_new_n19510__, new_new_n19511__, new_new_n19512__,
    new_new_n19513__, new_new_n19514__, new_new_n19515__, new_new_n19516__,
    new_new_n19517__, new_new_n19518__, new_new_n19519__, new_new_n19520__,
    new_new_n19521__, new_new_n19522__, new_new_n19523__, new_new_n19524__,
    new_new_n19525__, new_new_n19526__, new_new_n19527__, new_new_n19528__,
    new_new_n19529__, new_new_n19530__, new_new_n19531__, new_new_n19532__,
    new_new_n19533__, new_new_n19534__, new_new_n19535__, new_new_n19536__,
    new_new_n19537__, new_new_n19538__, new_new_n19539__, new_new_n19540__,
    new_new_n19541__, new_new_n19542__, new_new_n19543__, new_new_n19544__,
    new_new_n19545__, new_new_n19546__, new_new_n19547__, new_new_n19548__,
    new_new_n19549__, new_new_n19550__, new_new_n19551__, new_new_n19552__,
    new_new_n19553__, new_new_n19554__, new_new_n19555__, new_new_n19556__,
    new_new_n19557__, new_new_n19558__, new_new_n19559__, new_new_n19560__,
    new_new_n19561__, new_new_n19562__, new_new_n19563__, new_new_n19564__,
    new_new_n19565__, new_new_n19566__, new_new_n19567__, new_new_n19568__,
    new_new_n19569__, new_new_n19570__, new_new_n19571__, new_new_n19572__,
    new_new_n19573__, new_new_n19574__, new_new_n19575__, new_new_n19576__,
    new_new_n19577__, new_new_n19578__, new_new_n19579__, new_new_n19580__,
    new_new_n19581__, new_new_n19582__, new_new_n19583__, new_new_n19584__,
    new_new_n19585__, new_new_n19586__, new_new_n19587__, new_new_n19588__,
    new_new_n19589__, new_new_n19590__, new_new_n19591__, new_new_n19592__,
    new_new_n19593__, new_new_n19594__, new_new_n19595__, new_new_n19596__,
    new_new_n19597__, new_new_n19598__, new_new_n19599__, new_new_n19600__,
    new_new_n19601__, new_new_n19602__, new_new_n19603__, new_new_n19604__,
    new_new_n19605__, new_new_n19606__, new_new_n19607__, new_new_n19608__,
    new_new_n19609__, new_new_n19610__, new_new_n19611__, new_new_n19612__,
    new_new_n19613__, new_new_n19614__, new_new_n19615__, new_new_n19616__,
    new_new_n19617__, new_new_n19618__, new_new_n19619__, new_new_n19620__,
    new_new_n19621__, new_new_n19622__, new_new_n19623__, new_new_n19624__,
    new_new_n19625__, new_new_n19626__, new_new_n19627__, new_new_n19628__,
    new_new_n19629__, new_new_n19630__, new_new_n19631__, new_new_n19632__,
    new_new_n19633__, new_new_n19634__, new_new_n19635__, new_new_n19636__,
    new_new_n19637__, new_new_n19638__, new_new_n19639__, new_new_n19640__,
    new_new_n19641__, new_new_n19642__, new_new_n19643__, new_new_n19644__,
    new_new_n19645__, new_new_n19646__, new_new_n19647__, new_new_n19648__,
    new_new_n19649__, new_new_n19650__, new_new_n19651__, new_new_n19652__,
    new_new_n19653__, new_new_n19654__, new_new_n19655__, new_new_n19656__,
    new_new_n19657__, new_new_n19658__, new_new_n19659__, new_new_n19660__,
    new_new_n19661__, new_new_n19662__, new_new_n19663__, new_new_n19664__,
    new_new_n19665__, new_new_n19666__, new_new_n19667__, new_new_n19668__,
    new_new_n19669__, new_new_n19670__, new_new_n19671__, new_new_n19672__,
    new_new_n19673__, new_new_n19674__, new_new_n19675__, new_new_n19676__,
    new_new_n19677__, new_new_n19678__, new_new_n19679__, new_new_n19680__,
    new_new_n19681__, new_new_n19682__, new_new_n19683__, new_new_n19684__,
    new_new_n19685__, new_new_n19686__, new_new_n19687__, new_new_n19688__,
    new_new_n19689__, new_new_n19690__, new_new_n19691__, new_new_n19692__,
    new_new_n19693__, new_new_n19694__, new_new_n19695__, new_new_n19696__,
    new_new_n19697__, new_new_n19698__, new_new_n19699__, new_new_n19700__,
    new_new_n19701__, new_new_n19702__, new_new_n19703__, new_new_n19704__,
    new_new_n19705__, new_new_n19706__, new_new_n19707__, new_new_n19708__,
    new_new_n19709__, new_new_n19710__, new_new_n19711__, new_new_n19712__,
    new_new_n19713__, new_new_n19714__, new_new_n19715__, new_new_n19716__,
    new_new_n19717__, new_new_n19718__, new_new_n19719__, new_new_n19720__,
    new_new_n19721__, new_new_n19722__, new_new_n19723__, new_new_n19724__,
    new_new_n19725__, new_new_n19726__, new_new_n19727__, new_new_n19728__,
    new_new_n19729__, new_new_n19730__, new_new_n19731__, new_new_n19732__,
    new_new_n19733__, new_new_n19734__, new_new_n19735__, new_new_n19736__,
    new_new_n19737__, new_new_n19738__, new_new_n19739__, new_new_n19740__,
    new_new_n19741__, new_new_n19742__, new_new_n19743__, new_new_n19744__,
    new_new_n19745__, new_new_n19746__, new_new_n19747__, new_new_n19748__,
    new_new_n19749__, new_new_n19750__, new_new_n19751__, new_new_n19752__,
    new_new_n19753__, new_new_n19754__, new_new_n19755__, new_new_n19756__,
    new_new_n19757__, new_new_n19758__, new_new_n19759__, new_new_n19760__,
    new_new_n19761__, new_new_n19762__, new_new_n19763__, new_new_n19764__,
    new_new_n19765__, new_new_n19766__, new_new_n19767__, new_new_n19768__,
    new_new_n19769__, new_new_n19770__, new_new_n19771__, new_new_n19772__,
    new_new_n19773__, new_new_n19774__, new_new_n19775__, new_new_n19776__,
    new_new_n19777__, new_new_n19778__, new_new_n19779__, new_new_n19780__,
    new_new_n19781__, new_new_n19782__, new_new_n19783__, new_new_n19784__,
    new_new_n19785__, new_new_n19786__, new_new_n19787__, new_new_n19788__,
    new_new_n19789__, new_new_n19790__, new_new_n19791__, new_new_n19792__,
    new_new_n19793__, new_new_n19794__, new_new_n19795__, new_new_n19796__,
    new_new_n19797__, new_new_n19798__, new_new_n19799__, new_new_n19800__,
    new_new_n19801__, new_new_n19802__, new_new_n19803__, new_new_n19804__,
    new_new_n19805__, new_new_n19806__, new_new_n19807__, new_new_n19808__,
    new_new_n19809__, new_new_n19810__, new_new_n19811__, new_new_n19812__,
    new_new_n19813__, new_new_n19814__, new_new_n19815__, new_new_n19816__,
    new_new_n19817__, new_new_n19818__, new_new_n19819__, new_new_n19820__,
    new_new_n19821__, new_new_n19822__, new_new_n19823__, new_new_n19824__,
    new_new_n19825__, new_new_n19826__, new_new_n19827__, new_new_n19828__,
    new_new_n19829__, new_new_n19830__, new_new_n19831__, new_new_n19832__,
    new_new_n19833__, new_new_n19834__, new_new_n19835__, new_new_n19836__,
    new_new_n19837__, new_new_n19838__, new_new_n19839__, new_new_n19840__,
    new_new_n19841__, new_new_n19842__, new_new_n19843__, new_new_n19844__,
    new_new_n19845__, new_new_n19846__, new_new_n19847__, new_new_n19848__,
    new_new_n19849__, new_new_n19850__, new_new_n19851__, new_new_n19852__,
    new_new_n19853__, new_new_n19854__, new_new_n19855__, new_new_n19856__,
    new_new_n19857__, new_new_n19858__, new_new_n19859__, new_new_n19860__,
    new_new_n19861__, new_new_n19862__, new_new_n19863__, new_new_n19864__,
    new_new_n19865__, new_new_n19866__, new_new_n19867__, new_new_n19868__,
    new_new_n19869__, new_new_n19870__, new_new_n19871__, new_new_n19872__,
    new_new_n19873__, new_new_n19874__, new_new_n19875__, new_new_n19876__,
    new_new_n19877__, new_new_n19878__, new_new_n19879__, new_new_n19880__,
    new_new_n19881__, new_new_n19882__, new_new_n19883__, new_new_n19884__,
    new_new_n19885__, new_new_n19886__, new_new_n19887__, new_new_n19888__,
    new_new_n19889__, new_new_n19890__, new_new_n19891__, new_new_n19892__,
    new_new_n19893__, new_new_n19894__, new_new_n19895__, new_new_n19896__,
    new_new_n19897__, new_new_n19898__, new_new_n19899__, new_new_n19900__,
    new_new_n19901__, new_new_n19902__, new_new_n19903__, new_new_n19904__,
    new_new_n19905__, new_new_n19906__, new_new_n19907__, new_new_n19908__,
    new_new_n19909__, new_new_n19910__, new_new_n19911__, new_new_n19912__,
    new_new_n19913__, new_new_n19914__, new_new_n19915__, new_new_n19916__,
    new_new_n19917__, new_new_n19918__, new_new_n19919__, new_new_n19920__,
    new_new_n19921__, new_new_n19922__, new_new_n19923__, new_new_n19924__,
    new_new_n19925__, new_new_n19926__, new_new_n19927__, new_new_n19928__,
    new_new_n19929__, new_new_n19930__, new_new_n19931__, new_new_n19932__,
    new_new_n19933__, new_new_n19934__, new_new_n19935__, new_new_n19936__,
    new_new_n19937__, new_new_n19938__, new_new_n19939__, new_new_n19940__,
    new_new_n19941__, new_new_n19942__, new_new_n19943__, new_new_n19944__,
    new_new_n19945__, new_new_n19946__, new_new_n19947__, new_new_n19948__,
    new_new_n19949__, new_new_n19950__, new_new_n19951__, new_new_n19952__,
    new_new_n19953__, new_new_n19954__, new_new_n19955__, new_new_n19956__,
    new_new_n19957__, new_new_n19958__, new_new_n19959__, new_new_n19960__,
    new_new_n19961__, new_new_n19962__, new_new_n19963__, new_new_n19964__,
    new_new_n19965__, new_new_n19966__, new_new_n19967__, new_new_n19968__,
    new_new_n19969__, new_new_n19970__, new_new_n19971__, new_new_n19972__,
    new_new_n19973__, new_new_n19974__, new_new_n19975__, new_new_n19976__,
    new_new_n19977__, new_new_n19978__, new_new_n19979__, new_new_n19980__,
    new_new_n19981__, new_new_n19982__, new_new_n19983__, new_new_n19984__,
    new_new_n19985__, new_new_n19986__, new_new_n19987__, new_new_n19988__,
    new_new_n19989__, new_new_n19990__, new_new_n19991__, new_new_n19992__,
    new_new_n19993__, new_new_n19994__, new_new_n19995__, new_new_n19996__,
    new_new_n19997__, new_new_n19998__, new_new_n19999__, new_new_n20000__,
    new_new_n20001__, new_new_n20002__, new_new_n20003__, new_new_n20004__,
    new_new_n20005__, new_new_n20006__, new_new_n20007__, new_new_n20008__,
    new_new_n20009__, new_new_n20010__, new_new_n20011__, new_new_n20012__,
    new_new_n20013__, new_new_n20014__, new_new_n20016__, new_new_n20017__,
    new_new_n20018__, new_new_n20019__, new_new_n20020__, new_new_n20021__,
    new_new_n20022__, new_new_n20023__, new_new_n20024__, new_new_n20025__,
    new_new_n20026__, new_new_n20027__, new_new_n20028__, new_new_n20029__,
    new_new_n20030__, new_new_n20031__, new_new_n20032__, new_new_n20033__,
    new_new_n20034__, new_new_n20035__, new_new_n20036__, new_new_n20037__,
    new_new_n20038__, new_new_n20039__, new_new_n20040__, new_new_n20041__,
    new_new_n20042__, new_new_n20043__, new_new_n20044__, new_new_n20045__,
    new_new_n20046__, new_new_n20047__, new_new_n20048__, new_new_n20049__,
    new_new_n20050__, new_new_n20051__, new_new_n20052__, new_new_n20053__,
    new_new_n20054__, new_new_n20055__, new_new_n20056__, new_new_n20057__,
    new_new_n20058__, new_new_n20059__, new_new_n20060__, new_new_n20061__,
    new_new_n20062__, new_new_n20063__, new_new_n20064__, new_new_n20065__,
    new_new_n20066__, new_new_n20067__, new_new_n20068__, new_new_n20069__,
    new_new_n20070__, new_new_n20071__, new_new_n20072__, new_new_n20073__,
    new_new_n20074__, new_new_n20075__, new_new_n20076__, new_new_n20077__,
    new_new_n20078__, new_new_n20079__, new_new_n20080__, new_new_n20081__,
    new_new_n20082__, new_new_n20083__, new_new_n20084__, new_new_n20085__,
    new_new_n20086__, new_new_n20087__, new_new_n20088__, new_new_n20089__,
    new_new_n20090__, new_new_n20091__, new_new_n20092__, new_new_n20093__,
    new_new_n20094__, new_new_n20095__, new_new_n20096__, new_new_n20097__,
    new_new_n20098__, new_new_n20099__, new_new_n20100__, new_new_n20101__,
    new_new_n20102__, new_new_n20103__, new_new_n20104__, new_new_n20105__,
    new_new_n20106__, new_new_n20107__, new_new_n20108__, new_new_n20109__,
    new_new_n20110__, new_new_n20111__, new_new_n20112__, new_new_n20113__,
    new_new_n20114__, new_new_n20115__, new_new_n20116__, new_new_n20117__,
    new_new_n20118__, new_new_n20119__, new_new_n20120__, new_new_n20121__,
    new_new_n20122__, new_new_n20123__, new_new_n20124__, new_new_n20125__,
    new_new_n20126__, new_new_n20127__, new_new_n20128__, new_new_n20129__,
    new_new_n20130__, new_new_n20131__, new_new_n20132__, new_new_n20133__,
    new_new_n20134__, new_new_n20135__, new_new_n20136__, new_new_n20137__,
    new_new_n20138__, new_new_n20139__, new_new_n20140__, new_new_n20141__,
    new_new_n20142__, new_new_n20143__, new_new_n20144__, new_new_n20145__,
    new_new_n20146__, new_new_n20147__, new_new_n20148__, new_new_n20149__,
    new_new_n20150__, new_new_n20151__, new_new_n20152__, new_new_n20153__,
    new_new_n20154__, new_new_n20155__, new_new_n20156__, new_new_n20157__,
    new_new_n20158__, new_new_n20159__, new_new_n20160__, new_new_n20161__,
    new_new_n20162__, new_new_n20163__, new_new_n20164__, new_new_n20165__,
    new_new_n20166__, new_new_n20167__, new_new_n20168__, new_new_n20169__,
    new_new_n20170__, new_new_n20171__, new_new_n20172__, new_new_n20173__,
    new_new_n20174__, new_new_n20175__, new_new_n20176__, new_new_n20177__,
    new_new_n20178__, new_new_n20179__, new_new_n20180__, new_new_n20181__,
    new_new_n20182__, new_new_n20183__, new_new_n20184__, new_new_n20185__,
    new_new_n20186__, new_new_n20187__, new_new_n20188__, new_new_n20189__,
    new_new_n20190__, new_new_n20191__, new_new_n20192__, new_new_n20193__,
    new_new_n20194__, new_new_n20195__, new_new_n20196__, new_new_n20197__,
    new_new_n20198__, new_new_n20199__, new_new_n20200__, new_new_n20201__,
    new_new_n20202__, new_new_n20203__, new_new_n20204__, new_new_n20205__,
    new_new_n20206__, new_new_n20207__, new_new_n20208__, new_new_n20209__,
    new_new_n20210__, new_new_n20211__, new_new_n20212__, new_new_n20213__,
    new_new_n20214__, new_new_n20215__, new_new_n20216__, new_new_n20217__,
    new_new_n20218__, new_new_n20219__, new_new_n20220__, new_new_n20221__,
    new_new_n20222__, new_new_n20223__, new_new_n20224__, new_new_n20225__,
    new_new_n20226__, new_new_n20227__, new_new_n20228__, new_new_n20229__,
    new_new_n20230__, new_new_n20231__, new_new_n20232__, new_new_n20233__,
    new_new_n20234__, new_new_n20235__, new_new_n20236__, new_new_n20237__,
    new_new_n20238__, new_new_n20239__, new_new_n20240__, new_new_n20241__,
    new_new_n20242__, new_new_n20243__, new_new_n20244__, new_new_n20245__,
    new_new_n20246__, new_new_n20247__, new_new_n20248__, new_new_n20249__,
    new_new_n20250__, new_new_n20251__, new_new_n20252__, new_new_n20253__,
    new_new_n20254__, new_new_n20255__, new_new_n20256__, new_new_n20257__,
    new_new_n20258__, new_new_n20259__, new_new_n20260__, new_new_n20261__,
    new_new_n20262__, new_new_n20263__, new_new_n20264__, new_new_n20265__,
    new_new_n20266__, new_new_n20267__, new_new_n20268__, new_new_n20269__,
    new_new_n20270__, new_new_n20271__, new_new_n20272__, new_new_n20273__,
    new_new_n20274__, new_new_n20275__, new_new_n20276__, new_new_n20277__,
    new_new_n20278__, new_new_n20279__, new_new_n20280__, new_new_n20281__,
    new_new_n20282__, new_new_n20283__, new_new_n20284__, new_new_n20285__,
    new_new_n20286__, new_new_n20287__, new_new_n20288__, new_new_n20289__,
    new_new_n20290__, new_new_n20291__, new_new_n20292__, new_new_n20293__,
    new_new_n20294__, new_new_n20295__, new_new_n20296__, new_new_n20297__,
    new_new_n20298__, new_new_n20299__, new_new_n20300__, new_new_n20301__,
    new_new_n20302__, new_new_n20303__, new_new_n20304__, new_new_n20305__,
    new_new_n20306__, new_new_n20307__, new_new_n20308__, new_new_n20309__,
    new_new_n20310__, new_new_n20311__, new_new_n20312__, new_new_n20313__,
    new_new_n20314__, new_new_n20315__, new_new_n20316__, new_new_n20317__,
    new_new_n20318__, new_new_n20319__, new_new_n20320__, new_new_n20321__,
    new_new_n20322__, new_new_n20323__, new_new_n20324__, new_new_n20325__,
    new_new_n20326__, new_new_n20327__, new_new_n20328__, new_new_n20329__,
    new_new_n20330__, new_new_n20331__, new_new_n20332__, new_new_n20333__,
    new_new_n20334__, new_new_n20335__, new_new_n20336__, new_new_n20337__,
    new_new_n20338__, new_new_n20339__, new_new_n20340__, new_new_n20341__,
    new_new_n20342__, new_new_n20343__, new_new_n20344__, new_new_n20345__,
    new_new_n20346__, new_new_n20347__, new_new_n20348__, new_new_n20349__,
    new_new_n20350__, new_new_n20351__, new_new_n20352__, new_new_n20353__,
    new_new_n20354__, new_new_n20355__, new_new_n20356__, new_new_n20357__,
    new_new_n20358__, new_new_n20359__, new_new_n20360__, new_new_n20361__,
    new_new_n20362__, new_new_n20363__, new_new_n20364__, new_new_n20365__,
    new_new_n20366__, new_new_n20367__, new_new_n20368__, new_new_n20369__,
    new_new_n20370__, new_new_n20371__, new_new_n20372__, new_new_n20373__,
    new_new_n20374__, new_new_n20375__, new_new_n20376__, new_new_n20377__,
    new_new_n20378__, new_new_n20379__, new_new_n20380__, new_new_n20381__,
    new_new_n20382__, new_new_n20383__, new_new_n20384__, new_new_n20385__,
    new_new_n20386__, new_new_n20387__, new_new_n20388__, new_new_n20389__,
    new_new_n20390__, new_new_n20391__, new_new_n20392__, new_new_n20393__,
    new_new_n20394__, new_new_n20395__, new_new_n20396__, new_new_n20397__,
    new_new_n20398__, new_new_n20399__, new_new_n20400__, new_new_n20401__,
    new_new_n20402__, new_new_n20403__, new_new_n20404__, new_new_n20405__,
    new_new_n20406__, new_new_n20407__, new_new_n20408__, new_new_n20409__,
    new_new_n20410__, new_new_n20411__, new_new_n20412__, new_new_n20413__,
    new_new_n20414__, new_new_n20415__, new_new_n20416__, new_new_n20417__,
    new_new_n20418__, new_new_n20419__, new_new_n20420__, new_new_n20421__,
    new_new_n20422__, new_new_n20423__, new_new_n20424__, new_new_n20425__,
    new_new_n20426__, new_new_n20427__, new_new_n20428__, new_new_n20429__,
    new_new_n20430__, new_new_n20431__, new_new_n20432__, new_new_n20433__,
    new_new_n20434__, new_new_n20435__, new_new_n20436__, new_new_n20437__,
    new_new_n20438__, new_new_n20439__, new_new_n20440__, new_new_n20441__,
    new_new_n20442__, new_new_n20443__, new_new_n20444__, new_new_n20445__,
    new_new_n20446__, new_new_n20447__, new_new_n20448__, new_new_n20449__,
    new_new_n20450__, new_new_n20451__, new_new_n20452__, new_new_n20453__,
    new_new_n20454__, new_new_n20455__, new_new_n20456__, new_new_n20457__,
    new_new_n20458__, new_new_n20459__, new_new_n20460__, new_new_n20461__,
    new_new_n20462__, new_new_n20463__, new_new_n20464__, new_new_n20465__,
    new_new_n20466__, new_new_n20467__, new_new_n20468__, new_new_n20469__,
    new_new_n20470__, new_new_n20471__, new_new_n20472__, new_new_n20473__,
    new_new_n20474__, new_new_n20475__, new_new_n20476__, new_new_n20477__,
    new_new_n20478__, new_new_n20479__, new_new_n20480__, new_new_n20481__,
    new_new_n20482__, new_new_n20483__, new_new_n20484__, new_new_n20485__,
    new_new_n20486__, new_new_n20487__, new_new_n20488__, new_new_n20489__,
    new_new_n20490__, new_new_n20491__, new_new_n20492__, new_new_n20493__,
    new_new_n20494__, new_new_n20495__, new_new_n20496__, new_new_n20497__,
    new_new_n20498__, new_new_n20499__, new_new_n20500__, new_new_n20501__,
    new_new_n20502__, new_new_n20503__, new_new_n20504__, new_new_n20505__,
    new_new_n20506__, new_new_n20507__, new_new_n20508__, new_new_n20509__,
    new_new_n20510__, new_new_n20511__, new_new_n20512__, new_new_n20513__,
    new_new_n20514__, new_new_n20515__, new_new_n20516__, new_new_n20517__,
    new_new_n20518__, new_new_n20519__, new_new_n20520__, new_new_n20521__,
    new_new_n20522__, new_new_n20523__, new_new_n20524__, new_new_n20525__,
    new_new_n20526__, new_new_n20527__, new_new_n20528__, new_new_n20529__,
    new_new_n20530__, new_new_n20531__, new_new_n20532__, new_new_n20533__,
    new_new_n20534__, new_new_n20535__, new_new_n20536__, new_new_n20537__,
    new_new_n20538__, new_new_n20539__, new_new_n20540__, new_new_n20541__,
    new_new_n20542__, new_new_n20543__, new_new_n20544__, new_new_n20545__,
    new_new_n20546__, new_new_n20547__, new_new_n20548__, new_new_n20549__,
    new_new_n20550__, new_new_n20551__, new_new_n20552__, new_new_n20553__,
    new_new_n20554__, new_new_n20555__, new_new_n20556__, new_new_n20557__,
    new_new_n20558__, new_new_n20559__, new_new_n20560__, new_new_n20561__,
    new_new_n20562__, new_new_n20563__, new_new_n20564__, new_new_n20565__,
    new_new_n20566__, new_new_n20567__, new_new_n20568__, new_new_n20569__,
    new_new_n20570__, new_new_n20571__, new_new_n20572__, new_new_n20573__,
    new_new_n20574__, new_new_n20575__, new_new_n20576__, new_new_n20577__,
    new_new_n20578__, new_new_n20579__, new_new_n20580__, new_new_n20581__,
    new_new_n20582__, new_new_n20583__, new_new_n20584__, new_new_n20585__,
    new_new_n20586__, new_new_n20587__, new_new_n20588__, new_new_n20589__,
    new_new_n20590__, new_new_n20591__, new_new_n20592__, new_new_n20593__,
    new_new_n20594__, new_new_n20595__, new_new_n20596__, new_new_n20597__,
    new_new_n20598__, new_new_n20599__, new_new_n20600__, new_new_n20601__,
    new_new_n20602__, new_new_n20603__, new_new_n20604__, new_new_n20605__,
    new_new_n20606__, new_new_n20607__, new_new_n20608__, new_new_n20609__,
    new_new_n20610__, new_new_n20611__, new_new_n20612__, new_new_n20613__,
    new_new_n20614__, new_new_n20615__, new_new_n20616__, new_new_n20617__,
    new_new_n20618__, new_new_n20619__, new_new_n20620__, new_new_n20621__,
    new_new_n20622__, new_new_n20623__, new_new_n20624__, new_new_n20625__,
    new_new_n20626__, new_new_n20627__, new_new_n20628__, new_new_n20629__,
    new_new_n20630__, new_new_n20631__, new_new_n20632__, new_new_n20633__,
    new_new_n20634__, new_new_n20635__, new_new_n20636__, new_new_n20637__,
    new_new_n20638__, new_new_n20639__, new_new_n20640__, new_new_n20641__,
    new_new_n20642__, new_new_n20643__, new_new_n20644__, new_new_n20645__,
    new_new_n20646__, new_new_n20647__, new_new_n20648__, new_new_n20649__,
    new_new_n20650__, new_new_n20651__, new_new_n20652__, new_new_n20653__,
    new_new_n20654__, new_new_n20655__, new_new_n20656__, new_new_n20657__,
    new_new_n20658__, new_new_n20659__, new_new_n20660__, new_new_n20661__,
    new_new_n20662__, new_new_n20663__, new_new_n20664__, new_new_n20665__,
    new_new_n20666__, new_new_n20667__, new_new_n20668__, new_new_n20669__,
    new_new_n20670__, new_new_n20671__, new_new_n20672__, new_new_n20673__,
    new_new_n20674__, new_new_n20675__, new_new_n20676__, new_new_n20677__,
    new_new_n20679__, new_new_n20680__, new_new_n20681__, new_new_n20682__,
    new_new_n20683__, new_new_n20684__, new_new_n20685__, new_new_n20686__,
    new_new_n20687__, new_new_n20688__, new_new_n20689__, new_new_n20690__,
    new_new_n20691__, new_new_n20692__, new_new_n20693__, new_new_n20694__,
    new_new_n20695__, new_new_n20696__, new_new_n20697__, new_new_n20698__,
    new_new_n20699__, new_new_n20700__, new_new_n20701__, new_new_n20702__,
    new_new_n20703__, new_new_n20704__, new_new_n20705__, new_new_n20706__,
    new_new_n20707__, new_new_n20708__, new_new_n20709__, new_new_n20710__,
    new_new_n20711__, new_new_n20712__, new_new_n20713__, new_new_n20714__,
    new_new_n20715__, new_new_n20716__, new_new_n20717__, new_new_n20718__,
    new_new_n20719__, new_new_n20720__, new_new_n20721__, new_new_n20722__,
    new_new_n20723__, new_new_n20724__, new_new_n20725__, new_new_n20726__,
    new_new_n20727__, new_new_n20728__, new_new_n20729__, new_new_n20730__,
    new_new_n20731__, new_new_n20732__, new_new_n20733__, new_new_n20734__,
    new_new_n20735__, new_new_n20736__, new_new_n20737__, new_new_n20738__,
    new_new_n20739__, new_new_n20740__, new_new_n20741__, new_new_n20742__,
    new_new_n20743__, new_new_n20744__, new_new_n20745__, new_new_n20746__,
    new_new_n20747__, new_new_n20748__, new_new_n20749__, new_new_n20750__,
    new_new_n20751__, new_new_n20752__, new_new_n20753__, new_new_n20754__,
    new_new_n20755__, new_new_n20756__, new_new_n20757__, new_new_n20758__,
    new_new_n20759__, new_new_n20760__, new_new_n20761__, new_new_n20762__,
    new_new_n20763__, new_new_n20764__, new_new_n20765__, new_new_n20766__,
    new_new_n20767__, new_new_n20768__, new_new_n20769__, new_new_n20770__,
    new_new_n20771__, new_new_n20772__, new_new_n20773__, new_new_n20774__,
    new_new_n20775__, new_new_n20776__, new_new_n20777__, new_new_n20778__,
    new_new_n20779__, new_new_n20780__, new_new_n20781__, new_new_n20782__,
    new_new_n20783__, new_new_n20784__, new_new_n20785__, new_new_n20786__,
    new_new_n20787__, new_new_n20788__, new_new_n20789__, new_new_n20790__,
    new_new_n20791__, new_new_n20792__, new_new_n20793__, new_new_n20794__,
    new_new_n20795__, new_new_n20796__, new_new_n20797__, new_new_n20798__,
    new_new_n20799__, new_new_n20800__, new_new_n20801__, new_new_n20802__,
    new_new_n20803__, new_new_n20804__, new_new_n20805__, new_new_n20806__,
    new_new_n20807__, new_new_n20808__, new_new_n20809__, new_new_n20810__,
    new_new_n20811__, new_new_n20812__, new_new_n20813__, new_new_n20814__,
    new_new_n20815__, new_new_n20816__, new_new_n20817__, new_new_n20818__,
    new_new_n20819__, new_new_n20820__, new_new_n20821__, new_new_n20822__,
    new_new_n20823__, new_new_n20824__, new_new_n20825__, new_new_n20826__,
    new_new_n20827__, new_new_n20828__, new_new_n20829__, new_new_n20830__,
    new_new_n20831__, new_new_n20832__, new_new_n20833__, new_new_n20834__,
    new_new_n20835__, new_new_n20836__, new_new_n20837__, new_new_n20838__,
    new_new_n20839__, new_new_n20840__, new_new_n20841__, new_new_n20842__,
    new_new_n20843__, new_new_n20844__, new_new_n20845__, new_new_n20846__,
    new_new_n20847__, new_new_n20848__, new_new_n20849__, new_new_n20850__,
    new_new_n20851__, new_new_n20852__, new_new_n20853__, new_new_n20854__,
    new_new_n20855__, new_new_n20856__, new_new_n20857__, new_new_n20858__,
    new_new_n20859__, new_new_n20860__, new_new_n20861__, new_new_n20862__,
    new_new_n20863__, new_new_n20864__, new_new_n20865__, new_new_n20866__,
    new_new_n20867__, new_new_n20868__, new_new_n20869__, new_new_n20870__,
    new_new_n20871__, new_new_n20872__, new_new_n20873__, new_new_n20874__,
    new_new_n20875__, new_new_n20876__, new_new_n20877__, new_new_n20878__,
    new_new_n20879__, new_new_n20880__, new_new_n20881__, new_new_n20882__,
    new_new_n20883__, new_new_n20884__, new_new_n20885__, new_new_n20886__,
    new_new_n20887__, new_new_n20888__, new_new_n20889__, new_new_n20890__,
    new_new_n20891__, new_new_n20892__, new_new_n20893__, new_new_n20894__,
    new_new_n20895__, new_new_n20896__, new_new_n20897__, new_new_n20898__,
    new_new_n20899__, new_new_n20900__, new_new_n20901__, new_new_n20902__,
    new_new_n20903__, new_new_n20904__, new_new_n20905__, new_new_n20906__,
    new_new_n20907__, new_new_n20908__, new_new_n20909__, new_new_n20910__,
    new_new_n20911__, new_new_n20912__, new_new_n20913__, new_new_n20914__,
    new_new_n20915__, new_new_n20916__, new_new_n20917__, new_new_n20918__,
    new_new_n20919__, new_new_n20920__, new_new_n20921__, new_new_n20922__,
    new_new_n20923__, new_new_n20924__, new_new_n20925__, new_new_n20926__,
    new_new_n20927__, new_new_n20928__, new_new_n20929__, new_new_n20930__,
    new_new_n20931__, new_new_n20932__, new_new_n20933__, new_new_n20934__,
    new_new_n20935__, new_new_n20936__, new_new_n20937__, new_new_n20938__,
    new_new_n20939__, new_new_n20940__, new_new_n20941__, new_new_n20942__,
    new_new_n20943__, new_new_n20944__, new_new_n20945__, new_new_n20946__,
    new_new_n20947__, new_new_n20948__, new_new_n20949__, new_new_n20950__,
    new_new_n20951__, new_new_n20952__, new_new_n20953__, new_new_n20954__,
    new_new_n20955__, new_new_n20956__, new_new_n20957__, new_new_n20958__,
    new_new_n20959__, new_new_n20960__, new_new_n20961__, new_new_n20962__,
    new_new_n20963__, new_new_n20964__, new_new_n20965__, new_new_n20966__,
    new_new_n20967__, new_new_n20968__, new_new_n20969__, new_new_n20970__,
    new_new_n20971__, new_new_n20972__, new_new_n20973__, new_new_n20974__,
    new_new_n20975__, new_new_n20976__, new_new_n20977__, new_new_n20978__,
    new_new_n20979__, new_new_n20980__, new_new_n20981__, new_new_n20982__,
    new_new_n20983__, new_new_n20984__, new_new_n20985__, new_new_n20986__,
    new_new_n20987__, new_new_n20988__, new_new_n20989__, new_new_n20990__,
    new_new_n20991__, new_new_n20992__, new_new_n20993__, new_new_n20994__,
    new_new_n20995__, new_new_n20996__, new_new_n20997__, new_new_n20998__,
    new_new_n20999__, new_new_n21000__, new_new_n21001__, new_new_n21002__,
    new_new_n21003__, new_new_n21004__, new_new_n21005__, new_new_n21006__,
    new_new_n21007__, new_new_n21008__, new_new_n21009__, new_new_n21010__,
    new_new_n21011__, new_new_n21012__, new_new_n21013__, new_new_n21014__,
    new_new_n21015__, new_new_n21016__, new_new_n21017__, new_new_n21018__,
    new_new_n21019__, new_new_n21020__, new_new_n21021__, new_new_n21022__,
    new_new_n21023__, new_new_n21024__, new_new_n21025__, new_new_n21026__,
    new_new_n21027__, new_new_n21028__, new_new_n21029__, new_new_n21030__,
    new_new_n21031__, new_new_n21032__, new_new_n21033__, new_new_n21034__,
    new_new_n21035__, new_new_n21036__, new_new_n21037__, new_new_n21038__,
    new_new_n21039__, new_new_n21040__, new_new_n21041__, new_new_n21042__,
    new_new_n21043__, new_new_n21044__, new_new_n21045__, new_new_n21046__,
    new_new_n21047__, new_new_n21048__, new_new_n21049__, new_new_n21050__,
    new_new_n21051__, new_new_n21052__, new_new_n21053__, new_new_n21054__,
    new_new_n21055__, new_new_n21056__, new_new_n21057__, new_new_n21058__,
    new_new_n21059__, new_new_n21060__, new_new_n21061__, new_new_n21062__,
    new_new_n21063__, new_new_n21064__, new_new_n21065__, new_new_n21066__,
    new_new_n21067__, new_new_n21068__, new_new_n21069__, new_new_n21070__,
    new_new_n21071__, new_new_n21072__, new_new_n21073__, new_new_n21074__,
    new_new_n21075__, new_new_n21076__, new_new_n21077__, new_new_n21078__,
    new_new_n21079__, new_new_n21080__, new_new_n21081__, new_new_n21082__,
    new_new_n21083__, new_new_n21084__, new_new_n21085__, new_new_n21086__,
    new_new_n21087__, new_new_n21088__, new_new_n21089__, new_new_n21090__,
    new_new_n21091__, new_new_n21092__, new_new_n21093__, new_new_n21094__,
    new_new_n21095__, new_new_n21096__, new_new_n21097__, new_new_n21098__,
    new_new_n21099__, new_new_n21100__, new_new_n21101__, new_new_n21102__,
    new_new_n21103__, new_new_n21104__, new_new_n21105__, new_new_n21106__,
    new_new_n21107__, new_new_n21108__, new_new_n21109__, new_new_n21110__,
    new_new_n21111__, new_new_n21112__, new_new_n21113__, new_new_n21114__,
    new_new_n21115__, new_new_n21116__, new_new_n21117__, new_new_n21118__,
    new_new_n21119__, new_new_n21120__, new_new_n21121__, new_new_n21122__,
    new_new_n21123__, new_new_n21124__, new_new_n21125__, new_new_n21126__,
    new_new_n21127__, new_new_n21128__, new_new_n21129__, new_new_n21130__,
    new_new_n21131__, new_new_n21132__, new_new_n21133__, new_new_n21134__,
    new_new_n21135__, new_new_n21136__, new_new_n21137__, new_new_n21138__,
    new_new_n21139__, new_new_n21140__, new_new_n21141__, new_new_n21142__,
    new_new_n21143__, new_new_n21144__, new_new_n21145__, new_new_n21146__,
    new_new_n21147__, new_new_n21148__, new_new_n21149__, new_new_n21150__,
    new_new_n21151__, new_new_n21152__, new_new_n21153__, new_new_n21154__,
    new_new_n21155__, new_new_n21156__, new_new_n21157__, new_new_n21158__,
    new_new_n21159__, new_new_n21160__, new_new_n21161__, new_new_n21162__,
    new_new_n21163__, new_new_n21164__, new_new_n21165__, new_new_n21166__,
    new_new_n21167__, new_new_n21168__, new_new_n21169__, new_new_n21170__,
    new_new_n21171__, new_new_n21172__, new_new_n21173__, new_new_n21174__,
    new_new_n21175__, new_new_n21176__, new_new_n21177__, new_new_n21178__,
    new_new_n21179__, new_new_n21180__, new_new_n21181__, new_new_n21182__,
    new_new_n21183__, new_new_n21184__, new_new_n21185__, new_new_n21186__,
    new_new_n21187__, new_new_n21188__, new_new_n21189__, new_new_n21190__,
    new_new_n21191__, new_new_n21192__, new_new_n21193__, new_new_n21194__,
    new_new_n21195__, new_new_n21196__, new_new_n21197__, new_new_n21198__,
    new_new_n21199__, new_new_n21200__, new_new_n21201__, new_new_n21202__,
    new_new_n21203__, new_new_n21204__, new_new_n21205__, new_new_n21206__,
    new_new_n21207__, new_new_n21208__, new_new_n21209__, new_new_n21210__,
    new_new_n21211__, new_new_n21212__, new_new_n21213__, new_new_n21214__,
    new_new_n21215__, new_new_n21216__, new_new_n21217__, new_new_n21218__,
    new_new_n21219__, new_new_n21220__, new_new_n21221__, new_new_n21222__,
    new_new_n21223__, new_new_n21224__, new_new_n21225__, new_new_n21226__,
    new_new_n21227__, new_new_n21228__, new_new_n21229__, new_new_n21230__,
    new_new_n21231__, new_new_n21232__, new_new_n21233__, new_new_n21234__,
    new_new_n21235__, new_new_n21236__, new_new_n21237__, new_new_n21238__,
    new_new_n21239__, new_new_n21240__, new_new_n21241__, new_new_n21242__,
    new_new_n21243__, new_new_n21244__, new_new_n21245__, new_new_n21246__,
    new_new_n21247__, new_new_n21248__, new_new_n21249__, new_new_n21250__,
    new_new_n21251__, new_new_n21252__, new_new_n21253__, new_new_n21254__,
    new_new_n21255__, new_new_n21256__, new_new_n21257__, new_new_n21258__,
    new_new_n21259__, new_new_n21260__, new_new_n21261__, new_new_n21262__,
    new_new_n21263__, new_new_n21264__, new_new_n21265__, new_new_n21266__,
    new_new_n21267__, new_new_n21268__, new_new_n21269__, new_new_n21270__,
    new_new_n21271__, new_new_n21272__, new_new_n21273__, new_new_n21274__,
    new_new_n21275__, new_new_n21276__, new_new_n21277__, new_new_n21278__,
    new_new_n21279__, new_new_n21280__, new_new_n21281__, new_new_n21282__,
    new_new_n21283__, new_new_n21284__, new_new_n21285__, new_new_n21286__,
    new_new_n21287__, new_new_n21288__, new_new_n21289__, new_new_n21290__,
    new_new_n21291__, new_new_n21292__, new_new_n21293__, new_new_n21294__,
    new_new_n21295__, new_new_n21296__, new_new_n21297__, new_new_n21298__,
    new_new_n21299__, new_new_n21300__, new_new_n21301__, new_new_n21302__,
    new_new_n21303__, new_new_n21304__, new_new_n21305__, new_new_n21306__,
    new_new_n21307__, new_new_n21308__, new_new_n21309__, new_new_n21310__,
    new_new_n21311__, new_new_n21312__, new_new_n21313__, new_new_n21314__,
    new_new_n21315__, new_new_n21316__, new_new_n21317__, new_new_n21318__,
    new_new_n21319__, new_new_n21320__, new_new_n21321__, new_new_n21322__,
    new_new_n21323__, new_new_n21324__, new_new_n21325__, new_new_n21326__,
    new_new_n21327__, new_new_n21328__, new_new_n21329__, new_new_n21330__,
    new_new_n21331__, new_new_n21332__, new_new_n21333__, new_new_n21334__,
    new_new_n21335__, new_new_n21336__, new_new_n21337__, new_new_n21338__,
    new_new_n21339__, new_new_n21340__, new_new_n21341__, new_new_n21342__,
    new_new_n21344__, new_new_n21345__, new_new_n21346__, new_new_n21347__,
    new_new_n21348__, new_new_n21349__, new_new_n21350__, new_new_n21351__,
    new_new_n21352__, new_new_n21353__, new_new_n21354__, new_new_n21355__,
    new_new_n21356__, new_new_n21357__, new_new_n21358__, new_new_n21359__,
    new_new_n21360__, new_new_n21361__, new_new_n21362__, new_new_n21363__,
    new_new_n21364__, new_new_n21365__, new_new_n21366__, new_new_n21367__,
    new_new_n21368__, new_new_n21369__, new_new_n21370__, new_new_n21371__,
    new_new_n21372__, new_new_n21373__, new_new_n21374__, new_new_n21375__,
    new_new_n21376__, new_new_n21377__, new_new_n21378__, new_new_n21379__,
    new_new_n21380__, new_new_n21381__, new_new_n21382__, new_new_n21383__,
    new_new_n21384__, new_new_n21385__, new_new_n21386__, new_new_n21387__,
    new_new_n21388__, new_new_n21389__, new_new_n21390__, new_new_n21391__,
    new_new_n21392__, new_new_n21393__, new_new_n21394__, new_new_n21395__,
    new_new_n21396__, new_new_n21397__, new_new_n21398__, new_new_n21399__,
    new_new_n21400__, new_new_n21401__, new_new_n21402__, new_new_n21403__,
    new_new_n21404__, new_new_n21405__, new_new_n21406__, new_new_n21407__,
    new_new_n21408__, new_new_n21409__, new_new_n21410__, new_new_n21411__,
    new_new_n21412__, new_new_n21413__, new_new_n21414__, new_new_n21415__,
    new_new_n21416__, new_new_n21417__, new_new_n21418__, new_new_n21419__,
    new_new_n21420__, new_new_n21421__, new_new_n21422__, new_new_n21423__,
    new_new_n21424__, new_new_n21425__, new_new_n21426__, new_new_n21427__,
    new_new_n21428__, new_new_n21429__, new_new_n21430__, new_new_n21431__,
    new_new_n21432__, new_new_n21433__, new_new_n21434__, new_new_n21435__,
    new_new_n21436__, new_new_n21437__, new_new_n21438__, new_new_n21439__,
    new_new_n21440__, new_new_n21441__, new_new_n21442__, new_new_n21443__,
    new_new_n21444__, new_new_n21445__, new_new_n21446__, new_new_n21447__,
    new_new_n21448__, new_new_n21449__, new_new_n21450__, new_new_n21451__,
    new_new_n21452__, new_new_n21453__, new_new_n21454__, new_new_n21455__,
    new_new_n21456__, new_new_n21457__, new_new_n21458__, new_new_n21459__,
    new_new_n21460__, new_new_n21461__, new_new_n21462__, new_new_n21463__,
    new_new_n21464__, new_new_n21465__, new_new_n21466__, new_new_n21467__,
    new_new_n21468__, new_new_n21469__, new_new_n21470__, new_new_n21471__,
    new_new_n21472__, new_new_n21473__, new_new_n21474__, new_new_n21475__,
    new_new_n21476__, new_new_n21477__, new_new_n21478__, new_new_n21479__,
    new_new_n21480__, new_new_n21481__, new_new_n21482__, new_new_n21483__,
    new_new_n21484__, new_new_n21485__, new_new_n21486__, new_new_n21487__,
    new_new_n21488__, new_new_n21489__, new_new_n21490__, new_new_n21491__,
    new_new_n21492__, new_new_n21493__, new_new_n21494__, new_new_n21495__,
    new_new_n21496__, new_new_n21497__, new_new_n21498__, new_new_n21499__,
    new_new_n21500__, new_new_n21501__, new_new_n21502__, new_new_n21503__,
    new_new_n21504__, new_new_n21505__, new_new_n21506__, new_new_n21507__,
    new_new_n21508__, new_new_n21509__, new_new_n21510__, new_new_n21511__,
    new_new_n21512__, new_new_n21513__, new_new_n21514__, new_new_n21515__,
    new_new_n21516__, new_new_n21517__, new_new_n21518__, new_new_n21519__,
    new_new_n21520__, new_new_n21521__, new_new_n21522__, new_new_n21523__,
    new_new_n21524__, new_new_n21525__, new_new_n21526__, new_new_n21527__,
    new_new_n21528__, new_new_n21529__, new_new_n21530__, new_new_n21531__,
    new_new_n21532__, new_new_n21533__, new_new_n21534__, new_new_n21535__,
    new_new_n21536__, new_new_n21537__, new_new_n21538__, new_new_n21539__,
    new_new_n21540__, new_new_n21541__, new_new_n21542__, new_new_n21543__,
    new_new_n21544__, new_new_n21545__, new_new_n21546__, new_new_n21547__,
    new_new_n21548__, new_new_n21549__, new_new_n21550__, new_new_n21551__,
    new_new_n21552__, new_new_n21553__, new_new_n21554__, new_new_n21555__,
    new_new_n21556__, new_new_n21557__, new_new_n21558__, new_new_n21559__,
    new_new_n21560__, new_new_n21561__, new_new_n21562__, new_new_n21563__,
    new_new_n21564__, new_new_n21565__, new_new_n21566__, new_new_n21567__,
    new_new_n21568__, new_new_n21569__, new_new_n21570__, new_new_n21571__,
    new_new_n21572__, new_new_n21573__, new_new_n21574__, new_new_n21575__,
    new_new_n21576__, new_new_n21577__, new_new_n21578__, new_new_n21579__,
    new_new_n21580__, new_new_n21581__, new_new_n21582__, new_new_n21583__,
    new_new_n21584__, new_new_n21585__, new_new_n21586__, new_new_n21587__,
    new_new_n21588__, new_new_n21589__, new_new_n21590__, new_new_n21591__,
    new_new_n21592__, new_new_n21593__, new_new_n21594__, new_new_n21595__,
    new_new_n21596__, new_new_n21597__, new_new_n21598__, new_new_n21599__,
    new_new_n21600__, new_new_n21601__, new_new_n21602__, new_new_n21603__,
    new_new_n21604__, new_new_n21605__, new_new_n21606__, new_new_n21607__,
    new_new_n21608__, new_new_n21609__, new_new_n21610__, new_new_n21611__,
    new_new_n21612__, new_new_n21613__, new_new_n21614__, new_new_n21615__,
    new_new_n21616__, new_new_n21617__, new_new_n21618__, new_new_n21619__,
    new_new_n21620__, new_new_n21621__, new_new_n21622__, new_new_n21623__,
    new_new_n21624__, new_new_n21625__, new_new_n21626__, new_new_n21627__,
    new_new_n21628__, new_new_n21629__, new_new_n21630__, new_new_n21631__,
    new_new_n21632__, new_new_n21633__, new_new_n21634__, new_new_n21635__,
    new_new_n21636__, new_new_n21637__, new_new_n21638__, new_new_n21639__,
    new_new_n21640__, new_new_n21641__, new_new_n21642__, new_new_n21643__,
    new_new_n21644__, new_new_n21645__, new_new_n21646__, new_new_n21647__,
    new_new_n21648__, new_new_n21649__, new_new_n21650__, new_new_n21651__,
    new_new_n21652__, new_new_n21653__, new_new_n21654__, new_new_n21655__,
    new_new_n21656__, new_new_n21657__, new_new_n21658__, new_new_n21659__,
    new_new_n21660__, new_new_n21661__, new_new_n21662__, new_new_n21663__,
    new_new_n21664__, new_new_n21665__, new_new_n21666__, new_new_n21667__,
    new_new_n21668__, new_new_n21669__, new_new_n21670__, new_new_n21671__,
    new_new_n21672__, new_new_n21673__, new_new_n21674__, new_new_n21675__,
    new_new_n21676__, new_new_n21677__, new_new_n21678__, new_new_n21679__,
    new_new_n21680__, new_new_n21681__, new_new_n21682__, new_new_n21683__,
    new_new_n21684__, new_new_n21685__, new_new_n21686__, new_new_n21687__,
    new_new_n21688__, new_new_n21689__, new_new_n21690__, new_new_n21691__,
    new_new_n21692__, new_new_n21693__, new_new_n21694__, new_new_n21695__,
    new_new_n21696__, new_new_n21697__, new_new_n21698__, new_new_n21699__,
    new_new_n21700__, new_new_n21701__, new_new_n21702__, new_new_n21703__,
    new_new_n21704__, new_new_n21705__, new_new_n21706__, new_new_n21707__,
    new_new_n21708__, new_new_n21709__, new_new_n21710__, new_new_n21711__,
    new_new_n21712__, new_new_n21713__, new_new_n21714__, new_new_n21715__,
    new_new_n21716__, new_new_n21717__, new_new_n21718__, new_new_n21719__,
    new_new_n21720__, new_new_n21721__, new_new_n21722__, new_new_n21723__,
    new_new_n21724__, new_new_n21725__, new_new_n21726__, new_new_n21727__,
    new_new_n21728__, new_new_n21729__, new_new_n21730__, new_new_n21731__,
    new_new_n21732__, new_new_n21733__, new_new_n21734__, new_new_n21735__,
    new_new_n21736__, new_new_n21737__, new_new_n21738__, new_new_n21739__,
    new_new_n21740__, new_new_n21741__, new_new_n21742__, new_new_n21743__,
    new_new_n21744__, new_new_n21745__, new_new_n21746__, new_new_n21747__,
    new_new_n21748__, new_new_n21749__, new_new_n21750__, new_new_n21751__,
    new_new_n21752__, new_new_n21753__, new_new_n21754__, new_new_n21755__,
    new_new_n21756__, new_new_n21757__, new_new_n21758__, new_new_n21759__,
    new_new_n21760__, new_new_n21761__, new_new_n21762__, new_new_n21763__,
    new_new_n21764__, new_new_n21765__, new_new_n21766__, new_new_n21767__,
    new_new_n21768__, new_new_n21769__, new_new_n21770__, new_new_n21771__,
    new_new_n21772__, new_new_n21773__, new_new_n21774__, new_new_n21775__,
    new_new_n21776__, new_new_n21777__, new_new_n21778__, new_new_n21779__,
    new_new_n21780__, new_new_n21781__, new_new_n21782__, new_new_n21783__,
    new_new_n21784__, new_new_n21785__, new_new_n21786__, new_new_n21787__,
    new_new_n21788__, new_new_n21789__, new_new_n21790__, new_new_n21791__,
    new_new_n21792__, new_new_n21793__, new_new_n21794__, new_new_n21795__,
    new_new_n21796__, new_new_n21797__, new_new_n21798__, new_new_n21799__,
    new_new_n21800__, new_new_n21801__, new_new_n21802__, new_new_n21803__,
    new_new_n21804__, new_new_n21805__, new_new_n21806__, new_new_n21807__,
    new_new_n21808__, new_new_n21809__, new_new_n21810__, new_new_n21811__,
    new_new_n21812__, new_new_n21813__, new_new_n21814__, new_new_n21815__,
    new_new_n21816__, new_new_n21817__, new_new_n21818__, new_new_n21819__,
    new_new_n21820__, new_new_n21821__, new_new_n21822__, new_new_n21823__,
    new_new_n21824__, new_new_n21825__, new_new_n21826__, new_new_n21827__,
    new_new_n21828__, new_new_n21829__, new_new_n21830__, new_new_n21831__,
    new_new_n21832__, new_new_n21833__, new_new_n21834__, new_new_n21835__,
    new_new_n21836__, new_new_n21837__, new_new_n21838__, new_new_n21839__,
    new_new_n21840__, new_new_n21841__, new_new_n21842__, new_new_n21843__,
    new_new_n21844__, new_new_n21845__, new_new_n21846__, new_new_n21847__,
    new_new_n21848__, new_new_n21849__, new_new_n21850__, new_new_n21851__,
    new_new_n21852__, new_new_n21853__, new_new_n21854__, new_new_n21855__,
    new_new_n21856__, new_new_n21857__, new_new_n21858__, new_new_n21859__,
    new_new_n21860__, new_new_n21861__, new_new_n21862__, new_new_n21863__,
    new_new_n21864__, new_new_n21865__, new_new_n21866__, new_new_n21867__,
    new_new_n21868__, new_new_n21869__, new_new_n21870__, new_new_n21871__,
    new_new_n21872__, new_new_n21873__, new_new_n21874__, new_new_n21875__,
    new_new_n21876__, new_new_n21877__, new_new_n21878__, new_new_n21879__,
    new_new_n21880__, new_new_n21881__, new_new_n21882__, new_new_n21883__,
    new_new_n21884__, new_new_n21885__, new_new_n21886__, new_new_n21887__,
    new_new_n21888__, new_new_n21889__, new_new_n21890__, new_new_n21891__,
    new_new_n21892__, new_new_n21893__, new_new_n21894__, new_new_n21895__,
    new_new_n21896__, new_new_n21897__, new_new_n21898__, new_new_n21899__,
    new_new_n21900__, new_new_n21901__, new_new_n21902__, new_new_n21903__,
    new_new_n21904__, new_new_n21905__, new_new_n21906__, new_new_n21907__,
    new_new_n21908__, new_new_n21909__, new_new_n21910__, new_new_n21911__,
    new_new_n21912__, new_new_n21913__, new_new_n21914__, new_new_n21915__,
    new_new_n21916__, new_new_n21917__, new_new_n21918__, new_new_n21919__,
    new_new_n21920__, new_new_n21921__, new_new_n21922__, new_new_n21923__,
    new_new_n21924__, new_new_n21925__, new_new_n21926__, new_new_n21927__,
    new_new_n21928__, new_new_n21929__, new_new_n21930__, new_new_n21931__,
    new_new_n21932__, new_new_n21933__, new_new_n21934__, new_new_n21935__,
    new_new_n21936__, new_new_n21937__, new_new_n21938__, new_new_n21939__,
    new_new_n21940__, new_new_n21941__, new_new_n21942__, new_new_n21943__,
    new_new_n21944__, new_new_n21945__, new_new_n21946__, new_new_n21947__,
    new_new_n21948__, new_new_n21949__, new_new_n21950__, new_new_n21951__,
    new_new_n21952__, new_new_n21953__, new_new_n21954__, new_new_n21955__,
    new_new_n21956__, new_new_n21957__, new_new_n21958__, new_new_n21959__,
    new_new_n21960__, new_new_n21961__, new_new_n21962__, new_new_n21963__,
    new_new_n21964__, new_new_n21965__, new_new_n21966__, new_new_n21967__,
    new_new_n21968__, new_new_n21969__, new_new_n21970__, new_new_n21971__,
    new_new_n21972__, new_new_n21973__, new_new_n21974__, new_new_n21975__,
    new_new_n21976__, new_new_n21977__, new_new_n21978__, new_new_n21979__,
    new_new_n21980__, new_new_n21981__, new_new_n21982__, new_new_n21983__,
    new_new_n21984__, new_new_n21985__, new_new_n21986__, new_new_n21987__,
    new_new_n21988__, new_new_n21989__, new_new_n21990__, new_new_n21991__,
    new_new_n21992__, new_new_n21993__, new_new_n21994__, new_new_n21995__,
    new_new_n21996__, new_new_n21997__, new_new_n21998__, new_new_n21999__,
    new_new_n22000__, new_new_n22001__, new_new_n22002__, new_new_n22003__,
    new_new_n22004__, new_new_n22005__, new_new_n22006__, new_new_n22007__,
    new_new_n22008__, new_new_n22009__, new_new_n22010__, new_new_n22011__,
    new_new_n22012__, new_new_n22013__, new_new_n22014__, new_new_n22015__,
    new_new_n22016__, new_new_n22017__, new_new_n22018__, new_new_n22019__,
    new_new_n22020__, new_new_n22021__, new_new_n22022__, new_new_n22023__,
    new_new_n22024__, new_new_n22025__, new_new_n22026__, new_new_n22027__,
    new_new_n22028__, new_new_n22029__, new_new_n22030__, new_new_n22031__,
    new_new_n22032__, new_new_n22033__, new_new_n22034__, new_new_n22035__,
    new_new_n22037__, new_new_n22038__, new_new_n22039__, new_new_n22040__,
    new_new_n22041__, new_new_n22042__, new_new_n22043__, new_new_n22044__,
    new_new_n22045__, new_new_n22046__, new_new_n22047__, new_new_n22048__,
    new_new_n22049__, new_new_n22050__, new_new_n22051__, new_new_n22052__,
    new_new_n22053__, new_new_n22054__, new_new_n22055__, new_new_n22056__,
    new_new_n22057__, new_new_n22058__, new_new_n22059__, new_new_n22060__,
    new_new_n22061__, new_new_n22062__, new_new_n22063__, new_new_n22064__,
    new_new_n22065__, new_new_n22066__, new_new_n22067__, new_new_n22068__,
    new_new_n22069__, new_new_n22070__, new_new_n22071__, new_new_n22072__,
    new_new_n22073__, new_new_n22074__, new_new_n22075__, new_new_n22076__,
    new_new_n22077__, new_new_n22078__, new_new_n22079__, new_new_n22080__,
    new_new_n22081__, new_new_n22082__, new_new_n22083__, new_new_n22084__,
    new_new_n22085__, new_new_n22086__, new_new_n22087__, new_new_n22088__,
    new_new_n22089__, new_new_n22090__, new_new_n22091__, new_new_n22092__,
    new_new_n22093__, new_new_n22094__, new_new_n22095__, new_new_n22096__,
    new_new_n22097__, new_new_n22098__, new_new_n22099__, new_new_n22100__,
    new_new_n22101__, new_new_n22102__, new_new_n22103__, new_new_n22104__,
    new_new_n22105__, new_new_n22106__, new_new_n22107__, new_new_n22108__,
    new_new_n22109__, new_new_n22110__, new_new_n22111__, new_new_n22112__,
    new_new_n22113__, new_new_n22114__, new_new_n22115__, new_new_n22116__,
    new_new_n22117__, new_new_n22118__, new_new_n22119__, new_new_n22120__,
    new_new_n22121__, new_new_n22122__, new_new_n22123__, new_new_n22124__,
    new_new_n22125__, new_new_n22126__, new_new_n22127__, new_new_n22128__,
    new_new_n22129__, new_new_n22130__, new_new_n22131__, new_new_n22132__,
    new_new_n22133__, new_new_n22134__, new_new_n22135__, new_new_n22136__,
    new_new_n22137__, new_new_n22138__, new_new_n22139__, new_new_n22140__,
    new_new_n22141__, new_new_n22142__, new_new_n22143__, new_new_n22144__,
    new_new_n22145__, new_new_n22146__, new_new_n22147__, new_new_n22148__,
    new_new_n22149__, new_new_n22150__, new_new_n22151__, new_new_n22152__,
    new_new_n22153__, new_new_n22154__, new_new_n22155__, new_new_n22156__,
    new_new_n22157__, new_new_n22158__, new_new_n22159__, new_new_n22160__,
    new_new_n22161__, new_new_n22162__, new_new_n22163__, new_new_n22164__,
    new_new_n22165__, new_new_n22166__, new_new_n22167__, new_new_n22168__,
    new_new_n22169__, new_new_n22170__, new_new_n22171__, new_new_n22172__,
    new_new_n22173__, new_new_n22174__, new_new_n22175__, new_new_n22176__,
    new_new_n22177__, new_new_n22178__, new_new_n22179__, new_new_n22180__,
    new_new_n22181__, new_new_n22182__, new_new_n22183__, new_new_n22184__,
    new_new_n22185__, new_new_n22186__, new_new_n22187__, new_new_n22188__,
    new_new_n22189__, new_new_n22190__, new_new_n22191__, new_new_n22192__,
    new_new_n22193__, new_new_n22194__, new_new_n22195__, new_new_n22196__,
    new_new_n22197__, new_new_n22198__, new_new_n22199__, new_new_n22200__,
    new_new_n22201__, new_new_n22202__, new_new_n22203__, new_new_n22204__,
    new_new_n22205__, new_new_n22206__, new_new_n22207__, new_new_n22208__,
    new_new_n22209__, new_new_n22210__, new_new_n22211__, new_new_n22212__,
    new_new_n22213__, new_new_n22214__, new_new_n22215__, new_new_n22216__,
    new_new_n22217__, new_new_n22218__, new_new_n22219__, new_new_n22220__,
    new_new_n22221__, new_new_n22222__, new_new_n22223__, new_new_n22224__,
    new_new_n22225__, new_new_n22226__, new_new_n22227__, new_new_n22228__,
    new_new_n22229__, new_new_n22230__, new_new_n22231__, new_new_n22232__,
    new_new_n22233__, new_new_n22234__, new_new_n22235__, new_new_n22236__,
    new_new_n22237__, new_new_n22238__, new_new_n22239__, new_new_n22240__,
    new_new_n22241__, new_new_n22242__, new_new_n22243__, new_new_n22244__,
    new_new_n22245__, new_new_n22246__, new_new_n22247__, new_new_n22248__,
    new_new_n22249__, new_new_n22250__, new_new_n22251__, new_new_n22252__,
    new_new_n22253__, new_new_n22254__, new_new_n22255__, new_new_n22256__,
    new_new_n22257__, new_new_n22258__, new_new_n22259__, new_new_n22260__,
    new_new_n22261__, new_new_n22262__, new_new_n22263__, new_new_n22264__,
    new_new_n22265__, new_new_n22266__, new_new_n22267__, new_new_n22268__,
    new_new_n22269__, new_new_n22270__, new_new_n22271__, new_new_n22272__,
    new_new_n22273__, new_new_n22274__, new_new_n22275__, new_new_n22276__,
    new_new_n22277__, new_new_n22278__, new_new_n22279__, new_new_n22280__,
    new_new_n22281__, new_new_n22282__, new_new_n22283__, new_new_n22284__,
    new_new_n22285__, new_new_n22286__, new_new_n22287__, new_new_n22288__,
    new_new_n22289__, new_new_n22290__, new_new_n22291__, new_new_n22292__,
    new_new_n22293__, new_new_n22294__, new_new_n22295__, new_new_n22296__,
    new_new_n22297__, new_new_n22298__, new_new_n22299__, new_new_n22300__,
    new_new_n22301__, new_new_n22302__, new_new_n22303__, new_new_n22304__,
    new_new_n22305__, new_new_n22306__, new_new_n22307__, new_new_n22308__,
    new_new_n22309__, new_new_n22310__, new_new_n22311__, new_new_n22312__,
    new_new_n22313__, new_new_n22314__, new_new_n22315__, new_new_n22316__,
    new_new_n22317__, new_new_n22318__, new_new_n22319__, new_new_n22320__,
    new_new_n22321__, new_new_n22322__, new_new_n22323__, new_new_n22324__,
    new_new_n22325__, new_new_n22326__, new_new_n22327__, new_new_n22328__,
    new_new_n22329__, new_new_n22330__, new_new_n22331__, new_new_n22332__,
    new_new_n22333__, new_new_n22334__, new_new_n22335__, new_new_n22336__,
    new_new_n22337__, new_new_n22338__, new_new_n22339__, new_new_n22340__,
    new_new_n22341__, new_new_n22342__, new_new_n22343__, new_new_n22344__,
    new_new_n22345__, new_new_n22346__, new_new_n22347__, new_new_n22348__,
    new_new_n22349__, new_new_n22350__, new_new_n22351__, new_new_n22352__,
    new_new_n22353__, new_new_n22354__, new_new_n22355__, new_new_n22356__,
    new_new_n22357__, new_new_n22358__, new_new_n22359__, new_new_n22360__,
    new_new_n22361__, new_new_n22362__, new_new_n22363__, new_new_n22364__,
    new_new_n22365__, new_new_n22366__, new_new_n22367__, new_new_n22368__,
    new_new_n22369__, new_new_n22370__, new_new_n22371__, new_new_n22372__,
    new_new_n22373__, new_new_n22374__, new_new_n22375__, new_new_n22376__,
    new_new_n22377__, new_new_n22378__, new_new_n22379__, new_new_n22380__,
    new_new_n22381__, new_new_n22382__, new_new_n22383__, new_new_n22384__,
    new_new_n22385__, new_new_n22386__, new_new_n22387__, new_new_n22388__,
    new_new_n22389__, new_new_n22390__, new_new_n22391__, new_new_n22392__,
    new_new_n22393__, new_new_n22394__, new_new_n22395__, new_new_n22396__,
    new_new_n22397__, new_new_n22398__, new_new_n22399__, new_new_n22400__,
    new_new_n22401__, new_new_n22402__, new_new_n22403__, new_new_n22404__,
    new_new_n22405__, new_new_n22406__, new_new_n22407__, new_new_n22408__,
    new_new_n22409__, new_new_n22410__, new_new_n22411__, new_new_n22412__,
    new_new_n22413__, new_new_n22414__, new_new_n22415__, new_new_n22416__,
    new_new_n22417__, new_new_n22418__, new_new_n22419__, new_new_n22420__,
    new_new_n22421__, new_new_n22422__, new_new_n22423__, new_new_n22424__,
    new_new_n22425__, new_new_n22426__, new_new_n22427__, new_new_n22428__,
    new_new_n22429__, new_new_n22430__, new_new_n22431__, new_new_n22432__,
    new_new_n22433__, new_new_n22434__, new_new_n22435__, new_new_n22436__,
    new_new_n22437__, new_new_n22438__, new_new_n22439__, new_new_n22440__,
    new_new_n22441__, new_new_n22442__, new_new_n22443__, new_new_n22444__,
    new_new_n22445__, new_new_n22446__, new_new_n22447__, new_new_n22448__,
    new_new_n22449__, new_new_n22450__, new_new_n22451__, new_new_n22452__,
    new_new_n22453__, new_new_n22454__, new_new_n22455__, new_new_n22456__,
    new_new_n22457__, new_new_n22458__, new_new_n22459__, new_new_n22460__,
    new_new_n22461__, new_new_n22462__, new_new_n22463__, new_new_n22464__,
    new_new_n22465__, new_new_n22466__, new_new_n22467__, new_new_n22468__,
    new_new_n22469__, new_new_n22470__, new_new_n22471__, new_new_n22472__,
    new_new_n22473__, new_new_n22474__, new_new_n22475__, new_new_n22476__,
    new_new_n22477__, new_new_n22478__, new_new_n22479__, new_new_n22480__,
    new_new_n22481__, new_new_n22482__, new_new_n22483__, new_new_n22484__,
    new_new_n22485__, new_new_n22486__, new_new_n22487__, new_new_n22488__,
    new_new_n22489__, new_new_n22490__, new_new_n22491__, new_new_n22492__,
    new_new_n22493__, new_new_n22494__, new_new_n22495__, new_new_n22496__,
    new_new_n22497__, new_new_n22498__, new_new_n22499__, new_new_n22500__,
    new_new_n22501__, new_new_n22502__, new_new_n22503__, new_new_n22504__,
    new_new_n22505__, new_new_n22506__, new_new_n22507__, new_new_n22508__,
    new_new_n22509__, new_new_n22510__, new_new_n22511__, new_new_n22512__,
    new_new_n22513__, new_new_n22514__, new_new_n22515__, new_new_n22516__,
    new_new_n22517__, new_new_n22518__, new_new_n22519__, new_new_n22520__,
    new_new_n22521__, new_new_n22522__, new_new_n22523__, new_new_n22524__,
    new_new_n22525__, new_new_n22526__, new_new_n22527__, new_new_n22528__,
    new_new_n22529__, new_new_n22530__, new_new_n22531__, new_new_n22532__,
    new_new_n22533__, new_new_n22534__, new_new_n22535__, new_new_n22536__,
    new_new_n22537__, new_new_n22538__, new_new_n22539__, new_new_n22540__,
    new_new_n22541__, new_new_n22542__, new_new_n22543__, new_new_n22544__,
    new_new_n22545__, new_new_n22546__, new_new_n22547__, new_new_n22548__,
    new_new_n22549__, new_new_n22550__, new_new_n22551__, new_new_n22552__,
    new_new_n22553__, new_new_n22554__, new_new_n22555__, new_new_n22556__,
    new_new_n22557__, new_new_n22558__, new_new_n22559__, new_new_n22560__,
    new_new_n22561__, new_new_n22562__, new_new_n22563__, new_new_n22564__,
    new_new_n22565__, new_new_n22566__, new_new_n22567__, new_new_n22568__,
    new_new_n22569__, new_new_n22570__, new_new_n22571__, new_new_n22572__,
    new_new_n22573__, new_new_n22574__, new_new_n22575__, new_new_n22576__,
    new_new_n22577__, new_new_n22578__, new_new_n22579__, new_new_n22580__,
    new_new_n22581__, new_new_n22582__, new_new_n22583__, new_new_n22584__,
    new_new_n22585__, new_new_n22586__, new_new_n22587__, new_new_n22588__,
    new_new_n22589__, new_new_n22590__, new_new_n22591__, new_new_n22592__,
    new_new_n22593__, new_new_n22594__, new_new_n22595__, new_new_n22596__,
    new_new_n22597__, new_new_n22598__, new_new_n22599__, new_new_n22600__,
    new_new_n22601__, new_new_n22602__, new_new_n22603__, new_new_n22604__,
    new_new_n22605__, new_new_n22606__, new_new_n22607__, new_new_n22608__,
    new_new_n22609__, new_new_n22610__, new_new_n22611__, new_new_n22612__,
    new_new_n22613__, new_new_n22614__, new_new_n22615__, new_new_n22616__,
    new_new_n22617__, new_new_n22618__, new_new_n22619__, new_new_n22620__,
    new_new_n22621__, new_new_n22622__, new_new_n22623__, new_new_n22624__,
    new_new_n22625__, new_new_n22626__, new_new_n22627__, new_new_n22628__,
    new_new_n22629__, new_new_n22630__, new_new_n22631__, new_new_n22632__,
    new_new_n22633__, new_new_n22634__, new_new_n22635__, new_new_n22636__,
    new_new_n22637__, new_new_n22638__, new_new_n22639__, new_new_n22640__,
    new_new_n22641__, new_new_n22642__, new_new_n22643__, new_new_n22644__,
    new_new_n22645__, new_new_n22646__, new_new_n22647__, new_new_n22648__,
    new_new_n22649__, new_new_n22650__, new_new_n22651__, new_new_n22652__,
    new_new_n22653__, new_new_n22654__, new_new_n22655__, new_new_n22656__,
    new_new_n22657__, new_new_n22658__, new_new_n22659__, new_new_n22660__,
    new_new_n22661__, new_new_n22662__, new_new_n22663__, new_new_n22664__,
    new_new_n22665__, new_new_n22666__, new_new_n22667__, new_new_n22668__,
    new_new_n22669__, new_new_n22670__, new_new_n22671__, new_new_n22672__,
    new_new_n22673__, new_new_n22674__, new_new_n22675__, new_new_n22676__,
    new_new_n22677__, new_new_n22678__, new_new_n22679__, new_new_n22680__,
    new_new_n22681__, new_new_n22682__, new_new_n22683__, new_new_n22684__,
    new_new_n22685__, new_new_n22686__, new_new_n22687__, new_new_n22688__,
    new_new_n22689__, new_new_n22690__, new_new_n22691__, new_new_n22692__,
    new_new_n22693__, new_new_n22694__, new_new_n22695__, new_new_n22696__,
    new_new_n22697__, new_new_n22698__, new_new_n22699__, new_new_n22700__,
    new_new_n22701__, new_new_n22702__, new_new_n22703__, new_new_n22704__,
    new_new_n22705__, new_new_n22706__, new_new_n22707__, new_new_n22708__,
    new_new_n22709__, new_new_n22710__, new_new_n22711__, new_new_n22712__,
    new_new_n22713__, new_new_n22714__, new_new_n22715__, new_new_n22716__,
    new_new_n22717__, new_new_n22718__, new_new_n22719__, new_new_n22720__,
    new_new_n22721__, new_new_n22722__, new_new_n22723__, new_new_n22724__,
    new_new_n22725__, new_new_n22726__, new_new_n22727__, new_new_n22728__,
    new_new_n22729__, new_new_n22730__, new_new_n22731__, new_new_n22732__,
    new_new_n22733__, new_new_n22734__, new_new_n22735__, new_new_n22736__,
    new_new_n22737__, new_new_n22738__, new_new_n22739__, new_new_n22740__,
    new_new_n22741__, new_new_n22742__, new_new_n22743__, new_new_n22744__,
    new_new_n22745__, new_new_n22746__, new_new_n22747__, new_new_n22748__,
    new_new_n22749__, new_new_n22750__, new_new_n22751__, new_new_n22752__,
    new_new_n22753__, new_new_n22754__, new_new_n22755__, new_new_n22756__,
    new_new_n22757__, new_new_n22758__, new_new_n22759__, new_new_n22760__,
    new_new_n22761__, new_new_n22762__, new_new_n22763__, new_new_n22764__,
    new_new_n22765__, new_new_n22766__, new_new_n22767__, new_new_n22768__,
    new_new_n22770__, new_new_n22771__, new_new_n22772__, new_new_n22773__,
    new_new_n22774__, new_new_n22775__, new_new_n22776__, new_new_n22777__,
    new_new_n22778__, new_new_n22779__, new_new_n22780__, new_new_n22781__,
    new_new_n22782__, new_new_n22783__, new_new_n22784__, new_new_n22785__,
    new_new_n22786__, new_new_n22787__, new_new_n22788__, new_new_n22789__,
    new_new_n22790__, new_new_n22791__, new_new_n22792__, new_new_n22793__,
    new_new_n22794__, new_new_n22795__, new_new_n22796__, new_new_n22797__,
    new_new_n22798__, new_new_n22799__, new_new_n22800__, new_new_n22801__,
    new_new_n22802__, new_new_n22803__, new_new_n22804__, new_new_n22805__,
    new_new_n22806__, new_new_n22807__, new_new_n22808__, new_new_n22809__,
    new_new_n22810__, new_new_n22811__, new_new_n22812__, new_new_n22813__,
    new_new_n22814__, new_new_n22815__, new_new_n22816__, new_new_n22817__,
    new_new_n22818__, new_new_n22819__, new_new_n22820__, new_new_n22821__,
    new_new_n22822__, new_new_n22823__, new_new_n22824__, new_new_n22825__,
    new_new_n22826__, new_new_n22827__, new_new_n22828__, new_new_n22829__,
    new_new_n22830__, new_new_n22831__, new_new_n22832__, new_new_n22833__,
    new_new_n22834__, new_new_n22835__, new_new_n22836__, new_new_n22837__,
    new_new_n22838__, new_new_n22839__, new_new_n22840__, new_new_n22841__,
    new_new_n22842__, new_new_n22843__, new_new_n22844__, new_new_n22845__,
    new_new_n22846__, new_new_n22847__, new_new_n22848__, new_new_n22849__,
    new_new_n22850__, new_new_n22851__, new_new_n22852__, new_new_n22853__,
    new_new_n22854__, new_new_n22855__, new_new_n22856__, new_new_n22857__,
    new_new_n22858__, new_new_n22859__, new_new_n22860__, new_new_n22861__,
    new_new_n22862__, new_new_n22863__, new_new_n22864__, new_new_n22865__,
    new_new_n22866__, new_new_n22867__, new_new_n22868__, new_new_n22869__,
    new_new_n22870__, new_new_n22871__, new_new_n22872__, new_new_n22873__,
    new_new_n22874__, new_new_n22875__, new_new_n22876__, new_new_n22877__,
    new_new_n22878__, new_new_n22879__, new_new_n22880__, new_new_n22881__,
    new_new_n22882__, new_new_n22883__, new_new_n22884__, new_new_n22885__,
    new_new_n22886__, new_new_n22887__, new_new_n22888__, new_new_n22889__,
    new_new_n22890__, new_new_n22891__, new_new_n22892__, new_new_n22893__,
    new_new_n22894__, new_new_n22895__, new_new_n22896__, new_new_n22897__,
    new_new_n22898__, new_new_n22899__, new_new_n22900__, new_new_n22901__,
    new_new_n22902__, new_new_n22903__, new_new_n22904__, new_new_n22905__,
    new_new_n22906__, new_new_n22907__, new_new_n22908__, new_new_n22909__,
    new_new_n22910__, new_new_n22911__, new_new_n22912__, new_new_n22913__,
    new_new_n22914__, new_new_n22915__, new_new_n22916__, new_new_n22917__,
    new_new_n22918__, new_new_n22919__, new_new_n22920__, new_new_n22921__,
    new_new_n22922__, new_new_n22923__, new_new_n22924__, new_new_n22925__,
    new_new_n22926__, new_new_n22927__, new_new_n22928__, new_new_n22929__,
    new_new_n22930__, new_new_n22931__, new_new_n22932__, new_new_n22933__,
    new_new_n22934__, new_new_n22935__, new_new_n22936__, new_new_n22937__,
    new_new_n22938__, new_new_n22939__, new_new_n22940__, new_new_n22941__,
    new_new_n22942__, new_new_n22943__, new_new_n22944__, new_new_n22945__,
    new_new_n22946__, new_new_n22947__, new_new_n22948__, new_new_n22949__,
    new_new_n22950__, new_new_n22951__, new_new_n22952__, new_new_n22953__,
    new_new_n22954__, new_new_n22955__, new_new_n22956__, new_new_n22957__,
    new_new_n22958__, new_new_n22959__, new_new_n22960__, new_new_n22961__,
    new_new_n22962__, new_new_n22963__, new_new_n22964__, new_new_n22965__,
    new_new_n22966__, new_new_n22967__, new_new_n22968__, new_new_n22969__,
    new_new_n22970__, new_new_n22971__, new_new_n22972__, new_new_n22973__,
    new_new_n22974__, new_new_n22975__, new_new_n22976__, new_new_n22977__,
    new_new_n22978__, new_new_n22979__, new_new_n22980__, new_new_n22981__,
    new_new_n22982__, new_new_n22983__, new_new_n22984__, new_new_n22985__,
    new_new_n22986__, new_new_n22987__, new_new_n22988__, new_new_n22989__,
    new_new_n22990__, new_new_n22991__, new_new_n22992__, new_new_n22993__,
    new_new_n22994__, new_new_n22995__, new_new_n22996__, new_new_n22997__,
    new_new_n22998__, new_new_n22999__, new_new_n23000__, new_new_n23001__,
    new_new_n23002__, new_new_n23003__, new_new_n23004__, new_new_n23005__,
    new_new_n23006__, new_new_n23007__, new_new_n23008__, new_new_n23009__,
    new_new_n23010__, new_new_n23011__, new_new_n23012__, new_new_n23013__,
    new_new_n23014__, new_new_n23015__, new_new_n23016__, new_new_n23017__,
    new_new_n23018__, new_new_n23019__, new_new_n23020__, new_new_n23021__,
    new_new_n23022__, new_new_n23023__, new_new_n23024__, new_new_n23025__,
    new_new_n23026__, new_new_n23027__, new_new_n23028__, new_new_n23029__,
    new_new_n23030__, new_new_n23031__, new_new_n23032__, new_new_n23033__,
    new_new_n23034__, new_new_n23035__, new_new_n23036__, new_new_n23037__,
    new_new_n23038__, new_new_n23039__, new_new_n23040__, new_new_n23041__,
    new_new_n23042__, new_new_n23043__, new_new_n23044__, new_new_n23045__,
    new_new_n23046__, new_new_n23047__, new_new_n23048__, new_new_n23049__,
    new_new_n23050__, new_new_n23051__, new_new_n23052__, new_new_n23053__,
    new_new_n23054__, new_new_n23055__, new_new_n23056__, new_new_n23057__,
    new_new_n23058__, new_new_n23059__, new_new_n23060__, new_new_n23061__,
    new_new_n23062__, new_new_n23063__, new_new_n23064__, new_new_n23065__,
    new_new_n23066__, new_new_n23067__, new_new_n23068__, new_new_n23069__,
    new_new_n23070__, new_new_n23071__, new_new_n23072__, new_new_n23073__,
    new_new_n23074__, new_new_n23075__, new_new_n23076__, new_new_n23077__,
    new_new_n23078__, new_new_n23079__, new_new_n23080__, new_new_n23081__,
    new_new_n23082__, new_new_n23083__, new_new_n23084__, new_new_n23085__,
    new_new_n23086__, new_new_n23087__, new_new_n23088__, new_new_n23089__,
    new_new_n23090__, new_new_n23091__, new_new_n23092__, new_new_n23093__,
    new_new_n23094__, new_new_n23095__, new_new_n23096__, new_new_n23097__,
    new_new_n23098__, new_new_n23099__, new_new_n23100__, new_new_n23101__,
    new_new_n23102__, new_new_n23103__, new_new_n23104__, new_new_n23105__,
    new_new_n23106__, new_new_n23107__, new_new_n23108__, new_new_n23109__,
    new_new_n23110__, new_new_n23111__, new_new_n23112__, new_new_n23113__,
    new_new_n23114__, new_new_n23115__, new_new_n23116__, new_new_n23117__,
    new_new_n23118__, new_new_n23119__, new_new_n23120__, new_new_n23121__,
    new_new_n23122__, new_new_n23123__, new_new_n23124__, new_new_n23125__,
    new_new_n23126__, new_new_n23127__, new_new_n23128__, new_new_n23129__,
    new_new_n23130__, new_new_n23131__, new_new_n23132__, new_new_n23133__,
    new_new_n23134__, new_new_n23135__, new_new_n23136__, new_new_n23137__,
    new_new_n23138__, new_new_n23139__, new_new_n23140__, new_new_n23141__,
    new_new_n23142__, new_new_n23143__, new_new_n23144__, new_new_n23145__,
    new_new_n23146__, new_new_n23147__, new_new_n23148__, new_new_n23149__,
    new_new_n23150__, new_new_n23151__, new_new_n23152__, new_new_n23153__,
    new_new_n23154__, new_new_n23155__, new_new_n23156__, new_new_n23157__,
    new_new_n23158__, new_new_n23159__, new_new_n23160__, new_new_n23161__,
    new_new_n23162__, new_new_n23163__, new_new_n23164__, new_new_n23165__,
    new_new_n23166__, new_new_n23167__, new_new_n23168__, new_new_n23169__,
    new_new_n23170__, new_new_n23171__, new_new_n23172__, new_new_n23173__,
    new_new_n23174__, new_new_n23175__, new_new_n23176__, new_new_n23177__,
    new_new_n23178__, new_new_n23179__, new_new_n23180__, new_new_n23181__,
    new_new_n23182__, new_new_n23183__, new_new_n23184__, new_new_n23185__,
    new_new_n23186__, new_new_n23187__, new_new_n23188__, new_new_n23189__,
    new_new_n23190__, new_new_n23191__, new_new_n23192__, new_new_n23193__,
    new_new_n23194__, new_new_n23195__, new_new_n23196__, new_new_n23197__,
    new_new_n23198__, new_new_n23199__, new_new_n23200__, new_new_n23201__,
    new_new_n23202__, new_new_n23203__, new_new_n23204__, new_new_n23205__,
    new_new_n23206__, new_new_n23207__, new_new_n23208__, new_new_n23209__,
    new_new_n23210__, new_new_n23211__, new_new_n23212__, new_new_n23213__,
    new_new_n23214__, new_new_n23215__, new_new_n23216__, new_new_n23217__,
    new_new_n23218__, new_new_n23219__, new_new_n23220__, new_new_n23221__,
    new_new_n23222__, new_new_n23223__, new_new_n23224__, new_new_n23225__,
    new_new_n23226__, new_new_n23227__, new_new_n23228__, new_new_n23229__,
    new_new_n23230__, new_new_n23231__, new_new_n23232__, new_new_n23233__,
    new_new_n23234__, new_new_n23235__, new_new_n23236__, new_new_n23237__,
    new_new_n23238__, new_new_n23239__, new_new_n23240__, new_new_n23241__,
    new_new_n23242__, new_new_n23243__, new_new_n23244__, new_new_n23245__,
    new_new_n23246__, new_new_n23247__, new_new_n23248__, new_new_n23249__,
    new_new_n23250__, new_new_n23251__, new_new_n23252__, new_new_n23253__,
    new_new_n23254__, new_new_n23255__, new_new_n23256__, new_new_n23257__,
    new_new_n23258__, new_new_n23259__, new_new_n23260__, new_new_n23261__,
    new_new_n23262__, new_new_n23263__, new_new_n23264__, new_new_n23265__,
    new_new_n23266__, new_new_n23267__, new_new_n23268__, new_new_n23269__,
    new_new_n23270__, new_new_n23271__, new_new_n23272__, new_new_n23273__,
    new_new_n23274__, new_new_n23275__, new_new_n23276__, new_new_n23277__,
    new_new_n23278__, new_new_n23279__, new_new_n23280__, new_new_n23281__,
    new_new_n23282__, new_new_n23283__, new_new_n23284__, new_new_n23285__,
    new_new_n23286__, new_new_n23287__, new_new_n23288__, new_new_n23289__,
    new_new_n23290__, new_new_n23291__, new_new_n23292__, new_new_n23293__,
    new_new_n23294__, new_new_n23295__, new_new_n23296__, new_new_n23297__,
    new_new_n23298__, new_new_n23299__, new_new_n23300__, new_new_n23301__,
    new_new_n23302__, new_new_n23303__, new_new_n23304__, new_new_n23305__,
    new_new_n23306__, new_new_n23307__, new_new_n23308__, new_new_n23309__,
    new_new_n23310__, new_new_n23311__, new_new_n23312__, new_new_n23313__,
    new_new_n23314__, new_new_n23315__, new_new_n23316__, new_new_n23317__,
    new_new_n23318__, new_new_n23319__, new_new_n23320__, new_new_n23321__,
    new_new_n23322__, new_new_n23323__, new_new_n23324__, new_new_n23325__,
    new_new_n23326__, new_new_n23327__, new_new_n23328__, new_new_n23329__,
    new_new_n23330__, new_new_n23331__, new_new_n23332__, new_new_n23333__,
    new_new_n23334__, new_new_n23335__, new_new_n23336__, new_new_n23337__,
    new_new_n23338__, new_new_n23339__, new_new_n23340__, new_new_n23341__,
    new_new_n23342__, new_new_n23343__, new_new_n23344__, new_new_n23345__,
    new_new_n23346__, new_new_n23347__, new_new_n23348__, new_new_n23349__,
    new_new_n23350__, new_new_n23351__, new_new_n23352__, new_new_n23353__,
    new_new_n23354__, new_new_n23355__, new_new_n23356__, new_new_n23357__,
    new_new_n23358__, new_new_n23359__, new_new_n23360__, new_new_n23361__,
    new_new_n23362__, new_new_n23363__, new_new_n23364__, new_new_n23365__,
    new_new_n23366__, new_new_n23367__, new_new_n23368__, new_new_n23369__,
    new_new_n23370__, new_new_n23371__, new_new_n23372__, new_new_n23373__,
    new_new_n23374__, new_new_n23375__, new_new_n23376__, new_new_n23377__,
    new_new_n23378__, new_new_n23379__, new_new_n23380__, new_new_n23381__,
    new_new_n23382__, new_new_n23383__, new_new_n23384__, new_new_n23385__,
    new_new_n23386__, new_new_n23387__, new_new_n23388__, new_new_n23389__,
    new_new_n23390__, new_new_n23391__, new_new_n23392__, new_new_n23393__,
    new_new_n23394__, new_new_n23395__, new_new_n23396__, new_new_n23397__,
    new_new_n23398__, new_new_n23399__, new_new_n23400__, new_new_n23401__,
    new_new_n23402__, new_new_n23403__, new_new_n23404__, new_new_n23405__,
    new_new_n23406__, new_new_n23407__, new_new_n23408__, new_new_n23409__,
    new_new_n23410__, new_new_n23411__, new_new_n23412__, new_new_n23413__,
    new_new_n23414__, new_new_n23415__, new_new_n23416__, new_new_n23417__,
    new_new_n23418__, new_new_n23419__, new_new_n23420__, new_new_n23421__,
    new_new_n23422__, new_new_n23423__, new_new_n23424__, new_new_n23425__,
    new_new_n23426__, new_new_n23427__, new_new_n23428__, new_new_n23429__,
    new_new_n23430__, new_new_n23431__, new_new_n23432__, new_new_n23433__,
    new_new_n23434__, new_new_n23435__, new_new_n23436__, new_new_n23437__,
    new_new_n23438__, new_new_n23439__, new_new_n23440__, new_new_n23441__,
    new_new_n23442__, new_new_n23443__, new_new_n23444__, new_new_n23445__,
    new_new_n23446__, new_new_n23447__, new_new_n23448__, new_new_n23449__,
    new_new_n23450__, new_new_n23451__, new_new_n23452__, new_new_n23453__,
    new_new_n23454__, new_new_n23455__, new_new_n23456__, new_new_n23457__,
    new_new_n23458__, new_new_n23459__, new_new_n23460__, new_new_n23461__,
    new_new_n23464__, new_new_n23465__, new_new_n23466__, new_new_n23468__,
    new_new_n23469__, new_new_n23470__, new_new_n23472__, new_new_n23473__,
    new_new_n23474__, new_new_n23475__, new_new_n23476__, new_new_n23477__,
    new_new_n23478__, new_new_n23479__, new_new_n23480__, new_new_n23481__,
    new_new_n23482__, new_new_n23483__, new_new_n23484__, new_new_n23485__,
    new_new_n23486__, new_new_n23487__, new_new_n23488__, new_new_n23489__,
    new_new_n23490__, new_new_n23491__, new_new_n23492__, new_new_n23493__,
    new_new_n23494__, new_new_n23495__, new_new_n23497__, new_new_n23498__,
    new_new_n23499__, new_new_n23500__, new_new_n23502__, new_new_n23503__,
    new_new_n23504__, new_new_n23505__, new_new_n23506__, new_new_n23507__,
    new_new_n23509__, new_new_n23510__, new_new_n23511__, new_new_n23512__,
    new_new_n23514__, new_new_n23515__, new_new_n23516__, new_new_n23517__,
    new_new_n23518__, new_new_n23519__, new_new_n23521__, new_new_n23522__,
    new_new_n23523__, new_new_n23524__, new_new_n23525__, new_new_n23526__,
    new_new_n23528__, new_new_n23529__, new_new_n23530__, new_new_n23531__,
    new_new_n23532__, new_new_n23533__, new_new_n23535__, new_new_n23536__,
    new_new_n23537__, new_new_n23538__, new_new_n23539__, new_new_n23540__,
    new_new_n23542__, new_new_n23543__, new_new_n23544__, new_new_n23545__,
    new_new_n23546__, new_new_n23547__, new_new_n23549__, new_new_n23550__,
    new_new_n23551__, new_new_n23552__, new_new_n23553__, new_new_n23554__,
    new_new_n23556__, new_new_n23557__, new_new_n23558__, new_new_n23559__,
    new_new_n23560__, new_new_n23561__, new_new_n23563__, new_new_n23564__,
    new_new_n23565__, new_new_n23566__, new_new_n23567__, new_new_n23568__,
    new_new_n23570__, new_new_n23571__, new_new_n23572__, new_new_n23573__,
    new_new_n23574__, new_new_n23575__, new_new_n23577__, new_new_n23578__,
    new_new_n23579__, new_new_n23580__, new_new_n23581__, new_new_n23582__,
    new_new_n23584__, new_new_n23585__, new_new_n23586__, new_new_n23587__,
    new_new_n23588__, new_new_n23589__, new_new_n23591__, new_new_n23592__,
    new_new_n23593__, new_new_n23594__, new_new_n23595__, new_new_n23596__,
    new_new_n23598__, new_new_n23599__, new_new_n23600__, new_new_n23601__,
    new_new_n23602__, new_new_n23603__, new_new_n23605__, new_new_n23606__,
    new_new_n23607__, new_new_n23608__, new_new_n23609__, new_new_n23610__,
    new_new_n23612__, new_new_n23613__, new_new_n23614__, new_new_n23615__,
    new_new_n23616__, new_new_n23617__, new_new_n23619__, new_new_n23620__,
    new_new_n23621__, new_new_n23622__, new_new_n23623__, new_new_n23624__,
    new_new_n23626__, new_new_n23627__, new_new_n23628__, new_new_n23629__,
    new_new_n23630__, new_new_n23631__, new_new_n23633__, new_new_n23634__,
    new_new_n23635__, new_new_n23636__, new_new_n23637__, new_new_n23638__,
    new_new_n23640__, new_new_n23641__, new_new_n23642__, new_new_n23643__,
    new_new_n23644__, new_new_n23645__, new_new_n23647__, new_new_n23648__,
    new_new_n23649__, new_new_n23650__, new_new_n23651__, new_new_n23652__,
    new_new_n23654__, new_new_n23655__, new_new_n23656__, new_new_n23657__,
    new_new_n23658__, new_new_n23659__, new_new_n23661__, new_new_n23662__,
    new_new_n23663__, new_new_n23664__, new_new_n23665__, new_new_n23666__,
    new_new_n23668__, new_new_n23669__, new_new_n23670__, new_new_n23671__,
    new_new_n23672__, new_new_n23673__, new_new_n23675__, new_new_n23676__,
    new_new_n23677__, new_new_n23678__, new_new_n23679__, new_new_n23680__,
    new_new_n23682__, new_new_n23683__, new_new_n23684__, new_new_n23685__,
    new_new_n23686__, new_new_n23687__, new_new_n23689__, new_new_n23690__,
    new_new_n23691__, new_new_n23692__, new_new_n23693__, new_new_n23694__,
    new_new_n23696__, new_new_n23697__, new_new_n23698__, new_new_n23699__,
    new_new_n23700__, new_new_n23701__, new_new_n23703__, new_new_n23704__,
    new_new_n23705__, new_new_n23706__, new_new_n23707__, new_new_n23708__,
    new_new_n23710__, new_new_n23711__, new_new_n23712__, new_new_n23713__,
    new_new_n23714__, new_new_n23715__, new_new_n23717__, new_new_n23718__,
    new_new_n23719__, new_new_n23720__, new_new_n23721__, new_new_n23722__,
    new_new_n23724__, new_new_n23725__, new_new_n23726__, new_new_n23727__,
    new_new_n23728__, new_new_n23729__, new_new_n23731__, new_new_n23732__,
    new_new_n23733__, new_new_n23734__, new_new_n23735__, new_new_n23736__,
    new_new_n23738__, new_new_n23739__, new_new_n23740__, new_new_n23741__,
    new_new_n23742__, new_new_n23743__, new_new_n23745__, new_new_n23746__,
    new_new_n23747__, new_new_n23748__, new_new_n23749__, new_new_n23750__,
    new_new_n23752__, new_new_n23753__, new_new_n23754__, new_new_n23755__,
    new_new_n23756__, new_new_n23757__, new_new_n23759__, new_new_n23760__,
    new_new_n23761__, new_new_n23762__, new_new_n23763__, new_new_n23764__,
    new_new_n23766__, new_new_n23767__, new_new_n23768__, new_new_n23769__,
    new_new_n23770__, new_new_n23771__, new_new_n23773__, new_new_n23774__,
    new_new_n23775__, new_new_n23776__, new_new_n23777__, new_new_n23778__,
    new_new_n23780__, new_new_n23781__, new_new_n23782__, new_new_n23783__,
    new_new_n23784__, new_new_n23785__, new_new_n23787__, new_new_n23788__,
    new_new_n23789__, new_new_n23790__, new_new_n23791__, new_new_n23792__,
    new_new_n23794__, new_new_n23795__, new_new_n23796__, new_new_n23797__,
    new_new_n23798__, new_new_n23799__, new_new_n23801__, new_new_n23802__,
    new_new_n23803__, new_new_n23804__, new_new_n23805__, new_new_n23806__,
    new_new_n23808__, new_new_n23809__, new_new_n23810__, new_new_n23811__,
    new_new_n23812__, new_new_n23813__, new_new_n23815__, new_new_n23816__,
    new_new_n23817__, new_new_n23818__, new_new_n23819__, new_new_n23820__,
    new_new_n23822__, new_new_n23823__, new_new_n23824__, new_new_n23825__,
    new_new_n23826__, new_new_n23827__, new_new_n23829__, new_new_n23830__,
    new_new_n23831__, new_new_n23832__, new_new_n23833__, new_new_n23834__,
    new_new_n23836__, new_new_n23837__, new_new_n23838__, new_new_n23839__,
    new_new_n23840__, new_new_n23841__, new_new_n23843__, new_new_n23844__,
    new_new_n23845__, new_new_n23846__, new_new_n23847__, new_new_n23848__,
    new_new_n23850__, new_new_n23851__, new_new_n23852__, new_new_n23853__,
    new_new_n23854__, new_new_n23855__, new_new_n23857__, new_new_n23858__,
    new_new_n23859__, new_new_n23860__, new_new_n23861__, new_new_n23862__,
    new_new_n23864__, new_new_n23865__, new_new_n23866__, new_new_n23867__,
    new_new_n23868__, new_new_n23869__, new_new_n23871__, new_new_n23872__,
    new_new_n23873__, new_new_n23874__, new_new_n23875__, new_new_n23876__,
    new_new_n23878__, new_new_n23879__, new_new_n23880__, new_new_n23881__,
    new_new_n23882__, new_new_n23883__, new_new_n23885__, new_new_n23886__,
    new_new_n23887__, new_new_n23888__, new_new_n23889__, new_new_n23890__,
    new_new_n23892__, new_new_n23893__, new_new_n23894__, new_new_n23895__,
    new_new_n23896__, new_new_n23897__, new_new_n23899__, new_new_n23900__,
    new_new_n23901__, new_new_n23902__, new_new_n23903__, new_new_n23904__,
    new_new_n23906__, new_new_n23907__, new_new_n23908__, new_new_n23909__,
    new_new_n23910__, new_new_n23911__, new_new_n23913__, new_new_n23914__,
    new_new_n23915__, new_new_n23916__, new_new_n23917__, new_new_n23918__,
    new_new_n23920__, new_new_n23921__, new_new_n23922__;
  assign new_new_n257__ = ~pi089 & ~pi090;
  assign new_new_n258__ = ~pi088 & new_new_n257__;
  assign new_new_n259__ = ~pi097 & ~pi098;
  assign new_new_n260__ = ~pi126 & ~pi127;
  assign new_new_n261__ = ~pi124 & ~pi125;
  assign new_new_n262__ = new_new_n260__ & new_new_n261__;
  assign new_new_n263__ = ~pi122 & ~pi123;
  assign new_new_n264__ = new_new_n262__ & new_new_n263__;
  assign new_new_n265__ = ~pi117 & ~pi118;
  assign new_new_n266__ = ~pi119 & ~pi120;
  assign new_new_n267__ = ~pi121 & new_new_n266__;
  assign new_new_n268__ = new_new_n265__ & new_new_n267__;
  assign new_new_n269__ = new_new_n264__ & new_new_n268__;
  assign new_new_n270__ = ~pi112 & ~pi113;
  assign new_new_n271__ = ~pi114 & ~pi115;
  assign new_new_n272__ = ~pi116 & new_new_n271__;
  assign new_new_n273__ = new_new_n270__ & new_new_n272__;
  assign new_new_n274__ = new_new_n269__ & new_new_n273__;
  assign new_new_n275__ = ~pi107 & ~pi108;
  assign new_new_n276__ = ~pi109 & new_new_n275__;
  assign new_new_n277__ = ~pi110 & ~pi111;
  assign new_new_n278__ = new_new_n276__ & new_new_n277__;
  assign new_new_n279__ = new_new_n274__ & new_new_n278__;
  assign new_new_n280__ = ~pi105 & ~pi106;
  assign new_new_n281__ = ~pi102 & ~pi103;
  assign new_new_n282__ = ~pi104 & new_new_n281__;
  assign new_new_n283__ = new_new_n280__ & new_new_n282__;
  assign new_new_n284__ = new_new_n279__ & new_new_n283__;
  assign new_new_n285__ = ~pi099 & ~pi100;
  assign new_new_n286__ = ~pi101 & new_new_n285__;
  assign new_new_n287__ = new_new_n284__ & new_new_n286__;
  assign new_new_n288__ = ~pi096 & new_new_n259__;
  assign new_new_n289__ = new_new_n287__ & new_new_n288__;
  assign new_new_n290__ = ~pi091 & ~pi092;
  assign new_new_n291__ = ~pi093 & ~pi094;
  assign new_new_n292__ = new_new_n290__ & new_new_n291__;
  assign new_new_n293__ = ~pi095 & new_new_n292__;
  assign new_new_n294__ = new_new_n289__ & new_new_n293__;
  assign new_new_n295__ = ~pi086 & ~pi087;
  assign new_new_n296__ = new_new_n258__ & new_new_n295__;
  assign new_new_n297__ = new_new_n294__ & new_new_n296__;
  assign new_new_n298__ = ~pi083 & ~pi084;
  assign new_new_n299__ = ~pi085 & new_new_n298__;
  assign new_new_n300__ = ~pi081 & ~pi082;
  assign new_new_n301__ = new_new_n299__ & new_new_n300__;
  assign new_new_n302__ = new_new_n297__ & new_new_n301__;
  assign new_new_n303__ = ~pi078 & ~pi079;
  assign new_new_n304__ = ~pi080 & new_new_n303__;
  assign new_new_n305__ = new_new_n302__ & new_new_n304__;
  assign new_new_n306__ = ~pi077 & new_new_n305__;
  assign new_new_n307__ = ~pi074 & ~pi075;
  assign new_new_n308__ = ~pi076 & new_new_n307__;
  assign new_new_n309__ = new_new_n306__ & new_new_n308__;
  assign new_new_n310__ = ~pi071 & ~pi072;
  assign new_new_n311__ = ~pi073 & new_new_n310__;
  assign new_new_n312__ = new_new_n309__ & new_new_n311__;
  assign new_new_n313__ = ~pi068 & ~pi069;
  assign new_new_n314__ = ~pi070 & new_new_n313__;
  assign new_new_n315__ = new_new_n312__ & new_new_n314__;
  assign new_new_n316__ = ~pi067 & new_new_n315__;
  assign new_new_n317__ = ~pi061 & pi064;
  assign new_new_n318__ = ~pi065 & ~new_new_n317__;
  assign new_new_n319__ = ~pi066 & ~pi067;
  assign new_new_n320__ = ~pi063 & pi065;
  assign new_new_n321__ = new_new_n319__ & ~new_new_n320__;
  assign new_new_n322__ = new_new_n315__ & new_new_n321__;
  assign new_new_n323__ = ~pi061 & pi065;
  assign new_new_n324__ = ~new_new_n322__ & ~new_new_n323__;
  assign new_new_n325__ = pi064 & ~new_new_n324__;
  assign new_new_n326__ = pi062 & ~new_new_n325__;
  assign new_new_n327__ = ~new_new_n318__ & ~new_new_n326__;
  assign new_new_n328__ = ~pi066 & ~new_new_n327__;
  assign new_new_n329__ = pi066 & new_new_n327__;
  assign new_new_n330__ = new_new_n316__ & ~new_new_n329__;
  assign new_new_n331__ = ~new_new_n328__ & new_new_n330__;
  assign new_new_n332__ = ~pi064 & ~pi065;
  assign new_new_n333__ = ~pi062 & pi064;
  assign new_new_n334__ = pi065 & new_new_n333__;
  assign new_new_n335__ = ~pi066 & ~new_new_n332__;
  assign new_new_n336__ = ~new_new_n334__ & new_new_n335__;
  assign new_new_n337__ = new_new_n316__ & new_new_n336__;
  assign new_new_n338__ = pi063 & ~new_new_n337__;
  assign new_new_n339__ = ~new_new_n331__ & new_new_n338__;
  assign new_new_n340__ = ~new_new_n328__ & ~new_new_n338__;
  assign po061 = new_new_n330__ & ~new_new_n340__;
  assign new_new_n342__ = pi060 & ~pi065;
  assign new_new_n343__ = pi061 & ~new_new_n342__;
  assign new_new_n344__ = po061 & new_new_n343__;
  assign new_new_n345__ = ~pi061 & ~po061;
  assign new_new_n346__ = ~pi065 & ~new_new_n345__;
  assign new_new_n347__ = ~pi060 & ~new_new_n346__;
  assign new_new_n348__ = ~new_new_n344__ & ~new_new_n347__;
  assign new_new_n349__ = pi064 & ~new_new_n348__;
  assign new_new_n350__ = pi064 & po061;
  assign new_new_n351__ = new_new_n323__ & ~new_new_n350__;
  assign new_new_n352__ = ~new_new_n349__ & ~new_new_n351__;
  assign new_new_n353__ = pi066 & ~new_new_n352__;
  assign new_new_n354__ = ~pi066 & new_new_n352__;
  assign new_new_n355__ = ~pi062 & new_new_n332__;
  assign new_new_n356__ = pi061 & ~pi065;
  assign new_new_n357__ = po061 & ~new_new_n356__;
  assign new_new_n358__ = pi064 & new_new_n322__;
  assign new_new_n359__ = pi062 & ~new_new_n358__;
  assign new_new_n360__ = ~new_new_n357__ & ~new_new_n359__;
  assign new_new_n361__ = ~new_new_n318__ & new_new_n326__;
  assign new_new_n362__ = po061 & new_new_n361__;
  assign new_new_n363__ = pi062 & ~new_new_n322__;
  assign new_new_n364__ = pi065 & new_new_n317__;
  assign new_new_n365__ = ~new_new_n363__ & new_new_n364__;
  assign new_new_n366__ = ~new_new_n355__ & ~new_new_n365__;
  assign new_new_n367__ = ~new_new_n362__ & new_new_n366__;
  assign new_new_n368__ = ~new_new_n360__ & new_new_n367__;
  assign new_new_n369__ = ~new_new_n354__ & ~new_new_n368__;
  assign new_new_n370__ = ~new_new_n353__ & ~new_new_n369__;
  assign new_new_n371__ = pi067 & ~new_new_n370__;
  assign new_new_n372__ = ~pi067 & new_new_n370__;
  assign new_new_n373__ = new_new_n315__ & ~new_new_n371__;
  assign new_new_n374__ = ~new_new_n372__ & new_new_n373__;
  assign new_new_n375__ = new_new_n339__ & ~new_new_n374__;
  assign new_new_n376__ = new_new_n316__ & new_new_n375__;
  assign new_new_n377__ = ~pi068 & new_new_n375__;
  assign new_new_n378__ = ~new_new_n339__ & ~new_new_n370__;
  assign new_new_n379__ = ~pi067 & ~new_new_n378__;
  assign new_new_n380__ = pi063 & new_new_n370__;
  assign new_new_n381__ = ~new_new_n379__ & ~new_new_n380__;
  assign po060 = new_new_n315__ & ~new_new_n381__;
  assign new_new_n383__ = ~new_new_n353__ & ~new_new_n354__;
  assign new_new_n384__ = po060 & new_new_n383__;
  assign new_new_n385__ = new_new_n368__ & ~new_new_n384__;
  assign new_new_n386__ = ~new_new_n368__ & new_new_n384__;
  assign new_new_n387__ = ~new_new_n385__ & ~new_new_n386__;
  assign new_new_n388__ = pi067 & new_new_n387__;
  assign new_new_n389__ = ~pi067 & ~new_new_n387__;
  assign new_new_n390__ = ~pi060 & ~po060;
  assign new_new_n391__ = ~pi065 & ~new_new_n390__;
  assign new_new_n392__ = ~pi059 & ~new_new_n391__;
  assign new_new_n393__ = pi059 & ~pi065;
  assign new_new_n394__ = pi060 & ~new_new_n393__;
  assign new_new_n395__ = po060 & new_new_n394__;
  assign new_new_n396__ = ~new_new_n392__ & ~new_new_n395__;
  assign new_new_n397__ = pi064 & ~new_new_n396__;
  assign new_new_n398__ = ~pi060 & pi065;
  assign new_new_n399__ = pi064 & po060;
  assign new_new_n400__ = new_new_n398__ & ~new_new_n399__;
  assign new_new_n401__ = ~new_new_n397__ & ~new_new_n400__;
  assign new_new_n402__ = pi066 & ~new_new_n401__;
  assign new_new_n403__ = ~pi064 & pi065;
  assign new_new_n404__ = ~new_new_n342__ & ~new_new_n398__;
  assign new_new_n405__ = ~new_new_n332__ & new_new_n404__;
  assign new_new_n406__ = ~po061 & new_new_n405__;
  assign new_new_n407__ = ~new_new_n403__ & ~new_new_n406__;
  assign new_new_n408__ = po060 & ~new_new_n407__;
  assign new_new_n409__ = po060 & new_new_n404__;
  assign new_new_n410__ = new_new_n350__ & ~new_new_n409__;
  assign new_new_n411__ = ~new_new_n408__ & ~new_new_n410__;
  assign new_new_n412__ = ~pi061 & ~new_new_n411__;
  assign new_new_n413__ = pi061 & new_new_n411__;
  assign new_new_n414__ = ~new_new_n412__ & ~new_new_n413__;
  assign new_new_n415__ = ~pi066 & new_new_n401__;
  assign new_new_n416__ = new_new_n414__ & ~new_new_n415__;
  assign new_new_n417__ = ~new_new_n402__ & ~new_new_n416__;
  assign new_new_n418__ = ~new_new_n389__ & ~new_new_n417__;
  assign new_new_n419__ = ~new_new_n388__ & ~new_new_n418__;
  assign new_new_n420__ = ~new_new_n377__ & ~new_new_n419__;
  assign new_new_n421__ = pi068 & ~new_new_n375__;
  assign new_new_n422__ = ~pi070 & new_new_n312__;
  assign new_new_n423__ = ~pi069 & new_new_n422__;
  assign new_new_n424__ = ~new_new_n421__ & new_new_n423__;
  assign po059 = ~new_new_n420__ & new_new_n424__;
  assign new_new_n426__ = pi064 & pi065;
  assign new_new_n427__ = ~po059 & new_new_n426__;
  assign new_new_n428__ = ~pi065 & po059;
  assign new_new_n429__ = pi068 & ~new_new_n419__;
  assign new_new_n430__ = ~pi068 & new_new_n419__;
  assign new_new_n431__ = new_new_n423__ & ~new_new_n429__;
  assign new_new_n432__ = ~new_new_n430__ & new_new_n431__;
  assign new_new_n433__ = new_new_n375__ & ~new_new_n432__;
  assign new_new_n434__ = ~pi069 & new_new_n433__;
  assign new_new_n435__ = pi069 & ~new_new_n433__;
  assign new_new_n436__ = ~new_new_n402__ & ~new_new_n415__;
  assign new_new_n437__ = po059 & new_new_n436__;
  assign new_new_n438__ = ~new_new_n414__ & ~new_new_n437__;
  assign new_new_n439__ = new_new_n414__ & new_new_n437__;
  assign new_new_n440__ = ~new_new_n438__ & ~new_new_n439__;
  assign new_new_n441__ = ~pi067 & ~new_new_n440__;
  assign new_new_n442__ = pi067 & new_new_n440__;
  assign new_new_n443__ = pi059 & po059;
  assign new_new_n444__ = ~pi059 & ~po059;
  assign new_new_n445__ = ~pi065 & ~new_new_n443__;
  assign new_new_n446__ = ~new_new_n444__ & new_new_n445__;
  assign new_new_n447__ = ~pi058 & ~new_new_n446__;
  assign new_new_n448__ = pi065 & new_new_n443__;
  assign new_new_n449__ = ~new_new_n447__ & ~new_new_n448__;
  assign new_new_n450__ = pi064 & ~new_new_n449__;
  assign new_new_n451__ = pi064 & po059;
  assign new_new_n452__ = ~pi059 & pi065;
  assign new_new_n453__ = ~new_new_n451__ & new_new_n452__;
  assign new_new_n454__ = ~new_new_n450__ & ~new_new_n453__;
  assign new_new_n455__ = ~po060 & new_new_n426__;
  assign new_new_n456__ = po060 & new_new_n428__;
  assign new_new_n457__ = ~new_new_n455__ & ~new_new_n456__;
  assign new_new_n458__ = ~pi059 & ~new_new_n457__;
  assign new_new_n459__ = ~new_new_n332__ & po059;
  assign new_new_n460__ = ~new_new_n399__ & ~new_new_n459__;
  assign new_new_n461__ = pi065 & po059;
  assign new_new_n462__ = po060 & ~new_new_n461__;
  assign new_new_n463__ = pi065 & ~new_new_n399__;
  assign new_new_n464__ = pi059 & ~new_new_n463__;
  assign new_new_n465__ = ~new_new_n462__ & new_new_n464__;
  assign new_new_n466__ = ~new_new_n460__ & ~new_new_n465__;
  assign new_new_n467__ = ~new_new_n458__ & new_new_n466__;
  assign new_new_n468__ = ~pi060 & ~new_new_n467__;
  assign new_new_n469__ = ~new_new_n399__ & ~new_new_n461__;
  assign new_new_n470__ = pi065 & po060;
  assign new_new_n471__ = pi059 & ~new_new_n470__;
  assign new_new_n472__ = pi064 & ~new_new_n471__;
  assign new_new_n473__ = ~new_new_n469__ & ~new_new_n472__;
  assign new_new_n474__ = ~po060 & ~new_new_n428__;
  assign new_new_n475__ = pi064 & ~new_new_n443__;
  assign new_new_n476__ = ~new_new_n456__ & new_new_n475__;
  assign new_new_n477__ = ~new_new_n474__ & new_new_n476__;
  assign new_new_n478__ = ~new_new_n473__ & ~new_new_n477__;
  assign new_new_n479__ = pi060 & ~new_new_n478__;
  assign new_new_n480__ = ~new_new_n468__ & ~new_new_n479__;
  assign new_new_n481__ = ~pi066 & new_new_n480__;
  assign new_new_n482__ = ~new_new_n454__ & ~new_new_n481__;
  assign new_new_n483__ = pi066 & ~new_new_n480__;
  assign new_new_n484__ = ~new_new_n482__ & ~new_new_n483__;
  assign new_new_n485__ = ~new_new_n442__ & new_new_n484__;
  assign new_new_n486__ = ~new_new_n441__ & ~new_new_n485__;
  assign new_new_n487__ = ~pi068 & ~new_new_n486__;
  assign new_new_n488__ = ~new_new_n388__ & ~new_new_n389__;
  assign new_new_n489__ = ~new_new_n417__ & po059;
  assign new_new_n490__ = pi067 & ~po059;
  assign new_new_n491__ = ~new_new_n489__ & ~new_new_n490__;
  assign new_new_n492__ = new_new_n488__ & ~new_new_n491__;
  assign new_new_n493__ = ~new_new_n488__ & new_new_n491__;
  assign new_new_n494__ = ~new_new_n492__ & ~new_new_n493__;
  assign new_new_n495__ = pi068 & new_new_n486__;
  assign new_new_n496__ = ~new_new_n494__ & ~new_new_n495__;
  assign new_new_n497__ = ~new_new_n487__ & ~new_new_n496__;
  assign new_new_n498__ = ~new_new_n435__ & ~new_new_n497__;
  assign new_new_n499__ = ~new_new_n434__ & ~new_new_n498__;
  assign po058 = new_new_n422__ & ~new_new_n499__;
  assign new_new_n501__ = new_new_n428__ & po058;
  assign new_new_n502__ = ~new_new_n427__ & ~new_new_n501__;
  assign new_new_n503__ = ~pi058 & ~new_new_n502__;
  assign new_new_n504__ = ~new_new_n332__ & po058;
  assign new_new_n505__ = ~new_new_n451__ & ~new_new_n504__;
  assign new_new_n506__ = pi065 & po058;
  assign new_new_n507__ = po059 & ~new_new_n506__;
  assign new_new_n508__ = pi065 & ~new_new_n451__;
  assign new_new_n509__ = pi058 & ~new_new_n508__;
  assign new_new_n510__ = ~new_new_n507__ & new_new_n509__;
  assign new_new_n511__ = ~new_new_n503__ & ~new_new_n505__;
  assign new_new_n512__ = ~new_new_n510__ & new_new_n511__;
  assign new_new_n513__ = ~pi059 & ~new_new_n512__;
  assign new_new_n514__ = ~new_new_n451__ & ~new_new_n506__;
  assign new_new_n515__ = pi058 & ~new_new_n461__;
  assign new_new_n516__ = pi064 & ~new_new_n515__;
  assign new_new_n517__ = ~new_new_n514__ & ~new_new_n516__;
  assign new_new_n518__ = ~pi065 & po058;
  assign new_new_n519__ = ~po059 & ~new_new_n518__;
  assign new_new_n520__ = pi058 & po058;
  assign new_new_n521__ = pi064 & ~new_new_n501__;
  assign new_new_n522__ = ~new_new_n520__ & new_new_n521__;
  assign new_new_n523__ = ~new_new_n519__ & new_new_n522__;
  assign new_new_n524__ = ~new_new_n517__ & ~new_new_n523__;
  assign new_new_n525__ = pi059 & ~new_new_n524__;
  assign new_new_n526__ = ~new_new_n513__ & ~new_new_n525__;
  assign new_new_n527__ = pi057 & ~pi065;
  assign new_new_n528__ = new_new_n520__ & ~new_new_n527__;
  assign new_new_n529__ = ~pi058 & ~po058;
  assign new_new_n530__ = ~pi065 & ~new_new_n529__;
  assign new_new_n531__ = ~pi057 & ~new_new_n530__;
  assign new_new_n532__ = ~new_new_n528__ & ~new_new_n531__;
  assign new_new_n533__ = pi064 & ~new_new_n532__;
  assign new_new_n534__ = pi064 & po058;
  assign new_new_n535__ = ~pi058 & pi065;
  assign new_new_n536__ = ~new_new_n534__ & new_new_n535__;
  assign new_new_n537__ = ~new_new_n533__ & ~new_new_n536__;
  assign new_new_n538__ = ~pi066 & new_new_n537__;
  assign new_new_n539__ = pi066 & ~new_new_n537__;
  assign new_new_n540__ = pi070 & ~new_new_n433__;
  assign new_new_n541__ = ~new_new_n487__ & ~new_new_n495__;
  assign new_new_n542__ = po058 & new_new_n541__;
  assign new_new_n543__ = new_new_n494__ & ~new_new_n542__;
  assign new_new_n544__ = ~new_new_n494__ & new_new_n542__;
  assign new_new_n545__ = ~new_new_n543__ & ~new_new_n544__;
  assign new_new_n546__ = ~pi069 & new_new_n545__;
  assign new_new_n547__ = pi069 & ~new_new_n545__;
  assign new_new_n548__ = ~new_new_n441__ & ~new_new_n442__;
  assign new_new_n549__ = new_new_n484__ & po058;
  assign new_new_n550__ = ~pi067 & ~po058;
  assign new_new_n551__ = ~new_new_n549__ & ~new_new_n550__;
  assign new_new_n552__ = ~new_new_n548__ & ~new_new_n551__;
  assign new_new_n553__ = new_new_n548__ & new_new_n551__;
  assign new_new_n554__ = ~new_new_n552__ & ~new_new_n553__;
  assign new_new_n555__ = ~pi068 & ~new_new_n554__;
  assign new_new_n556__ = pi068 & new_new_n554__;
  assign new_new_n557__ = pi066 & ~new_new_n454__;
  assign new_new_n558__ = ~pi066 & new_new_n454__;
  assign new_new_n559__ = ~new_new_n557__ & ~new_new_n558__;
  assign new_new_n560__ = po058 & new_new_n559__;
  assign new_new_n561__ = new_new_n480__ & ~new_new_n560__;
  assign new_new_n562__ = ~new_new_n480__ & new_new_n560__;
  assign new_new_n563__ = ~new_new_n561__ & ~new_new_n562__;
  assign new_new_n564__ = ~pi067 & ~new_new_n563__;
  assign new_new_n565__ = pi067 & new_new_n563__;
  assign new_new_n566__ = ~new_new_n526__ & ~new_new_n538__;
  assign new_new_n567__ = ~new_new_n539__ & ~new_new_n566__;
  assign new_new_n568__ = ~new_new_n565__ & new_new_n567__;
  assign new_new_n569__ = ~new_new_n564__ & ~new_new_n568__;
  assign new_new_n570__ = ~new_new_n556__ & ~new_new_n569__;
  assign new_new_n571__ = ~new_new_n555__ & ~new_new_n570__;
  assign new_new_n572__ = ~new_new_n547__ & ~new_new_n571__;
  assign new_new_n573__ = ~new_new_n546__ & ~new_new_n572__;
  assign new_new_n574__ = ~new_new_n540__ & ~new_new_n573__;
  assign new_new_n575__ = new_new_n433__ & new_new_n499__;
  assign new_new_n576__ = ~new_new_n376__ & ~new_new_n575__;
  assign new_new_n577__ = ~new_new_n574__ & new_new_n576__;
  assign new_new_n578__ = pi070 & new_new_n573__;
  assign new_new_n579__ = new_new_n312__ & ~new_new_n578__;
  assign po057 = ~new_new_n577__ & new_new_n579__;
  assign new_new_n581__ = ~new_new_n539__ & po057;
  assign new_new_n582__ = ~new_new_n538__ & new_new_n581__;
  assign new_new_n583__ = new_new_n526__ & ~new_new_n582__;
  assign new_new_n584__ = new_new_n566__ & new_new_n581__;
  assign new_new_n585__ = ~new_new_n583__ & ~new_new_n584__;
  assign new_new_n586__ = pi057 & po057;
  assign new_new_n587__ = ~pi057 & ~po057;
  assign new_new_n588__ = ~pi065 & ~new_new_n586__;
  assign new_new_n589__ = ~new_new_n587__ & new_new_n588__;
  assign new_new_n590__ = ~pi056 & ~new_new_n589__;
  assign new_new_n591__ = pi065 & new_new_n586__;
  assign new_new_n592__ = ~new_new_n590__ & ~new_new_n591__;
  assign new_new_n593__ = pi064 & ~new_new_n592__;
  assign new_new_n594__ = pi064 & po057;
  assign new_new_n595__ = ~pi057 & pi065;
  assign new_new_n596__ = ~new_new_n594__ & new_new_n595__;
  assign new_new_n597__ = ~new_new_n593__ & ~new_new_n596__;
  assign new_new_n598__ = pi066 & ~new_new_n597__;
  assign new_new_n599__ = ~pi066 & new_new_n597__;
  assign new_new_n600__ = new_new_n426__ & ~po058;
  assign new_new_n601__ = new_new_n518__ & po057;
  assign new_new_n602__ = ~new_new_n600__ & ~new_new_n601__;
  assign new_new_n603__ = ~pi057 & ~new_new_n602__;
  assign new_new_n604__ = pi065 & po057;
  assign new_new_n605__ = po058 & ~new_new_n604__;
  assign new_new_n606__ = pi065 & ~new_new_n534__;
  assign new_new_n607__ = pi057 & ~new_new_n606__;
  assign new_new_n608__ = ~new_new_n605__ & new_new_n607__;
  assign new_new_n609__ = ~new_new_n332__ & po057;
  assign new_new_n610__ = ~new_new_n534__ & ~new_new_n609__;
  assign new_new_n611__ = ~new_new_n603__ & ~new_new_n610__;
  assign new_new_n612__ = ~new_new_n608__ & new_new_n611__;
  assign new_new_n613__ = pi058 & ~new_new_n612__;
  assign new_new_n614__ = ~pi064 & ~new_new_n604__;
  assign new_new_n615__ = ~pi065 & po057;
  assign new_new_n616__ = ~po058 & ~new_new_n615__;
  assign new_new_n617__ = ~new_new_n586__ & ~new_new_n601__;
  assign new_new_n618__ = ~new_new_n616__ & new_new_n617__;
  assign new_new_n619__ = pi064 & ~new_new_n618__;
  assign new_new_n620__ = ~new_new_n614__ & ~new_new_n619__;
  assign new_new_n621__ = ~new_new_n534__ & ~new_new_n604__;
  assign new_new_n622__ = pi057 & ~new_new_n506__;
  assign new_new_n623__ = ~new_new_n621__ & new_new_n622__;
  assign new_new_n624__ = ~new_new_n620__ & ~new_new_n623__;
  assign new_new_n625__ = ~pi058 & ~new_new_n624__;
  assign new_new_n626__ = ~new_new_n613__ & ~new_new_n625__;
  assign new_new_n627__ = ~new_new_n599__ & new_new_n626__;
  assign new_new_n628__ = ~new_new_n598__ & ~new_new_n627__;
  assign new_new_n629__ = pi067 & ~new_new_n628__;
  assign new_new_n630__ = ~pi067 & new_new_n628__;
  assign new_new_n631__ = ~pi073 & new_new_n309__;
  assign new_new_n632__ = ~pi072 & new_new_n631__;
  assign new_new_n633__ = ~new_new_n546__ & ~new_new_n547__;
  assign new_new_n634__ = ~new_new_n571__ & po057;
  assign new_new_n635__ = ~pi069 & ~po057;
  assign new_new_n636__ = ~new_new_n634__ & ~new_new_n635__;
  assign new_new_n637__ = new_new_n633__ & ~new_new_n636__;
  assign new_new_n638__ = ~new_new_n633__ & new_new_n636__;
  assign new_new_n639__ = ~new_new_n637__ & ~new_new_n638__;
  assign new_new_n640__ = ~new_new_n555__ & ~new_new_n556__;
  assign new_new_n641__ = ~new_new_n569__ & po057;
  assign new_new_n642__ = ~pi068 & ~po057;
  assign new_new_n643__ = ~new_new_n641__ & ~new_new_n642__;
  assign new_new_n644__ = new_new_n640__ & ~new_new_n643__;
  assign new_new_n645__ = ~new_new_n640__ & new_new_n643__;
  assign new_new_n646__ = ~new_new_n644__ & ~new_new_n645__;
  assign new_new_n647__ = pi069 & ~new_new_n646__;
  assign new_new_n648__ = ~pi069 & new_new_n646__;
  assign new_new_n649__ = ~new_new_n585__ & ~new_new_n629__;
  assign new_new_n650__ = ~new_new_n630__ & ~new_new_n649__;
  assign new_new_n651__ = ~pi068 & ~new_new_n650__;
  assign new_new_n652__ = pi068 & new_new_n650__;
  assign new_new_n653__ = ~new_new_n564__ & ~new_new_n565__;
  assign new_new_n654__ = new_new_n567__ & po057;
  assign new_new_n655__ = ~pi067 & ~po057;
  assign new_new_n656__ = ~new_new_n654__ & ~new_new_n655__;
  assign new_new_n657__ = ~new_new_n653__ & ~new_new_n656__;
  assign new_new_n658__ = new_new_n653__ & new_new_n656__;
  assign new_new_n659__ = ~new_new_n657__ & ~new_new_n658__;
  assign new_new_n660__ = ~new_new_n652__ & ~new_new_n659__;
  assign new_new_n661__ = ~new_new_n651__ & ~new_new_n660__;
  assign new_new_n662__ = ~new_new_n648__ & new_new_n661__;
  assign new_new_n663__ = ~new_new_n647__ & ~new_new_n662__;
  assign new_new_n664__ = ~pi070 & new_new_n663__;
  assign new_new_n665__ = ~new_new_n639__ & ~new_new_n664__;
  assign new_new_n666__ = pi070 & ~new_new_n663__;
  assign new_new_n667__ = new_new_n433__ & ~po058;
  assign new_new_n668__ = ~new_new_n376__ & ~new_new_n667__;
  assign new_new_n669__ = pi071 & new_new_n668__;
  assign new_new_n670__ = ~new_new_n666__ & ~new_new_n669__;
  assign new_new_n671__ = ~new_new_n665__ & new_new_n670__;
  assign new_new_n672__ = ~pi071 & ~new_new_n668__;
  assign new_new_n673__ = new_new_n578__ & new_new_n672__;
  assign new_new_n674__ = ~new_new_n671__ & ~new_new_n673__;
  assign po056 = new_new_n632__ & ~new_new_n674__;
  assign new_new_n676__ = ~new_new_n629__ & ~new_new_n630__;
  assign new_new_n677__ = po056 & new_new_n676__;
  assign new_new_n678__ = new_new_n585__ & ~new_new_n677__;
  assign new_new_n679__ = ~new_new_n585__ & new_new_n677__;
  assign new_new_n680__ = ~new_new_n678__ & ~new_new_n679__;
  assign new_new_n681__ = ~new_new_n598__ & ~new_new_n599__;
  assign new_new_n682__ = po056 & new_new_n681__;
  assign new_new_n683__ = new_new_n626__ & ~new_new_n682__;
  assign new_new_n684__ = ~new_new_n626__ & new_new_n682__;
  assign new_new_n685__ = ~new_new_n683__ & ~new_new_n684__;
  assign new_new_n686__ = pi067 & ~new_new_n685__;
  assign new_new_n687__ = ~pi067 & new_new_n685__;
  assign new_new_n688__ = ~pi056 & ~po056;
  assign new_new_n689__ = ~pi065 & ~new_new_n688__;
  assign new_new_n690__ = ~pi055 & ~new_new_n689__;
  assign new_new_n691__ = pi055 & ~pi065;
  assign new_new_n692__ = pi056 & ~new_new_n691__;
  assign new_new_n693__ = po056 & new_new_n692__;
  assign new_new_n694__ = ~new_new_n690__ & ~new_new_n693__;
  assign new_new_n695__ = pi064 & ~new_new_n694__;
  assign new_new_n696__ = pi064 & po056;
  assign new_new_n697__ = ~pi056 & pi065;
  assign new_new_n698__ = ~new_new_n696__ & new_new_n697__;
  assign new_new_n699__ = ~new_new_n695__ & ~new_new_n698__;
  assign new_new_n700__ = pi066 & ~new_new_n699__;
  assign new_new_n701__ = ~pi066 & new_new_n699__;
  assign new_new_n702__ = ~pi065 & po056;
  assign new_new_n703__ = ~po057 & ~new_new_n702__;
  assign new_new_n704__ = ~pi056 & ~new_new_n615__;
  assign new_new_n705__ = po056 & ~new_new_n704__;
  assign new_new_n706__ = pi064 & ~new_new_n705__;
  assign new_new_n707__ = ~new_new_n703__ & new_new_n706__;
  assign new_new_n708__ = pi065 & po056;
  assign new_new_n709__ = ~pi064 & new_new_n708__;
  assign new_new_n710__ = ~new_new_n594__ & ~new_new_n708__;
  assign new_new_n711__ = pi056 & ~new_new_n604__;
  assign new_new_n712__ = ~new_new_n710__ & new_new_n711__;
  assign new_new_n713__ = ~new_new_n707__ & ~new_new_n709__;
  assign new_new_n714__ = ~new_new_n712__ & new_new_n713__;
  assign new_new_n715__ = ~pi057 & ~new_new_n714__;
  assign new_new_n716__ = pi057 & new_new_n714__;
  assign new_new_n717__ = ~new_new_n715__ & ~new_new_n716__;
  assign new_new_n718__ = ~new_new_n701__ & new_new_n717__;
  assign new_new_n719__ = ~new_new_n700__ & ~new_new_n718__;
  assign new_new_n720__ = ~new_new_n687__ & ~new_new_n719__;
  assign new_new_n721__ = ~new_new_n686__ & ~new_new_n720__;
  assign new_new_n722__ = ~pi068 & new_new_n721__;
  assign new_new_n723__ = pi068 & ~new_new_n721__;
  assign new_new_n724__ = ~new_new_n664__ & ~new_new_n666__;
  assign new_new_n725__ = po056 & new_new_n724__;
  assign new_new_n726__ = new_new_n639__ & new_new_n725__;
  assign new_new_n727__ = ~new_new_n639__ & ~new_new_n725__;
  assign new_new_n728__ = ~new_new_n726__ & ~new_new_n727__;
  assign new_new_n729__ = ~pi071 & new_new_n728__;
  assign new_new_n730__ = ~new_new_n647__ & ~new_new_n648__;
  assign new_new_n731__ = ~new_new_n661__ & po056;
  assign new_new_n732__ = ~pi069 & ~po056;
  assign new_new_n733__ = ~new_new_n731__ & ~new_new_n732__;
  assign new_new_n734__ = new_new_n730__ & ~new_new_n733__;
  assign new_new_n735__ = ~new_new_n730__ & new_new_n733__;
  assign new_new_n736__ = ~new_new_n734__ & ~new_new_n735__;
  assign new_new_n737__ = ~pi070 & new_new_n736__;
  assign new_new_n738__ = pi070 & ~new_new_n736__;
  assign new_new_n739__ = ~new_new_n651__ & ~new_new_n652__;
  assign new_new_n740__ = po056 & new_new_n739__;
  assign new_new_n741__ = ~new_new_n659__ & ~new_new_n740__;
  assign new_new_n742__ = new_new_n659__ & new_new_n740__;
  assign new_new_n743__ = ~new_new_n741__ & ~new_new_n742__;
  assign new_new_n744__ = ~pi069 & ~new_new_n743__;
  assign new_new_n745__ = pi069 & new_new_n743__;
  assign new_new_n746__ = new_new_n680__ & ~new_new_n723__;
  assign new_new_n747__ = ~new_new_n722__ & ~new_new_n746__;
  assign new_new_n748__ = ~new_new_n745__ & ~new_new_n747__;
  assign new_new_n749__ = ~new_new_n744__ & ~new_new_n748__;
  assign new_new_n750__ = ~new_new_n738__ & ~new_new_n749__;
  assign new_new_n751__ = ~new_new_n737__ & ~new_new_n750__;
  assign new_new_n752__ = ~new_new_n729__ & new_new_n751__;
  assign new_new_n753__ = pi071 & ~new_new_n728__;
  assign new_new_n754__ = ~pi063 & pi072;
  assign new_new_n755__ = new_new_n631__ & ~new_new_n754__;
  assign new_new_n756__ = ~new_new_n753__ & new_new_n755__;
  assign new_new_n757__ = ~new_new_n752__ & new_new_n756__;
  assign new_new_n758__ = ~new_new_n376__ & ~new_new_n674__;
  assign new_new_n759__ = ~new_new_n376__ & po057;
  assign new_new_n760__ = ~new_new_n668__ & ~new_new_n759__;
  assign new_new_n761__ = new_new_n632__ & new_new_n760__;
  assign new_new_n762__ = ~new_new_n758__ & new_new_n761__;
  assign po055 = new_new_n757__ | new_new_n762__;
  assign new_new_n764__ = ~new_new_n722__ & ~new_new_n723__;
  assign new_new_n765__ = po055 & new_new_n764__;
  assign new_new_n766__ = new_new_n680__ & new_new_n765__;
  assign new_new_n767__ = ~new_new_n680__ & ~new_new_n765__;
  assign new_new_n768__ = ~new_new_n766__ & ~new_new_n767__;
  assign new_new_n769__ = pi069 & ~new_new_n768__;
  assign new_new_n770__ = ~pi069 & new_new_n768__;
  assign new_new_n771__ = ~new_new_n769__ & ~new_new_n770__;
  assign new_new_n772__ = ~new_new_n686__ & ~new_new_n687__;
  assign new_new_n773__ = new_new_n719__ & po055;
  assign new_new_n774__ = ~pi067 & ~po055;
  assign new_new_n775__ = ~new_new_n773__ & ~new_new_n774__;
  assign new_new_n776__ = new_new_n772__ & new_new_n775__;
  assign new_new_n777__ = ~new_new_n772__ & ~new_new_n775__;
  assign new_new_n778__ = ~new_new_n776__ & ~new_new_n777__;
  assign new_new_n779__ = pi068 & new_new_n778__;
  assign new_new_n780__ = ~pi068 & ~new_new_n778__;
  assign new_new_n781__ = ~new_new_n700__ & ~new_new_n701__;
  assign new_new_n782__ = po055 & new_new_n781__;
  assign new_new_n783__ = new_new_n717__ & ~new_new_n782__;
  assign new_new_n784__ = ~new_new_n717__ & new_new_n782__;
  assign new_new_n785__ = ~new_new_n783__ & ~new_new_n784__;
  assign new_new_n786__ = pi067 & ~new_new_n785__;
  assign new_new_n787__ = ~pi067 & new_new_n785__;
  assign new_new_n788__ = pi055 & po055;
  assign new_new_n789__ = pi054 & ~pi065;
  assign new_new_n790__ = new_new_n788__ & ~new_new_n789__;
  assign new_new_n791__ = ~pi055 & ~po055;
  assign new_new_n792__ = ~pi065 & ~new_new_n791__;
  assign new_new_n793__ = ~pi054 & ~new_new_n792__;
  assign new_new_n794__ = ~new_new_n790__ & ~new_new_n793__;
  assign new_new_n795__ = pi064 & ~new_new_n794__;
  assign new_new_n796__ = pi064 & po055;
  assign new_new_n797__ = ~pi055 & pi065;
  assign new_new_n798__ = ~new_new_n796__ & new_new_n797__;
  assign new_new_n799__ = ~new_new_n795__ & ~new_new_n798__;
  assign new_new_n800__ = pi066 & ~new_new_n799__;
  assign new_new_n801__ = pi065 & po055;
  assign new_new_n802__ = ~new_new_n696__ & ~new_new_n801__;
  assign new_new_n803__ = ~new_new_n796__ & new_new_n802__;
  assign new_new_n804__ = new_new_n426__ & ~po056;
  assign new_new_n805__ = new_new_n702__ & po055;
  assign new_new_n806__ = ~new_new_n804__ & ~new_new_n805__;
  assign new_new_n807__ = ~pi055 & ~new_new_n806__;
  assign new_new_n808__ = po056 & ~new_new_n801__;
  assign new_new_n809__ = pi065 & ~new_new_n696__;
  assign new_new_n810__ = pi055 & ~new_new_n809__;
  assign new_new_n811__ = ~new_new_n808__ & new_new_n810__;
  assign new_new_n812__ = ~new_new_n803__ & ~new_new_n807__;
  assign new_new_n813__ = ~new_new_n811__ & new_new_n812__;
  assign new_new_n814__ = ~pi056 & ~new_new_n813__;
  assign new_new_n815__ = pi055 & ~new_new_n708__;
  assign new_new_n816__ = pi064 & ~new_new_n815__;
  assign new_new_n817__ = ~new_new_n802__ & ~new_new_n816__;
  assign new_new_n818__ = ~pi065 & po055;
  assign new_new_n819__ = ~po056 & ~new_new_n818__;
  assign new_new_n820__ = pi064 & ~new_new_n788__;
  assign new_new_n821__ = ~new_new_n805__ & new_new_n820__;
  assign new_new_n822__ = ~new_new_n819__ & new_new_n821__;
  assign new_new_n823__ = ~new_new_n817__ & ~new_new_n822__;
  assign new_new_n824__ = pi056 & ~new_new_n823__;
  assign new_new_n825__ = ~new_new_n814__ & ~new_new_n824__;
  assign new_new_n826__ = ~pi066 & new_new_n799__;
  assign new_new_n827__ = ~new_new_n825__ & ~new_new_n826__;
  assign new_new_n828__ = ~new_new_n800__ & ~new_new_n827__;
  assign new_new_n829__ = ~new_new_n787__ & ~new_new_n828__;
  assign new_new_n830__ = ~new_new_n786__ & ~new_new_n829__;
  assign new_new_n831__ = ~new_new_n780__ & ~new_new_n830__;
  assign new_new_n832__ = ~new_new_n779__ & ~new_new_n831__;
  assign new_new_n833__ = ~new_new_n757__ & new_new_n760__;
  assign new_new_n834__ = ~new_new_n632__ & new_new_n833__;
  assign new_new_n835__ = ~pi073 & new_new_n834__;
  assign new_new_n836__ = ~new_new_n737__ & ~new_new_n738__;
  assign new_new_n837__ = ~pi070 & ~po055;
  assign new_new_n838__ = ~new_new_n749__ & po055;
  assign new_new_n839__ = ~new_new_n837__ & ~new_new_n838__;
  assign new_new_n840__ = new_new_n836__ & ~new_new_n839__;
  assign new_new_n841__ = ~new_new_n836__ & new_new_n839__;
  assign new_new_n842__ = ~new_new_n840__ & ~new_new_n841__;
  assign new_new_n843__ = pi071 & ~new_new_n842__;
  assign new_new_n844__ = ~pi071 & new_new_n842__;
  assign new_new_n845__ = ~new_new_n744__ & ~new_new_n745__;
  assign new_new_n846__ = ~pi069 & ~po055;
  assign new_new_n847__ = ~new_new_n747__ & po055;
  assign new_new_n848__ = ~new_new_n846__ & ~new_new_n847__;
  assign new_new_n849__ = new_new_n845__ & ~new_new_n848__;
  assign new_new_n850__ = ~new_new_n845__ & new_new_n848__;
  assign new_new_n851__ = ~new_new_n849__ & ~new_new_n850__;
  assign new_new_n852__ = pi070 & ~new_new_n851__;
  assign new_new_n853__ = ~pi070 & new_new_n851__;
  assign new_new_n854__ = ~new_new_n770__ & ~new_new_n832__;
  assign new_new_n855__ = ~new_new_n769__ & ~new_new_n854__;
  assign new_new_n856__ = ~new_new_n853__ & ~new_new_n855__;
  assign new_new_n857__ = ~new_new_n852__ & ~new_new_n856__;
  assign new_new_n858__ = ~new_new_n844__ & ~new_new_n857__;
  assign new_new_n859__ = ~new_new_n843__ & ~new_new_n858__;
  assign new_new_n860__ = pi072 & ~new_new_n859__;
  assign new_new_n861__ = pi073 & ~new_new_n833__;
  assign new_new_n862__ = ~new_new_n860__ & ~new_new_n861__;
  assign new_new_n863__ = ~new_new_n729__ & ~new_new_n753__;
  assign new_new_n864__ = ~new_new_n751__ & po055;
  assign new_new_n865__ = ~pi071 & ~po055;
  assign new_new_n866__ = ~new_new_n864__ & ~new_new_n865__;
  assign new_new_n867__ = new_new_n863__ & ~new_new_n866__;
  assign new_new_n868__ = ~new_new_n863__ & new_new_n866__;
  assign new_new_n869__ = ~new_new_n867__ & ~new_new_n868__;
  assign new_new_n870__ = ~pi072 & new_new_n859__;
  assign new_new_n871__ = ~new_new_n869__ & ~new_new_n870__;
  assign new_new_n872__ = new_new_n862__ & ~new_new_n871__;
  assign new_new_n873__ = ~new_new_n835__ & ~new_new_n872__;
  assign po054 = new_new_n309__ & ~new_new_n873__;
  assign new_new_n875__ = ~new_new_n832__ & po054;
  assign new_new_n876__ = pi069 & ~po054;
  assign new_new_n877__ = ~new_new_n875__ & ~new_new_n876__;
  assign new_new_n878__ = new_new_n771__ & new_new_n877__;
  assign new_new_n879__ = ~new_new_n771__ & ~new_new_n877__;
  assign new_new_n880__ = ~new_new_n878__ & ~new_new_n879__;
  assign new_new_n881__ = new_new_n830__ & po054;
  assign new_new_n882__ = ~pi068 & ~po054;
  assign new_new_n883__ = ~new_new_n881__ & ~new_new_n882__;
  assign new_new_n884__ = ~new_new_n779__ & ~new_new_n780__;
  assign new_new_n885__ = ~new_new_n883__ & ~new_new_n884__;
  assign new_new_n886__ = new_new_n883__ & new_new_n884__;
  assign new_new_n887__ = ~new_new_n885__ & ~new_new_n886__;
  assign new_new_n888__ = ~pi069 & ~new_new_n887__;
  assign new_new_n889__ = ~pi067 & ~new_new_n828__;
  assign new_new_n890__ = pi067 & new_new_n828__;
  assign new_new_n891__ = ~new_new_n889__ & ~new_new_n890__;
  assign new_new_n892__ = po054 & ~new_new_n891__;
  assign new_new_n893__ = new_new_n785__ & new_new_n892__;
  assign new_new_n894__ = ~new_new_n785__ & ~new_new_n892__;
  assign new_new_n895__ = ~new_new_n893__ & ~new_new_n894__;
  assign new_new_n896__ = pi068 & ~new_new_n895__;
  assign new_new_n897__ = ~pi068 & new_new_n895__;
  assign new_new_n898__ = ~new_new_n800__ & ~new_new_n826__;
  assign new_new_n899__ = po054 & new_new_n898__;
  assign new_new_n900__ = new_new_n825__ & ~new_new_n899__;
  assign new_new_n901__ = ~new_new_n825__ & new_new_n899__;
  assign new_new_n902__ = ~new_new_n900__ & ~new_new_n901__;
  assign new_new_n903__ = pi067 & new_new_n902__;
  assign new_new_n904__ = ~pi067 & ~new_new_n902__;
  assign new_new_n905__ = pi054 & po054;
  assign new_new_n906__ = pi053 & ~pi065;
  assign new_new_n907__ = new_new_n905__ & ~new_new_n906__;
  assign new_new_n908__ = ~pi054 & ~po054;
  assign new_new_n909__ = ~pi065 & ~new_new_n908__;
  assign new_new_n910__ = ~pi053 & ~new_new_n909__;
  assign new_new_n911__ = ~new_new_n907__ & ~new_new_n910__;
  assign new_new_n912__ = pi064 & ~new_new_n911__;
  assign new_new_n913__ = pi064 & po054;
  assign new_new_n914__ = ~pi054 & pi065;
  assign new_new_n915__ = ~new_new_n913__ & new_new_n914__;
  assign new_new_n916__ = ~new_new_n912__ & ~new_new_n915__;
  assign new_new_n917__ = pi066 & ~new_new_n916__;
  assign new_new_n918__ = ~pi066 & new_new_n916__;
  assign new_new_n919__ = new_new_n426__ & ~po055;
  assign new_new_n920__ = new_new_n818__ & po054;
  assign new_new_n921__ = ~new_new_n919__ & ~new_new_n920__;
  assign new_new_n922__ = ~pi054 & ~new_new_n921__;
  assign new_new_n923__ = ~new_new_n332__ & po054;
  assign new_new_n924__ = ~new_new_n796__ & ~new_new_n923__;
  assign new_new_n925__ = pi065 & ~new_new_n796__;
  assign new_new_n926__ = pi065 & po054;
  assign new_new_n927__ = po055 & ~new_new_n926__;
  assign new_new_n928__ = pi054 & ~new_new_n925__;
  assign new_new_n929__ = ~new_new_n927__ & new_new_n928__;
  assign new_new_n930__ = ~new_new_n922__ & ~new_new_n924__;
  assign new_new_n931__ = ~new_new_n929__ & new_new_n930__;
  assign new_new_n932__ = pi055 & ~new_new_n931__;
  assign new_new_n933__ = ~new_new_n796__ & ~new_new_n926__;
  assign new_new_n934__ = pi054 & ~new_new_n801__;
  assign new_new_n935__ = pi064 & ~new_new_n934__;
  assign new_new_n936__ = ~new_new_n933__ & ~new_new_n935__;
  assign new_new_n937__ = ~pi065 & po054;
  assign new_new_n938__ = ~po055 & ~new_new_n937__;
  assign new_new_n939__ = pi064 & ~new_new_n905__;
  assign new_new_n940__ = ~new_new_n920__ & new_new_n939__;
  assign new_new_n941__ = ~new_new_n938__ & new_new_n940__;
  assign new_new_n942__ = ~new_new_n936__ & ~new_new_n941__;
  assign new_new_n943__ = ~pi055 & ~new_new_n942__;
  assign new_new_n944__ = ~new_new_n932__ & ~new_new_n943__;
  assign new_new_n945__ = ~new_new_n918__ & new_new_n944__;
  assign new_new_n946__ = ~new_new_n917__ & ~new_new_n945__;
  assign new_new_n947__ = ~new_new_n904__ & ~new_new_n946__;
  assign new_new_n948__ = ~new_new_n903__ & ~new_new_n947__;
  assign new_new_n949__ = ~new_new_n897__ & ~new_new_n948__;
  assign new_new_n950__ = ~new_new_n896__ & ~new_new_n949__;
  assign new_new_n951__ = pi069 & new_new_n887__;
  assign new_new_n952__ = new_new_n950__ & ~new_new_n951__;
  assign new_new_n953__ = ~new_new_n888__ & ~new_new_n952__;
  assign new_new_n954__ = pi070 & new_new_n953__;
  assign new_new_n955__ = ~pi070 & ~new_new_n953__;
  assign new_new_n956__ = new_new_n309__ & ~new_new_n870__;
  assign new_new_n957__ = new_new_n862__ & new_new_n956__;
  assign new_new_n958__ = new_new_n869__ & ~new_new_n957__;
  assign new_new_n959__ = new_new_n631__ & new_new_n834__;
  assign new_new_n960__ = ~new_new_n860__ & new_new_n959__;
  assign new_new_n961__ = new_new_n871__ & new_new_n960__;
  assign new_new_n962__ = ~new_new_n958__ & ~new_new_n961__;
  assign new_new_n963__ = ~pi073 & ~new_new_n962__;
  assign new_new_n964__ = pi073 & ~new_new_n958__;
  assign new_new_n965__ = pi071 & ~new_new_n857__;
  assign new_new_n966__ = ~pi071 & new_new_n857__;
  assign new_new_n967__ = ~new_new_n965__ & ~new_new_n966__;
  assign new_new_n968__ = po054 & new_new_n967__;
  assign new_new_n969__ = new_new_n842__ & new_new_n968__;
  assign new_new_n970__ = ~new_new_n842__ & ~new_new_n968__;
  assign new_new_n971__ = ~new_new_n969__ & ~new_new_n970__;
  assign new_new_n972__ = pi072 & ~new_new_n971__;
  assign new_new_n973__ = ~pi072 & new_new_n971__;
  assign new_new_n974__ = ~new_new_n855__ & po054;
  assign new_new_n975__ = pi070 & ~po054;
  assign new_new_n976__ = ~new_new_n974__ & ~new_new_n975__;
  assign new_new_n977__ = ~new_new_n852__ & ~new_new_n853__;
  assign new_new_n978__ = ~new_new_n976__ & new_new_n977__;
  assign new_new_n979__ = new_new_n976__ & ~new_new_n977__;
  assign new_new_n980__ = ~new_new_n978__ & ~new_new_n979__;
  assign new_new_n981__ = ~pi071 & ~new_new_n980__;
  assign new_new_n982__ = pi071 & new_new_n980__;
  assign new_new_n983__ = ~new_new_n880__ & ~new_new_n955__;
  assign new_new_n984__ = ~new_new_n954__ & ~new_new_n983__;
  assign new_new_n985__ = ~new_new_n982__ & new_new_n984__;
  assign new_new_n986__ = ~new_new_n981__ & ~new_new_n985__;
  assign new_new_n987__ = ~new_new_n973__ & new_new_n986__;
  assign new_new_n988__ = ~new_new_n972__ & ~new_new_n987__;
  assign new_new_n989__ = ~new_new_n964__ & new_new_n988__;
  assign new_new_n990__ = ~new_new_n963__ & ~new_new_n989__;
  assign new_new_n991__ = pi074 & new_new_n990__;
  assign new_new_n992__ = ~pi076 & new_new_n306__;
  assign new_new_n993__ = ~pi075 & new_new_n992__;
  assign new_new_n994__ = ~new_new_n991__ & new_new_n993__;
  assign new_new_n995__ = ~pi074 & ~new_new_n990__;
  assign new_new_n996__ = new_new_n834__ & ~po054;
  assign new_new_n997__ = ~new_new_n376__ & ~new_new_n996__;
  assign new_new_n998__ = ~new_new_n995__ & new_new_n997__;
  assign po053 = new_new_n994__ & ~new_new_n998__;
  assign new_new_n1000__ = ~new_new_n954__ & ~new_new_n955__;
  assign new_new_n1001__ = po053 & new_new_n1000__;
  assign new_new_n1002__ = ~new_new_n880__ & ~new_new_n1001__;
  assign new_new_n1003__ = new_new_n880__ & new_new_n1001__;
  assign new_new_n1004__ = ~new_new_n1002__ & ~new_new_n1003__;
  assign new_new_n1005__ = ~pi071 & new_new_n1004__;
  assign new_new_n1006__ = pi071 & ~new_new_n1004__;
  assign new_new_n1007__ = ~new_new_n1005__ & ~new_new_n1006__;
  assign new_new_n1008__ = ~new_new_n888__ & ~new_new_n951__;
  assign new_new_n1009__ = new_new_n950__ & po053;
  assign new_new_n1010__ = ~pi069 & ~po053;
  assign new_new_n1011__ = ~new_new_n1009__ & ~new_new_n1010__;
  assign new_new_n1012__ = ~new_new_n1008__ & ~new_new_n1011__;
  assign new_new_n1013__ = new_new_n1008__ & new_new_n1011__;
  assign new_new_n1014__ = ~new_new_n1012__ & ~new_new_n1013__;
  assign new_new_n1015__ = ~pi070 & ~new_new_n1014__;
  assign new_new_n1016__ = pi070 & new_new_n1014__;
  assign new_new_n1017__ = ~new_new_n948__ & po053;
  assign new_new_n1018__ = pi068 & ~po053;
  assign new_new_n1019__ = ~new_new_n1017__ & ~new_new_n1018__;
  assign new_new_n1020__ = ~new_new_n896__ & ~new_new_n897__;
  assign new_new_n1021__ = ~new_new_n1019__ & new_new_n1020__;
  assign new_new_n1022__ = new_new_n1019__ & ~new_new_n1020__;
  assign new_new_n1023__ = ~new_new_n1021__ & ~new_new_n1022__;
  assign new_new_n1024__ = ~pi069 & ~new_new_n1023__;
  assign new_new_n1025__ = pi069 & new_new_n1023__;
  assign new_new_n1026__ = ~new_new_n917__ & ~new_new_n918__;
  assign new_new_n1027__ = po053 & new_new_n1026__;
  assign new_new_n1028__ = new_new_n944__ & ~new_new_n1027__;
  assign new_new_n1029__ = ~new_new_n944__ & new_new_n1027__;
  assign new_new_n1030__ = ~new_new_n1028__ & ~new_new_n1029__;
  assign new_new_n1031__ = pi067 & ~new_new_n1030__;
  assign new_new_n1032__ = ~pi067 & new_new_n1030__;
  assign new_new_n1033__ = pi053 & po053;
  assign new_new_n1034__ = ~pi053 & ~po053;
  assign new_new_n1035__ = ~pi065 & ~new_new_n1033__;
  assign new_new_n1036__ = ~new_new_n1034__ & new_new_n1035__;
  assign new_new_n1037__ = ~pi052 & ~new_new_n1036__;
  assign new_new_n1038__ = pi065 & new_new_n1033__;
  assign new_new_n1039__ = ~new_new_n1037__ & ~new_new_n1038__;
  assign new_new_n1040__ = pi064 & ~new_new_n1039__;
  assign new_new_n1041__ = pi064 & po053;
  assign new_new_n1042__ = ~pi053 & pi065;
  assign new_new_n1043__ = ~new_new_n1041__ & new_new_n1042__;
  assign new_new_n1044__ = ~new_new_n1040__ & ~new_new_n1043__;
  assign new_new_n1045__ = pi066 & ~new_new_n1044__;
  assign new_new_n1046__ = ~pi066 & new_new_n1044__;
  assign new_new_n1047__ = new_new_n426__ & ~po054;
  assign new_new_n1048__ = new_new_n937__ & po053;
  assign new_new_n1049__ = ~new_new_n1047__ & ~new_new_n1048__;
  assign new_new_n1050__ = ~pi053 & ~new_new_n1049__;
  assign new_new_n1051__ = ~new_new_n332__ & po053;
  assign new_new_n1052__ = ~new_new_n913__ & ~new_new_n1051__;
  assign new_new_n1053__ = pi065 & po053;
  assign new_new_n1054__ = po054 & ~new_new_n1053__;
  assign new_new_n1055__ = pi065 & ~new_new_n913__;
  assign new_new_n1056__ = pi053 & ~new_new_n1055__;
  assign new_new_n1057__ = ~new_new_n1054__ & new_new_n1056__;
  assign new_new_n1058__ = ~new_new_n1050__ & ~new_new_n1052__;
  assign new_new_n1059__ = ~new_new_n1057__ & new_new_n1058__;
  assign new_new_n1060__ = pi054 & ~new_new_n1059__;
  assign new_new_n1061__ = ~pi064 & ~new_new_n1053__;
  assign new_new_n1062__ = ~pi065 & po053;
  assign new_new_n1063__ = ~po054 & ~new_new_n1062__;
  assign new_new_n1064__ = ~new_new_n1033__ & ~new_new_n1048__;
  assign new_new_n1065__ = ~new_new_n1063__ & new_new_n1064__;
  assign new_new_n1066__ = pi064 & ~new_new_n1065__;
  assign new_new_n1067__ = ~new_new_n1061__ & ~new_new_n1066__;
  assign new_new_n1068__ = ~new_new_n913__ & ~new_new_n1053__;
  assign new_new_n1069__ = pi053 & ~new_new_n926__;
  assign new_new_n1070__ = ~new_new_n1068__ & new_new_n1069__;
  assign new_new_n1071__ = ~new_new_n1067__ & ~new_new_n1070__;
  assign new_new_n1072__ = ~pi054 & ~new_new_n1071__;
  assign new_new_n1073__ = ~new_new_n1060__ & ~new_new_n1072__;
  assign new_new_n1074__ = ~new_new_n1046__ & new_new_n1073__;
  assign new_new_n1075__ = ~new_new_n1045__ & ~new_new_n1074__;
  assign new_new_n1076__ = ~new_new_n1032__ & ~new_new_n1075__;
  assign new_new_n1077__ = ~new_new_n1031__ & ~new_new_n1076__;
  assign new_new_n1078__ = ~pi068 & new_new_n1077__;
  assign new_new_n1079__ = pi068 & ~new_new_n1077__;
  assign new_new_n1080__ = ~new_new_n903__ & ~new_new_n904__;
  assign new_new_n1081__ = ~new_new_n946__ & po053;
  assign new_new_n1082__ = pi067 & ~po053;
  assign new_new_n1083__ = ~new_new_n1081__ & ~new_new_n1082__;
  assign new_new_n1084__ = new_new_n1080__ & ~new_new_n1083__;
  assign new_new_n1085__ = ~new_new_n1080__ & new_new_n1083__;
  assign new_new_n1086__ = ~new_new_n1084__ & ~new_new_n1085__;
  assign new_new_n1087__ = ~new_new_n1079__ & ~new_new_n1086__;
  assign new_new_n1088__ = ~new_new_n1078__ & ~new_new_n1087__;
  assign new_new_n1089__ = ~new_new_n1025__ & ~new_new_n1088__;
  assign new_new_n1090__ = ~new_new_n1024__ & ~new_new_n1089__;
  assign new_new_n1091__ = ~new_new_n1016__ & ~new_new_n1090__;
  assign new_new_n1092__ = ~new_new_n1015__ & ~new_new_n1091__;
  assign new_new_n1093__ = pi073 & ~new_new_n988__;
  assign new_new_n1094__ = ~pi073 & new_new_n988__;
  assign new_new_n1095__ = ~new_new_n1093__ & ~new_new_n1094__;
  assign new_new_n1096__ = po053 & new_new_n1095__;
  assign new_new_n1097__ = ~new_new_n962__ & new_new_n1096__;
  assign new_new_n1098__ = new_new_n962__ & ~new_new_n1096__;
  assign new_new_n1099__ = ~new_new_n1097__ & ~new_new_n1098__;
  assign new_new_n1100__ = pi074 & ~new_new_n1099__;
  assign new_new_n1101__ = ~pi074 & new_new_n1099__;
  assign new_new_n1102__ = new_new_n986__ & po053;
  assign new_new_n1103__ = pi072 & ~po053;
  assign new_new_n1104__ = ~new_new_n1102__ & ~new_new_n1103__;
  assign new_new_n1105__ = ~new_new_n972__ & ~new_new_n973__;
  assign new_new_n1106__ = ~new_new_n1104__ & ~new_new_n1105__;
  assign new_new_n1107__ = new_new_n1104__ & new_new_n1105__;
  assign new_new_n1108__ = ~new_new_n1106__ & ~new_new_n1107__;
  assign new_new_n1109__ = pi073 & ~new_new_n1108__;
  assign new_new_n1110__ = ~pi073 & new_new_n1108__;
  assign new_new_n1111__ = ~new_new_n981__ & ~new_new_n982__;
  assign new_new_n1112__ = ~new_new_n984__ & po053;
  assign new_new_n1113__ = pi071 & ~po053;
  assign new_new_n1114__ = ~new_new_n1112__ & ~new_new_n1113__;
  assign new_new_n1115__ = new_new_n1111__ & ~new_new_n1114__;
  assign new_new_n1116__ = ~new_new_n1111__ & new_new_n1114__;
  assign new_new_n1117__ = ~new_new_n1115__ & ~new_new_n1116__;
  assign new_new_n1118__ = ~pi072 & ~new_new_n1117__;
  assign new_new_n1119__ = pi072 & new_new_n1117__;
  assign new_new_n1120__ = ~new_new_n1006__ & ~new_new_n1092__;
  assign new_new_n1121__ = ~new_new_n1005__ & ~new_new_n1120__;
  assign new_new_n1122__ = ~new_new_n1119__ & ~new_new_n1121__;
  assign new_new_n1123__ = ~new_new_n1118__ & ~new_new_n1122__;
  assign new_new_n1124__ = ~new_new_n1110__ & new_new_n1123__;
  assign new_new_n1125__ = ~new_new_n1109__ & ~new_new_n1124__;
  assign new_new_n1126__ = ~new_new_n1101__ & ~new_new_n1125__;
  assign new_new_n1127__ = ~new_new_n1100__ & ~new_new_n1126__;
  assign new_new_n1128__ = pi075 & ~new_new_n1127__;
  assign new_new_n1129__ = new_new_n992__ & ~new_new_n1128__;
  assign new_new_n1130__ = ~pi075 & new_new_n1127__;
  assign new_new_n1131__ = ~new_new_n994__ & new_new_n996__;
  assign new_new_n1132__ = ~new_new_n376__ & ~new_new_n1131__;
  assign new_new_n1133__ = ~new_new_n1130__ & new_new_n1132__;
  assign po052 = new_new_n1129__ & ~new_new_n1133__;
  assign new_new_n1135__ = ~new_new_n1092__ & po052;
  assign new_new_n1136__ = ~pi071 & ~po052;
  assign new_new_n1137__ = ~new_new_n1135__ & ~new_new_n1136__;
  assign new_new_n1138__ = new_new_n1007__ & ~new_new_n1137__;
  assign new_new_n1139__ = ~new_new_n1007__ & new_new_n1137__;
  assign new_new_n1140__ = ~new_new_n1138__ & ~new_new_n1139__;
  assign new_new_n1141__ = ~pi072 & new_new_n1140__;
  assign new_new_n1142__ = pi072 & ~new_new_n1140__;
  assign new_new_n1143__ = ~new_new_n1141__ & ~new_new_n1142__;
  assign new_new_n1144__ = ~new_new_n1015__ & ~new_new_n1016__;
  assign new_new_n1145__ = ~new_new_n1090__ & po052;
  assign new_new_n1146__ = ~pi070 & ~po052;
  assign new_new_n1147__ = ~new_new_n1145__ & ~new_new_n1146__;
  assign new_new_n1148__ = new_new_n1144__ & ~new_new_n1147__;
  assign new_new_n1149__ = ~new_new_n1144__ & new_new_n1147__;
  assign new_new_n1150__ = ~new_new_n1148__ & ~new_new_n1149__;
  assign new_new_n1151__ = ~pi071 & new_new_n1150__;
  assign new_new_n1152__ = pi071 & ~new_new_n1150__;
  assign new_new_n1153__ = ~new_new_n1024__ & ~new_new_n1025__;
  assign new_new_n1154__ = ~new_new_n1088__ & po052;
  assign new_new_n1155__ = ~pi069 & ~po052;
  assign new_new_n1156__ = ~new_new_n1154__ & ~new_new_n1155__;
  assign new_new_n1157__ = ~new_new_n1153__ & ~new_new_n1156__;
  assign new_new_n1158__ = new_new_n1153__ & new_new_n1156__;
  assign new_new_n1159__ = ~new_new_n1157__ & ~new_new_n1158__;
  assign new_new_n1160__ = ~pi070 & ~new_new_n1159__;
  assign new_new_n1161__ = pi070 & new_new_n1159__;
  assign new_new_n1162__ = ~new_new_n1078__ & ~new_new_n1079__;
  assign new_new_n1163__ = po052 & new_new_n1162__;
  assign new_new_n1164__ = new_new_n1086__ & new_new_n1163__;
  assign new_new_n1165__ = ~new_new_n1086__ & ~new_new_n1163__;
  assign new_new_n1166__ = ~new_new_n1164__ & ~new_new_n1165__;
  assign new_new_n1167__ = ~pi069 & ~new_new_n1166__;
  assign new_new_n1168__ = pi069 & new_new_n1166__;
  assign new_new_n1169__ = ~new_new_n1045__ & ~new_new_n1046__;
  assign new_new_n1170__ = po052 & new_new_n1169__;
  assign new_new_n1171__ = new_new_n1073__ & ~new_new_n1170__;
  assign new_new_n1172__ = ~new_new_n1073__ & new_new_n1170__;
  assign new_new_n1173__ = ~new_new_n1171__ & ~new_new_n1172__;
  assign new_new_n1174__ = pi067 & ~new_new_n1173__;
  assign new_new_n1175__ = ~pi067 & new_new_n1173__;
  assign new_new_n1176__ = pi052 & po052;
  assign new_new_n1177__ = ~pi052 & ~po052;
  assign new_new_n1178__ = ~pi065 & ~new_new_n1176__;
  assign new_new_n1179__ = ~new_new_n1177__ & new_new_n1178__;
  assign new_new_n1180__ = ~pi051 & ~new_new_n1179__;
  assign new_new_n1181__ = pi065 & new_new_n1176__;
  assign new_new_n1182__ = ~new_new_n1180__ & ~new_new_n1181__;
  assign new_new_n1183__ = pi064 & ~new_new_n1182__;
  assign new_new_n1184__ = pi064 & po052;
  assign new_new_n1185__ = ~pi052 & pi065;
  assign new_new_n1186__ = ~new_new_n1184__ & new_new_n1185__;
  assign new_new_n1187__ = ~new_new_n1183__ & ~new_new_n1186__;
  assign new_new_n1188__ = pi066 & ~new_new_n1187__;
  assign new_new_n1189__ = new_new_n426__ & ~po053;
  assign new_new_n1190__ = new_new_n1062__ & po052;
  assign new_new_n1191__ = ~new_new_n1189__ & ~new_new_n1190__;
  assign new_new_n1192__ = ~pi052 & ~new_new_n1191__;
  assign new_new_n1193__ = ~new_new_n332__ & po052;
  assign new_new_n1194__ = ~new_new_n1041__ & ~new_new_n1193__;
  assign new_new_n1195__ = pi065 & po052;
  assign new_new_n1196__ = po053 & ~new_new_n1195__;
  assign new_new_n1197__ = pi065 & ~new_new_n1041__;
  assign new_new_n1198__ = pi052 & ~new_new_n1197__;
  assign new_new_n1199__ = ~new_new_n1196__ & new_new_n1198__;
  assign new_new_n1200__ = ~new_new_n1192__ & ~new_new_n1194__;
  assign new_new_n1201__ = ~new_new_n1199__ & new_new_n1200__;
  assign new_new_n1202__ = ~pi053 & ~new_new_n1201__;
  assign new_new_n1203__ = ~pi064 & ~new_new_n1195__;
  assign new_new_n1204__ = ~pi065 & po052;
  assign new_new_n1205__ = ~po053 & ~new_new_n1204__;
  assign new_new_n1206__ = ~new_new_n1176__ & ~new_new_n1190__;
  assign new_new_n1207__ = ~new_new_n1205__ & new_new_n1206__;
  assign new_new_n1208__ = pi064 & ~new_new_n1207__;
  assign new_new_n1209__ = ~new_new_n1203__ & ~new_new_n1208__;
  assign new_new_n1210__ = ~new_new_n1041__ & ~new_new_n1195__;
  assign new_new_n1211__ = pi052 & ~new_new_n1053__;
  assign new_new_n1212__ = ~new_new_n1210__ & new_new_n1211__;
  assign new_new_n1213__ = ~new_new_n1209__ & ~new_new_n1212__;
  assign new_new_n1214__ = pi053 & ~new_new_n1213__;
  assign new_new_n1215__ = ~new_new_n1202__ & ~new_new_n1214__;
  assign new_new_n1216__ = ~pi066 & new_new_n1187__;
  assign new_new_n1217__ = ~new_new_n1215__ & ~new_new_n1216__;
  assign new_new_n1218__ = ~new_new_n1188__ & ~new_new_n1217__;
  assign new_new_n1219__ = ~new_new_n1175__ & ~new_new_n1218__;
  assign new_new_n1220__ = ~new_new_n1174__ & ~new_new_n1219__;
  assign new_new_n1221__ = ~pi068 & new_new_n1220__;
  assign new_new_n1222__ = pi068 & ~new_new_n1220__;
  assign new_new_n1223__ = ~new_new_n1075__ & po052;
  assign new_new_n1224__ = pi067 & ~po052;
  assign new_new_n1225__ = ~new_new_n1223__ & ~new_new_n1224__;
  assign new_new_n1226__ = ~new_new_n1031__ & ~new_new_n1032__;
  assign new_new_n1227__ = ~new_new_n1225__ & new_new_n1226__;
  assign new_new_n1228__ = new_new_n1225__ & ~new_new_n1226__;
  assign new_new_n1229__ = ~new_new_n1227__ & ~new_new_n1228__;
  assign new_new_n1230__ = ~new_new_n1222__ & ~new_new_n1229__;
  assign new_new_n1231__ = ~new_new_n1221__ & ~new_new_n1230__;
  assign new_new_n1232__ = ~new_new_n1168__ & ~new_new_n1231__;
  assign new_new_n1233__ = ~new_new_n1167__ & ~new_new_n1232__;
  assign new_new_n1234__ = ~new_new_n1161__ & ~new_new_n1233__;
  assign new_new_n1235__ = ~new_new_n1160__ & ~new_new_n1234__;
  assign new_new_n1236__ = ~new_new_n1152__ & ~new_new_n1235__;
  assign new_new_n1237__ = ~new_new_n1151__ & ~new_new_n1236__;
  assign new_new_n1238__ = ~new_new_n1129__ & ~new_new_n1132__;
  assign new_new_n1239__ = ~pi076 & new_new_n1238__;
  assign new_new_n1240__ = new_new_n1123__ & po052;
  assign new_new_n1241__ = pi073 & ~po052;
  assign new_new_n1242__ = ~new_new_n1240__ & ~new_new_n1241__;
  assign new_new_n1243__ = ~new_new_n1109__ & ~new_new_n1110__;
  assign new_new_n1244__ = ~new_new_n1242__ & ~new_new_n1243__;
  assign new_new_n1245__ = new_new_n1242__ & new_new_n1243__;
  assign new_new_n1246__ = ~new_new_n1244__ & ~new_new_n1245__;
  assign new_new_n1247__ = pi074 & ~new_new_n1246__;
  assign new_new_n1248__ = ~pi074 & new_new_n1246__;
  assign new_new_n1249__ = ~pi072 & ~new_new_n1121__;
  assign new_new_n1250__ = pi072 & new_new_n1121__;
  assign new_new_n1251__ = ~new_new_n1249__ & ~new_new_n1250__;
  assign new_new_n1252__ = po052 & new_new_n1251__;
  assign new_new_n1253__ = new_new_n1117__ & new_new_n1252__;
  assign new_new_n1254__ = ~new_new_n1117__ & ~new_new_n1252__;
  assign new_new_n1255__ = ~new_new_n1253__ & ~new_new_n1254__;
  assign new_new_n1256__ = ~pi073 & ~new_new_n1255__;
  assign new_new_n1257__ = pi073 & new_new_n1255__;
  assign new_new_n1258__ = ~new_new_n1142__ & ~new_new_n1237__;
  assign new_new_n1259__ = ~new_new_n1141__ & ~new_new_n1258__;
  assign new_new_n1260__ = ~new_new_n1257__ & ~new_new_n1259__;
  assign new_new_n1261__ = ~new_new_n1256__ & ~new_new_n1260__;
  assign new_new_n1262__ = ~new_new_n1248__ & new_new_n1261__;
  assign new_new_n1263__ = ~new_new_n1247__ & ~new_new_n1262__;
  assign new_new_n1264__ = pi075 & ~new_new_n1263__;
  assign new_new_n1265__ = pi076 & new_new_n1132__;
  assign new_new_n1266__ = ~new_new_n1264__ & ~new_new_n1265__;
  assign new_new_n1267__ = ~new_new_n1100__ & ~new_new_n1101__;
  assign new_new_n1268__ = ~new_new_n1125__ & po052;
  assign new_new_n1269__ = pi074 & ~po052;
  assign new_new_n1270__ = ~new_new_n1268__ & ~new_new_n1269__;
  assign new_new_n1271__ = new_new_n1267__ & ~new_new_n1270__;
  assign new_new_n1272__ = ~new_new_n1267__ & new_new_n1270__;
  assign new_new_n1273__ = ~new_new_n1271__ & ~new_new_n1272__;
  assign new_new_n1274__ = ~pi075 & new_new_n1263__;
  assign new_new_n1275__ = new_new_n1273__ & ~new_new_n1274__;
  assign new_new_n1276__ = new_new_n1266__ & ~new_new_n1275__;
  assign new_new_n1277__ = ~new_new_n1239__ & ~new_new_n1276__;
  assign po051 = new_new_n306__ & ~new_new_n1277__;
  assign new_new_n1279__ = ~new_new_n1237__ & po051;
  assign new_new_n1280__ = ~pi072 & ~po051;
  assign new_new_n1281__ = ~new_new_n1279__ & ~new_new_n1280__;
  assign new_new_n1282__ = new_new_n1143__ & ~new_new_n1281__;
  assign new_new_n1283__ = ~new_new_n1143__ & new_new_n1281__;
  assign new_new_n1284__ = ~new_new_n1282__ & ~new_new_n1283__;
  assign new_new_n1285__ = new_new_n1238__ & ~po051;
  assign new_new_n1286__ = ~new_new_n376__ & ~new_new_n1285__;
  assign new_new_n1287__ = ~pi077 & ~new_new_n1286__;
  assign new_new_n1288__ = pi077 & new_new_n1286__;
  assign new_new_n1289__ = new_new_n1261__ & po051;
  assign new_new_n1290__ = pi074 & ~po051;
  assign new_new_n1291__ = ~new_new_n1289__ & ~new_new_n1290__;
  assign new_new_n1292__ = ~new_new_n1247__ & ~new_new_n1248__;
  assign new_new_n1293__ = ~new_new_n1291__ & ~new_new_n1292__;
  assign new_new_n1294__ = new_new_n1291__ & new_new_n1292__;
  assign new_new_n1295__ = ~new_new_n1293__ & ~new_new_n1294__;
  assign new_new_n1296__ = pi075 & ~new_new_n1295__;
  assign new_new_n1297__ = ~pi075 & new_new_n1295__;
  assign new_new_n1298__ = ~new_new_n1256__ & ~new_new_n1257__;
  assign new_new_n1299__ = ~new_new_n1259__ & po051;
  assign new_new_n1300__ = ~pi073 & ~po051;
  assign new_new_n1301__ = ~new_new_n1299__ & ~new_new_n1300__;
  assign new_new_n1302__ = new_new_n1298__ & ~new_new_n1301__;
  assign new_new_n1303__ = ~new_new_n1298__ & new_new_n1301__;
  assign new_new_n1304__ = ~new_new_n1302__ & ~new_new_n1303__;
  assign new_new_n1305__ = pi074 & ~new_new_n1304__;
  assign new_new_n1306__ = ~pi074 & new_new_n1304__;
  assign new_new_n1307__ = pi073 & ~new_new_n1284__;
  assign new_new_n1308__ = ~pi073 & new_new_n1284__;
  assign new_new_n1309__ = ~new_new_n1151__ & ~new_new_n1152__;
  assign new_new_n1310__ = ~new_new_n1235__ & po051;
  assign new_new_n1311__ = ~pi071 & ~po051;
  assign new_new_n1312__ = ~new_new_n1310__ & ~new_new_n1311__;
  assign new_new_n1313__ = new_new_n1309__ & ~new_new_n1312__;
  assign new_new_n1314__ = ~new_new_n1309__ & new_new_n1312__;
  assign new_new_n1315__ = ~new_new_n1313__ & ~new_new_n1314__;
  assign new_new_n1316__ = pi072 & ~new_new_n1315__;
  assign new_new_n1317__ = ~pi072 & new_new_n1315__;
  assign new_new_n1318__ = ~pi070 & ~new_new_n1233__;
  assign new_new_n1319__ = pi070 & new_new_n1233__;
  assign new_new_n1320__ = ~new_new_n1318__ & ~new_new_n1319__;
  assign new_new_n1321__ = po051 & new_new_n1320__;
  assign new_new_n1322__ = new_new_n1159__ & ~new_new_n1321__;
  assign new_new_n1323__ = ~new_new_n1159__ & new_new_n1321__;
  assign new_new_n1324__ = ~new_new_n1322__ & ~new_new_n1323__;
  assign new_new_n1325__ = pi071 & ~new_new_n1324__;
  assign new_new_n1326__ = ~pi071 & new_new_n1324__;
  assign new_new_n1327__ = ~new_new_n1167__ & ~new_new_n1168__;
  assign new_new_n1328__ = ~new_new_n1231__ & po051;
  assign new_new_n1329__ = ~pi069 & ~po051;
  assign new_new_n1330__ = ~new_new_n1328__ & ~new_new_n1329__;
  assign new_new_n1331__ = new_new_n1327__ & ~new_new_n1330__;
  assign new_new_n1332__ = ~new_new_n1327__ & new_new_n1330__;
  assign new_new_n1333__ = ~new_new_n1331__ & ~new_new_n1332__;
  assign new_new_n1334__ = pi070 & ~new_new_n1333__;
  assign new_new_n1335__ = ~pi070 & new_new_n1333__;
  assign new_new_n1336__ = ~new_new_n1221__ & ~new_new_n1222__;
  assign new_new_n1337__ = po051 & new_new_n1336__;
  assign new_new_n1338__ = new_new_n1229__ & new_new_n1337__;
  assign new_new_n1339__ = ~new_new_n1229__ & ~new_new_n1337__;
  assign new_new_n1340__ = ~new_new_n1338__ & ~new_new_n1339__;
  assign new_new_n1341__ = ~pi069 & ~new_new_n1340__;
  assign new_new_n1342__ = pi069 & new_new_n1340__;
  assign new_new_n1343__ = ~pi067 & ~new_new_n1218__;
  assign new_new_n1344__ = pi067 & new_new_n1218__;
  assign new_new_n1345__ = ~new_new_n1343__ & ~new_new_n1344__;
  assign new_new_n1346__ = po051 & ~new_new_n1345__;
  assign new_new_n1347__ = new_new_n1173__ & new_new_n1346__;
  assign new_new_n1348__ = ~new_new_n1173__ & ~new_new_n1346__;
  assign new_new_n1349__ = ~new_new_n1347__ & ~new_new_n1348__;
  assign new_new_n1350__ = pi068 & ~new_new_n1349__;
  assign new_new_n1351__ = ~pi068 & new_new_n1349__;
  assign new_new_n1352__ = ~new_new_n1188__ & po051;
  assign new_new_n1353__ = ~new_new_n1216__ & new_new_n1352__;
  assign new_new_n1354__ = new_new_n1215__ & ~new_new_n1353__;
  assign new_new_n1355__ = new_new_n1217__ & new_new_n1352__;
  assign new_new_n1356__ = ~new_new_n1354__ & ~new_new_n1355__;
  assign new_new_n1357__ = ~pi067 & ~new_new_n1356__;
  assign new_new_n1358__ = pi067 & new_new_n1356__;
  assign new_new_n1359__ = pi051 & po051;
  assign new_new_n1360__ = pi050 & ~pi065;
  assign new_new_n1361__ = new_new_n1359__ & ~new_new_n1360__;
  assign new_new_n1362__ = ~pi051 & ~po051;
  assign new_new_n1363__ = ~pi065 & ~new_new_n1362__;
  assign new_new_n1364__ = ~pi050 & ~new_new_n1363__;
  assign new_new_n1365__ = ~new_new_n1361__ & ~new_new_n1364__;
  assign new_new_n1366__ = pi064 & ~new_new_n1365__;
  assign new_new_n1367__ = pi064 & po051;
  assign new_new_n1368__ = ~pi051 & pi065;
  assign new_new_n1369__ = ~new_new_n1367__ & new_new_n1368__;
  assign new_new_n1370__ = ~new_new_n1366__ & ~new_new_n1369__;
  assign new_new_n1371__ = pi066 & ~new_new_n1370__;
  assign new_new_n1372__ = new_new_n426__ & ~po052;
  assign new_new_n1373__ = new_new_n1204__ & po051;
  assign new_new_n1374__ = ~new_new_n1372__ & ~new_new_n1373__;
  assign new_new_n1375__ = ~pi051 & ~new_new_n1374__;
  assign new_new_n1376__ = ~new_new_n332__ & po051;
  assign new_new_n1377__ = ~new_new_n1184__ & ~new_new_n1376__;
  assign new_new_n1378__ = pi065 & po051;
  assign new_new_n1379__ = po052 & ~new_new_n1378__;
  assign new_new_n1380__ = pi065 & ~new_new_n1184__;
  assign new_new_n1381__ = pi051 & ~new_new_n1380__;
  assign new_new_n1382__ = ~new_new_n1379__ & new_new_n1381__;
  assign new_new_n1383__ = ~new_new_n1375__ & ~new_new_n1377__;
  assign new_new_n1384__ = ~new_new_n1382__ & new_new_n1383__;
  assign new_new_n1385__ = ~pi052 & ~new_new_n1384__;
  assign new_new_n1386__ = ~new_new_n1184__ & ~new_new_n1378__;
  assign new_new_n1387__ = pi051 & ~new_new_n1195__;
  assign new_new_n1388__ = pi064 & ~new_new_n1387__;
  assign new_new_n1389__ = ~new_new_n1386__ & ~new_new_n1388__;
  assign new_new_n1390__ = ~pi065 & po051;
  assign new_new_n1391__ = ~po052 & ~new_new_n1390__;
  assign new_new_n1392__ = pi064 & ~new_new_n1359__;
  assign new_new_n1393__ = ~new_new_n1373__ & new_new_n1392__;
  assign new_new_n1394__ = ~new_new_n1391__ & new_new_n1393__;
  assign new_new_n1395__ = ~new_new_n1389__ & ~new_new_n1394__;
  assign new_new_n1396__ = pi052 & ~new_new_n1395__;
  assign new_new_n1397__ = ~new_new_n1385__ & ~new_new_n1396__;
  assign new_new_n1398__ = ~pi066 & new_new_n1370__;
  assign new_new_n1399__ = ~new_new_n1397__ & ~new_new_n1398__;
  assign new_new_n1400__ = ~new_new_n1371__ & ~new_new_n1399__;
  assign new_new_n1401__ = ~new_new_n1358__ & new_new_n1400__;
  assign new_new_n1402__ = ~new_new_n1357__ & ~new_new_n1401__;
  assign new_new_n1403__ = ~new_new_n1351__ & new_new_n1402__;
  assign new_new_n1404__ = ~new_new_n1350__ & ~new_new_n1403__;
  assign new_new_n1405__ = ~new_new_n1342__ & new_new_n1404__;
  assign new_new_n1406__ = ~new_new_n1341__ & ~new_new_n1405__;
  assign new_new_n1407__ = ~new_new_n1335__ & new_new_n1406__;
  assign new_new_n1408__ = ~new_new_n1334__ & ~new_new_n1407__;
  assign new_new_n1409__ = ~new_new_n1326__ & ~new_new_n1408__;
  assign new_new_n1410__ = ~new_new_n1325__ & ~new_new_n1409__;
  assign new_new_n1411__ = ~new_new_n1317__ & ~new_new_n1410__;
  assign new_new_n1412__ = ~new_new_n1316__ & ~new_new_n1411__;
  assign new_new_n1413__ = ~new_new_n1308__ & ~new_new_n1412__;
  assign new_new_n1414__ = ~new_new_n1307__ & ~new_new_n1413__;
  assign new_new_n1415__ = ~new_new_n1306__ & ~new_new_n1414__;
  assign new_new_n1416__ = ~new_new_n1305__ & ~new_new_n1415__;
  assign new_new_n1417__ = ~new_new_n1297__ & ~new_new_n1416__;
  assign new_new_n1418__ = ~new_new_n1296__ & ~new_new_n1417__;
  assign new_new_n1419__ = pi076 & ~new_new_n1418__;
  assign new_new_n1420__ = ~new_new_n1288__ & ~new_new_n1419__;
  assign new_new_n1421__ = new_new_n306__ & ~new_new_n1274__;
  assign new_new_n1422__ = new_new_n1266__ & new_new_n1421__;
  assign new_new_n1423__ = ~new_new_n1273__ & ~new_new_n1422__;
  assign new_new_n1424__ = new_new_n992__ & new_new_n1238__;
  assign new_new_n1425__ = ~new_new_n1264__ & new_new_n1424__;
  assign new_new_n1426__ = new_new_n1275__ & new_new_n1425__;
  assign new_new_n1427__ = ~new_new_n1423__ & ~new_new_n1426__;
  assign new_new_n1428__ = ~pi076 & new_new_n1418__;
  assign new_new_n1429__ = new_new_n1427__ & ~new_new_n1428__;
  assign new_new_n1430__ = new_new_n1420__ & ~new_new_n1429__;
  assign new_new_n1431__ = ~new_new_n1287__ & ~new_new_n1430__;
  assign po050 = new_new_n305__ & ~new_new_n1431__;
  assign new_new_n1433__ = ~pi073 & ~new_new_n1412__;
  assign new_new_n1434__ = pi073 & new_new_n1412__;
  assign new_new_n1435__ = ~new_new_n1433__ & ~new_new_n1434__;
  assign new_new_n1436__ = po050 & ~new_new_n1435__;
  assign new_new_n1437__ = new_new_n1284__ & new_new_n1436__;
  assign new_new_n1438__ = ~new_new_n1284__ & ~new_new_n1436__;
  assign new_new_n1439__ = ~new_new_n1437__ & ~new_new_n1438__;
  assign new_new_n1440__ = pi074 & ~new_new_n1439__;
  assign new_new_n1441__ = ~pi074 & new_new_n1439__;
  assign new_new_n1442__ = ~new_new_n1440__ & ~new_new_n1441__;
  assign new_new_n1443__ = ~pi080 & new_new_n302__;
  assign new_new_n1444__ = ~pi079 & new_new_n1443__;
  assign new_new_n1445__ = ~new_new_n376__ & po050;
  assign new_new_n1446__ = ~new_new_n1286__ & ~new_new_n1445__;
  assign new_new_n1447__ = ~pi078 & new_new_n1446__;
  assign new_new_n1448__ = new_new_n1444__ & new_new_n1447__;
  assign new_new_n1449__ = new_new_n305__ & ~new_new_n1428__;
  assign new_new_n1450__ = new_new_n1420__ & new_new_n1449__;
  assign new_new_n1451__ = ~new_new_n1427__ & ~new_new_n1450__;
  assign new_new_n1452__ = new_new_n305__ & new_new_n1287__;
  assign new_new_n1453__ = ~new_new_n1419__ & new_new_n1452__;
  assign new_new_n1454__ = new_new_n1429__ & new_new_n1453__;
  assign new_new_n1455__ = ~new_new_n1451__ & ~new_new_n1454__;
  assign new_new_n1456__ = ~new_new_n1416__ & po050;
  assign new_new_n1457__ = pi075 & ~po050;
  assign new_new_n1458__ = ~new_new_n1456__ & ~new_new_n1457__;
  assign new_new_n1459__ = ~new_new_n1296__ & ~new_new_n1297__;
  assign new_new_n1460__ = ~new_new_n1458__ & new_new_n1459__;
  assign new_new_n1461__ = new_new_n1458__ & ~new_new_n1459__;
  assign new_new_n1462__ = ~new_new_n1460__ & ~new_new_n1461__;
  assign new_new_n1463__ = pi076 & new_new_n1462__;
  assign new_new_n1464__ = ~pi076 & ~new_new_n1462__;
  assign new_new_n1465__ = pi074 & ~new_new_n1414__;
  assign new_new_n1466__ = ~pi074 & new_new_n1414__;
  assign new_new_n1467__ = ~new_new_n1465__ & ~new_new_n1466__;
  assign new_new_n1468__ = po050 & new_new_n1467__;
  assign new_new_n1469__ = new_new_n1304__ & new_new_n1468__;
  assign new_new_n1470__ = ~new_new_n1304__ & ~new_new_n1468__;
  assign new_new_n1471__ = ~new_new_n1469__ & ~new_new_n1470__;
  assign new_new_n1472__ = pi075 & ~new_new_n1471__;
  assign new_new_n1473__ = ~pi075 & new_new_n1471__;
  assign new_new_n1474__ = ~new_new_n1316__ & ~new_new_n1317__;
  assign new_new_n1475__ = pi072 & ~po050;
  assign new_new_n1476__ = ~new_new_n1410__ & po050;
  assign new_new_n1477__ = ~new_new_n1475__ & ~new_new_n1476__;
  assign new_new_n1478__ = new_new_n1474__ & new_new_n1477__;
  assign new_new_n1479__ = ~new_new_n1474__ & ~new_new_n1477__;
  assign new_new_n1480__ = ~new_new_n1478__ & ~new_new_n1479__;
  assign new_new_n1481__ = pi073 & ~new_new_n1480__;
  assign new_new_n1482__ = ~pi073 & new_new_n1480__;
  assign new_new_n1483__ = ~new_new_n1408__ & po050;
  assign new_new_n1484__ = pi071 & ~po050;
  assign new_new_n1485__ = ~new_new_n1483__ & ~new_new_n1484__;
  assign new_new_n1486__ = ~new_new_n1325__ & ~new_new_n1326__;
  assign new_new_n1487__ = ~new_new_n1485__ & new_new_n1486__;
  assign new_new_n1488__ = new_new_n1485__ & ~new_new_n1486__;
  assign new_new_n1489__ = ~new_new_n1487__ & ~new_new_n1488__;
  assign new_new_n1490__ = pi072 & new_new_n1489__;
  assign new_new_n1491__ = ~pi072 & ~new_new_n1489__;
  assign new_new_n1492__ = ~new_new_n1334__ & ~new_new_n1335__;
  assign new_new_n1493__ = ~new_new_n1406__ & po050;
  assign new_new_n1494__ = ~pi070 & ~po050;
  assign new_new_n1495__ = ~new_new_n1493__ & ~new_new_n1494__;
  assign new_new_n1496__ = new_new_n1492__ & ~new_new_n1495__;
  assign new_new_n1497__ = ~new_new_n1492__ & new_new_n1495__;
  assign new_new_n1498__ = ~new_new_n1496__ & ~new_new_n1497__;
  assign new_new_n1499__ = pi071 & ~new_new_n1498__;
  assign new_new_n1500__ = ~pi071 & new_new_n1498__;
  assign new_new_n1501__ = ~new_new_n1341__ & ~new_new_n1342__;
  assign new_new_n1502__ = new_new_n1404__ & po050;
  assign new_new_n1503__ = ~pi069 & ~po050;
  assign new_new_n1504__ = ~new_new_n1502__ & ~new_new_n1503__;
  assign new_new_n1505__ = ~new_new_n1501__ & ~new_new_n1504__;
  assign new_new_n1506__ = new_new_n1501__ & new_new_n1504__;
  assign new_new_n1507__ = ~new_new_n1505__ & ~new_new_n1506__;
  assign new_new_n1508__ = ~pi070 & ~new_new_n1507__;
  assign new_new_n1509__ = pi070 & new_new_n1507__;
  assign new_new_n1510__ = new_new_n1402__ & po050;
  assign new_new_n1511__ = pi068 & ~po050;
  assign new_new_n1512__ = ~new_new_n1510__ & ~new_new_n1511__;
  assign new_new_n1513__ = ~new_new_n1350__ & ~new_new_n1351__;
  assign new_new_n1514__ = ~new_new_n1512__ & ~new_new_n1513__;
  assign new_new_n1515__ = new_new_n1512__ & new_new_n1513__;
  assign new_new_n1516__ = ~new_new_n1514__ & ~new_new_n1515__;
  assign new_new_n1517__ = pi069 & ~new_new_n1516__;
  assign new_new_n1518__ = ~pi069 & new_new_n1516__;
  assign new_new_n1519__ = ~new_new_n1357__ & ~new_new_n1358__;
  assign new_new_n1520__ = ~new_new_n1400__ & po050;
  assign new_new_n1521__ = pi067 & ~po050;
  assign new_new_n1522__ = ~new_new_n1520__ & ~new_new_n1521__;
  assign new_new_n1523__ = new_new_n1519__ & ~new_new_n1522__;
  assign new_new_n1524__ = ~new_new_n1519__ & new_new_n1522__;
  assign new_new_n1525__ = ~new_new_n1523__ & ~new_new_n1524__;
  assign new_new_n1526__ = ~pi068 & ~new_new_n1525__;
  assign new_new_n1527__ = pi068 & new_new_n1525__;
  assign new_new_n1528__ = pi050 & po050;
  assign new_new_n1529__ = ~pi050 & ~po050;
  assign new_new_n1530__ = ~pi065 & ~new_new_n1528__;
  assign new_new_n1531__ = ~new_new_n1529__ & new_new_n1530__;
  assign new_new_n1532__ = ~pi049 & ~new_new_n1531__;
  assign new_new_n1533__ = pi065 & new_new_n1528__;
  assign new_new_n1534__ = ~new_new_n1532__ & ~new_new_n1533__;
  assign new_new_n1535__ = pi064 & ~new_new_n1534__;
  assign new_new_n1536__ = pi064 & po050;
  assign new_new_n1537__ = ~pi050 & pi065;
  assign new_new_n1538__ = ~new_new_n1536__ & new_new_n1537__;
  assign new_new_n1539__ = ~new_new_n1535__ & ~new_new_n1538__;
  assign new_new_n1540__ = pi066 & ~new_new_n1539__;
  assign new_new_n1541__ = ~pi066 & new_new_n1539__;
  assign new_new_n1542__ = new_new_n426__ & ~po051;
  assign new_new_n1543__ = new_new_n1390__ & po050;
  assign new_new_n1544__ = ~new_new_n1542__ & ~new_new_n1543__;
  assign new_new_n1545__ = ~pi050 & ~new_new_n1544__;
  assign new_new_n1546__ = ~new_new_n332__ & po050;
  assign new_new_n1547__ = ~new_new_n1367__ & ~new_new_n1546__;
  assign new_new_n1548__ = pi065 & po050;
  assign new_new_n1549__ = po051 & ~new_new_n1548__;
  assign new_new_n1550__ = pi065 & ~new_new_n1367__;
  assign new_new_n1551__ = pi050 & ~new_new_n1550__;
  assign new_new_n1552__ = ~new_new_n1549__ & new_new_n1551__;
  assign new_new_n1553__ = ~new_new_n1545__ & ~new_new_n1547__;
  assign new_new_n1554__ = ~new_new_n1552__ & new_new_n1553__;
  assign new_new_n1555__ = pi051 & ~new_new_n1554__;
  assign new_new_n1556__ = ~pi064 & ~new_new_n1548__;
  assign new_new_n1557__ = ~pi065 & po050;
  assign new_new_n1558__ = ~po051 & ~new_new_n1557__;
  assign new_new_n1559__ = ~new_new_n1528__ & ~new_new_n1543__;
  assign new_new_n1560__ = ~new_new_n1558__ & new_new_n1559__;
  assign new_new_n1561__ = pi064 & ~new_new_n1560__;
  assign new_new_n1562__ = ~new_new_n1556__ & ~new_new_n1561__;
  assign new_new_n1563__ = ~new_new_n1367__ & ~new_new_n1548__;
  assign new_new_n1564__ = pi050 & ~new_new_n1378__;
  assign new_new_n1565__ = ~new_new_n1563__ & new_new_n1564__;
  assign new_new_n1566__ = ~new_new_n1562__ & ~new_new_n1565__;
  assign new_new_n1567__ = ~pi051 & ~new_new_n1566__;
  assign new_new_n1568__ = ~new_new_n1555__ & ~new_new_n1567__;
  assign new_new_n1569__ = ~new_new_n1541__ & new_new_n1568__;
  assign new_new_n1570__ = ~new_new_n1540__ & ~new_new_n1569__;
  assign new_new_n1571__ = pi067 & ~new_new_n1570__;
  assign new_new_n1572__ = ~new_new_n1371__ & po050;
  assign new_new_n1573__ = ~new_new_n1398__ & new_new_n1572__;
  assign new_new_n1574__ = new_new_n1397__ & ~new_new_n1573__;
  assign new_new_n1575__ = new_new_n1399__ & new_new_n1572__;
  assign new_new_n1576__ = ~new_new_n1574__ & ~new_new_n1575__;
  assign new_new_n1577__ = ~new_new_n1571__ & ~new_new_n1576__;
  assign new_new_n1578__ = ~pi067 & new_new_n1570__;
  assign new_new_n1579__ = ~new_new_n1577__ & ~new_new_n1578__;
  assign new_new_n1580__ = ~new_new_n1527__ & ~new_new_n1579__;
  assign new_new_n1581__ = ~new_new_n1526__ & ~new_new_n1580__;
  assign new_new_n1582__ = ~new_new_n1518__ & new_new_n1581__;
  assign new_new_n1583__ = ~new_new_n1517__ & ~new_new_n1582__;
  assign new_new_n1584__ = ~new_new_n1509__ & new_new_n1583__;
  assign new_new_n1585__ = ~new_new_n1508__ & ~new_new_n1584__;
  assign new_new_n1586__ = ~new_new_n1500__ & new_new_n1585__;
  assign new_new_n1587__ = ~new_new_n1499__ & ~new_new_n1586__;
  assign new_new_n1588__ = ~new_new_n1491__ & ~new_new_n1587__;
  assign new_new_n1589__ = ~new_new_n1490__ & ~new_new_n1588__;
  assign new_new_n1590__ = ~new_new_n1482__ & ~new_new_n1589__;
  assign new_new_n1591__ = ~new_new_n1481__ & ~new_new_n1590__;
  assign new_new_n1592__ = ~new_new_n1441__ & ~new_new_n1591__;
  assign new_new_n1593__ = ~new_new_n1440__ & ~new_new_n1592__;
  assign new_new_n1594__ = ~new_new_n1473__ & ~new_new_n1593__;
  assign new_new_n1595__ = ~new_new_n1472__ & ~new_new_n1594__;
  assign new_new_n1596__ = ~new_new_n1464__ & ~new_new_n1595__;
  assign new_new_n1597__ = ~new_new_n1463__ & ~new_new_n1596__;
  assign new_new_n1598__ = ~pi077 & new_new_n1597__;
  assign new_new_n1599__ = new_new_n1455__ & ~new_new_n1598__;
  assign new_new_n1600__ = pi077 & ~new_new_n1597__;
  assign new_new_n1601__ = pi078 & ~new_new_n1446__;
  assign new_new_n1602__ = new_new_n1444__ & ~new_new_n1601__;
  assign new_new_n1603__ = ~new_new_n1447__ & new_new_n1602__;
  assign new_new_n1604__ = ~new_new_n1600__ & new_new_n1603__;
  assign new_new_n1605__ = ~new_new_n1599__ & new_new_n1604__;
  assign po049 = new_new_n1448__ | new_new_n1605__;
  assign new_new_n1607__ = ~pi074 & ~po049;
  assign new_new_n1608__ = new_new_n1591__ & po049;
  assign new_new_n1609__ = ~new_new_n1607__ & ~new_new_n1608__;
  assign new_new_n1610__ = new_new_n1442__ & ~new_new_n1609__;
  assign new_new_n1611__ = ~new_new_n1442__ & new_new_n1609__;
  assign new_new_n1612__ = ~new_new_n1610__ & ~new_new_n1611__;
  assign new_new_n1613__ = pi075 & ~new_new_n1612__;
  assign new_new_n1614__ = ~pi075 & new_new_n1612__;
  assign new_new_n1615__ = ~new_new_n1613__ & ~new_new_n1614__;
  assign new_new_n1616__ = ~new_new_n1481__ & ~new_new_n1482__;
  assign new_new_n1617__ = ~pi073 & ~po049;
  assign new_new_n1618__ = new_new_n1589__ & po049;
  assign new_new_n1619__ = ~new_new_n1617__ & ~new_new_n1618__;
  assign new_new_n1620__ = new_new_n1616__ & ~new_new_n1619__;
  assign new_new_n1621__ = ~new_new_n1616__ & new_new_n1619__;
  assign new_new_n1622__ = ~new_new_n1620__ & ~new_new_n1621__;
  assign new_new_n1623__ = pi074 & ~new_new_n1622__;
  assign new_new_n1624__ = ~pi074 & new_new_n1622__;
  assign new_new_n1625__ = ~new_new_n1490__ & ~new_new_n1491__;
  assign new_new_n1626__ = new_new_n1587__ & po049;
  assign new_new_n1627__ = ~pi072 & ~po049;
  assign new_new_n1628__ = ~new_new_n1626__ & ~new_new_n1627__;
  assign new_new_n1629__ = ~new_new_n1625__ & ~new_new_n1628__;
  assign new_new_n1630__ = new_new_n1625__ & new_new_n1628__;
  assign new_new_n1631__ = ~new_new_n1629__ & ~new_new_n1630__;
  assign new_new_n1632__ = ~pi073 & ~new_new_n1631__;
  assign new_new_n1633__ = pi073 & new_new_n1631__;
  assign new_new_n1634__ = ~new_new_n1499__ & ~new_new_n1500__;
  assign new_new_n1635__ = ~new_new_n1585__ & po049;
  assign new_new_n1636__ = ~pi071 & ~po049;
  assign new_new_n1637__ = ~new_new_n1635__ & ~new_new_n1636__;
  assign new_new_n1638__ = new_new_n1634__ & new_new_n1637__;
  assign new_new_n1639__ = ~new_new_n1634__ & ~new_new_n1637__;
  assign new_new_n1640__ = ~new_new_n1638__ & ~new_new_n1639__;
  assign new_new_n1641__ = ~pi072 & ~new_new_n1640__;
  assign new_new_n1642__ = pi072 & new_new_n1640__;
  assign new_new_n1643__ = new_new_n1583__ & po049;
  assign new_new_n1644__ = ~pi070 & ~po049;
  assign new_new_n1645__ = ~new_new_n1643__ & ~new_new_n1644__;
  assign new_new_n1646__ = ~new_new_n1508__ & ~new_new_n1509__;
  assign new_new_n1647__ = ~new_new_n1645__ & ~new_new_n1646__;
  assign new_new_n1648__ = new_new_n1645__ & new_new_n1646__;
  assign new_new_n1649__ = ~new_new_n1647__ & ~new_new_n1648__;
  assign new_new_n1650__ = ~pi071 & ~new_new_n1649__;
  assign new_new_n1651__ = pi071 & new_new_n1649__;
  assign new_new_n1652__ = ~new_new_n1517__ & ~new_new_n1518__;
  assign new_new_n1653__ = ~new_new_n1581__ & po049;
  assign new_new_n1654__ = ~pi069 & ~po049;
  assign new_new_n1655__ = ~new_new_n1653__ & ~new_new_n1654__;
  assign new_new_n1656__ = new_new_n1652__ & ~new_new_n1655__;
  assign new_new_n1657__ = ~new_new_n1652__ & new_new_n1655__;
  assign new_new_n1658__ = ~new_new_n1656__ & ~new_new_n1657__;
  assign new_new_n1659__ = pi070 & ~new_new_n1658__;
  assign new_new_n1660__ = ~pi070 & new_new_n1658__;
  assign new_new_n1661__ = ~new_new_n1571__ & ~new_new_n1578__;
  assign new_new_n1662__ = po049 & new_new_n1661__;
  assign new_new_n1663__ = new_new_n1576__ & ~new_new_n1662__;
  assign new_new_n1664__ = ~new_new_n1576__ & new_new_n1662__;
  assign new_new_n1665__ = ~new_new_n1663__ & ~new_new_n1664__;
  assign new_new_n1666__ = pi068 & ~new_new_n1665__;
  assign new_new_n1667__ = ~pi068 & new_new_n1665__;
  assign new_new_n1668__ = ~new_new_n1540__ & ~new_new_n1541__;
  assign new_new_n1669__ = po049 & new_new_n1668__;
  assign new_new_n1670__ = new_new_n1568__ & ~new_new_n1669__;
  assign new_new_n1671__ = ~new_new_n1568__ & new_new_n1669__;
  assign new_new_n1672__ = ~new_new_n1670__ & ~new_new_n1671__;
  assign new_new_n1673__ = pi067 & ~new_new_n1672__;
  assign new_new_n1674__ = ~pi067 & new_new_n1672__;
  assign new_new_n1675__ = pi049 & po049;
  assign new_new_n1676__ = pi048 & ~pi065;
  assign new_new_n1677__ = new_new_n1675__ & ~new_new_n1676__;
  assign new_new_n1678__ = ~pi049 & ~po049;
  assign new_new_n1679__ = ~pi065 & ~new_new_n1678__;
  assign new_new_n1680__ = ~pi048 & ~new_new_n1679__;
  assign new_new_n1681__ = ~new_new_n1677__ & ~new_new_n1680__;
  assign new_new_n1682__ = pi064 & ~new_new_n1681__;
  assign new_new_n1683__ = pi064 & po049;
  assign new_new_n1684__ = ~pi049 & pi065;
  assign new_new_n1685__ = ~new_new_n1683__ & new_new_n1684__;
  assign new_new_n1686__ = ~new_new_n1682__ & ~new_new_n1685__;
  assign new_new_n1687__ = pi066 & ~new_new_n1686__;
  assign new_new_n1688__ = pi065 & po049;
  assign new_new_n1689__ = ~new_new_n1536__ & ~new_new_n1688__;
  assign new_new_n1690__ = ~new_new_n1683__ & new_new_n1689__;
  assign new_new_n1691__ = new_new_n426__ & ~po050;
  assign new_new_n1692__ = new_new_n1557__ & po049;
  assign new_new_n1693__ = ~new_new_n1691__ & ~new_new_n1692__;
  assign new_new_n1694__ = ~pi049 & ~new_new_n1693__;
  assign new_new_n1695__ = po050 & ~new_new_n1688__;
  assign new_new_n1696__ = pi065 & ~new_new_n1536__;
  assign new_new_n1697__ = pi049 & ~new_new_n1696__;
  assign new_new_n1698__ = ~new_new_n1695__ & new_new_n1697__;
  assign new_new_n1699__ = ~new_new_n1690__ & ~new_new_n1694__;
  assign new_new_n1700__ = ~new_new_n1698__ & new_new_n1699__;
  assign new_new_n1701__ = ~pi050 & ~new_new_n1700__;
  assign new_new_n1702__ = pi049 & ~new_new_n1548__;
  assign new_new_n1703__ = pi064 & ~new_new_n1702__;
  assign new_new_n1704__ = ~new_new_n1689__ & ~new_new_n1703__;
  assign new_new_n1705__ = ~pi065 & po049;
  assign new_new_n1706__ = ~po050 & ~new_new_n1705__;
  assign new_new_n1707__ = pi064 & ~new_new_n1675__;
  assign new_new_n1708__ = ~new_new_n1692__ & new_new_n1707__;
  assign new_new_n1709__ = ~new_new_n1706__ & new_new_n1708__;
  assign new_new_n1710__ = ~new_new_n1704__ & ~new_new_n1709__;
  assign new_new_n1711__ = pi050 & ~new_new_n1710__;
  assign new_new_n1712__ = ~new_new_n1701__ & ~new_new_n1711__;
  assign new_new_n1713__ = ~pi066 & new_new_n1686__;
  assign new_new_n1714__ = ~new_new_n1712__ & ~new_new_n1713__;
  assign new_new_n1715__ = ~new_new_n1687__ & ~new_new_n1714__;
  assign new_new_n1716__ = ~new_new_n1674__ & ~new_new_n1715__;
  assign new_new_n1717__ = ~new_new_n1673__ & ~new_new_n1716__;
  assign new_new_n1718__ = ~new_new_n1667__ & ~new_new_n1717__;
  assign new_new_n1719__ = ~new_new_n1666__ & ~new_new_n1718__;
  assign new_new_n1720__ = pi069 & ~new_new_n1719__;
  assign new_new_n1721__ = ~pi069 & new_new_n1719__;
  assign new_new_n1722__ = ~pi068 & ~new_new_n1579__;
  assign new_new_n1723__ = pi068 & new_new_n1579__;
  assign new_new_n1724__ = ~new_new_n1722__ & ~new_new_n1723__;
  assign new_new_n1725__ = po049 & new_new_n1724__;
  assign new_new_n1726__ = ~new_new_n1525__ & ~new_new_n1725__;
  assign new_new_n1727__ = new_new_n1525__ & new_new_n1725__;
  assign new_new_n1728__ = ~new_new_n1726__ & ~new_new_n1727__;
  assign new_new_n1729__ = ~new_new_n1721__ & new_new_n1728__;
  assign new_new_n1730__ = ~new_new_n1720__ & ~new_new_n1729__;
  assign new_new_n1731__ = ~new_new_n1660__ & ~new_new_n1730__;
  assign new_new_n1732__ = ~new_new_n1659__ & ~new_new_n1731__;
  assign new_new_n1733__ = ~new_new_n1651__ & new_new_n1732__;
  assign new_new_n1734__ = ~new_new_n1650__ & ~new_new_n1733__;
  assign new_new_n1735__ = ~new_new_n1642__ & ~new_new_n1734__;
  assign new_new_n1736__ = ~new_new_n1641__ & ~new_new_n1735__;
  assign new_new_n1737__ = ~new_new_n1633__ & ~new_new_n1736__;
  assign new_new_n1738__ = ~new_new_n1632__ & ~new_new_n1737__;
  assign new_new_n1739__ = ~new_new_n1624__ & new_new_n1738__;
  assign new_new_n1740__ = ~new_new_n1623__ & ~new_new_n1739__;
  assign new_new_n1741__ = ~new_new_n1598__ & ~new_new_n1600__;
  assign new_new_n1742__ = new_new_n1602__ & new_new_n1741__;
  assign new_new_n1743__ = ~new_new_n1455__ & ~new_new_n1742__;
  assign new_new_n1744__ = new_new_n1448__ & new_new_n1455__;
  assign new_new_n1745__ = new_new_n1741__ & new_new_n1744__;
  assign new_new_n1746__ = ~new_new_n1743__ & ~new_new_n1745__;
  assign new_new_n1747__ = pi078 & new_new_n1746__;
  assign new_new_n1748__ = ~pi078 & ~new_new_n1746__;
  assign new_new_n1749__ = ~new_new_n1463__ & ~new_new_n1464__;
  assign new_new_n1750__ = new_new_n1595__ & po049;
  assign new_new_n1751__ = ~pi076 & ~po049;
  assign new_new_n1752__ = ~new_new_n1750__ & ~new_new_n1751__;
  assign new_new_n1753__ = ~new_new_n1749__ & ~new_new_n1752__;
  assign new_new_n1754__ = new_new_n1749__ & new_new_n1752__;
  assign new_new_n1755__ = ~new_new_n1753__ & ~new_new_n1754__;
  assign new_new_n1756__ = pi077 & new_new_n1755__;
  assign new_new_n1757__ = ~pi077 & ~new_new_n1755__;
  assign new_new_n1758__ = pi075 & ~new_new_n1593__;
  assign new_new_n1759__ = ~pi075 & new_new_n1593__;
  assign new_new_n1760__ = ~new_new_n1758__ & ~new_new_n1759__;
  assign new_new_n1761__ = po049 & new_new_n1760__;
  assign new_new_n1762__ = new_new_n1471__ & new_new_n1761__;
  assign new_new_n1763__ = ~new_new_n1471__ & ~new_new_n1761__;
  assign new_new_n1764__ = ~new_new_n1762__ & ~new_new_n1763__;
  assign new_new_n1765__ = pi076 & ~new_new_n1764__;
  assign new_new_n1766__ = ~pi076 & new_new_n1764__;
  assign new_new_n1767__ = ~new_new_n1614__ & ~new_new_n1740__;
  assign new_new_n1768__ = ~new_new_n1613__ & ~new_new_n1767__;
  assign new_new_n1769__ = ~new_new_n1766__ & ~new_new_n1768__;
  assign new_new_n1770__ = ~new_new_n1765__ & ~new_new_n1769__;
  assign new_new_n1771__ = ~new_new_n1757__ & ~new_new_n1770__;
  assign new_new_n1772__ = ~new_new_n1756__ & ~new_new_n1771__;
  assign new_new_n1773__ = ~new_new_n1748__ & ~new_new_n1772__;
  assign new_new_n1774__ = ~new_new_n1747__ & ~new_new_n1773__;
  assign new_new_n1775__ = pi079 & ~new_new_n1774__;
  assign new_new_n1776__ = new_new_n1443__ & ~new_new_n1775__;
  assign new_new_n1777__ = new_new_n1446__ & ~po049;
  assign new_new_n1778__ = ~pi079 & new_new_n1774__;
  assign new_new_n1779__ = ~new_new_n376__ & ~new_new_n1777__;
  assign new_new_n1780__ = ~new_new_n1778__ & new_new_n1779__;
  assign po048 = new_new_n1776__ & ~new_new_n1780__;
  assign new_new_n1782__ = ~new_new_n1740__ & po048;
  assign new_new_n1783__ = pi075 & ~po048;
  assign new_new_n1784__ = ~new_new_n1782__ & ~new_new_n1783__;
  assign new_new_n1785__ = new_new_n1615__ & new_new_n1784__;
  assign new_new_n1786__ = ~new_new_n1615__ & ~new_new_n1784__;
  assign new_new_n1787__ = ~new_new_n1785__ & ~new_new_n1786__;
  assign new_new_n1788__ = pi076 & ~new_new_n1787__;
  assign new_new_n1789__ = ~pi076 & new_new_n1787__;
  assign new_new_n1790__ = ~new_new_n1788__ & ~new_new_n1789__;
  assign new_new_n1791__ = ~new_new_n1776__ & new_new_n1777__;
  assign new_new_n1792__ = ~new_new_n376__ & ~new_new_n1791__;
  assign new_new_n1793__ = ~pi080 & ~new_new_n1792__;
  assign new_new_n1794__ = pi080 & new_new_n1792__;
  assign new_new_n1795__ = ~new_new_n1770__ & po048;
  assign new_new_n1796__ = pi077 & ~po048;
  assign new_new_n1797__ = ~new_new_n1795__ & ~new_new_n1796__;
  assign new_new_n1798__ = ~new_new_n1756__ & ~new_new_n1757__;
  assign new_new_n1799__ = ~new_new_n1797__ & new_new_n1798__;
  assign new_new_n1800__ = new_new_n1797__ & ~new_new_n1798__;
  assign new_new_n1801__ = ~new_new_n1799__ & ~new_new_n1800__;
  assign new_new_n1802__ = ~pi078 & ~new_new_n1801__;
  assign new_new_n1803__ = pi078 & new_new_n1801__;
  assign new_new_n1804__ = ~new_new_n1765__ & ~new_new_n1766__;
  assign new_new_n1805__ = pi076 & ~po048;
  assign new_new_n1806__ = ~new_new_n1768__ & po048;
  assign new_new_n1807__ = ~new_new_n1805__ & ~new_new_n1806__;
  assign new_new_n1808__ = new_new_n1804__ & new_new_n1807__;
  assign new_new_n1809__ = ~new_new_n1804__ & ~new_new_n1807__;
  assign new_new_n1810__ = ~new_new_n1808__ & ~new_new_n1809__;
  assign new_new_n1811__ = pi077 & ~new_new_n1810__;
  assign new_new_n1812__ = ~pi077 & new_new_n1810__;
  assign new_new_n1813__ = new_new_n1738__ & po048;
  assign new_new_n1814__ = pi074 & ~po048;
  assign new_new_n1815__ = ~new_new_n1813__ & ~new_new_n1814__;
  assign new_new_n1816__ = ~new_new_n1623__ & ~new_new_n1624__;
  assign new_new_n1817__ = ~new_new_n1815__ & ~new_new_n1816__;
  assign new_new_n1818__ = new_new_n1815__ & new_new_n1816__;
  assign new_new_n1819__ = ~new_new_n1817__ & ~new_new_n1818__;
  assign new_new_n1820__ = pi075 & ~new_new_n1819__;
  assign new_new_n1821__ = ~pi075 & new_new_n1819__;
  assign new_new_n1822__ = ~pi073 & ~new_new_n1736__;
  assign new_new_n1823__ = pi073 & new_new_n1736__;
  assign new_new_n1824__ = ~new_new_n1822__ & ~new_new_n1823__;
  assign new_new_n1825__ = po048 & new_new_n1824__;
  assign new_new_n1826__ = new_new_n1631__ & ~new_new_n1825__;
  assign new_new_n1827__ = ~new_new_n1631__ & new_new_n1825__;
  assign new_new_n1828__ = ~new_new_n1826__ & ~new_new_n1827__;
  assign new_new_n1829__ = pi074 & ~new_new_n1828__;
  assign new_new_n1830__ = ~pi074 & new_new_n1828__;
  assign new_new_n1831__ = ~new_new_n1641__ & ~new_new_n1642__;
  assign new_new_n1832__ = ~new_new_n1734__ & po048;
  assign new_new_n1833__ = ~pi072 & ~po048;
  assign new_new_n1834__ = ~new_new_n1832__ & ~new_new_n1833__;
  assign new_new_n1835__ = ~new_new_n1831__ & ~new_new_n1834__;
  assign new_new_n1836__ = new_new_n1831__ & new_new_n1834__;
  assign new_new_n1837__ = ~new_new_n1835__ & ~new_new_n1836__;
  assign new_new_n1838__ = ~pi073 & ~new_new_n1837__;
  assign new_new_n1839__ = pi073 & new_new_n1837__;
  assign new_new_n1840__ = new_new_n1732__ & po048;
  assign new_new_n1841__ = ~pi071 & ~po048;
  assign new_new_n1842__ = ~new_new_n1840__ & ~new_new_n1841__;
  assign new_new_n1843__ = ~new_new_n1650__ & ~new_new_n1651__;
  assign new_new_n1844__ = ~new_new_n1842__ & ~new_new_n1843__;
  assign new_new_n1845__ = new_new_n1842__ & new_new_n1843__;
  assign new_new_n1846__ = ~new_new_n1844__ & ~new_new_n1845__;
  assign new_new_n1847__ = ~pi072 & ~new_new_n1846__;
  assign new_new_n1848__ = pi072 & new_new_n1846__;
  assign new_new_n1849__ = pi070 & ~new_new_n1730__;
  assign new_new_n1850__ = ~pi070 & new_new_n1730__;
  assign new_new_n1851__ = ~new_new_n1849__ & ~new_new_n1850__;
  assign new_new_n1852__ = po048 & new_new_n1851__;
  assign new_new_n1853__ = new_new_n1658__ & new_new_n1852__;
  assign new_new_n1854__ = ~new_new_n1658__ & ~new_new_n1852__;
  assign new_new_n1855__ = ~new_new_n1853__ & ~new_new_n1854__;
  assign new_new_n1856__ = pi071 & ~new_new_n1855__;
  assign new_new_n1857__ = ~pi071 & new_new_n1855__;
  assign new_new_n1858__ = pi068 & ~new_new_n1717__;
  assign new_new_n1859__ = ~pi068 & new_new_n1717__;
  assign new_new_n1860__ = ~new_new_n1858__ & ~new_new_n1859__;
  assign new_new_n1861__ = po048 & new_new_n1860__;
  assign new_new_n1862__ = new_new_n1665__ & new_new_n1861__;
  assign new_new_n1863__ = ~new_new_n1665__ & ~new_new_n1861__;
  assign new_new_n1864__ = ~new_new_n1862__ & ~new_new_n1863__;
  assign new_new_n1865__ = pi069 & ~new_new_n1864__;
  assign new_new_n1866__ = ~pi069 & new_new_n1864__;
  assign new_new_n1867__ = ~new_new_n1687__ & ~new_new_n1713__;
  assign new_new_n1868__ = po048 & new_new_n1867__;
  assign new_new_n1869__ = new_new_n1712__ & ~new_new_n1868__;
  assign new_new_n1870__ = ~new_new_n1712__ & new_new_n1868__;
  assign new_new_n1871__ = ~new_new_n1869__ & ~new_new_n1870__;
  assign new_new_n1872__ = pi067 & new_new_n1871__;
  assign new_new_n1873__ = ~pi067 & ~new_new_n1871__;
  assign new_new_n1874__ = pi048 & po048;
  assign new_new_n1875__ = pi047 & ~pi065;
  assign new_new_n1876__ = new_new_n1874__ & ~new_new_n1875__;
  assign new_new_n1877__ = ~pi048 & ~po048;
  assign new_new_n1878__ = ~pi065 & ~new_new_n1877__;
  assign new_new_n1879__ = ~pi047 & ~new_new_n1878__;
  assign new_new_n1880__ = ~new_new_n1876__ & ~new_new_n1879__;
  assign new_new_n1881__ = pi064 & ~new_new_n1880__;
  assign new_new_n1882__ = pi064 & po048;
  assign new_new_n1883__ = ~pi048 & pi065;
  assign new_new_n1884__ = ~new_new_n1882__ & new_new_n1883__;
  assign new_new_n1885__ = ~new_new_n1881__ & ~new_new_n1884__;
  assign new_new_n1886__ = pi066 & ~new_new_n1885__;
  assign new_new_n1887__ = new_new_n426__ & ~po049;
  assign new_new_n1888__ = new_new_n1705__ & po048;
  assign new_new_n1889__ = ~new_new_n1887__ & ~new_new_n1888__;
  assign new_new_n1890__ = ~pi048 & ~new_new_n1889__;
  assign new_new_n1891__ = ~new_new_n332__ & po048;
  assign new_new_n1892__ = ~new_new_n1683__ & ~new_new_n1891__;
  assign new_new_n1893__ = pi065 & ~new_new_n1683__;
  assign new_new_n1894__ = pi065 & po048;
  assign new_new_n1895__ = po049 & ~new_new_n1894__;
  assign new_new_n1896__ = pi048 & ~new_new_n1893__;
  assign new_new_n1897__ = ~new_new_n1895__ & new_new_n1896__;
  assign new_new_n1898__ = ~new_new_n1890__ & ~new_new_n1892__;
  assign new_new_n1899__ = ~new_new_n1897__ & new_new_n1898__;
  assign new_new_n1900__ = ~pi049 & ~new_new_n1899__;
  assign new_new_n1901__ = ~new_new_n1683__ & ~new_new_n1894__;
  assign new_new_n1902__ = pi048 & ~new_new_n1688__;
  assign new_new_n1903__ = pi064 & ~new_new_n1902__;
  assign new_new_n1904__ = ~new_new_n1901__ & ~new_new_n1903__;
  assign new_new_n1905__ = ~pi065 & po048;
  assign new_new_n1906__ = ~po049 & ~new_new_n1905__;
  assign new_new_n1907__ = pi064 & ~new_new_n1874__;
  assign new_new_n1908__ = ~new_new_n1888__ & new_new_n1907__;
  assign new_new_n1909__ = ~new_new_n1906__ & new_new_n1908__;
  assign new_new_n1910__ = ~new_new_n1904__ & ~new_new_n1909__;
  assign new_new_n1911__ = pi049 & ~new_new_n1910__;
  assign new_new_n1912__ = ~new_new_n1900__ & ~new_new_n1911__;
  assign new_new_n1913__ = ~pi066 & new_new_n1885__;
  assign new_new_n1914__ = ~new_new_n1912__ & ~new_new_n1913__;
  assign new_new_n1915__ = ~new_new_n1886__ & ~new_new_n1914__;
  assign new_new_n1916__ = ~new_new_n1873__ & ~new_new_n1915__;
  assign new_new_n1917__ = ~new_new_n1872__ & ~new_new_n1916__;
  assign new_new_n1918__ = pi068 & ~new_new_n1917__;
  assign new_new_n1919__ = ~pi068 & new_new_n1917__;
  assign new_new_n1920__ = ~pi067 & ~new_new_n1715__;
  assign new_new_n1921__ = pi067 & new_new_n1715__;
  assign new_new_n1922__ = ~new_new_n1920__ & ~new_new_n1921__;
  assign new_new_n1923__ = po048 & ~new_new_n1922__;
  assign new_new_n1924__ = new_new_n1672__ & new_new_n1923__;
  assign new_new_n1925__ = ~new_new_n1672__ & ~new_new_n1923__;
  assign new_new_n1926__ = ~new_new_n1924__ & ~new_new_n1925__;
  assign new_new_n1927__ = ~new_new_n1919__ & ~new_new_n1926__;
  assign new_new_n1928__ = ~new_new_n1918__ & ~new_new_n1927__;
  assign new_new_n1929__ = ~new_new_n1866__ & ~new_new_n1928__;
  assign new_new_n1930__ = ~new_new_n1865__ & ~new_new_n1929__;
  assign new_new_n1931__ = pi070 & ~new_new_n1930__;
  assign new_new_n1932__ = ~pi070 & new_new_n1930__;
  assign new_new_n1933__ = ~new_new_n1720__ & ~new_new_n1721__;
  assign new_new_n1934__ = po048 & new_new_n1933__;
  assign new_new_n1935__ = new_new_n1728__ & new_new_n1934__;
  assign new_new_n1936__ = ~new_new_n1728__ & ~new_new_n1934__;
  assign new_new_n1937__ = ~new_new_n1935__ & ~new_new_n1936__;
  assign new_new_n1938__ = ~new_new_n1932__ & new_new_n1937__;
  assign new_new_n1939__ = ~new_new_n1931__ & ~new_new_n1938__;
  assign new_new_n1940__ = ~new_new_n1857__ & ~new_new_n1939__;
  assign new_new_n1941__ = ~new_new_n1856__ & ~new_new_n1940__;
  assign new_new_n1942__ = ~new_new_n1848__ & new_new_n1941__;
  assign new_new_n1943__ = ~new_new_n1847__ & ~new_new_n1942__;
  assign new_new_n1944__ = ~new_new_n1839__ & ~new_new_n1943__;
  assign new_new_n1945__ = ~new_new_n1838__ & ~new_new_n1944__;
  assign new_new_n1946__ = ~new_new_n1830__ & new_new_n1945__;
  assign new_new_n1947__ = ~new_new_n1829__ & ~new_new_n1946__;
  assign new_new_n1948__ = ~new_new_n1821__ & ~new_new_n1947__;
  assign new_new_n1949__ = ~new_new_n1820__ & ~new_new_n1948__;
  assign new_new_n1950__ = ~new_new_n1789__ & ~new_new_n1949__;
  assign new_new_n1951__ = ~new_new_n1788__ & ~new_new_n1950__;
  assign new_new_n1952__ = ~new_new_n1812__ & ~new_new_n1951__;
  assign new_new_n1953__ = ~new_new_n1811__ & ~new_new_n1952__;
  assign new_new_n1954__ = ~new_new_n1803__ & new_new_n1953__;
  assign new_new_n1955__ = ~new_new_n1802__ & ~new_new_n1954__;
  assign new_new_n1956__ = pi079 & new_new_n1955__;
  assign new_new_n1957__ = ~new_new_n1794__ & ~new_new_n1956__;
  assign new_new_n1958__ = ~new_new_n1747__ & ~new_new_n1748__;
  assign new_new_n1959__ = ~new_new_n1772__ & po048;
  assign new_new_n1960__ = pi078 & ~po048;
  assign new_new_n1961__ = ~new_new_n1959__ & ~new_new_n1960__;
  assign new_new_n1962__ = new_new_n1958__ & ~new_new_n1961__;
  assign new_new_n1963__ = ~new_new_n1958__ & new_new_n1961__;
  assign new_new_n1964__ = ~new_new_n1962__ & ~new_new_n1963__;
  assign new_new_n1965__ = ~pi079 & ~new_new_n1955__;
  assign new_new_n1966__ = new_new_n1964__ & ~new_new_n1965__;
  assign new_new_n1967__ = new_new_n1957__ & ~new_new_n1966__;
  assign new_new_n1968__ = ~new_new_n1793__ & ~new_new_n1967__;
  assign po047 = new_new_n302__ & ~new_new_n1968__;
  assign new_new_n1970__ = pi076 & ~po047;
  assign new_new_n1971__ = ~new_new_n1949__ & po047;
  assign new_new_n1972__ = ~new_new_n1970__ & ~new_new_n1971__;
  assign new_new_n1973__ = new_new_n1790__ & new_new_n1972__;
  assign new_new_n1974__ = ~new_new_n1790__ & ~new_new_n1972__;
  assign new_new_n1975__ = ~new_new_n1973__ & ~new_new_n1974__;
  assign new_new_n1976__ = pi077 & ~new_new_n1975__;
  assign new_new_n1977__ = ~pi077 & new_new_n1975__;
  assign new_new_n1978__ = ~new_new_n1976__ & ~new_new_n1977__;
  assign new_new_n1979__ = new_new_n302__ & ~new_new_n1965__;
  assign new_new_n1980__ = new_new_n1957__ & new_new_n1979__;
  assign new_new_n1981__ = ~new_new_n1964__ & ~new_new_n1980__;
  assign new_new_n1982__ = new_new_n1443__ & ~new_new_n1792__;
  assign new_new_n1983__ = ~new_new_n1956__ & new_new_n1982__;
  assign new_new_n1984__ = new_new_n1966__ & new_new_n1983__;
  assign new_new_n1985__ = ~new_new_n1981__ & ~new_new_n1984__;
  assign new_new_n1986__ = ~pi080 & ~new_new_n1985__;
  assign new_new_n1987__ = ~new_new_n1953__ & po047;
  assign new_new_n1988__ = pi078 & ~po047;
  assign new_new_n1989__ = ~new_new_n1987__ & ~new_new_n1988__;
  assign new_new_n1990__ = ~new_new_n1802__ & ~new_new_n1803__;
  assign new_new_n1991__ = ~new_new_n1989__ & new_new_n1990__;
  assign new_new_n1992__ = new_new_n1989__ & ~new_new_n1990__;
  assign new_new_n1993__ = ~new_new_n1991__ & ~new_new_n1992__;
  assign new_new_n1994__ = ~pi079 & ~new_new_n1993__;
  assign new_new_n1995__ = pi079 & new_new_n1993__;
  assign new_new_n1996__ = ~new_new_n1811__ & ~new_new_n1812__;
  assign new_new_n1997__ = ~new_new_n1951__ & po047;
  assign new_new_n1998__ = pi077 & ~po047;
  assign new_new_n1999__ = ~new_new_n1997__ & ~new_new_n1998__;
  assign new_new_n2000__ = new_new_n1996__ & ~new_new_n1999__;
  assign new_new_n2001__ = ~new_new_n1996__ & new_new_n1999__;
  assign new_new_n2002__ = ~new_new_n2000__ & ~new_new_n2001__;
  assign new_new_n2003__ = pi078 & new_new_n2002__;
  assign new_new_n2004__ = ~pi078 & ~new_new_n2002__;
  assign new_new_n2005__ = ~new_new_n1820__ & ~new_new_n1821__;
  assign new_new_n2006__ = ~new_new_n1947__ & po047;
  assign new_new_n2007__ = pi075 & ~po047;
  assign new_new_n2008__ = ~new_new_n2006__ & ~new_new_n2007__;
  assign new_new_n2009__ = new_new_n2005__ & new_new_n2008__;
  assign new_new_n2010__ = ~new_new_n2005__ & ~new_new_n2008__;
  assign new_new_n2011__ = ~new_new_n2009__ & ~new_new_n2010__;
  assign new_new_n2012__ = ~pi076 & new_new_n2011__;
  assign new_new_n2013__ = pi076 & ~new_new_n2011__;
  assign new_new_n2014__ = new_new_n1945__ & po047;
  assign new_new_n2015__ = pi074 & ~po047;
  assign new_new_n2016__ = ~new_new_n2014__ & ~new_new_n2015__;
  assign new_new_n2017__ = ~new_new_n1829__ & ~new_new_n1830__;
  assign new_new_n2018__ = ~new_new_n2016__ & ~new_new_n2017__;
  assign new_new_n2019__ = new_new_n2016__ & new_new_n2017__;
  assign new_new_n2020__ = ~new_new_n2018__ & ~new_new_n2019__;
  assign new_new_n2021__ = ~pi075 & new_new_n2020__;
  assign new_new_n2022__ = pi075 & ~new_new_n2020__;
  assign new_new_n2023__ = ~new_new_n1838__ & ~new_new_n1839__;
  assign new_new_n2024__ = ~new_new_n1943__ & po047;
  assign new_new_n2025__ = ~pi073 & ~po047;
  assign new_new_n2026__ = ~new_new_n2024__ & ~new_new_n2025__;
  assign new_new_n2027__ = ~new_new_n2023__ & ~new_new_n2026__;
  assign new_new_n2028__ = new_new_n2023__ & new_new_n2026__;
  assign new_new_n2029__ = ~new_new_n2027__ & ~new_new_n2028__;
  assign new_new_n2030__ = ~pi074 & ~new_new_n2029__;
  assign new_new_n2031__ = pi074 & new_new_n2029__;
  assign new_new_n2032__ = new_new_n1941__ & po047;
  assign new_new_n2033__ = ~pi072 & ~po047;
  assign new_new_n2034__ = ~new_new_n2032__ & ~new_new_n2033__;
  assign new_new_n2035__ = ~new_new_n1847__ & ~new_new_n1848__;
  assign new_new_n2036__ = ~new_new_n2034__ & ~new_new_n2035__;
  assign new_new_n2037__ = new_new_n2034__ & new_new_n2035__;
  assign new_new_n2038__ = ~new_new_n2036__ & ~new_new_n2037__;
  assign new_new_n2039__ = ~pi073 & ~new_new_n2038__;
  assign new_new_n2040__ = pi073 & new_new_n2038__;
  assign new_new_n2041__ = ~new_new_n1856__ & ~new_new_n1857__;
  assign new_new_n2042__ = ~new_new_n1939__ & po047;
  assign new_new_n2043__ = pi071 & ~po047;
  assign new_new_n2044__ = ~new_new_n2042__ & ~new_new_n2043__;
  assign new_new_n2045__ = new_new_n2041__ & ~new_new_n2044__;
  assign new_new_n2046__ = ~new_new_n2041__ & new_new_n2044__;
  assign new_new_n2047__ = ~new_new_n2045__ & ~new_new_n2046__;
  assign new_new_n2048__ = ~pi072 & ~new_new_n2047__;
  assign new_new_n2049__ = pi072 & new_new_n2047__;
  assign new_new_n2050__ = ~new_new_n1931__ & ~new_new_n1932__;
  assign new_new_n2051__ = po047 & new_new_n2050__;
  assign new_new_n2052__ = ~new_new_n1937__ & ~new_new_n2051__;
  assign new_new_n2053__ = new_new_n1937__ & new_new_n2051__;
  assign new_new_n2054__ = ~new_new_n2052__ & ~new_new_n2053__;
  assign new_new_n2055__ = ~pi071 & ~new_new_n2054__;
  assign new_new_n2056__ = pi071 & new_new_n2054__;
  assign new_new_n2057__ = ~new_new_n1865__ & ~new_new_n1866__;
  assign new_new_n2058__ = ~new_new_n1928__ & po047;
  assign new_new_n2059__ = pi069 & ~po047;
  assign new_new_n2060__ = ~new_new_n2058__ & ~new_new_n2059__;
  assign new_new_n2061__ = new_new_n2057__ & new_new_n2060__;
  assign new_new_n2062__ = ~new_new_n2057__ & ~new_new_n2060__;
  assign new_new_n2063__ = ~new_new_n2061__ & ~new_new_n2062__;
  assign new_new_n2064__ = pi070 & ~new_new_n2063__;
  assign new_new_n2065__ = ~pi070 & new_new_n2063__;
  assign new_new_n2066__ = ~new_new_n1918__ & ~new_new_n1919__;
  assign new_new_n2067__ = po047 & new_new_n2066__;
  assign new_new_n2068__ = new_new_n1926__ & new_new_n2067__;
  assign new_new_n2069__ = ~new_new_n1926__ & ~new_new_n2067__;
  assign new_new_n2070__ = ~new_new_n2068__ & ~new_new_n2069__;
  assign new_new_n2071__ = pi069 & ~new_new_n2070__;
  assign new_new_n2072__ = ~pi069 & new_new_n2070__;
  assign new_new_n2073__ = ~new_new_n1886__ & ~new_new_n1913__;
  assign new_new_n2074__ = po047 & new_new_n2073__;
  assign new_new_n2075__ = new_new_n1912__ & ~new_new_n2074__;
  assign new_new_n2076__ = ~new_new_n1912__ & new_new_n2074__;
  assign new_new_n2077__ = ~new_new_n2075__ & ~new_new_n2076__;
  assign new_new_n2078__ = pi067 & new_new_n2077__;
  assign new_new_n2079__ = ~pi067 & ~new_new_n2077__;
  assign new_new_n2080__ = pi047 & po047;
  assign new_new_n2081__ = ~pi047 & ~po047;
  assign new_new_n2082__ = ~new_new_n2080__ & ~new_new_n2081__;
  assign new_new_n2083__ = ~pi046 & ~new_new_n2082__;
  assign new_new_n2084__ = ~pi046 & pi065;
  assign new_new_n2085__ = pi065 & new_new_n2080__;
  assign new_new_n2086__ = ~new_new_n2084__ & ~new_new_n2085__;
  assign new_new_n2087__ = ~new_new_n2083__ & new_new_n2086__;
  assign new_new_n2088__ = pi064 & ~new_new_n2087__;
  assign new_new_n2089__ = pi064 & po047;
  assign new_new_n2090__ = ~pi047 & pi065;
  assign new_new_n2091__ = ~new_new_n2089__ & new_new_n2090__;
  assign new_new_n2092__ = ~new_new_n2088__ & ~new_new_n2091__;
  assign new_new_n2093__ = pi066 & ~new_new_n2092__;
  assign new_new_n2094__ = new_new_n426__ & ~po048;
  assign new_new_n2095__ = new_new_n1905__ & po047;
  assign new_new_n2096__ = ~new_new_n2094__ & ~new_new_n2095__;
  assign new_new_n2097__ = ~pi047 & ~new_new_n2096__;
  assign new_new_n2098__ = ~new_new_n332__ & po047;
  assign new_new_n2099__ = ~new_new_n1882__ & ~new_new_n2098__;
  assign new_new_n2100__ = pi065 & po047;
  assign new_new_n2101__ = po048 & ~new_new_n2100__;
  assign new_new_n2102__ = pi065 & ~new_new_n1882__;
  assign new_new_n2103__ = pi047 & ~new_new_n2102__;
  assign new_new_n2104__ = ~new_new_n2101__ & new_new_n2103__;
  assign new_new_n2105__ = ~new_new_n2097__ & ~new_new_n2099__;
  assign new_new_n2106__ = ~new_new_n2104__ & new_new_n2105__;
  assign new_new_n2107__ = ~pi048 & ~new_new_n2106__;
  assign new_new_n2108__ = ~new_new_n1882__ & ~new_new_n2100__;
  assign new_new_n2109__ = pi047 & ~new_new_n1894__;
  assign new_new_n2110__ = pi064 & ~new_new_n2109__;
  assign new_new_n2111__ = ~new_new_n2108__ & ~new_new_n2110__;
  assign new_new_n2112__ = ~pi065 & po047;
  assign new_new_n2113__ = ~po048 & ~new_new_n2112__;
  assign new_new_n2114__ = pi064 & ~new_new_n2080__;
  assign new_new_n2115__ = ~new_new_n2095__ & new_new_n2114__;
  assign new_new_n2116__ = ~new_new_n2113__ & new_new_n2115__;
  assign new_new_n2117__ = ~new_new_n2111__ & ~new_new_n2116__;
  assign new_new_n2118__ = pi048 & ~new_new_n2117__;
  assign new_new_n2119__ = ~new_new_n2107__ & ~new_new_n2118__;
  assign new_new_n2120__ = ~pi066 & new_new_n2092__;
  assign new_new_n2121__ = ~new_new_n2119__ & ~new_new_n2120__;
  assign new_new_n2122__ = ~new_new_n2093__ & ~new_new_n2121__;
  assign new_new_n2123__ = ~new_new_n2079__ & ~new_new_n2122__;
  assign new_new_n2124__ = ~new_new_n2078__ & ~new_new_n2123__;
  assign new_new_n2125__ = pi068 & ~new_new_n2124__;
  assign new_new_n2126__ = ~pi068 & new_new_n2124__;
  assign new_new_n2127__ = ~new_new_n1872__ & ~new_new_n1873__;
  assign new_new_n2128__ = new_new_n1915__ & po047;
  assign new_new_n2129__ = ~pi067 & ~po047;
  assign new_new_n2130__ = ~new_new_n2128__ & ~new_new_n2129__;
  assign new_new_n2131__ = ~new_new_n2127__ & ~new_new_n2130__;
  assign new_new_n2132__ = new_new_n2127__ & new_new_n2130__;
  assign new_new_n2133__ = ~new_new_n2131__ & ~new_new_n2132__;
  assign new_new_n2134__ = ~new_new_n2126__ & new_new_n2133__;
  assign new_new_n2135__ = ~new_new_n2125__ & ~new_new_n2134__;
  assign new_new_n2136__ = ~new_new_n2072__ & ~new_new_n2135__;
  assign new_new_n2137__ = ~new_new_n2071__ & ~new_new_n2136__;
  assign new_new_n2138__ = ~new_new_n2065__ & ~new_new_n2137__;
  assign new_new_n2139__ = ~new_new_n2064__ & ~new_new_n2138__;
  assign new_new_n2140__ = ~new_new_n2056__ & new_new_n2139__;
  assign new_new_n2141__ = ~new_new_n2055__ & ~new_new_n2140__;
  assign new_new_n2142__ = ~new_new_n2049__ & ~new_new_n2141__;
  assign new_new_n2143__ = ~new_new_n2048__ & ~new_new_n2142__;
  assign new_new_n2144__ = ~new_new_n2040__ & ~new_new_n2143__;
  assign new_new_n2145__ = ~new_new_n2039__ & ~new_new_n2144__;
  assign new_new_n2146__ = ~new_new_n2031__ & ~new_new_n2145__;
  assign new_new_n2147__ = ~new_new_n2030__ & ~new_new_n2146__;
  assign new_new_n2148__ = ~new_new_n2022__ & ~new_new_n2147__;
  assign new_new_n2149__ = ~new_new_n2021__ & ~new_new_n2148__;
  assign new_new_n2150__ = ~new_new_n2013__ & ~new_new_n2149__;
  assign new_new_n2151__ = ~new_new_n2012__ & ~new_new_n2150__;
  assign new_new_n2152__ = ~new_new_n1977__ & new_new_n2151__;
  assign new_new_n2153__ = ~new_new_n1976__ & ~new_new_n2152__;
  assign new_new_n2154__ = ~new_new_n2004__ & ~new_new_n2153__;
  assign new_new_n2155__ = ~new_new_n2003__ & ~new_new_n2154__;
  assign new_new_n2156__ = ~new_new_n1995__ & new_new_n2155__;
  assign new_new_n2157__ = ~new_new_n1994__ & ~new_new_n2156__;
  assign new_new_n2158__ = ~new_new_n1986__ & new_new_n2157__;
  assign new_new_n2159__ = ~pi085 & new_new_n297__;
  assign new_new_n2160__ = pi080 & new_new_n1985__;
  assign new_new_n2161__ = ~new_new_n376__ & po047;
  assign new_new_n2162__ = ~new_new_n1792__ & ~new_new_n2161__;
  assign new_new_n2163__ = ~pi081 & new_new_n2162__;
  assign new_new_n2164__ = pi081 & ~new_new_n2162__;
  assign new_new_n2165__ = ~pi082 & new_new_n298__;
  assign new_new_n2166__ = new_new_n2159__ & new_new_n2165__;
  assign new_new_n2167__ = ~new_new_n2160__ & new_new_n2166__;
  assign new_new_n2168__ = ~new_new_n2163__ & new_new_n2167__;
  assign new_new_n2169__ = ~new_new_n2164__ & new_new_n2168__;
  assign new_new_n2170__ = ~new_new_n2158__ & new_new_n2169__;
  assign new_new_n2171__ = new_new_n302__ & new_new_n2162__;
  assign po046 = new_new_n2170__ | new_new_n2171__;
  assign new_new_n2173__ = ~pi077 & ~po046;
  assign new_new_n2174__ = ~new_new_n2151__ & po046;
  assign new_new_n2175__ = ~new_new_n2173__ & ~new_new_n2174__;
  assign new_new_n2176__ = new_new_n1978__ & ~new_new_n2175__;
  assign new_new_n2177__ = ~new_new_n1978__ & new_new_n2175__;
  assign new_new_n2178__ = ~new_new_n2176__ & ~new_new_n2177__;
  assign new_new_n2179__ = new_new_n297__ & new_new_n299__;
  assign new_new_n2180__ = ~new_new_n302__ & ~new_new_n1792__;
  assign new_new_n2181__ = ~new_new_n2170__ & new_new_n2180__;
  assign new_new_n2182__ = ~new_new_n376__ & ~new_new_n2181__;
  assign new_new_n2183__ = ~pi082 & ~new_new_n2182__;
  assign new_new_n2184__ = pi082 & new_new_n2182__;
  assign new_new_n2185__ = ~new_new_n1994__ & ~new_new_n1995__;
  assign new_new_n2186__ = ~pi079 & ~po046;
  assign new_new_n2187__ = new_new_n2155__ & po046;
  assign new_new_n2188__ = ~new_new_n2186__ & ~new_new_n2187__;
  assign new_new_n2189__ = new_new_n2185__ & ~new_new_n2188__;
  assign new_new_n2190__ = ~new_new_n2185__ & new_new_n2188__;
  assign new_new_n2191__ = ~new_new_n2189__ & ~new_new_n2190__;
  assign new_new_n2192__ = pi080 & ~new_new_n2191__;
  assign new_new_n2193__ = ~pi080 & new_new_n2191__;
  assign new_new_n2194__ = ~new_new_n2003__ & ~new_new_n2004__;
  assign new_new_n2195__ = new_new_n2153__ & po046;
  assign new_new_n2196__ = ~pi078 & ~po046;
  assign new_new_n2197__ = ~new_new_n2195__ & ~new_new_n2196__;
  assign new_new_n2198__ = ~new_new_n2194__ & ~new_new_n2197__;
  assign new_new_n2199__ = new_new_n2194__ & new_new_n2197__;
  assign new_new_n2200__ = ~new_new_n2198__ & ~new_new_n2199__;
  assign new_new_n2201__ = ~pi079 & ~new_new_n2200__;
  assign new_new_n2202__ = pi079 & new_new_n2200__;
  assign new_new_n2203__ = pi078 & ~new_new_n2178__;
  assign new_new_n2204__ = ~pi078 & new_new_n2178__;
  assign new_new_n2205__ = ~new_new_n2012__ & ~new_new_n2013__;
  assign new_new_n2206__ = ~pi076 & ~po046;
  assign new_new_n2207__ = ~new_new_n2149__ & po046;
  assign new_new_n2208__ = ~new_new_n2206__ & ~new_new_n2207__;
  assign new_new_n2209__ = new_new_n2205__ & ~new_new_n2208__;
  assign new_new_n2210__ = ~new_new_n2205__ & new_new_n2208__;
  assign new_new_n2211__ = ~new_new_n2209__ & ~new_new_n2210__;
  assign new_new_n2212__ = pi077 & ~new_new_n2211__;
  assign new_new_n2213__ = ~pi077 & new_new_n2211__;
  assign new_new_n2214__ = ~new_new_n2021__ & ~new_new_n2022__;
  assign new_new_n2215__ = ~pi075 & ~po046;
  assign new_new_n2216__ = ~new_new_n2147__ & po046;
  assign new_new_n2217__ = ~new_new_n2215__ & ~new_new_n2216__;
  assign new_new_n2218__ = new_new_n2214__ & ~new_new_n2217__;
  assign new_new_n2219__ = ~new_new_n2214__ & new_new_n2217__;
  assign new_new_n2220__ = ~new_new_n2218__ & ~new_new_n2219__;
  assign new_new_n2221__ = ~pi076 & new_new_n2220__;
  assign new_new_n2222__ = pi076 & ~new_new_n2220__;
  assign new_new_n2223__ = ~pi074 & ~new_new_n2145__;
  assign new_new_n2224__ = pi074 & new_new_n2145__;
  assign new_new_n2225__ = ~new_new_n2223__ & ~new_new_n2224__;
  assign new_new_n2226__ = po046 & new_new_n2225__;
  assign new_new_n2227__ = new_new_n2029__ & ~new_new_n2226__;
  assign new_new_n2228__ = ~new_new_n2029__ & new_new_n2226__;
  assign new_new_n2229__ = ~new_new_n2227__ & ~new_new_n2228__;
  assign new_new_n2230__ = ~pi075 & new_new_n2229__;
  assign new_new_n2231__ = pi075 & ~new_new_n2229__;
  assign new_new_n2232__ = ~new_new_n2039__ & ~new_new_n2040__;
  assign new_new_n2233__ = ~pi073 & ~po046;
  assign new_new_n2234__ = ~new_new_n2143__ & po046;
  assign new_new_n2235__ = ~new_new_n2233__ & ~new_new_n2234__;
  assign new_new_n2236__ = new_new_n2232__ & ~new_new_n2235__;
  assign new_new_n2237__ = ~new_new_n2232__ & new_new_n2235__;
  assign new_new_n2238__ = ~new_new_n2236__ & ~new_new_n2237__;
  assign new_new_n2239__ = ~pi074 & new_new_n2238__;
  assign new_new_n2240__ = pi074 & ~new_new_n2238__;
  assign new_new_n2241__ = ~new_new_n2048__ & ~new_new_n2049__;
  assign new_new_n2242__ = ~new_new_n2141__ & po046;
  assign new_new_n2243__ = ~pi072 & ~po046;
  assign new_new_n2244__ = ~new_new_n2242__ & ~new_new_n2243__;
  assign new_new_n2245__ = ~new_new_n2241__ & ~new_new_n2244__;
  assign new_new_n2246__ = new_new_n2241__ & new_new_n2244__;
  assign new_new_n2247__ = ~new_new_n2245__ & ~new_new_n2246__;
  assign new_new_n2248__ = ~pi073 & ~new_new_n2247__;
  assign new_new_n2249__ = pi073 & new_new_n2247__;
  assign new_new_n2250__ = new_new_n2139__ & po046;
  assign new_new_n2251__ = ~pi071 & ~po046;
  assign new_new_n2252__ = ~new_new_n2250__ & ~new_new_n2251__;
  assign new_new_n2253__ = ~new_new_n2055__ & ~new_new_n2056__;
  assign new_new_n2254__ = ~new_new_n2252__ & ~new_new_n2253__;
  assign new_new_n2255__ = new_new_n2252__ & new_new_n2253__;
  assign new_new_n2256__ = ~new_new_n2254__ & ~new_new_n2255__;
  assign new_new_n2257__ = pi072 & new_new_n2256__;
  assign new_new_n2258__ = ~pi072 & ~new_new_n2256__;
  assign new_new_n2259__ = ~new_new_n2064__ & ~new_new_n2065__;
  assign new_new_n2260__ = ~pi070 & ~po046;
  assign new_new_n2261__ = new_new_n2137__ & po046;
  assign new_new_n2262__ = ~new_new_n2260__ & ~new_new_n2261__;
  assign new_new_n2263__ = new_new_n2259__ & ~new_new_n2262__;
  assign new_new_n2264__ = ~new_new_n2259__ & new_new_n2262__;
  assign new_new_n2265__ = ~new_new_n2263__ & ~new_new_n2264__;
  assign new_new_n2266__ = pi071 & ~new_new_n2265__;
  assign new_new_n2267__ = ~pi071 & new_new_n2265__;
  assign new_new_n2268__ = ~new_new_n2071__ & ~new_new_n2072__;
  assign new_new_n2269__ = new_new_n2135__ & po046;
  assign new_new_n2270__ = ~pi069 & ~po046;
  assign new_new_n2271__ = ~new_new_n2269__ & ~new_new_n2270__;
  assign new_new_n2272__ = new_new_n2268__ & new_new_n2271__;
  assign new_new_n2273__ = ~new_new_n2268__ & ~new_new_n2271__;
  assign new_new_n2274__ = ~new_new_n2272__ & ~new_new_n2273__;
  assign new_new_n2275__ = ~pi070 & ~new_new_n2274__;
  assign new_new_n2276__ = pi070 & new_new_n2274__;
  assign new_new_n2277__ = ~new_new_n2125__ & ~new_new_n2126__;
  assign new_new_n2278__ = po046 & new_new_n2277__;
  assign new_new_n2279__ = ~new_new_n2133__ & ~new_new_n2278__;
  assign new_new_n2280__ = new_new_n2133__ & new_new_n2278__;
  assign new_new_n2281__ = ~new_new_n2279__ & ~new_new_n2280__;
  assign new_new_n2282__ = ~pi069 & ~new_new_n2281__;
  assign new_new_n2283__ = pi069 & new_new_n2281__;
  assign new_new_n2284__ = ~new_new_n2078__ & ~new_new_n2079__;
  assign new_new_n2285__ = ~pi067 & ~po046;
  assign new_new_n2286__ = new_new_n2122__ & po046;
  assign new_new_n2287__ = ~new_new_n2285__ & ~new_new_n2286__;
  assign new_new_n2288__ = ~new_new_n2284__ & ~new_new_n2287__;
  assign new_new_n2289__ = new_new_n2284__ & new_new_n2287__;
  assign new_new_n2290__ = ~new_new_n2288__ & ~new_new_n2289__;
  assign new_new_n2291__ = ~pi068 & ~new_new_n2290__;
  assign new_new_n2292__ = pi068 & new_new_n2290__;
  assign new_new_n2293__ = ~new_new_n2093__ & po046;
  assign new_new_n2294__ = ~new_new_n2120__ & new_new_n2293__;
  assign new_new_n2295__ = new_new_n2119__ & ~new_new_n2294__;
  assign new_new_n2296__ = new_new_n2121__ & new_new_n2293__;
  assign new_new_n2297__ = ~new_new_n2295__ & ~new_new_n2296__;
  assign new_new_n2298__ = ~pi067 & ~new_new_n2297__;
  assign new_new_n2299__ = pi067 & new_new_n2297__;
  assign new_new_n2300__ = pi046 & po046;
  assign new_new_n2301__ = pi045 & ~pi065;
  assign new_new_n2302__ = new_new_n2300__ & ~new_new_n2301__;
  assign new_new_n2303__ = ~pi046 & ~po046;
  assign new_new_n2304__ = ~pi065 & ~new_new_n2303__;
  assign new_new_n2305__ = ~pi045 & ~new_new_n2304__;
  assign new_new_n2306__ = ~new_new_n2302__ & ~new_new_n2305__;
  assign new_new_n2307__ = pi064 & ~new_new_n2306__;
  assign new_new_n2308__ = pi064 & po046;
  assign new_new_n2309__ = new_new_n2084__ & ~new_new_n2308__;
  assign new_new_n2310__ = ~new_new_n2307__ & ~new_new_n2309__;
  assign new_new_n2311__ = pi066 & ~new_new_n2310__;
  assign new_new_n2312__ = ~pi066 & new_new_n2310__;
  assign new_new_n2313__ = pi065 & po046;
  assign new_new_n2314__ = ~new_new_n2089__ & ~new_new_n2313__;
  assign new_new_n2315__ = ~new_new_n2308__ & new_new_n2314__;
  assign new_new_n2316__ = new_new_n426__ & ~po047;
  assign new_new_n2317__ = new_new_n2112__ & po046;
  assign new_new_n2318__ = ~new_new_n2316__ & ~new_new_n2317__;
  assign new_new_n2319__ = ~pi046 & ~new_new_n2318__;
  assign new_new_n2320__ = po047 & ~new_new_n2313__;
  assign new_new_n2321__ = pi065 & ~new_new_n2089__;
  assign new_new_n2322__ = pi046 & ~new_new_n2321__;
  assign new_new_n2323__ = ~new_new_n2320__ & new_new_n2322__;
  assign new_new_n2324__ = ~new_new_n2315__ & ~new_new_n2319__;
  assign new_new_n2325__ = ~new_new_n2323__ & new_new_n2324__;
  assign new_new_n2326__ = pi047 & ~new_new_n2325__;
  assign new_new_n2327__ = pi046 & ~new_new_n2100__;
  assign new_new_n2328__ = pi064 & ~new_new_n2327__;
  assign new_new_n2329__ = ~new_new_n2314__ & ~new_new_n2328__;
  assign new_new_n2330__ = ~pi065 & po046;
  assign new_new_n2331__ = ~po047 & ~new_new_n2330__;
  assign new_new_n2332__ = pi064 & ~new_new_n2300__;
  assign new_new_n2333__ = ~new_new_n2317__ & new_new_n2332__;
  assign new_new_n2334__ = ~new_new_n2331__ & new_new_n2333__;
  assign new_new_n2335__ = ~new_new_n2329__ & ~new_new_n2334__;
  assign new_new_n2336__ = ~pi047 & ~new_new_n2335__;
  assign new_new_n2337__ = ~new_new_n2326__ & ~new_new_n2336__;
  assign new_new_n2338__ = ~new_new_n2312__ & new_new_n2337__;
  assign new_new_n2339__ = ~new_new_n2311__ & ~new_new_n2338__;
  assign new_new_n2340__ = ~new_new_n2299__ & new_new_n2339__;
  assign new_new_n2341__ = ~new_new_n2298__ & ~new_new_n2340__;
  assign new_new_n2342__ = ~new_new_n2292__ & ~new_new_n2341__;
  assign new_new_n2343__ = ~new_new_n2291__ & ~new_new_n2342__;
  assign new_new_n2344__ = ~new_new_n2283__ & ~new_new_n2343__;
  assign new_new_n2345__ = ~new_new_n2282__ & ~new_new_n2344__;
  assign new_new_n2346__ = ~new_new_n2276__ & ~new_new_n2345__;
  assign new_new_n2347__ = ~new_new_n2275__ & ~new_new_n2346__;
  assign new_new_n2348__ = ~new_new_n2267__ & new_new_n2347__;
  assign new_new_n2349__ = ~new_new_n2266__ & ~new_new_n2348__;
  assign new_new_n2350__ = ~new_new_n2258__ & ~new_new_n2349__;
  assign new_new_n2351__ = ~new_new_n2257__ & ~new_new_n2350__;
  assign new_new_n2352__ = ~new_new_n2249__ & new_new_n2351__;
  assign new_new_n2353__ = ~new_new_n2248__ & ~new_new_n2352__;
  assign new_new_n2354__ = ~new_new_n2240__ & ~new_new_n2353__;
  assign new_new_n2355__ = ~new_new_n2239__ & ~new_new_n2354__;
  assign new_new_n2356__ = ~new_new_n2231__ & ~new_new_n2355__;
  assign new_new_n2357__ = ~new_new_n2230__ & ~new_new_n2356__;
  assign new_new_n2358__ = ~new_new_n2222__ & ~new_new_n2357__;
  assign new_new_n2359__ = ~new_new_n2221__ & ~new_new_n2358__;
  assign new_new_n2360__ = ~new_new_n2213__ & new_new_n2359__;
  assign new_new_n2361__ = ~new_new_n2212__ & ~new_new_n2360__;
  assign new_new_n2362__ = ~new_new_n2204__ & ~new_new_n2361__;
  assign new_new_n2363__ = ~new_new_n2203__ & ~new_new_n2362__;
  assign new_new_n2364__ = ~new_new_n2202__ & new_new_n2363__;
  assign new_new_n2365__ = ~new_new_n2201__ & ~new_new_n2364__;
  assign new_new_n2366__ = ~new_new_n2193__ & new_new_n2365__;
  assign new_new_n2367__ = ~new_new_n2192__ & ~new_new_n2366__;
  assign new_new_n2368__ = pi081 & ~new_new_n2367__;
  assign new_new_n2369__ = ~new_new_n2184__ & ~new_new_n2368__;
  assign new_new_n2370__ = ~pi081 & new_new_n2367__;
  assign new_new_n2371__ = ~new_new_n1986__ & ~new_new_n2160__;
  assign new_new_n2372__ = ~pi080 & ~po046;
  assign new_new_n2373__ = ~new_new_n2157__ & po046;
  assign new_new_n2374__ = ~new_new_n2372__ & ~new_new_n2373__;
  assign new_new_n2375__ = new_new_n2371__ & ~new_new_n2374__;
  assign new_new_n2376__ = ~new_new_n2371__ & new_new_n2374__;
  assign new_new_n2377__ = ~new_new_n2375__ & ~new_new_n2376__;
  assign new_new_n2378__ = ~new_new_n2370__ & ~new_new_n2377__;
  assign new_new_n2379__ = new_new_n2369__ & ~new_new_n2378__;
  assign new_new_n2380__ = ~new_new_n2183__ & ~new_new_n2379__;
  assign po045 = new_new_n2179__ & ~new_new_n2380__;
  assign new_new_n2382__ = pi078 & ~new_new_n2361__;
  assign new_new_n2383__ = ~pi078 & new_new_n2361__;
  assign new_new_n2384__ = ~new_new_n2382__ & ~new_new_n2383__;
  assign new_new_n2385__ = po045 & new_new_n2384__;
  assign new_new_n2386__ = new_new_n2178__ & new_new_n2385__;
  assign new_new_n2387__ = ~new_new_n2178__ & ~new_new_n2385__;
  assign new_new_n2388__ = ~new_new_n2386__ & ~new_new_n2387__;
  assign new_new_n2389__ = pi079 & ~new_new_n2388__;
  assign new_new_n2390__ = ~pi079 & new_new_n2388__;
  assign new_new_n2391__ = ~new_new_n2212__ & ~new_new_n2213__;
  assign new_new_n2392__ = ~new_new_n2359__ & po045;
  assign new_new_n2393__ = ~pi077 & ~po045;
  assign new_new_n2394__ = ~new_new_n2392__ & ~new_new_n2393__;
  assign new_new_n2395__ = new_new_n2391__ & ~new_new_n2394__;
  assign new_new_n2396__ = ~new_new_n2391__ & new_new_n2394__;
  assign new_new_n2397__ = ~new_new_n2395__ & ~new_new_n2396__;
  assign new_new_n2398__ = pi078 & ~new_new_n2397__;
  assign new_new_n2399__ = ~pi078 & new_new_n2397__;
  assign new_new_n2400__ = ~new_new_n2221__ & ~new_new_n2222__;
  assign new_new_n2401__ = ~new_new_n2357__ & po045;
  assign new_new_n2402__ = ~pi076 & ~po045;
  assign new_new_n2403__ = ~new_new_n2401__ & ~new_new_n2402__;
  assign new_new_n2404__ = new_new_n2400__ & ~new_new_n2403__;
  assign new_new_n2405__ = ~new_new_n2400__ & new_new_n2403__;
  assign new_new_n2406__ = ~new_new_n2404__ & ~new_new_n2405__;
  assign new_new_n2407__ = pi077 & ~new_new_n2406__;
  assign new_new_n2408__ = ~pi077 & new_new_n2406__;
  assign new_new_n2409__ = ~new_new_n2230__ & ~new_new_n2231__;
  assign new_new_n2410__ = ~new_new_n2355__ & po045;
  assign new_new_n2411__ = ~pi075 & ~po045;
  assign new_new_n2412__ = ~new_new_n2410__ & ~new_new_n2411__;
  assign new_new_n2413__ = new_new_n2409__ & ~new_new_n2412__;
  assign new_new_n2414__ = ~new_new_n2409__ & new_new_n2412__;
  assign new_new_n2415__ = ~new_new_n2413__ & ~new_new_n2414__;
  assign new_new_n2416__ = ~pi076 & new_new_n2415__;
  assign new_new_n2417__ = pi076 & ~new_new_n2415__;
  assign new_new_n2418__ = ~new_new_n2239__ & ~new_new_n2240__;
  assign new_new_n2419__ = ~new_new_n2353__ & po045;
  assign new_new_n2420__ = ~pi074 & ~po045;
  assign new_new_n2421__ = ~new_new_n2419__ & ~new_new_n2420__;
  assign new_new_n2422__ = new_new_n2418__ & ~new_new_n2421__;
  assign new_new_n2423__ = ~new_new_n2418__ & new_new_n2421__;
  assign new_new_n2424__ = ~new_new_n2422__ & ~new_new_n2423__;
  assign new_new_n2425__ = ~pi075 & new_new_n2424__;
  assign new_new_n2426__ = pi075 & ~new_new_n2424__;
  assign new_new_n2427__ = ~new_new_n2248__ & ~new_new_n2249__;
  assign new_new_n2428__ = ~new_new_n2351__ & po045;
  assign new_new_n2429__ = pi073 & ~po045;
  assign new_new_n2430__ = ~new_new_n2428__ & ~new_new_n2429__;
  assign new_new_n2431__ = new_new_n2427__ & ~new_new_n2430__;
  assign new_new_n2432__ = ~new_new_n2427__ & new_new_n2430__;
  assign new_new_n2433__ = ~new_new_n2431__ & ~new_new_n2432__;
  assign new_new_n2434__ = ~pi074 & ~new_new_n2433__;
  assign new_new_n2435__ = pi074 & new_new_n2433__;
  assign new_new_n2436__ = ~new_new_n2349__ & po045;
  assign new_new_n2437__ = pi072 & ~po045;
  assign new_new_n2438__ = ~new_new_n2436__ & ~new_new_n2437__;
  assign new_new_n2439__ = ~new_new_n2257__ & ~new_new_n2258__;
  assign new_new_n2440__ = ~new_new_n2438__ & new_new_n2439__;
  assign new_new_n2441__ = new_new_n2438__ & ~new_new_n2439__;
  assign new_new_n2442__ = ~new_new_n2440__ & ~new_new_n2441__;
  assign new_new_n2443__ = pi073 & new_new_n2442__;
  assign new_new_n2444__ = ~pi073 & ~new_new_n2442__;
  assign new_new_n2445__ = ~new_new_n2266__ & ~new_new_n2267__;
  assign new_new_n2446__ = ~new_new_n2347__ & po045;
  assign new_new_n2447__ = ~pi071 & ~po045;
  assign new_new_n2448__ = ~new_new_n2446__ & ~new_new_n2447__;
  assign new_new_n2449__ = new_new_n2445__ & ~new_new_n2448__;
  assign new_new_n2450__ = ~new_new_n2445__ & new_new_n2448__;
  assign new_new_n2451__ = ~new_new_n2449__ & ~new_new_n2450__;
  assign new_new_n2452__ = pi072 & ~new_new_n2451__;
  assign new_new_n2453__ = ~pi072 & new_new_n2451__;
  assign new_new_n2454__ = ~new_new_n2275__ & ~new_new_n2276__;
  assign new_new_n2455__ = ~new_new_n2345__ & po045;
  assign new_new_n2456__ = ~pi070 & ~po045;
  assign new_new_n2457__ = ~new_new_n2455__ & ~new_new_n2456__;
  assign new_new_n2458__ = ~new_new_n2454__ & ~new_new_n2457__;
  assign new_new_n2459__ = new_new_n2454__ & new_new_n2457__;
  assign new_new_n2460__ = ~new_new_n2458__ & ~new_new_n2459__;
  assign new_new_n2461__ = ~pi071 & ~new_new_n2460__;
  assign new_new_n2462__ = pi071 & new_new_n2460__;
  assign new_new_n2463__ = ~new_new_n2282__ & ~new_new_n2283__;
  assign new_new_n2464__ = ~new_new_n2343__ & po045;
  assign new_new_n2465__ = ~pi069 & ~po045;
  assign new_new_n2466__ = ~new_new_n2464__ & ~new_new_n2465__;
  assign new_new_n2467__ = new_new_n2463__ & ~new_new_n2466__;
  assign new_new_n2468__ = ~new_new_n2463__ & new_new_n2466__;
  assign new_new_n2469__ = ~new_new_n2467__ & ~new_new_n2468__;
  assign new_new_n2470__ = pi070 & ~new_new_n2469__;
  assign new_new_n2471__ = ~pi070 & new_new_n2469__;
  assign new_new_n2472__ = ~new_new_n2291__ & ~new_new_n2292__;
  assign new_new_n2473__ = ~new_new_n2341__ & po045;
  assign new_new_n2474__ = ~pi068 & ~po045;
  assign new_new_n2475__ = ~new_new_n2473__ & ~new_new_n2474__;
  assign new_new_n2476__ = ~new_new_n2472__ & ~new_new_n2475__;
  assign new_new_n2477__ = new_new_n2472__ & new_new_n2475__;
  assign new_new_n2478__ = ~new_new_n2476__ & ~new_new_n2477__;
  assign new_new_n2479__ = ~pi069 & ~new_new_n2478__;
  assign new_new_n2480__ = pi069 & new_new_n2478__;
  assign new_new_n2481__ = ~new_new_n2311__ & ~new_new_n2312__;
  assign new_new_n2482__ = po045 & new_new_n2481__;
  assign new_new_n2483__ = ~new_new_n2337__ & new_new_n2482__;
  assign new_new_n2484__ = new_new_n2337__ & ~new_new_n2482__;
  assign new_new_n2485__ = ~new_new_n2483__ & ~new_new_n2484__;
  assign new_new_n2486__ = pi067 & ~new_new_n2485__;
  assign new_new_n2487__ = pi045 & po045;
  assign new_new_n2488__ = ~pi045 & ~po045;
  assign new_new_n2489__ = ~pi065 & ~new_new_n2487__;
  assign new_new_n2490__ = ~new_new_n2488__ & new_new_n2489__;
  assign new_new_n2491__ = ~pi044 & ~new_new_n2490__;
  assign new_new_n2492__ = pi065 & new_new_n2487__;
  assign new_new_n2493__ = ~new_new_n2491__ & ~new_new_n2492__;
  assign new_new_n2494__ = pi064 & ~new_new_n2493__;
  assign new_new_n2495__ = pi064 & po045;
  assign new_new_n2496__ = ~pi045 & pi065;
  assign new_new_n2497__ = ~new_new_n2495__ & new_new_n2496__;
  assign new_new_n2498__ = ~new_new_n2494__ & ~new_new_n2497__;
  assign new_new_n2499__ = pi066 & ~new_new_n2498__;
  assign new_new_n2500__ = new_new_n426__ & ~po046;
  assign new_new_n2501__ = new_new_n2330__ & po045;
  assign new_new_n2502__ = ~new_new_n2500__ & ~new_new_n2501__;
  assign new_new_n2503__ = ~pi045 & ~new_new_n2502__;
  assign new_new_n2504__ = ~new_new_n332__ & po045;
  assign new_new_n2505__ = ~new_new_n2308__ & ~new_new_n2504__;
  assign new_new_n2506__ = pi065 & ~new_new_n2308__;
  assign new_new_n2507__ = pi065 & po045;
  assign new_new_n2508__ = po046 & ~new_new_n2507__;
  assign new_new_n2509__ = pi045 & ~new_new_n2506__;
  assign new_new_n2510__ = ~new_new_n2508__ & new_new_n2509__;
  assign new_new_n2511__ = ~new_new_n2503__ & ~new_new_n2505__;
  assign new_new_n2512__ = ~new_new_n2510__ & new_new_n2511__;
  assign new_new_n2513__ = ~pi046 & ~new_new_n2512__;
  assign new_new_n2514__ = ~pi064 & ~new_new_n2507__;
  assign new_new_n2515__ = ~pi065 & po045;
  assign new_new_n2516__ = ~po046 & ~new_new_n2515__;
  assign new_new_n2517__ = ~new_new_n2487__ & ~new_new_n2501__;
  assign new_new_n2518__ = ~new_new_n2516__ & new_new_n2517__;
  assign new_new_n2519__ = pi064 & ~new_new_n2518__;
  assign new_new_n2520__ = ~new_new_n2514__ & ~new_new_n2519__;
  assign new_new_n2521__ = ~new_new_n2308__ & ~new_new_n2507__;
  assign new_new_n2522__ = pi045 & ~new_new_n2313__;
  assign new_new_n2523__ = ~new_new_n2521__ & new_new_n2522__;
  assign new_new_n2524__ = ~new_new_n2520__ & ~new_new_n2523__;
  assign new_new_n2525__ = pi046 & ~new_new_n2524__;
  assign new_new_n2526__ = ~new_new_n2513__ & ~new_new_n2525__;
  assign new_new_n2527__ = ~pi066 & new_new_n2498__;
  assign new_new_n2528__ = ~new_new_n2526__ & ~new_new_n2527__;
  assign new_new_n2529__ = ~new_new_n2499__ & ~new_new_n2528__;
  assign new_new_n2530__ = ~pi067 & new_new_n2485__;
  assign new_new_n2531__ = ~new_new_n2529__ & ~new_new_n2530__;
  assign new_new_n2532__ = ~new_new_n2486__ & ~new_new_n2531__;
  assign new_new_n2533__ = ~pi068 & new_new_n2532__;
  assign new_new_n2534__ = pi068 & ~new_new_n2532__;
  assign new_new_n2535__ = new_new_n2339__ & po045;
  assign new_new_n2536__ = ~pi067 & ~po045;
  assign new_new_n2537__ = ~new_new_n2535__ & ~new_new_n2536__;
  assign new_new_n2538__ = ~new_new_n2298__ & ~new_new_n2299__;
  assign new_new_n2539__ = ~new_new_n2537__ & ~new_new_n2538__;
  assign new_new_n2540__ = new_new_n2537__ & new_new_n2538__;
  assign new_new_n2541__ = ~new_new_n2539__ & ~new_new_n2540__;
  assign new_new_n2542__ = ~new_new_n2534__ & ~new_new_n2541__;
  assign new_new_n2543__ = ~new_new_n2533__ & ~new_new_n2542__;
  assign new_new_n2544__ = ~new_new_n2480__ & ~new_new_n2543__;
  assign new_new_n2545__ = ~new_new_n2479__ & ~new_new_n2544__;
  assign new_new_n2546__ = ~new_new_n2471__ & new_new_n2545__;
  assign new_new_n2547__ = ~new_new_n2470__ & ~new_new_n2546__;
  assign new_new_n2548__ = ~new_new_n2462__ & new_new_n2547__;
  assign new_new_n2549__ = ~new_new_n2461__ & ~new_new_n2548__;
  assign new_new_n2550__ = ~new_new_n2453__ & new_new_n2549__;
  assign new_new_n2551__ = ~new_new_n2452__ & ~new_new_n2550__;
  assign new_new_n2552__ = ~new_new_n2444__ & ~new_new_n2551__;
  assign new_new_n2553__ = ~new_new_n2443__ & ~new_new_n2552__;
  assign new_new_n2554__ = ~new_new_n2435__ & new_new_n2553__;
  assign new_new_n2555__ = ~new_new_n2434__ & ~new_new_n2554__;
  assign new_new_n2556__ = ~new_new_n2426__ & ~new_new_n2555__;
  assign new_new_n2557__ = ~new_new_n2425__ & ~new_new_n2556__;
  assign new_new_n2558__ = ~new_new_n2417__ & ~new_new_n2557__;
  assign new_new_n2559__ = ~new_new_n2416__ & ~new_new_n2558__;
  assign new_new_n2560__ = ~new_new_n2408__ & new_new_n2559__;
  assign new_new_n2561__ = ~new_new_n2407__ & ~new_new_n2560__;
  assign new_new_n2562__ = ~new_new_n2399__ & ~new_new_n2561__;
  assign new_new_n2563__ = ~new_new_n2398__ & ~new_new_n2562__;
  assign new_new_n2564__ = ~new_new_n2390__ & ~new_new_n2563__;
  assign new_new_n2565__ = ~new_new_n2389__ & ~new_new_n2564__;
  assign new_new_n2566__ = ~pi084 & new_new_n2159__;
  assign new_new_n2567__ = new_new_n2181__ & ~po045;
  assign new_new_n2568__ = ~new_new_n376__ & ~new_new_n2567__;
  assign new_new_n2569__ = ~pi083 & ~new_new_n2568__;
  assign new_new_n2570__ = pi083 & new_new_n2568__;
  assign new_new_n2571__ = new_new_n2365__ & po045;
  assign new_new_n2572__ = pi080 & ~po045;
  assign new_new_n2573__ = ~new_new_n2571__ & ~new_new_n2572__;
  assign new_new_n2574__ = ~new_new_n2192__ & ~new_new_n2193__;
  assign new_new_n2575__ = ~new_new_n2573__ & ~new_new_n2574__;
  assign new_new_n2576__ = new_new_n2573__ & new_new_n2574__;
  assign new_new_n2577__ = ~new_new_n2575__ & ~new_new_n2576__;
  assign new_new_n2578__ = pi081 & ~new_new_n2577__;
  assign new_new_n2579__ = ~pi081 & new_new_n2577__;
  assign new_new_n2580__ = ~new_new_n2363__ & po045;
  assign new_new_n2581__ = pi079 & ~po045;
  assign new_new_n2582__ = ~new_new_n2580__ & ~new_new_n2581__;
  assign new_new_n2583__ = ~new_new_n2201__ & ~new_new_n2202__;
  assign new_new_n2584__ = ~new_new_n2582__ & new_new_n2583__;
  assign new_new_n2585__ = new_new_n2582__ & ~new_new_n2583__;
  assign new_new_n2586__ = ~new_new_n2584__ & ~new_new_n2585__;
  assign new_new_n2587__ = ~pi080 & ~new_new_n2586__;
  assign new_new_n2588__ = pi080 & new_new_n2586__;
  assign new_new_n2589__ = new_new_n2565__ & ~new_new_n2588__;
  assign new_new_n2590__ = ~new_new_n2587__ & ~new_new_n2589__;
  assign new_new_n2591__ = ~new_new_n2579__ & new_new_n2590__;
  assign new_new_n2592__ = ~new_new_n2578__ & ~new_new_n2591__;
  assign new_new_n2593__ = pi082 & ~new_new_n2592__;
  assign new_new_n2594__ = ~new_new_n2570__ & ~new_new_n2593__;
  assign new_new_n2595__ = new_new_n2179__ & ~new_new_n2370__;
  assign new_new_n2596__ = new_new_n2369__ & new_new_n2595__;
  assign new_new_n2597__ = new_new_n2377__ & ~new_new_n2596__;
  assign new_new_n2598__ = new_new_n2183__ & ~new_new_n2377__;
  assign new_new_n2599__ = ~new_new_n2368__ & new_new_n2598__;
  assign new_new_n2600__ = new_new_n2595__ & new_new_n2599__;
  assign new_new_n2601__ = ~new_new_n2597__ & ~new_new_n2600__;
  assign new_new_n2602__ = ~pi082 & new_new_n2592__;
  assign new_new_n2603__ = new_new_n2601__ & ~new_new_n2602__;
  assign new_new_n2604__ = new_new_n2594__ & ~new_new_n2603__;
  assign new_new_n2605__ = ~new_new_n2569__ & ~new_new_n2604__;
  assign po044 = new_new_n2566__ & ~new_new_n2605__;
  assign new_new_n2607__ = ~new_new_n2565__ & po044;
  assign new_new_n2608__ = pi080 & ~po044;
  assign new_new_n2609__ = ~new_new_n2607__ & ~new_new_n2608__;
  assign new_new_n2610__ = ~new_new_n2587__ & ~new_new_n2588__;
  assign new_new_n2611__ = ~new_new_n2609__ & new_new_n2610__;
  assign new_new_n2612__ = new_new_n2609__ & ~new_new_n2610__;
  assign new_new_n2613__ = ~new_new_n2611__ & ~new_new_n2612__;
  assign new_new_n2614__ = ~pi081 & ~new_new_n2613__;
  assign new_new_n2615__ = pi081 & new_new_n2613__;
  assign new_new_n2616__ = ~new_new_n2614__ & ~new_new_n2615__;
  assign new_new_n2617__ = ~new_new_n2389__ & ~new_new_n2390__;
  assign new_new_n2618__ = ~new_new_n2563__ & po044;
  assign new_new_n2619__ = pi079 & ~po044;
  assign new_new_n2620__ = ~new_new_n2618__ & ~new_new_n2619__;
  assign new_new_n2621__ = new_new_n2617__ & ~new_new_n2620__;
  assign new_new_n2622__ = ~new_new_n2617__ & new_new_n2620__;
  assign new_new_n2623__ = ~new_new_n2621__ & ~new_new_n2622__;
  assign new_new_n2624__ = pi080 & new_new_n2623__;
  assign new_new_n2625__ = ~pi080 & ~new_new_n2623__;
  assign new_new_n2626__ = pi078 & ~new_new_n2561__;
  assign new_new_n2627__ = ~pi078 & new_new_n2561__;
  assign new_new_n2628__ = ~new_new_n2626__ & ~new_new_n2627__;
  assign new_new_n2629__ = po044 & new_new_n2628__;
  assign new_new_n2630__ = new_new_n2397__ & new_new_n2629__;
  assign new_new_n2631__ = ~new_new_n2397__ & ~new_new_n2629__;
  assign new_new_n2632__ = ~new_new_n2630__ & ~new_new_n2631__;
  assign new_new_n2633__ = pi079 & ~new_new_n2632__;
  assign new_new_n2634__ = ~pi079 & new_new_n2632__;
  assign new_new_n2635__ = ~new_new_n2416__ & ~new_new_n2417__;
  assign new_new_n2636__ = ~new_new_n2557__ & po044;
  assign new_new_n2637__ = ~pi076 & ~po044;
  assign new_new_n2638__ = ~new_new_n2636__ & ~new_new_n2637__;
  assign new_new_n2639__ = new_new_n2635__ & ~new_new_n2638__;
  assign new_new_n2640__ = ~new_new_n2635__ & new_new_n2638__;
  assign new_new_n2641__ = ~new_new_n2639__ & ~new_new_n2640__;
  assign new_new_n2642__ = pi077 & ~new_new_n2641__;
  assign new_new_n2643__ = ~pi077 & new_new_n2641__;
  assign new_new_n2644__ = ~new_new_n2425__ & ~new_new_n2426__;
  assign new_new_n2645__ = ~new_new_n2555__ & po044;
  assign new_new_n2646__ = ~pi075 & ~po044;
  assign new_new_n2647__ = ~new_new_n2645__ & ~new_new_n2646__;
  assign new_new_n2648__ = new_new_n2644__ & ~new_new_n2647__;
  assign new_new_n2649__ = ~new_new_n2644__ & new_new_n2647__;
  assign new_new_n2650__ = ~new_new_n2648__ & ~new_new_n2649__;
  assign new_new_n2651__ = ~pi076 & new_new_n2650__;
  assign new_new_n2652__ = pi076 & ~new_new_n2650__;
  assign new_new_n2653__ = ~new_new_n2434__ & ~new_new_n2435__;
  assign new_new_n2654__ = ~new_new_n2553__ & po044;
  assign new_new_n2655__ = pi074 & ~po044;
  assign new_new_n2656__ = ~new_new_n2654__ & ~new_new_n2655__;
  assign new_new_n2657__ = new_new_n2653__ & ~new_new_n2656__;
  assign new_new_n2658__ = ~new_new_n2653__ & new_new_n2656__;
  assign new_new_n2659__ = ~new_new_n2657__ & ~new_new_n2658__;
  assign new_new_n2660__ = ~pi075 & ~new_new_n2659__;
  assign new_new_n2661__ = pi075 & new_new_n2659__;
  assign new_new_n2662__ = ~new_new_n2443__ & ~new_new_n2444__;
  assign new_new_n2663__ = ~new_new_n2551__ & po044;
  assign new_new_n2664__ = pi073 & ~po044;
  assign new_new_n2665__ = ~new_new_n2663__ & ~new_new_n2664__;
  assign new_new_n2666__ = new_new_n2662__ & ~new_new_n2665__;
  assign new_new_n2667__ = ~new_new_n2662__ & new_new_n2665__;
  assign new_new_n2668__ = ~new_new_n2666__ & ~new_new_n2667__;
  assign new_new_n2669__ = ~pi074 & ~new_new_n2668__;
  assign new_new_n2670__ = pi074 & new_new_n2668__;
  assign new_new_n2671__ = ~new_new_n2452__ & ~new_new_n2453__;
  assign new_new_n2672__ = ~new_new_n2549__ & po044;
  assign new_new_n2673__ = ~pi072 & ~po044;
  assign new_new_n2674__ = ~new_new_n2672__ & ~new_new_n2673__;
  assign new_new_n2675__ = new_new_n2671__ & ~new_new_n2674__;
  assign new_new_n2676__ = ~new_new_n2671__ & new_new_n2674__;
  assign new_new_n2677__ = ~new_new_n2675__ & ~new_new_n2676__;
  assign new_new_n2678__ = pi073 & ~new_new_n2677__;
  assign new_new_n2679__ = ~pi073 & new_new_n2677__;
  assign new_new_n2680__ = ~new_new_n2461__ & ~new_new_n2462__;
  assign new_new_n2681__ = new_new_n2547__ & po044;
  assign new_new_n2682__ = ~pi071 & ~po044;
  assign new_new_n2683__ = ~new_new_n2681__ & ~new_new_n2682__;
  assign new_new_n2684__ = ~new_new_n2680__ & ~new_new_n2683__;
  assign new_new_n2685__ = new_new_n2680__ & new_new_n2683__;
  assign new_new_n2686__ = ~new_new_n2684__ & ~new_new_n2685__;
  assign new_new_n2687__ = pi072 & new_new_n2686__;
  assign new_new_n2688__ = ~pi072 & ~new_new_n2686__;
  assign new_new_n2689__ = new_new_n2545__ & po044;
  assign new_new_n2690__ = pi070 & ~po044;
  assign new_new_n2691__ = ~new_new_n2689__ & ~new_new_n2690__;
  assign new_new_n2692__ = ~new_new_n2470__ & ~new_new_n2471__;
  assign new_new_n2693__ = ~new_new_n2691__ & ~new_new_n2692__;
  assign new_new_n2694__ = new_new_n2691__ & new_new_n2692__;
  assign new_new_n2695__ = ~new_new_n2693__ & ~new_new_n2694__;
  assign new_new_n2696__ = pi071 & ~new_new_n2695__;
  assign new_new_n2697__ = ~pi071 & new_new_n2695__;
  assign new_new_n2698__ = ~pi069 & ~new_new_n2543__;
  assign new_new_n2699__ = pi069 & new_new_n2543__;
  assign new_new_n2700__ = ~new_new_n2698__ & ~new_new_n2699__;
  assign new_new_n2701__ = po044 & new_new_n2700__;
  assign new_new_n2702__ = ~new_new_n2478__ & new_new_n2701__;
  assign new_new_n2703__ = new_new_n2478__ & ~new_new_n2701__;
  assign new_new_n2704__ = ~new_new_n2702__ & ~new_new_n2703__;
  assign new_new_n2705__ = pi070 & ~new_new_n2704__;
  assign new_new_n2706__ = ~pi070 & new_new_n2704__;
  assign new_new_n2707__ = ~new_new_n2533__ & ~new_new_n2534__;
  assign new_new_n2708__ = po044 & new_new_n2707__;
  assign new_new_n2709__ = ~new_new_n2541__ & ~new_new_n2708__;
  assign new_new_n2710__ = new_new_n2541__ & new_new_n2708__;
  assign new_new_n2711__ = ~new_new_n2709__ & ~new_new_n2710__;
  assign new_new_n2712__ = pi069 & new_new_n2711__;
  assign new_new_n2713__ = ~pi069 & ~new_new_n2711__;
  assign new_new_n2714__ = ~new_new_n2499__ & ~new_new_n2527__;
  assign new_new_n2715__ = po044 & new_new_n2714__;
  assign new_new_n2716__ = new_new_n2526__ & ~new_new_n2715__;
  assign new_new_n2717__ = ~new_new_n2526__ & new_new_n2715__;
  assign new_new_n2718__ = ~new_new_n2716__ & ~new_new_n2717__;
  assign new_new_n2719__ = pi067 & new_new_n2718__;
  assign new_new_n2720__ = ~pi067 & ~new_new_n2718__;
  assign new_new_n2721__ = pi044 & po044;
  assign new_new_n2722__ = ~pi044 & ~po044;
  assign new_new_n2723__ = ~pi065 & ~new_new_n2721__;
  assign new_new_n2724__ = ~new_new_n2722__ & new_new_n2723__;
  assign new_new_n2725__ = ~pi043 & ~new_new_n2724__;
  assign new_new_n2726__ = pi065 & new_new_n2721__;
  assign new_new_n2727__ = ~new_new_n2725__ & ~new_new_n2726__;
  assign new_new_n2728__ = pi064 & ~new_new_n2727__;
  assign new_new_n2729__ = pi064 & po044;
  assign new_new_n2730__ = ~pi044 & pi065;
  assign new_new_n2731__ = ~new_new_n2729__ & new_new_n2730__;
  assign new_new_n2732__ = ~new_new_n2728__ & ~new_new_n2731__;
  assign new_new_n2733__ = pi066 & ~new_new_n2732__;
  assign new_new_n2734__ = ~pi066 & new_new_n2732__;
  assign new_new_n2735__ = new_new_n426__ & ~po045;
  assign new_new_n2736__ = new_new_n2515__ & po044;
  assign new_new_n2737__ = ~new_new_n2735__ & ~new_new_n2736__;
  assign new_new_n2738__ = ~pi044 & ~new_new_n2737__;
  assign new_new_n2739__ = ~new_new_n332__ & po044;
  assign new_new_n2740__ = ~new_new_n2495__ & ~new_new_n2739__;
  assign new_new_n2741__ = pi065 & po044;
  assign new_new_n2742__ = po045 & ~new_new_n2741__;
  assign new_new_n2743__ = pi065 & ~new_new_n2495__;
  assign new_new_n2744__ = pi044 & ~new_new_n2743__;
  assign new_new_n2745__ = ~new_new_n2742__ & new_new_n2744__;
  assign new_new_n2746__ = ~new_new_n2738__ & ~new_new_n2740__;
  assign new_new_n2747__ = ~new_new_n2745__ & new_new_n2746__;
  assign new_new_n2748__ = pi045 & ~new_new_n2747__;
  assign new_new_n2749__ = ~pi064 & ~new_new_n2741__;
  assign new_new_n2750__ = ~pi065 & po044;
  assign new_new_n2751__ = ~po045 & ~new_new_n2750__;
  assign new_new_n2752__ = ~new_new_n2721__ & ~new_new_n2736__;
  assign new_new_n2753__ = ~new_new_n2751__ & new_new_n2752__;
  assign new_new_n2754__ = pi064 & ~new_new_n2753__;
  assign new_new_n2755__ = ~new_new_n2749__ & ~new_new_n2754__;
  assign new_new_n2756__ = ~new_new_n2495__ & ~new_new_n2741__;
  assign new_new_n2757__ = pi044 & ~new_new_n2507__;
  assign new_new_n2758__ = ~new_new_n2756__ & new_new_n2757__;
  assign new_new_n2759__ = ~new_new_n2755__ & ~new_new_n2758__;
  assign new_new_n2760__ = ~pi045 & ~new_new_n2759__;
  assign new_new_n2761__ = ~new_new_n2748__ & ~new_new_n2760__;
  assign new_new_n2762__ = ~new_new_n2734__ & new_new_n2761__;
  assign new_new_n2763__ = ~new_new_n2733__ & ~new_new_n2762__;
  assign new_new_n2764__ = ~new_new_n2720__ & ~new_new_n2763__;
  assign new_new_n2765__ = ~new_new_n2719__ & ~new_new_n2764__;
  assign new_new_n2766__ = pi068 & ~new_new_n2765__;
  assign new_new_n2767__ = ~pi068 & new_new_n2765__;
  assign new_new_n2768__ = ~new_new_n2486__ & ~new_new_n2530__;
  assign new_new_n2769__ = pi067 & ~po044;
  assign new_new_n2770__ = ~new_new_n2529__ & po044;
  assign new_new_n2771__ = ~new_new_n2769__ & ~new_new_n2770__;
  assign new_new_n2772__ = new_new_n2768__ & ~new_new_n2771__;
  assign new_new_n2773__ = ~new_new_n2768__ & new_new_n2771__;
  assign new_new_n2774__ = ~new_new_n2772__ & ~new_new_n2773__;
  assign new_new_n2775__ = ~new_new_n2767__ & new_new_n2774__;
  assign new_new_n2776__ = ~new_new_n2766__ & ~new_new_n2775__;
  assign new_new_n2777__ = ~new_new_n2713__ & ~new_new_n2776__;
  assign new_new_n2778__ = ~new_new_n2712__ & ~new_new_n2777__;
  assign new_new_n2779__ = ~new_new_n2706__ & ~new_new_n2778__;
  assign new_new_n2780__ = ~new_new_n2705__ & ~new_new_n2779__;
  assign new_new_n2781__ = ~new_new_n2697__ & ~new_new_n2780__;
  assign new_new_n2782__ = ~new_new_n2696__ & ~new_new_n2781__;
  assign new_new_n2783__ = ~new_new_n2688__ & ~new_new_n2782__;
  assign new_new_n2784__ = ~new_new_n2687__ & ~new_new_n2783__;
  assign new_new_n2785__ = ~new_new_n2679__ & ~new_new_n2784__;
  assign new_new_n2786__ = ~new_new_n2678__ & ~new_new_n2785__;
  assign new_new_n2787__ = ~new_new_n2670__ & new_new_n2786__;
  assign new_new_n2788__ = ~new_new_n2669__ & ~new_new_n2787__;
  assign new_new_n2789__ = ~new_new_n2661__ & ~new_new_n2788__;
  assign new_new_n2790__ = ~new_new_n2660__ & ~new_new_n2789__;
  assign new_new_n2791__ = ~new_new_n2652__ & ~new_new_n2790__;
  assign new_new_n2792__ = ~new_new_n2651__ & ~new_new_n2791__;
  assign new_new_n2793__ = ~new_new_n2643__ & new_new_n2792__;
  assign new_new_n2794__ = ~new_new_n2642__ & ~new_new_n2793__;
  assign new_new_n2795__ = ~pi078 & new_new_n2794__;
  assign new_new_n2796__ = pi078 & ~new_new_n2794__;
  assign new_new_n2797__ = ~new_new_n2407__ & ~new_new_n2408__;
  assign new_new_n2798__ = ~new_new_n2559__ & po044;
  assign new_new_n2799__ = ~pi077 & ~po044;
  assign new_new_n2800__ = ~new_new_n2798__ & ~new_new_n2799__;
  assign new_new_n2801__ = new_new_n2797__ & ~new_new_n2800__;
  assign new_new_n2802__ = ~new_new_n2797__ & new_new_n2800__;
  assign new_new_n2803__ = ~new_new_n2801__ & ~new_new_n2802__;
  assign new_new_n2804__ = ~new_new_n2796__ & new_new_n2803__;
  assign new_new_n2805__ = ~new_new_n2795__ & ~new_new_n2804__;
  assign new_new_n2806__ = ~new_new_n2634__ & new_new_n2805__;
  assign new_new_n2807__ = ~new_new_n2633__ & ~new_new_n2806__;
  assign new_new_n2808__ = ~new_new_n2625__ & ~new_new_n2807__;
  assign new_new_n2809__ = ~new_new_n2624__ & ~new_new_n2808__;
  assign new_new_n2810__ = new_new_n2566__ & ~new_new_n2602__;
  assign new_new_n2811__ = new_new_n2594__ & new_new_n2810__;
  assign new_new_n2812__ = ~new_new_n2601__ & ~new_new_n2811__;
  assign new_new_n2813__ = new_new_n2566__ & ~new_new_n2568__;
  assign new_new_n2814__ = ~new_new_n2593__ & new_new_n2813__;
  assign new_new_n2815__ = new_new_n2603__ & new_new_n2814__;
  assign new_new_n2816__ = ~new_new_n2812__ & ~new_new_n2815__;
  assign new_new_n2817__ = ~pi083 & ~new_new_n2816__;
  assign new_new_n2818__ = pi083 & ~new_new_n2812__;
  assign new_new_n2819__ = new_new_n2590__ & po044;
  assign new_new_n2820__ = pi081 & ~po044;
  assign new_new_n2821__ = ~new_new_n2819__ & ~new_new_n2820__;
  assign new_new_n2822__ = ~new_new_n2578__ & ~new_new_n2579__;
  assign new_new_n2823__ = ~new_new_n2821__ & ~new_new_n2822__;
  assign new_new_n2824__ = new_new_n2821__ & new_new_n2822__;
  assign new_new_n2825__ = ~new_new_n2823__ & ~new_new_n2824__;
  assign new_new_n2826__ = ~pi082 & new_new_n2825__;
  assign new_new_n2827__ = pi082 & ~new_new_n2825__;
  assign new_new_n2828__ = ~new_new_n2615__ & new_new_n2809__;
  assign new_new_n2829__ = ~new_new_n2614__ & ~new_new_n2828__;
  assign new_new_n2830__ = ~new_new_n2827__ & ~new_new_n2829__;
  assign new_new_n2831__ = ~new_new_n2826__ & ~new_new_n2830__;
  assign new_new_n2832__ = ~new_new_n2818__ & ~new_new_n2831__;
  assign new_new_n2833__ = ~new_new_n2817__ & ~new_new_n2832__;
  assign new_new_n2834__ = ~pi084 & ~new_new_n2833__;
  assign new_new_n2835__ = ~new_new_n376__ & po044;
  assign new_new_n2836__ = ~new_new_n2568__ & ~new_new_n2835__;
  assign new_new_n2837__ = ~new_new_n2834__ & ~new_new_n2836__;
  assign new_new_n2838__ = pi084 & new_new_n2833__;
  assign new_new_n2839__ = new_new_n2159__ & ~new_new_n2838__;
  assign po043 = ~new_new_n2837__ & new_new_n2839__;
  assign new_new_n2841__ = ~new_new_n2809__ & po043;
  assign new_new_n2842__ = pi081 & ~po043;
  assign new_new_n2843__ = ~new_new_n2841__ & ~new_new_n2842__;
  assign new_new_n2844__ = new_new_n2616__ & ~new_new_n2843__;
  assign new_new_n2845__ = ~new_new_n2616__ & new_new_n2843__;
  assign new_new_n2846__ = ~new_new_n2844__ & ~new_new_n2845__;
  assign new_new_n2847__ = new_new_n2836__ & ~new_new_n2839__;
  assign new_new_n2848__ = ~pi085 & new_new_n2847__;
  assign new_new_n2849__ = ~new_new_n2826__ & ~new_new_n2827__;
  assign new_new_n2850__ = ~new_new_n2829__ & po043;
  assign new_new_n2851__ = ~pi082 & ~po043;
  assign new_new_n2852__ = ~new_new_n2850__ & ~new_new_n2851__;
  assign new_new_n2853__ = new_new_n2849__ & ~new_new_n2852__;
  assign new_new_n2854__ = ~new_new_n2849__ & new_new_n2852__;
  assign new_new_n2855__ = ~new_new_n2853__ & ~new_new_n2854__;
  assign new_new_n2856__ = ~pi083 & new_new_n2855__;
  assign new_new_n2857__ = pi083 & ~new_new_n2855__;
  assign new_new_n2858__ = ~pi082 & ~new_new_n2846__;
  assign new_new_n2859__ = pi082 & new_new_n2846__;
  assign new_new_n2860__ = ~new_new_n2807__ & po043;
  assign new_new_n2861__ = pi080 & ~po043;
  assign new_new_n2862__ = ~new_new_n2860__ & ~new_new_n2861__;
  assign new_new_n2863__ = ~new_new_n2624__ & ~new_new_n2625__;
  assign new_new_n2864__ = ~new_new_n2862__ & new_new_n2863__;
  assign new_new_n2865__ = new_new_n2862__ & ~new_new_n2863__;
  assign new_new_n2866__ = ~new_new_n2864__ & ~new_new_n2865__;
  assign new_new_n2867__ = ~pi081 & ~new_new_n2866__;
  assign new_new_n2868__ = pi081 & new_new_n2866__;
  assign new_new_n2869__ = ~new_new_n2633__ & ~new_new_n2634__;
  assign new_new_n2870__ = ~new_new_n2805__ & po043;
  assign new_new_n2871__ = ~pi079 & ~po043;
  assign new_new_n2872__ = ~new_new_n2870__ & ~new_new_n2871__;
  assign new_new_n2873__ = new_new_n2869__ & ~new_new_n2872__;
  assign new_new_n2874__ = ~new_new_n2869__ & new_new_n2872__;
  assign new_new_n2875__ = ~new_new_n2873__ & ~new_new_n2874__;
  assign new_new_n2876__ = pi080 & ~new_new_n2875__;
  assign new_new_n2877__ = ~pi080 & new_new_n2875__;
  assign new_new_n2878__ = ~new_new_n2795__ & ~new_new_n2796__;
  assign new_new_n2879__ = po043 & new_new_n2878__;
  assign new_new_n2880__ = new_new_n2803__ & new_new_n2879__;
  assign new_new_n2881__ = ~new_new_n2803__ & ~new_new_n2879__;
  assign new_new_n2882__ = ~new_new_n2880__ & ~new_new_n2881__;
  assign new_new_n2883__ = pi079 & ~new_new_n2882__;
  assign new_new_n2884__ = ~pi079 & new_new_n2882__;
  assign new_new_n2885__ = ~new_new_n2642__ & ~new_new_n2643__;
  assign new_new_n2886__ = ~new_new_n2792__ & po043;
  assign new_new_n2887__ = ~pi077 & ~po043;
  assign new_new_n2888__ = ~new_new_n2886__ & ~new_new_n2887__;
  assign new_new_n2889__ = new_new_n2885__ & ~new_new_n2888__;
  assign new_new_n2890__ = ~new_new_n2885__ & new_new_n2888__;
  assign new_new_n2891__ = ~new_new_n2889__ & ~new_new_n2890__;
  assign new_new_n2892__ = pi078 & ~new_new_n2891__;
  assign new_new_n2893__ = ~pi078 & new_new_n2891__;
  assign new_new_n2894__ = new_new_n2790__ & po043;
  assign new_new_n2895__ = pi076 & ~po043;
  assign new_new_n2896__ = ~new_new_n2894__ & ~new_new_n2895__;
  assign new_new_n2897__ = ~new_new_n2651__ & ~new_new_n2652__;
  assign new_new_n2898__ = ~new_new_n2896__ & ~new_new_n2897__;
  assign new_new_n2899__ = new_new_n2896__ & new_new_n2897__;
  assign new_new_n2900__ = ~new_new_n2898__ & ~new_new_n2899__;
  assign new_new_n2901__ = ~pi077 & new_new_n2900__;
  assign new_new_n2902__ = pi077 & ~new_new_n2900__;
  assign new_new_n2903__ = ~pi075 & ~new_new_n2788__;
  assign new_new_n2904__ = pi075 & new_new_n2788__;
  assign new_new_n2905__ = ~new_new_n2903__ & ~new_new_n2904__;
  assign new_new_n2906__ = po043 & new_new_n2905__;
  assign new_new_n2907__ = new_new_n2659__ & new_new_n2906__;
  assign new_new_n2908__ = ~new_new_n2659__ & ~new_new_n2906__;
  assign new_new_n2909__ = ~new_new_n2907__ & ~new_new_n2908__;
  assign new_new_n2910__ = ~pi076 & ~new_new_n2909__;
  assign new_new_n2911__ = pi076 & new_new_n2909__;
  assign new_new_n2912__ = ~new_new_n2669__ & ~new_new_n2670__;
  assign new_new_n2913__ = ~new_new_n2786__ & po043;
  assign new_new_n2914__ = pi074 & ~po043;
  assign new_new_n2915__ = ~new_new_n2913__ & ~new_new_n2914__;
  assign new_new_n2916__ = new_new_n2912__ & ~new_new_n2915__;
  assign new_new_n2917__ = ~new_new_n2912__ & new_new_n2915__;
  assign new_new_n2918__ = ~new_new_n2916__ & ~new_new_n2917__;
  assign new_new_n2919__ = ~pi075 & ~new_new_n2918__;
  assign new_new_n2920__ = pi075 & new_new_n2918__;
  assign new_new_n2921__ = ~new_new_n2678__ & ~new_new_n2679__;
  assign new_new_n2922__ = ~new_new_n2784__ & po043;
  assign new_new_n2923__ = pi073 & ~po043;
  assign new_new_n2924__ = ~new_new_n2922__ & ~new_new_n2923__;
  assign new_new_n2925__ = new_new_n2921__ & ~new_new_n2924__;
  assign new_new_n2926__ = ~new_new_n2921__ & new_new_n2924__;
  assign new_new_n2927__ = ~new_new_n2925__ & ~new_new_n2926__;
  assign new_new_n2928__ = pi074 & new_new_n2927__;
  assign new_new_n2929__ = ~pi074 & ~new_new_n2927__;
  assign new_new_n2930__ = ~new_new_n2687__ & ~new_new_n2688__;
  assign new_new_n2931__ = new_new_n2782__ & po043;
  assign new_new_n2932__ = ~pi072 & ~po043;
  assign new_new_n2933__ = ~new_new_n2931__ & ~new_new_n2932__;
  assign new_new_n2934__ = ~new_new_n2930__ & ~new_new_n2933__;
  assign new_new_n2935__ = new_new_n2930__ & new_new_n2933__;
  assign new_new_n2936__ = ~new_new_n2934__ & ~new_new_n2935__;
  assign new_new_n2937__ = pi073 & new_new_n2936__;
  assign new_new_n2938__ = ~pi073 & ~new_new_n2936__;
  assign new_new_n2939__ = ~new_new_n2780__ & po043;
  assign new_new_n2940__ = pi071 & ~po043;
  assign new_new_n2941__ = ~new_new_n2939__ & ~new_new_n2940__;
  assign new_new_n2942__ = ~new_new_n2696__ & ~new_new_n2697__;
  assign new_new_n2943__ = new_new_n2941__ & new_new_n2942__;
  assign new_new_n2944__ = ~new_new_n2941__ & ~new_new_n2942__;
  assign new_new_n2945__ = ~new_new_n2943__ & ~new_new_n2944__;
  assign new_new_n2946__ = pi072 & ~new_new_n2945__;
  assign new_new_n2947__ = ~pi072 & new_new_n2945__;
  assign new_new_n2948__ = ~new_new_n2778__ & po043;
  assign new_new_n2949__ = pi070 & ~po043;
  assign new_new_n2950__ = ~new_new_n2948__ & ~new_new_n2949__;
  assign new_new_n2951__ = ~new_new_n2705__ & ~new_new_n2706__;
  assign new_new_n2952__ = ~new_new_n2950__ & new_new_n2951__;
  assign new_new_n2953__ = new_new_n2950__ & ~new_new_n2951__;
  assign new_new_n2954__ = ~new_new_n2952__ & ~new_new_n2953__;
  assign new_new_n2955__ = pi071 & new_new_n2954__;
  assign new_new_n2956__ = ~pi071 & ~new_new_n2954__;
  assign new_new_n2957__ = ~new_new_n2712__ & ~new_new_n2713__;
  assign new_new_n2958__ = ~new_new_n2776__ & po043;
  assign new_new_n2959__ = pi069 & ~po043;
  assign new_new_n2960__ = ~new_new_n2958__ & ~new_new_n2959__;
  assign new_new_n2961__ = new_new_n2957__ & ~new_new_n2960__;
  assign new_new_n2962__ = ~new_new_n2957__ & new_new_n2960__;
  assign new_new_n2963__ = ~new_new_n2961__ & ~new_new_n2962__;
  assign new_new_n2964__ = pi070 & new_new_n2963__;
  assign new_new_n2965__ = ~pi070 & ~new_new_n2963__;
  assign new_new_n2966__ = ~new_new_n2766__ & ~new_new_n2767__;
  assign new_new_n2967__ = po043 & new_new_n2966__;
  assign new_new_n2968__ = new_new_n2774__ & new_new_n2967__;
  assign new_new_n2969__ = ~new_new_n2774__ & ~new_new_n2967__;
  assign new_new_n2970__ = ~new_new_n2968__ & ~new_new_n2969__;
  assign new_new_n2971__ = pi069 & new_new_n2970__;
  assign new_new_n2972__ = ~pi069 & ~new_new_n2970__;
  assign new_new_n2973__ = ~new_new_n2719__ & ~new_new_n2720__;
  assign new_new_n2974__ = ~new_new_n2763__ & po043;
  assign new_new_n2975__ = pi067 & ~po043;
  assign new_new_n2976__ = ~new_new_n2974__ & ~new_new_n2975__;
  assign new_new_n2977__ = new_new_n2973__ & ~new_new_n2976__;
  assign new_new_n2978__ = ~new_new_n2973__ & new_new_n2976__;
  assign new_new_n2979__ = ~new_new_n2977__ & ~new_new_n2978__;
  assign new_new_n2980__ = pi068 & new_new_n2979__;
  assign new_new_n2981__ = ~pi068 & ~new_new_n2979__;
  assign new_new_n2982__ = ~new_new_n2733__ & ~new_new_n2734__;
  assign new_new_n2983__ = po043 & new_new_n2982__;
  assign new_new_n2984__ = ~new_new_n2761__ & new_new_n2983__;
  assign new_new_n2985__ = new_new_n2761__ & ~new_new_n2983__;
  assign new_new_n2986__ = ~new_new_n2984__ & ~new_new_n2985__;
  assign new_new_n2987__ = pi067 & ~new_new_n2986__;
  assign new_new_n2988__ = ~pi067 & new_new_n2986__;
  assign new_new_n2989__ = pi043 & po043;
  assign new_new_n2990__ = pi042 & ~pi065;
  assign new_new_n2991__ = new_new_n2989__ & ~new_new_n2990__;
  assign new_new_n2992__ = ~pi043 & ~po043;
  assign new_new_n2993__ = ~pi065 & ~new_new_n2992__;
  assign new_new_n2994__ = ~pi042 & ~new_new_n2993__;
  assign new_new_n2995__ = ~new_new_n2991__ & ~new_new_n2994__;
  assign new_new_n2996__ = pi064 & ~new_new_n2995__;
  assign new_new_n2997__ = pi064 & po043;
  assign new_new_n2998__ = ~pi043 & pi065;
  assign new_new_n2999__ = ~new_new_n2997__ & new_new_n2998__;
  assign new_new_n3000__ = ~new_new_n2996__ & ~new_new_n2999__;
  assign new_new_n3001__ = pi066 & ~new_new_n3000__;
  assign new_new_n3002__ = ~pi066 & new_new_n3000__;
  assign new_new_n3003__ = new_new_n426__ & ~po044;
  assign new_new_n3004__ = new_new_n2750__ & po043;
  assign new_new_n3005__ = ~new_new_n3003__ & ~new_new_n3004__;
  assign new_new_n3006__ = ~pi043 & ~new_new_n3005__;
  assign new_new_n3007__ = ~new_new_n332__ & po043;
  assign new_new_n3008__ = ~new_new_n2729__ & ~new_new_n3007__;
  assign new_new_n3009__ = pi065 & po043;
  assign new_new_n3010__ = po044 & ~new_new_n3009__;
  assign new_new_n3011__ = pi065 & ~new_new_n2729__;
  assign new_new_n3012__ = pi043 & ~new_new_n3011__;
  assign new_new_n3013__ = ~new_new_n3010__ & new_new_n3012__;
  assign new_new_n3014__ = ~new_new_n3006__ & ~new_new_n3008__;
  assign new_new_n3015__ = ~new_new_n3013__ & new_new_n3014__;
  assign new_new_n3016__ = pi044 & ~new_new_n3015__;
  assign new_new_n3017__ = ~new_new_n2729__ & ~new_new_n3009__;
  assign new_new_n3018__ = pi043 & ~new_new_n2741__;
  assign new_new_n3019__ = pi064 & ~new_new_n3018__;
  assign new_new_n3020__ = ~new_new_n3017__ & ~new_new_n3019__;
  assign new_new_n3021__ = ~pi065 & po043;
  assign new_new_n3022__ = ~po044 & ~new_new_n3021__;
  assign new_new_n3023__ = pi064 & ~new_new_n2989__;
  assign new_new_n3024__ = ~new_new_n3004__ & new_new_n3023__;
  assign new_new_n3025__ = ~new_new_n3022__ & new_new_n3024__;
  assign new_new_n3026__ = ~new_new_n3020__ & ~new_new_n3025__;
  assign new_new_n3027__ = ~pi044 & ~new_new_n3026__;
  assign new_new_n3028__ = ~new_new_n3016__ & ~new_new_n3027__;
  assign new_new_n3029__ = ~new_new_n3002__ & new_new_n3028__;
  assign new_new_n3030__ = ~new_new_n3001__ & ~new_new_n3029__;
  assign new_new_n3031__ = ~new_new_n2988__ & ~new_new_n3030__;
  assign new_new_n3032__ = ~new_new_n2987__ & ~new_new_n3031__;
  assign new_new_n3033__ = ~new_new_n2981__ & ~new_new_n3032__;
  assign new_new_n3034__ = ~new_new_n2980__ & ~new_new_n3033__;
  assign new_new_n3035__ = ~new_new_n2972__ & ~new_new_n3034__;
  assign new_new_n3036__ = ~new_new_n2971__ & ~new_new_n3035__;
  assign new_new_n3037__ = ~new_new_n2965__ & ~new_new_n3036__;
  assign new_new_n3038__ = ~new_new_n2964__ & ~new_new_n3037__;
  assign new_new_n3039__ = ~new_new_n2956__ & ~new_new_n3038__;
  assign new_new_n3040__ = ~new_new_n2955__ & ~new_new_n3039__;
  assign new_new_n3041__ = ~new_new_n2947__ & ~new_new_n3040__;
  assign new_new_n3042__ = ~new_new_n2946__ & ~new_new_n3041__;
  assign new_new_n3043__ = ~new_new_n2938__ & ~new_new_n3042__;
  assign new_new_n3044__ = ~new_new_n2937__ & ~new_new_n3043__;
  assign new_new_n3045__ = ~new_new_n2929__ & ~new_new_n3044__;
  assign new_new_n3046__ = ~new_new_n2928__ & ~new_new_n3045__;
  assign new_new_n3047__ = ~new_new_n2920__ & new_new_n3046__;
  assign new_new_n3048__ = ~new_new_n2919__ & ~new_new_n3047__;
  assign new_new_n3049__ = ~new_new_n2911__ & ~new_new_n3048__;
  assign new_new_n3050__ = ~new_new_n2910__ & ~new_new_n3049__;
  assign new_new_n3051__ = ~new_new_n2902__ & ~new_new_n3050__;
  assign new_new_n3052__ = ~new_new_n2901__ & ~new_new_n3051__;
  assign new_new_n3053__ = ~new_new_n2893__ & new_new_n3052__;
  assign new_new_n3054__ = ~new_new_n2892__ & ~new_new_n3053__;
  assign new_new_n3055__ = ~new_new_n2884__ & ~new_new_n3054__;
  assign new_new_n3056__ = ~new_new_n2883__ & ~new_new_n3055__;
  assign new_new_n3057__ = ~new_new_n2877__ & ~new_new_n3056__;
  assign new_new_n3058__ = ~new_new_n2876__ & ~new_new_n3057__;
  assign new_new_n3059__ = ~new_new_n2868__ & new_new_n3058__;
  assign new_new_n3060__ = ~new_new_n2867__ & ~new_new_n3059__;
  assign new_new_n3061__ = ~new_new_n2859__ & ~new_new_n3060__;
  assign new_new_n3062__ = ~new_new_n2858__ & ~new_new_n3061__;
  assign new_new_n3063__ = ~new_new_n2857__ & ~new_new_n3062__;
  assign new_new_n3064__ = ~new_new_n2856__ & ~new_new_n3063__;
  assign new_new_n3065__ = pi084 & new_new_n3064__;
  assign new_new_n3066__ = pi085 & ~new_new_n2836__;
  assign new_new_n3067__ = ~new_new_n3065__ & ~new_new_n3066__;
  assign new_new_n3068__ = ~new_new_n2817__ & ~new_new_n2818__;
  assign new_new_n3069__ = ~new_new_n2831__ & po043;
  assign new_new_n3070__ = ~pi083 & ~po043;
  assign new_new_n3071__ = ~new_new_n3069__ & ~new_new_n3070__;
  assign new_new_n3072__ = new_new_n3068__ & ~new_new_n3071__;
  assign new_new_n3073__ = ~new_new_n3068__ & new_new_n3071__;
  assign new_new_n3074__ = ~new_new_n3072__ & ~new_new_n3073__;
  assign new_new_n3075__ = ~pi084 & ~new_new_n3064__;
  assign new_new_n3076__ = ~new_new_n3074__ & ~new_new_n3075__;
  assign new_new_n3077__ = new_new_n3067__ & ~new_new_n3076__;
  assign new_new_n3078__ = ~new_new_n2848__ & ~new_new_n3077__;
  assign po042 = new_new_n297__ & ~new_new_n3078__;
  assign new_new_n3080__ = ~pi082 & ~new_new_n3060__;
  assign new_new_n3081__ = pi082 & new_new_n3060__;
  assign new_new_n3082__ = ~new_new_n3080__ & ~new_new_n3081__;
  assign new_new_n3083__ = po042 & new_new_n3082__;
  assign new_new_n3084__ = new_new_n2846__ & new_new_n3083__;
  assign new_new_n3085__ = ~new_new_n2846__ & ~new_new_n3083__;
  assign new_new_n3086__ = ~new_new_n3084__ & ~new_new_n3085__;
  assign new_new_n3087__ = ~pi083 & ~new_new_n3086__;
  assign new_new_n3088__ = pi083 & new_new_n3086__;
  assign new_new_n3089__ = ~new_new_n3087__ & ~new_new_n3088__;
  assign new_new_n3090__ = pi080 & ~new_new_n3056__;
  assign new_new_n3091__ = ~pi080 & new_new_n3056__;
  assign new_new_n3092__ = ~new_new_n3090__ & ~new_new_n3091__;
  assign new_new_n3093__ = po042 & new_new_n3092__;
  assign new_new_n3094__ = ~new_new_n2875__ & ~new_new_n3093__;
  assign new_new_n3095__ = new_new_n2875__ & new_new_n3093__;
  assign new_new_n3096__ = ~new_new_n3094__ & ~new_new_n3095__;
  assign new_new_n3097__ = pi081 & ~new_new_n3096__;
  assign new_new_n3098__ = ~pi081 & new_new_n3096__;
  assign new_new_n3099__ = ~new_new_n2883__ & ~new_new_n2884__;
  assign new_new_n3100__ = ~new_new_n3054__ & po042;
  assign new_new_n3101__ = pi079 & ~po042;
  assign new_new_n3102__ = ~new_new_n3100__ & ~new_new_n3101__;
  assign new_new_n3103__ = new_new_n3099__ & ~new_new_n3102__;
  assign new_new_n3104__ = ~new_new_n3099__ & new_new_n3102__;
  assign new_new_n3105__ = ~new_new_n3103__ & ~new_new_n3104__;
  assign new_new_n3106__ = ~pi080 & ~new_new_n3105__;
  assign new_new_n3107__ = pi080 & new_new_n3105__;
  assign new_new_n3108__ = ~new_new_n2892__ & ~new_new_n2893__;
  assign new_new_n3109__ = ~new_new_n3052__ & po042;
  assign new_new_n3110__ = ~pi078 & ~po042;
  assign new_new_n3111__ = ~new_new_n3109__ & ~new_new_n3110__;
  assign new_new_n3112__ = new_new_n3108__ & ~new_new_n3111__;
  assign new_new_n3113__ = ~new_new_n3108__ & new_new_n3111__;
  assign new_new_n3114__ = ~new_new_n3112__ & ~new_new_n3113__;
  assign new_new_n3115__ = pi079 & ~new_new_n3114__;
  assign new_new_n3116__ = ~pi079 & new_new_n3114__;
  assign new_new_n3117__ = ~new_new_n2901__ & ~new_new_n2902__;
  assign new_new_n3118__ = ~new_new_n3050__ & po042;
  assign new_new_n3119__ = ~pi077 & ~po042;
  assign new_new_n3120__ = ~new_new_n3118__ & ~new_new_n3119__;
  assign new_new_n3121__ = new_new_n3117__ & ~new_new_n3120__;
  assign new_new_n3122__ = ~new_new_n3117__ & new_new_n3120__;
  assign new_new_n3123__ = ~new_new_n3121__ & ~new_new_n3122__;
  assign new_new_n3124__ = pi078 & ~new_new_n3123__;
  assign new_new_n3125__ = ~pi078 & new_new_n3123__;
  assign new_new_n3126__ = ~pi076 & ~new_new_n3048__;
  assign new_new_n3127__ = pi076 & new_new_n3048__;
  assign new_new_n3128__ = ~new_new_n3126__ & ~new_new_n3127__;
  assign new_new_n3129__ = po042 & new_new_n3128__;
  assign new_new_n3130__ = new_new_n2909__ & new_new_n3129__;
  assign new_new_n3131__ = ~new_new_n2909__ & ~new_new_n3129__;
  assign new_new_n3132__ = ~new_new_n3130__ & ~new_new_n3131__;
  assign new_new_n3133__ = ~pi077 & ~new_new_n3132__;
  assign new_new_n3134__ = pi077 & new_new_n3132__;
  assign new_new_n3135__ = ~new_new_n3046__ & po042;
  assign new_new_n3136__ = pi075 & ~po042;
  assign new_new_n3137__ = ~new_new_n3135__ & ~new_new_n3136__;
  assign new_new_n3138__ = ~new_new_n2919__ & ~new_new_n2920__;
  assign new_new_n3139__ = ~new_new_n3137__ & new_new_n3138__;
  assign new_new_n3140__ = new_new_n3137__ & ~new_new_n3138__;
  assign new_new_n3141__ = ~new_new_n3139__ & ~new_new_n3140__;
  assign new_new_n3142__ = ~pi076 & ~new_new_n3141__;
  assign new_new_n3143__ = pi076 & new_new_n3141__;
  assign new_new_n3144__ = ~new_new_n3044__ & po042;
  assign new_new_n3145__ = pi074 & ~po042;
  assign new_new_n3146__ = ~new_new_n3144__ & ~new_new_n3145__;
  assign new_new_n3147__ = ~new_new_n2928__ & ~new_new_n2929__;
  assign new_new_n3148__ = ~new_new_n3146__ & new_new_n3147__;
  assign new_new_n3149__ = new_new_n3146__ & ~new_new_n3147__;
  assign new_new_n3150__ = ~new_new_n3148__ & ~new_new_n3149__;
  assign new_new_n3151__ = ~pi075 & ~new_new_n3150__;
  assign new_new_n3152__ = pi075 & new_new_n3150__;
  assign new_new_n3153__ = ~new_new_n2937__ & ~new_new_n2938__;
  assign new_new_n3154__ = new_new_n3042__ & po042;
  assign new_new_n3155__ = ~pi073 & ~po042;
  assign new_new_n3156__ = ~new_new_n3154__ & ~new_new_n3155__;
  assign new_new_n3157__ = ~new_new_n3153__ & ~new_new_n3156__;
  assign new_new_n3158__ = new_new_n3153__ & new_new_n3156__;
  assign new_new_n3159__ = ~new_new_n3157__ & ~new_new_n3158__;
  assign new_new_n3160__ = ~pi074 & ~new_new_n3159__;
  assign new_new_n3161__ = pi074 & new_new_n3159__;
  assign new_new_n3162__ = ~new_new_n2946__ & ~new_new_n2947__;
  assign new_new_n3163__ = ~new_new_n3040__ & po042;
  assign new_new_n3164__ = pi072 & ~po042;
  assign new_new_n3165__ = ~new_new_n3163__ & ~new_new_n3164__;
  assign new_new_n3166__ = new_new_n3162__ & new_new_n3165__;
  assign new_new_n3167__ = ~new_new_n3162__ & ~new_new_n3165__;
  assign new_new_n3168__ = ~new_new_n3166__ & ~new_new_n3167__;
  assign new_new_n3169__ = ~pi073 & new_new_n3168__;
  assign new_new_n3170__ = pi073 & ~new_new_n3168__;
  assign new_new_n3171__ = new_new_n3038__ & po042;
  assign new_new_n3172__ = ~pi071 & ~po042;
  assign new_new_n3173__ = ~new_new_n3171__ & ~new_new_n3172__;
  assign new_new_n3174__ = ~new_new_n2955__ & ~new_new_n2956__;
  assign new_new_n3175__ = ~new_new_n3173__ & ~new_new_n3174__;
  assign new_new_n3176__ = new_new_n3173__ & new_new_n3174__;
  assign new_new_n3177__ = ~new_new_n3175__ & ~new_new_n3176__;
  assign new_new_n3178__ = ~pi072 & ~new_new_n3177__;
  assign new_new_n3179__ = pi072 & new_new_n3177__;
  assign new_new_n3180__ = new_new_n3036__ & po042;
  assign new_new_n3181__ = ~pi070 & ~po042;
  assign new_new_n3182__ = ~new_new_n3180__ & ~new_new_n3181__;
  assign new_new_n3183__ = ~new_new_n2964__ & ~new_new_n2965__;
  assign new_new_n3184__ = ~new_new_n3182__ & ~new_new_n3183__;
  assign new_new_n3185__ = new_new_n3182__ & new_new_n3183__;
  assign new_new_n3186__ = ~new_new_n3184__ & ~new_new_n3185__;
  assign new_new_n3187__ = ~pi071 & ~new_new_n3186__;
  assign new_new_n3188__ = pi071 & new_new_n3186__;
  assign new_new_n3189__ = new_new_n3034__ & po042;
  assign new_new_n3190__ = ~pi069 & ~po042;
  assign new_new_n3191__ = ~new_new_n3189__ & ~new_new_n3190__;
  assign new_new_n3192__ = ~new_new_n2971__ & ~new_new_n2972__;
  assign new_new_n3193__ = ~new_new_n3191__ & ~new_new_n3192__;
  assign new_new_n3194__ = new_new_n3191__ & new_new_n3192__;
  assign new_new_n3195__ = ~new_new_n3193__ & ~new_new_n3194__;
  assign new_new_n3196__ = ~pi070 & ~new_new_n3195__;
  assign new_new_n3197__ = pi070 & new_new_n3195__;
  assign new_new_n3198__ = new_new_n3032__ & po042;
  assign new_new_n3199__ = ~pi068 & ~po042;
  assign new_new_n3200__ = ~new_new_n3198__ & ~new_new_n3199__;
  assign new_new_n3201__ = ~new_new_n2980__ & ~new_new_n2981__;
  assign new_new_n3202__ = ~new_new_n3200__ & ~new_new_n3201__;
  assign new_new_n3203__ = new_new_n3200__ & new_new_n3201__;
  assign new_new_n3204__ = ~new_new_n3202__ & ~new_new_n3203__;
  assign new_new_n3205__ = ~pi069 & ~new_new_n3204__;
  assign new_new_n3206__ = pi069 & new_new_n3204__;
  assign new_new_n3207__ = ~new_new_n3001__ & ~new_new_n3002__;
  assign new_new_n3208__ = po042 & new_new_n3207__;
  assign new_new_n3209__ = ~new_new_n3028__ & new_new_n3208__;
  assign new_new_n3210__ = new_new_n3028__ & ~new_new_n3208__;
  assign new_new_n3211__ = ~new_new_n3209__ & ~new_new_n3210__;
  assign new_new_n3212__ = pi067 & ~new_new_n3211__;
  assign new_new_n3213__ = ~pi067 & new_new_n3211__;
  assign new_new_n3214__ = pi042 & po042;
  assign new_new_n3215__ = ~pi042 & ~po042;
  assign new_new_n3216__ = ~pi065 & ~new_new_n3214__;
  assign new_new_n3217__ = ~new_new_n3215__ & new_new_n3216__;
  assign new_new_n3218__ = ~pi041 & ~new_new_n3217__;
  assign new_new_n3219__ = pi065 & new_new_n3214__;
  assign new_new_n3220__ = ~new_new_n3218__ & ~new_new_n3219__;
  assign new_new_n3221__ = pi064 & ~new_new_n3220__;
  assign new_new_n3222__ = pi064 & po042;
  assign new_new_n3223__ = ~pi042 & pi065;
  assign new_new_n3224__ = ~new_new_n3222__ & new_new_n3223__;
  assign new_new_n3225__ = ~new_new_n3221__ & ~new_new_n3224__;
  assign new_new_n3226__ = pi066 & ~new_new_n3225__;
  assign new_new_n3227__ = ~pi066 & new_new_n3225__;
  assign new_new_n3228__ = new_new_n426__ & ~po043;
  assign new_new_n3229__ = new_new_n3021__ & po042;
  assign new_new_n3230__ = ~new_new_n3228__ & ~new_new_n3229__;
  assign new_new_n3231__ = ~pi042 & ~new_new_n3230__;
  assign new_new_n3232__ = ~new_new_n332__ & po042;
  assign new_new_n3233__ = ~new_new_n2997__ & ~new_new_n3232__;
  assign new_new_n3234__ = pi065 & po042;
  assign new_new_n3235__ = po043 & ~new_new_n3234__;
  assign new_new_n3236__ = pi065 & ~new_new_n2997__;
  assign new_new_n3237__ = pi042 & ~new_new_n3236__;
  assign new_new_n3238__ = ~new_new_n3235__ & new_new_n3237__;
  assign new_new_n3239__ = ~new_new_n3231__ & ~new_new_n3233__;
  assign new_new_n3240__ = ~new_new_n3238__ & new_new_n3239__;
  assign new_new_n3241__ = pi043 & ~new_new_n3240__;
  assign new_new_n3242__ = ~pi064 & ~new_new_n3234__;
  assign new_new_n3243__ = ~pi065 & po042;
  assign new_new_n3244__ = ~po043 & ~new_new_n3243__;
  assign new_new_n3245__ = ~new_new_n3214__ & ~new_new_n3229__;
  assign new_new_n3246__ = ~new_new_n3244__ & new_new_n3245__;
  assign new_new_n3247__ = pi064 & ~new_new_n3246__;
  assign new_new_n3248__ = ~new_new_n3242__ & ~new_new_n3247__;
  assign new_new_n3249__ = ~new_new_n2997__ & ~new_new_n3234__;
  assign new_new_n3250__ = pi042 & ~new_new_n3009__;
  assign new_new_n3251__ = ~new_new_n3249__ & new_new_n3250__;
  assign new_new_n3252__ = ~new_new_n3248__ & ~new_new_n3251__;
  assign new_new_n3253__ = ~pi043 & ~new_new_n3252__;
  assign new_new_n3254__ = ~new_new_n3241__ & ~new_new_n3253__;
  assign new_new_n3255__ = ~new_new_n3227__ & new_new_n3254__;
  assign new_new_n3256__ = ~new_new_n3226__ & ~new_new_n3255__;
  assign new_new_n3257__ = ~new_new_n3213__ & ~new_new_n3256__;
  assign new_new_n3258__ = ~new_new_n3212__ & ~new_new_n3257__;
  assign new_new_n3259__ = pi068 & ~new_new_n3258__;
  assign new_new_n3260__ = ~pi068 & new_new_n3258__;
  assign new_new_n3261__ = ~new_new_n2987__ & ~new_new_n2988__;
  assign new_new_n3262__ = ~new_new_n3030__ & po042;
  assign new_new_n3263__ = pi067 & ~po042;
  assign new_new_n3264__ = ~new_new_n3262__ & ~new_new_n3263__;
  assign new_new_n3265__ = new_new_n3261__ & ~new_new_n3264__;
  assign new_new_n3266__ = ~new_new_n3261__ & new_new_n3264__;
  assign new_new_n3267__ = ~new_new_n3265__ & ~new_new_n3266__;
  assign new_new_n3268__ = ~new_new_n3260__ & new_new_n3267__;
  assign new_new_n3269__ = ~new_new_n3259__ & ~new_new_n3268__;
  assign new_new_n3270__ = ~new_new_n3206__ & new_new_n3269__;
  assign new_new_n3271__ = ~new_new_n3205__ & ~new_new_n3270__;
  assign new_new_n3272__ = ~new_new_n3197__ & ~new_new_n3271__;
  assign new_new_n3273__ = ~new_new_n3196__ & ~new_new_n3272__;
  assign new_new_n3274__ = ~new_new_n3188__ & ~new_new_n3273__;
  assign new_new_n3275__ = ~new_new_n3187__ & ~new_new_n3274__;
  assign new_new_n3276__ = ~new_new_n3179__ & ~new_new_n3275__;
  assign new_new_n3277__ = ~new_new_n3178__ & ~new_new_n3276__;
  assign new_new_n3278__ = ~new_new_n3170__ & ~new_new_n3277__;
  assign new_new_n3279__ = ~new_new_n3169__ & ~new_new_n3278__;
  assign new_new_n3280__ = ~new_new_n3161__ & ~new_new_n3279__;
  assign new_new_n3281__ = ~new_new_n3160__ & ~new_new_n3280__;
  assign new_new_n3282__ = ~new_new_n3152__ & ~new_new_n3281__;
  assign new_new_n3283__ = ~new_new_n3151__ & ~new_new_n3282__;
  assign new_new_n3284__ = ~new_new_n3143__ & ~new_new_n3283__;
  assign new_new_n3285__ = ~new_new_n3142__ & ~new_new_n3284__;
  assign new_new_n3286__ = ~new_new_n3134__ & ~new_new_n3285__;
  assign new_new_n3287__ = ~new_new_n3133__ & ~new_new_n3286__;
  assign new_new_n3288__ = ~new_new_n3125__ & new_new_n3287__;
  assign new_new_n3289__ = ~new_new_n3124__ & ~new_new_n3288__;
  assign new_new_n3290__ = ~new_new_n3116__ & ~new_new_n3289__;
  assign new_new_n3291__ = ~new_new_n3115__ & ~new_new_n3290__;
  assign new_new_n3292__ = ~new_new_n3107__ & new_new_n3291__;
  assign new_new_n3293__ = ~new_new_n3106__ & ~new_new_n3292__;
  assign new_new_n3294__ = ~new_new_n3098__ & new_new_n3293__;
  assign new_new_n3295__ = ~new_new_n3097__ & ~new_new_n3294__;
  assign new_new_n3296__ = ~pi082 & new_new_n3295__;
  assign new_new_n3297__ = pi082 & ~new_new_n3295__;
  assign new_new_n3298__ = ~new_new_n2867__ & ~new_new_n2868__;
  assign new_new_n3299__ = new_new_n3058__ & po042;
  assign new_new_n3300__ = ~pi081 & ~po042;
  assign new_new_n3301__ = ~new_new_n3299__ & ~new_new_n3300__;
  assign new_new_n3302__ = ~new_new_n3298__ & ~new_new_n3301__;
  assign new_new_n3303__ = new_new_n3298__ & new_new_n3301__;
  assign new_new_n3304__ = ~new_new_n3302__ & ~new_new_n3303__;
  assign new_new_n3305__ = ~new_new_n3297__ & ~new_new_n3304__;
  assign new_new_n3306__ = ~new_new_n3296__ & ~new_new_n3305__;
  assign new_new_n3307__ = new_new_n297__ & ~new_new_n3075__;
  assign new_new_n3308__ = new_new_n3067__ & new_new_n3307__;
  assign new_new_n3309__ = new_new_n3074__ & ~new_new_n3308__;
  assign new_new_n3310__ = new_new_n2159__ & new_new_n2847__;
  assign new_new_n3311__ = ~new_new_n3065__ & new_new_n3310__;
  assign new_new_n3312__ = new_new_n3076__ & new_new_n3311__;
  assign new_new_n3313__ = ~new_new_n3309__ & ~new_new_n3312__;
  assign new_new_n3314__ = pi085 & new_new_n3313__;
  assign new_new_n3315__ = ~pi085 & ~new_new_n3313__;
  assign new_new_n3316__ = ~new_new_n2856__ & ~new_new_n2857__;
  assign new_new_n3317__ = ~new_new_n3062__ & po042;
  assign new_new_n3318__ = ~pi083 & ~po042;
  assign new_new_n3319__ = ~new_new_n3317__ & ~new_new_n3318__;
  assign new_new_n3320__ = new_new_n3316__ & ~new_new_n3319__;
  assign new_new_n3321__ = ~new_new_n3316__ & new_new_n3319__;
  assign new_new_n3322__ = ~new_new_n3320__ & ~new_new_n3321__;
  assign new_new_n3323__ = pi084 & ~new_new_n3322__;
  assign new_new_n3324__ = ~pi084 & new_new_n3322__;
  assign new_new_n3325__ = ~new_new_n3088__ & ~new_new_n3306__;
  assign new_new_n3326__ = ~new_new_n3087__ & ~new_new_n3325__;
  assign new_new_n3327__ = ~new_new_n3324__ & new_new_n3326__;
  assign new_new_n3328__ = ~new_new_n3323__ & ~new_new_n3327__;
  assign new_new_n3329__ = ~new_new_n3315__ & ~new_new_n3328__;
  assign new_new_n3330__ = ~new_new_n3314__ & ~new_new_n3329__;
  assign new_new_n3331__ = pi086 & ~new_new_n3330__;
  assign new_new_n3332__ = ~pi095 & new_new_n289__;
  assign new_new_n3333__ = new_new_n292__ & new_new_n3332__;
  assign new_new_n3334__ = new_new_n258__ & new_new_n3333__;
  assign new_new_n3335__ = ~pi087 & new_new_n3334__;
  assign new_new_n3336__ = ~new_new_n3331__ & new_new_n3335__;
  assign new_new_n3337__ = ~pi086 & new_new_n3330__;
  assign new_new_n3338__ = new_new_n2847__ & ~po042;
  assign new_new_n3339__ = ~new_new_n376__ & ~new_new_n3338__;
  assign new_new_n3340__ = ~new_new_n3337__ & new_new_n3339__;
  assign po041 = new_new_n3336__ & ~new_new_n3340__;
  assign new_new_n3342__ = ~new_new_n3306__ & po041;
  assign new_new_n3343__ = ~pi083 & ~po041;
  assign new_new_n3344__ = ~new_new_n3342__ & ~new_new_n3343__;
  assign new_new_n3345__ = new_new_n3089__ & ~new_new_n3344__;
  assign new_new_n3346__ = ~new_new_n3089__ & new_new_n3344__;
  assign new_new_n3347__ = ~new_new_n3345__ & ~new_new_n3346__;
  assign new_new_n3348__ = ~pi084 & new_new_n3347__;
  assign new_new_n3349__ = pi084 & ~new_new_n3347__;
  assign new_new_n3350__ = ~new_new_n3348__ & ~new_new_n3349__;
  assign new_new_n3351__ = ~new_new_n3296__ & ~new_new_n3297__;
  assign new_new_n3352__ = po041 & new_new_n3351__;
  assign new_new_n3353__ = ~new_new_n3304__ & ~new_new_n3352__;
  assign new_new_n3354__ = new_new_n3304__ & new_new_n3352__;
  assign new_new_n3355__ = ~new_new_n3353__ & ~new_new_n3354__;
  assign new_new_n3356__ = ~pi083 & ~new_new_n3355__;
  assign new_new_n3357__ = pi083 & new_new_n3355__;
  assign new_new_n3358__ = new_new_n3293__ & po041;
  assign new_new_n3359__ = pi081 & ~po041;
  assign new_new_n3360__ = ~new_new_n3358__ & ~new_new_n3359__;
  assign new_new_n3361__ = ~new_new_n3097__ & ~new_new_n3098__;
  assign new_new_n3362__ = ~new_new_n3360__ & ~new_new_n3361__;
  assign new_new_n3363__ = new_new_n3360__ & new_new_n3361__;
  assign new_new_n3364__ = ~new_new_n3362__ & ~new_new_n3363__;
  assign new_new_n3365__ = ~pi082 & new_new_n3364__;
  assign new_new_n3366__ = pi082 & ~new_new_n3364__;
  assign new_new_n3367__ = ~new_new_n3106__ & ~new_new_n3107__;
  assign new_new_n3368__ = new_new_n3291__ & po041;
  assign new_new_n3369__ = ~pi080 & ~po041;
  assign new_new_n3370__ = ~new_new_n3368__ & ~new_new_n3369__;
  assign new_new_n3371__ = ~new_new_n3367__ & ~new_new_n3370__;
  assign new_new_n3372__ = new_new_n3367__ & new_new_n3370__;
  assign new_new_n3373__ = ~new_new_n3371__ & ~new_new_n3372__;
  assign new_new_n3374__ = ~pi081 & ~new_new_n3373__;
  assign new_new_n3375__ = pi081 & new_new_n3373__;
  assign new_new_n3376__ = pi079 & ~new_new_n3289__;
  assign new_new_n3377__ = ~pi079 & new_new_n3289__;
  assign new_new_n3378__ = ~new_new_n3376__ & ~new_new_n3377__;
  assign new_new_n3379__ = po041 & new_new_n3378__;
  assign new_new_n3380__ = new_new_n3114__ & new_new_n3379__;
  assign new_new_n3381__ = ~new_new_n3114__ & ~new_new_n3379__;
  assign new_new_n3382__ = ~new_new_n3380__ & ~new_new_n3381__;
  assign new_new_n3383__ = pi080 & ~new_new_n3382__;
  assign new_new_n3384__ = ~pi080 & new_new_n3382__;
  assign new_new_n3385__ = ~new_new_n3133__ & ~new_new_n3134__;
  assign new_new_n3386__ = ~new_new_n3285__ & po041;
  assign new_new_n3387__ = ~pi077 & ~po041;
  assign new_new_n3388__ = ~new_new_n3386__ & ~new_new_n3387__;
  assign new_new_n3389__ = ~new_new_n3385__ & ~new_new_n3388__;
  assign new_new_n3390__ = new_new_n3385__ & new_new_n3388__;
  assign new_new_n3391__ = ~new_new_n3389__ & ~new_new_n3390__;
  assign new_new_n3392__ = ~pi078 & ~new_new_n3391__;
  assign new_new_n3393__ = pi078 & new_new_n3391__;
  assign new_new_n3394__ = ~new_new_n3142__ & ~new_new_n3143__;
  assign new_new_n3395__ = ~new_new_n3283__ & po041;
  assign new_new_n3396__ = ~pi076 & ~po041;
  assign new_new_n3397__ = ~new_new_n3395__ & ~new_new_n3396__;
  assign new_new_n3398__ = ~new_new_n3394__ & ~new_new_n3397__;
  assign new_new_n3399__ = new_new_n3394__ & new_new_n3397__;
  assign new_new_n3400__ = ~new_new_n3398__ & ~new_new_n3399__;
  assign new_new_n3401__ = ~pi077 & ~new_new_n3400__;
  assign new_new_n3402__ = pi077 & new_new_n3400__;
  assign new_new_n3403__ = ~new_new_n3151__ & ~new_new_n3152__;
  assign new_new_n3404__ = ~new_new_n3281__ & po041;
  assign new_new_n3405__ = ~pi075 & ~po041;
  assign new_new_n3406__ = ~new_new_n3404__ & ~new_new_n3405__;
  assign new_new_n3407__ = ~new_new_n3403__ & ~new_new_n3406__;
  assign new_new_n3408__ = new_new_n3403__ & new_new_n3406__;
  assign new_new_n3409__ = ~new_new_n3407__ & ~new_new_n3408__;
  assign new_new_n3410__ = ~pi076 & ~new_new_n3409__;
  assign new_new_n3411__ = pi076 & new_new_n3409__;
  assign new_new_n3412__ = ~pi074 & ~new_new_n3279__;
  assign new_new_n3413__ = pi074 & new_new_n3279__;
  assign new_new_n3414__ = ~new_new_n3412__ & ~new_new_n3413__;
  assign new_new_n3415__ = po041 & new_new_n3414__;
  assign new_new_n3416__ = ~new_new_n3159__ & ~new_new_n3415__;
  assign new_new_n3417__ = new_new_n3159__ & new_new_n3415__;
  assign new_new_n3418__ = ~new_new_n3416__ & ~new_new_n3417__;
  assign new_new_n3419__ = pi075 & new_new_n3418__;
  assign new_new_n3420__ = ~pi075 & ~new_new_n3418__;
  assign new_new_n3421__ = new_new_n3277__ & po041;
  assign new_new_n3422__ = pi073 & ~po041;
  assign new_new_n3423__ = ~new_new_n3421__ & ~new_new_n3422__;
  assign new_new_n3424__ = ~new_new_n3169__ & ~new_new_n3170__;
  assign new_new_n3425__ = ~new_new_n3423__ & ~new_new_n3424__;
  assign new_new_n3426__ = new_new_n3423__ & new_new_n3424__;
  assign new_new_n3427__ = ~new_new_n3425__ & ~new_new_n3426__;
  assign new_new_n3428__ = pi074 & ~new_new_n3427__;
  assign new_new_n3429__ = ~pi074 & new_new_n3427__;
  assign new_new_n3430__ = ~new_new_n3178__ & ~new_new_n3179__;
  assign new_new_n3431__ = ~new_new_n3275__ & po041;
  assign new_new_n3432__ = ~pi072 & ~po041;
  assign new_new_n3433__ = ~new_new_n3431__ & ~new_new_n3432__;
  assign new_new_n3434__ = new_new_n3430__ & ~new_new_n3433__;
  assign new_new_n3435__ = ~new_new_n3430__ & new_new_n3433__;
  assign new_new_n3436__ = ~new_new_n3434__ & ~new_new_n3435__;
  assign new_new_n3437__ = pi073 & ~new_new_n3436__;
  assign new_new_n3438__ = ~pi073 & new_new_n3436__;
  assign new_new_n3439__ = ~new_new_n3187__ & ~new_new_n3188__;
  assign new_new_n3440__ = ~new_new_n3273__ & po041;
  assign new_new_n3441__ = ~pi071 & ~po041;
  assign new_new_n3442__ = ~new_new_n3440__ & ~new_new_n3441__;
  assign new_new_n3443__ = ~new_new_n3439__ & ~new_new_n3442__;
  assign new_new_n3444__ = new_new_n3439__ & new_new_n3442__;
  assign new_new_n3445__ = ~new_new_n3443__ & ~new_new_n3444__;
  assign new_new_n3446__ = pi072 & new_new_n3445__;
  assign new_new_n3447__ = ~pi072 & ~new_new_n3445__;
  assign new_new_n3448__ = ~new_new_n3196__ & ~new_new_n3197__;
  assign new_new_n3449__ = ~new_new_n3271__ & po041;
  assign new_new_n3450__ = ~pi070 & ~po041;
  assign new_new_n3451__ = ~new_new_n3449__ & ~new_new_n3450__;
  assign new_new_n3452__ = new_new_n3448__ & ~new_new_n3451__;
  assign new_new_n3453__ = ~new_new_n3448__ & new_new_n3451__;
  assign new_new_n3454__ = ~new_new_n3452__ & ~new_new_n3453__;
  assign new_new_n3455__ = pi071 & ~new_new_n3454__;
  assign new_new_n3456__ = ~pi071 & new_new_n3454__;
  assign new_new_n3457__ = ~new_new_n3205__ & ~new_new_n3206__;
  assign new_new_n3458__ = new_new_n3269__ & po041;
  assign new_new_n3459__ = ~pi069 & ~po041;
  assign new_new_n3460__ = ~new_new_n3458__ & ~new_new_n3459__;
  assign new_new_n3461__ = ~new_new_n3457__ & ~new_new_n3460__;
  assign new_new_n3462__ = new_new_n3457__ & new_new_n3460__;
  assign new_new_n3463__ = ~new_new_n3461__ & ~new_new_n3462__;
  assign new_new_n3464__ = ~pi070 & ~new_new_n3463__;
  assign new_new_n3465__ = pi070 & new_new_n3463__;
  assign new_new_n3466__ = ~new_new_n3259__ & ~new_new_n3260__;
  assign new_new_n3467__ = po041 & new_new_n3466__;
  assign new_new_n3468__ = ~new_new_n3267__ & ~new_new_n3467__;
  assign new_new_n3469__ = new_new_n3267__ & new_new_n3467__;
  assign new_new_n3470__ = ~new_new_n3468__ & ~new_new_n3469__;
  assign new_new_n3471__ = pi069 & new_new_n3470__;
  assign new_new_n3472__ = ~pi069 & ~new_new_n3470__;
  assign new_new_n3473__ = ~new_new_n3212__ & ~new_new_n3213__;
  assign new_new_n3474__ = ~new_new_n3256__ & po041;
  assign new_new_n3475__ = pi067 & ~po041;
  assign new_new_n3476__ = ~new_new_n3474__ & ~new_new_n3475__;
  assign new_new_n3477__ = new_new_n3473__ & ~new_new_n3476__;
  assign new_new_n3478__ = ~new_new_n3473__ & new_new_n3476__;
  assign new_new_n3479__ = ~new_new_n3477__ & ~new_new_n3478__;
  assign new_new_n3480__ = pi068 & new_new_n3479__;
  assign new_new_n3481__ = ~pi068 & ~new_new_n3479__;
  assign new_new_n3482__ = ~new_new_n3226__ & ~new_new_n3227__;
  assign new_new_n3483__ = po041 & new_new_n3482__;
  assign new_new_n3484__ = ~new_new_n3254__ & new_new_n3483__;
  assign new_new_n3485__ = new_new_n3254__ & ~new_new_n3483__;
  assign new_new_n3486__ = ~new_new_n3484__ & ~new_new_n3485__;
  assign new_new_n3487__ = pi067 & ~new_new_n3486__;
  assign new_new_n3488__ = ~pi067 & new_new_n3486__;
  assign new_new_n3489__ = pi041 & po041;
  assign new_new_n3490__ = pi040 & ~pi065;
  assign new_new_n3491__ = new_new_n3489__ & ~new_new_n3490__;
  assign new_new_n3492__ = ~pi041 & ~po041;
  assign new_new_n3493__ = ~pi065 & ~new_new_n3492__;
  assign new_new_n3494__ = ~pi040 & ~new_new_n3493__;
  assign new_new_n3495__ = ~new_new_n3491__ & ~new_new_n3494__;
  assign new_new_n3496__ = pi064 & ~new_new_n3495__;
  assign new_new_n3497__ = pi064 & po041;
  assign new_new_n3498__ = ~pi041 & pi065;
  assign new_new_n3499__ = ~new_new_n3497__ & new_new_n3498__;
  assign new_new_n3500__ = ~new_new_n3496__ & ~new_new_n3499__;
  assign new_new_n3501__ = ~pi066 & new_new_n3500__;
  assign new_new_n3502__ = pi066 & ~new_new_n3500__;
  assign new_new_n3503__ = new_new_n426__ & ~po042;
  assign new_new_n3504__ = new_new_n3243__ & po041;
  assign new_new_n3505__ = ~new_new_n3503__ & ~new_new_n3504__;
  assign new_new_n3506__ = ~pi041 & ~new_new_n3505__;
  assign new_new_n3507__ = ~new_new_n332__ & po041;
  assign new_new_n3508__ = ~new_new_n3222__ & ~new_new_n3507__;
  assign new_new_n3509__ = pi065 & po041;
  assign new_new_n3510__ = po042 & ~new_new_n3509__;
  assign new_new_n3511__ = pi065 & ~new_new_n3222__;
  assign new_new_n3512__ = pi041 & ~new_new_n3511__;
  assign new_new_n3513__ = ~new_new_n3510__ & new_new_n3512__;
  assign new_new_n3514__ = ~new_new_n3506__ & ~new_new_n3508__;
  assign new_new_n3515__ = ~new_new_n3513__ & new_new_n3514__;
  assign new_new_n3516__ = pi042 & ~new_new_n3515__;
  assign new_new_n3517__ = ~new_new_n3222__ & ~new_new_n3509__;
  assign new_new_n3518__ = pi041 & ~new_new_n3234__;
  assign new_new_n3519__ = pi064 & ~new_new_n3518__;
  assign new_new_n3520__ = ~new_new_n3517__ & ~new_new_n3519__;
  assign new_new_n3521__ = ~pi065 & po041;
  assign new_new_n3522__ = ~po042 & ~new_new_n3521__;
  assign new_new_n3523__ = pi064 & ~new_new_n3489__;
  assign new_new_n3524__ = ~new_new_n3504__ & new_new_n3523__;
  assign new_new_n3525__ = ~new_new_n3522__ & new_new_n3524__;
  assign new_new_n3526__ = ~new_new_n3520__ & ~new_new_n3525__;
  assign new_new_n3527__ = ~pi042 & ~new_new_n3526__;
  assign new_new_n3528__ = ~new_new_n3516__ & ~new_new_n3527__;
  assign new_new_n3529__ = ~new_new_n3502__ & ~new_new_n3528__;
  assign new_new_n3530__ = ~new_new_n3501__ & ~new_new_n3529__;
  assign new_new_n3531__ = ~new_new_n3488__ & new_new_n3530__;
  assign new_new_n3532__ = ~new_new_n3487__ & ~new_new_n3531__;
  assign new_new_n3533__ = ~new_new_n3481__ & ~new_new_n3532__;
  assign new_new_n3534__ = ~new_new_n3480__ & ~new_new_n3533__;
  assign new_new_n3535__ = ~new_new_n3472__ & ~new_new_n3534__;
  assign new_new_n3536__ = ~new_new_n3471__ & ~new_new_n3535__;
  assign new_new_n3537__ = ~new_new_n3465__ & new_new_n3536__;
  assign new_new_n3538__ = ~new_new_n3464__ & ~new_new_n3537__;
  assign new_new_n3539__ = ~new_new_n3456__ & new_new_n3538__;
  assign new_new_n3540__ = ~new_new_n3455__ & ~new_new_n3539__;
  assign new_new_n3541__ = ~new_new_n3447__ & ~new_new_n3540__;
  assign new_new_n3542__ = ~new_new_n3446__ & ~new_new_n3541__;
  assign new_new_n3543__ = ~new_new_n3438__ & ~new_new_n3542__;
  assign new_new_n3544__ = ~new_new_n3437__ & ~new_new_n3543__;
  assign new_new_n3545__ = ~new_new_n3429__ & ~new_new_n3544__;
  assign new_new_n3546__ = ~new_new_n3428__ & ~new_new_n3545__;
  assign new_new_n3547__ = ~new_new_n3420__ & ~new_new_n3546__;
  assign new_new_n3548__ = ~new_new_n3419__ & ~new_new_n3547__;
  assign new_new_n3549__ = ~new_new_n3411__ & new_new_n3548__;
  assign new_new_n3550__ = ~new_new_n3410__ & ~new_new_n3549__;
  assign new_new_n3551__ = ~new_new_n3402__ & ~new_new_n3550__;
  assign new_new_n3552__ = ~new_new_n3401__ & ~new_new_n3551__;
  assign new_new_n3553__ = ~new_new_n3393__ & ~new_new_n3552__;
  assign new_new_n3554__ = ~new_new_n3392__ & ~new_new_n3553__;
  assign new_new_n3555__ = pi079 & new_new_n3554__;
  assign new_new_n3556__ = ~pi079 & ~new_new_n3554__;
  assign new_new_n3557__ = ~new_new_n3124__ & ~new_new_n3125__;
  assign new_new_n3558__ = ~new_new_n3287__ & po041;
  assign new_new_n3559__ = ~pi078 & ~po041;
  assign new_new_n3560__ = ~new_new_n3558__ & ~new_new_n3559__;
  assign new_new_n3561__ = new_new_n3557__ & ~new_new_n3560__;
  assign new_new_n3562__ = ~new_new_n3557__ & new_new_n3560__;
  assign new_new_n3563__ = ~new_new_n3561__ & ~new_new_n3562__;
  assign new_new_n3564__ = ~new_new_n3556__ & ~new_new_n3563__;
  assign new_new_n3565__ = ~new_new_n3555__ & ~new_new_n3564__;
  assign new_new_n3566__ = ~new_new_n3384__ & ~new_new_n3565__;
  assign new_new_n3567__ = ~new_new_n3383__ & ~new_new_n3566__;
  assign new_new_n3568__ = ~new_new_n3375__ & new_new_n3567__;
  assign new_new_n3569__ = ~new_new_n3374__ & ~new_new_n3568__;
  assign new_new_n3570__ = ~new_new_n3366__ & ~new_new_n3569__;
  assign new_new_n3571__ = ~new_new_n3365__ & ~new_new_n3570__;
  assign new_new_n3572__ = ~new_new_n3357__ & ~new_new_n3571__;
  assign new_new_n3573__ = ~new_new_n3356__ & ~new_new_n3572__;
  assign new_new_n3574__ = ~new_new_n3336__ & new_new_n3338__;
  assign new_new_n3575__ = ~new_new_n376__ & ~new_new_n3574__;
  assign new_new_n3576__ = pi087 & new_new_n3575__;
  assign new_new_n3577__ = new_new_n3334__ & ~new_new_n3576__;
  assign new_new_n3578__ = ~new_new_n3314__ & ~new_new_n3315__;
  assign new_new_n3579__ = ~new_new_n3328__ & po041;
  assign new_new_n3580__ = pi085 & ~po041;
  assign new_new_n3581__ = ~new_new_n3579__ & ~new_new_n3580__;
  assign new_new_n3582__ = new_new_n3578__ & ~new_new_n3581__;
  assign new_new_n3583__ = ~new_new_n3578__ & new_new_n3581__;
  assign new_new_n3584__ = ~new_new_n3582__ & ~new_new_n3583__;
  assign new_new_n3585__ = pi086 & new_new_n3584__;
  assign new_new_n3586__ = ~pi086 & ~new_new_n3584__;
  assign new_new_n3587__ = ~new_new_n3323__ & ~new_new_n3324__;
  assign new_new_n3588__ = ~new_new_n3326__ & po041;
  assign new_new_n3589__ = ~pi084 & ~po041;
  assign new_new_n3590__ = ~new_new_n3588__ & ~new_new_n3589__;
  assign new_new_n3591__ = new_new_n3587__ & ~new_new_n3590__;
  assign new_new_n3592__ = ~new_new_n3587__ & new_new_n3590__;
  assign new_new_n3593__ = ~new_new_n3591__ & ~new_new_n3592__;
  assign new_new_n3594__ = pi085 & ~new_new_n3593__;
  assign new_new_n3595__ = ~pi085 & new_new_n3593__;
  assign new_new_n3596__ = ~new_new_n3349__ & ~new_new_n3573__;
  assign new_new_n3597__ = ~new_new_n3348__ & ~new_new_n3596__;
  assign new_new_n3598__ = ~new_new_n3595__ & new_new_n3597__;
  assign new_new_n3599__ = ~new_new_n3594__ & ~new_new_n3598__;
  assign new_new_n3600__ = ~new_new_n3586__ & ~new_new_n3599__;
  assign new_new_n3601__ = ~new_new_n3585__ & ~new_new_n3600__;
  assign new_new_n3602__ = ~pi087 & ~new_new_n3575__;
  assign new_new_n3603__ = ~new_new_n3601__ & ~new_new_n3602__;
  assign po040 = new_new_n3577__ & ~new_new_n3603__;
  assign new_new_n3605__ = ~new_new_n3573__ & po040;
  assign new_new_n3606__ = ~pi084 & ~po040;
  assign new_new_n3607__ = ~new_new_n3605__ & ~new_new_n3606__;
  assign new_new_n3608__ = new_new_n3350__ & ~new_new_n3607__;
  assign new_new_n3609__ = ~new_new_n3350__ & new_new_n3607__;
  assign new_new_n3610__ = ~new_new_n3608__ & ~new_new_n3609__;
  assign new_new_n3611__ = pi087 & ~new_new_n3601__;
  assign new_new_n3612__ = new_new_n3334__ & ~new_new_n3611__;
  assign new_new_n3613__ = ~new_new_n3575__ & ~new_new_n3612__;
  assign new_new_n3614__ = ~pi088 & new_new_n3613__;
  assign new_new_n3615__ = pi088 & ~new_new_n3613__;
  assign new_new_n3616__ = ~new_new_n3594__ & ~new_new_n3595__;
  assign new_new_n3617__ = ~new_new_n3597__ & po040;
  assign new_new_n3618__ = ~pi085 & ~po040;
  assign new_new_n3619__ = ~new_new_n3617__ & ~new_new_n3618__;
  assign new_new_n3620__ = new_new_n3616__ & ~new_new_n3619__;
  assign new_new_n3621__ = ~new_new_n3616__ & new_new_n3619__;
  assign new_new_n3622__ = ~new_new_n3620__ & ~new_new_n3621__;
  assign new_new_n3623__ = pi086 & ~new_new_n3622__;
  assign new_new_n3624__ = ~pi086 & new_new_n3622__;
  assign new_new_n3625__ = pi085 & ~new_new_n3610__;
  assign new_new_n3626__ = ~pi085 & new_new_n3610__;
  assign new_new_n3627__ = ~new_new_n3356__ & ~new_new_n3357__;
  assign new_new_n3628__ = ~new_new_n3571__ & po040;
  assign new_new_n3629__ = ~pi083 & ~po040;
  assign new_new_n3630__ = ~new_new_n3628__ & ~new_new_n3629__;
  assign new_new_n3631__ = new_new_n3627__ & ~new_new_n3630__;
  assign new_new_n3632__ = ~new_new_n3627__ & new_new_n3630__;
  assign new_new_n3633__ = ~new_new_n3631__ & ~new_new_n3632__;
  assign new_new_n3634__ = pi084 & ~new_new_n3633__;
  assign new_new_n3635__ = ~pi084 & new_new_n3633__;
  assign new_new_n3636__ = ~new_new_n3365__ & ~new_new_n3366__;
  assign new_new_n3637__ = ~new_new_n3569__ & po040;
  assign new_new_n3638__ = ~pi082 & ~po040;
  assign new_new_n3639__ = ~new_new_n3637__ & ~new_new_n3638__;
  assign new_new_n3640__ = new_new_n3636__ & new_new_n3639__;
  assign new_new_n3641__ = ~new_new_n3636__ & ~new_new_n3639__;
  assign new_new_n3642__ = ~new_new_n3640__ & ~new_new_n3641__;
  assign new_new_n3643__ = ~pi083 & ~new_new_n3642__;
  assign new_new_n3644__ = pi083 & new_new_n3642__;
  assign new_new_n3645__ = new_new_n3567__ & po040;
  assign new_new_n3646__ = ~pi081 & ~po040;
  assign new_new_n3647__ = ~new_new_n3645__ & ~new_new_n3646__;
  assign new_new_n3648__ = ~new_new_n3374__ & ~new_new_n3375__;
  assign new_new_n3649__ = ~new_new_n3647__ & ~new_new_n3648__;
  assign new_new_n3650__ = new_new_n3647__ & new_new_n3648__;
  assign new_new_n3651__ = ~new_new_n3649__ & ~new_new_n3650__;
  assign new_new_n3652__ = ~pi082 & ~new_new_n3651__;
  assign new_new_n3653__ = pi082 & new_new_n3651__;
  assign new_new_n3654__ = ~new_new_n3383__ & ~new_new_n3384__;
  assign new_new_n3655__ = ~new_new_n3565__ & po040;
  assign new_new_n3656__ = pi080 & ~po040;
  assign new_new_n3657__ = ~new_new_n3655__ & ~new_new_n3656__;
  assign new_new_n3658__ = new_new_n3654__ & ~new_new_n3657__;
  assign new_new_n3659__ = ~new_new_n3654__ & new_new_n3657__;
  assign new_new_n3660__ = ~new_new_n3658__ & ~new_new_n3659__;
  assign new_new_n3661__ = ~pi081 & ~new_new_n3660__;
  assign new_new_n3662__ = pi081 & new_new_n3660__;
  assign new_new_n3663__ = ~new_new_n3555__ & ~new_new_n3556__;
  assign new_new_n3664__ = po040 & new_new_n3663__;
  assign new_new_n3665__ = new_new_n3563__ & new_new_n3664__;
  assign new_new_n3666__ = ~new_new_n3563__ & ~new_new_n3664__;
  assign new_new_n3667__ = ~new_new_n3665__ & ~new_new_n3666__;
  assign new_new_n3668__ = pi080 & ~new_new_n3667__;
  assign new_new_n3669__ = ~pi080 & new_new_n3667__;
  assign new_new_n3670__ = ~pi078 & ~new_new_n3552__;
  assign new_new_n3671__ = pi078 & new_new_n3552__;
  assign new_new_n3672__ = ~new_new_n3670__ & ~new_new_n3671__;
  assign new_new_n3673__ = po040 & new_new_n3672__;
  assign new_new_n3674__ = ~new_new_n3391__ & new_new_n3673__;
  assign new_new_n3675__ = new_new_n3391__ & ~new_new_n3673__;
  assign new_new_n3676__ = ~new_new_n3674__ & ~new_new_n3675__;
  assign new_new_n3677__ = pi079 & ~new_new_n3676__;
  assign new_new_n3678__ = ~pi079 & new_new_n3676__;
  assign new_new_n3679__ = ~pi077 & ~new_new_n3550__;
  assign new_new_n3680__ = pi077 & new_new_n3550__;
  assign new_new_n3681__ = ~new_new_n3679__ & ~new_new_n3680__;
  assign new_new_n3682__ = po040 & new_new_n3681__;
  assign new_new_n3683__ = ~new_new_n3400__ & new_new_n3682__;
  assign new_new_n3684__ = new_new_n3400__ & ~new_new_n3682__;
  assign new_new_n3685__ = ~new_new_n3683__ & ~new_new_n3684__;
  assign new_new_n3686__ = pi078 & ~new_new_n3685__;
  assign new_new_n3687__ = ~pi078 & new_new_n3685__;
  assign new_new_n3688__ = ~new_new_n3410__ & ~new_new_n3411__;
  assign new_new_n3689__ = ~new_new_n3548__ & po040;
  assign new_new_n3690__ = pi076 & ~po040;
  assign new_new_n3691__ = ~new_new_n3689__ & ~new_new_n3690__;
  assign new_new_n3692__ = new_new_n3688__ & ~new_new_n3691__;
  assign new_new_n3693__ = ~new_new_n3688__ & new_new_n3691__;
  assign new_new_n3694__ = ~new_new_n3692__ & ~new_new_n3693__;
  assign new_new_n3695__ = ~pi077 & ~new_new_n3694__;
  assign new_new_n3696__ = pi077 & new_new_n3694__;
  assign new_new_n3697__ = ~new_new_n3419__ & ~new_new_n3420__;
  assign new_new_n3698__ = new_new_n3546__ & po040;
  assign new_new_n3699__ = ~pi075 & ~po040;
  assign new_new_n3700__ = ~new_new_n3698__ & ~new_new_n3699__;
  assign new_new_n3701__ = ~new_new_n3697__ & ~new_new_n3700__;
  assign new_new_n3702__ = new_new_n3697__ & new_new_n3700__;
  assign new_new_n3703__ = ~new_new_n3701__ & ~new_new_n3702__;
  assign new_new_n3704__ = ~pi076 & ~new_new_n3703__;
  assign new_new_n3705__ = pi076 & new_new_n3703__;
  assign new_new_n3706__ = pi074 & ~new_new_n3544__;
  assign new_new_n3707__ = ~pi074 & new_new_n3544__;
  assign new_new_n3708__ = ~new_new_n3706__ & ~new_new_n3707__;
  assign new_new_n3709__ = po040 & new_new_n3708__;
  assign new_new_n3710__ = new_new_n3427__ & new_new_n3709__;
  assign new_new_n3711__ = ~new_new_n3427__ & ~new_new_n3709__;
  assign new_new_n3712__ = ~new_new_n3710__ & ~new_new_n3711__;
  assign new_new_n3713__ = pi075 & ~new_new_n3712__;
  assign new_new_n3714__ = ~pi075 & new_new_n3712__;
  assign new_new_n3715__ = ~new_new_n3542__ & po040;
  assign new_new_n3716__ = pi073 & ~po040;
  assign new_new_n3717__ = ~new_new_n3715__ & ~new_new_n3716__;
  assign new_new_n3718__ = ~new_new_n3437__ & ~new_new_n3438__;
  assign new_new_n3719__ = ~new_new_n3717__ & new_new_n3718__;
  assign new_new_n3720__ = new_new_n3717__ & ~new_new_n3718__;
  assign new_new_n3721__ = ~new_new_n3719__ & ~new_new_n3720__;
  assign new_new_n3722__ = ~pi074 & ~new_new_n3721__;
  assign new_new_n3723__ = pi074 & new_new_n3721__;
  assign new_new_n3724__ = ~new_new_n3540__ & po040;
  assign new_new_n3725__ = pi072 & ~po040;
  assign new_new_n3726__ = ~new_new_n3724__ & ~new_new_n3725__;
  assign new_new_n3727__ = ~new_new_n3446__ & ~new_new_n3447__;
  assign new_new_n3728__ = ~new_new_n3726__ & new_new_n3727__;
  assign new_new_n3729__ = new_new_n3726__ & ~new_new_n3727__;
  assign new_new_n3730__ = ~new_new_n3728__ & ~new_new_n3729__;
  assign new_new_n3731__ = ~pi073 & ~new_new_n3730__;
  assign new_new_n3732__ = pi073 & new_new_n3730__;
  assign new_new_n3733__ = ~new_new_n3455__ & ~new_new_n3456__;
  assign new_new_n3734__ = ~new_new_n3538__ & po040;
  assign new_new_n3735__ = ~pi071 & ~po040;
  assign new_new_n3736__ = ~new_new_n3734__ & ~new_new_n3735__;
  assign new_new_n3737__ = new_new_n3733__ & new_new_n3736__;
  assign new_new_n3738__ = ~new_new_n3733__ & ~new_new_n3736__;
  assign new_new_n3739__ = ~new_new_n3737__ & ~new_new_n3738__;
  assign new_new_n3740__ = ~pi072 & ~new_new_n3739__;
  assign new_new_n3741__ = pi072 & new_new_n3739__;
  assign new_new_n3742__ = new_new_n3536__ & po040;
  assign new_new_n3743__ = ~pi070 & ~po040;
  assign new_new_n3744__ = ~new_new_n3742__ & ~new_new_n3743__;
  assign new_new_n3745__ = ~new_new_n3464__ & ~new_new_n3465__;
  assign new_new_n3746__ = ~new_new_n3744__ & ~new_new_n3745__;
  assign new_new_n3747__ = new_new_n3744__ & new_new_n3745__;
  assign new_new_n3748__ = ~new_new_n3746__ & ~new_new_n3747__;
  assign new_new_n3749__ = ~pi071 & ~new_new_n3748__;
  assign new_new_n3750__ = pi071 & new_new_n3748__;
  assign new_new_n3751__ = ~new_new_n3471__ & ~new_new_n3472__;
  assign new_new_n3752__ = new_new_n3534__ & po040;
  assign new_new_n3753__ = ~pi069 & ~po040;
  assign new_new_n3754__ = ~new_new_n3752__ & ~new_new_n3753__;
  assign new_new_n3755__ = ~new_new_n3751__ & ~new_new_n3754__;
  assign new_new_n3756__ = new_new_n3751__ & new_new_n3754__;
  assign new_new_n3757__ = ~new_new_n3755__ & ~new_new_n3756__;
  assign new_new_n3758__ = ~pi070 & ~new_new_n3757__;
  assign new_new_n3759__ = pi070 & new_new_n3757__;
  assign new_new_n3760__ = new_new_n3532__ & po040;
  assign new_new_n3761__ = ~pi068 & ~po040;
  assign new_new_n3762__ = ~new_new_n3760__ & ~new_new_n3761__;
  assign new_new_n3763__ = ~new_new_n3480__ & ~new_new_n3481__;
  assign new_new_n3764__ = ~new_new_n3762__ & ~new_new_n3763__;
  assign new_new_n3765__ = new_new_n3762__ & new_new_n3763__;
  assign new_new_n3766__ = ~new_new_n3764__ & ~new_new_n3765__;
  assign new_new_n3767__ = ~pi069 & ~new_new_n3766__;
  assign new_new_n3768__ = pi069 & new_new_n3766__;
  assign new_new_n3769__ = new_new_n3530__ & po040;
  assign new_new_n3770__ = pi067 & ~po040;
  assign new_new_n3771__ = ~new_new_n3769__ & ~new_new_n3770__;
  assign new_new_n3772__ = ~new_new_n3487__ & ~new_new_n3488__;
  assign new_new_n3773__ = ~new_new_n3771__ & ~new_new_n3772__;
  assign new_new_n3774__ = new_new_n3771__ & new_new_n3772__;
  assign new_new_n3775__ = ~new_new_n3773__ & ~new_new_n3774__;
  assign new_new_n3776__ = pi068 & ~new_new_n3775__;
  assign new_new_n3777__ = ~pi068 & new_new_n3775__;
  assign new_new_n3778__ = ~new_new_n3501__ & ~new_new_n3502__;
  assign new_new_n3779__ = po040 & new_new_n3778__;
  assign new_new_n3780__ = ~new_new_n3528__ & new_new_n3779__;
  assign new_new_n3781__ = new_new_n3528__ & ~new_new_n3779__;
  assign new_new_n3782__ = ~new_new_n3780__ & ~new_new_n3781__;
  assign new_new_n3783__ = pi067 & ~new_new_n3782__;
  assign new_new_n3784__ = ~pi067 & new_new_n3782__;
  assign new_new_n3785__ = pi040 & po040;
  assign new_new_n3786__ = pi039 & ~pi065;
  assign new_new_n3787__ = new_new_n3785__ & ~new_new_n3786__;
  assign new_new_n3788__ = ~pi040 & ~po040;
  assign new_new_n3789__ = ~pi065 & ~new_new_n3788__;
  assign new_new_n3790__ = ~pi039 & ~new_new_n3789__;
  assign new_new_n3791__ = ~new_new_n3787__ & ~new_new_n3790__;
  assign new_new_n3792__ = pi064 & ~new_new_n3791__;
  assign new_new_n3793__ = pi064 & po040;
  assign new_new_n3794__ = ~pi040 & pi065;
  assign new_new_n3795__ = ~new_new_n3793__ & new_new_n3794__;
  assign new_new_n3796__ = ~new_new_n3792__ & ~new_new_n3795__;
  assign new_new_n3797__ = pi066 & ~new_new_n3796__;
  assign new_new_n3798__ = ~pi066 & new_new_n3796__;
  assign new_new_n3799__ = new_new_n426__ & ~po041;
  assign new_new_n3800__ = new_new_n3521__ & po040;
  assign new_new_n3801__ = ~new_new_n3799__ & ~new_new_n3800__;
  assign new_new_n3802__ = ~pi040 & ~new_new_n3801__;
  assign new_new_n3803__ = ~new_new_n332__ & po040;
  assign new_new_n3804__ = ~new_new_n3497__ & ~new_new_n3803__;
  assign new_new_n3805__ = pi065 & po040;
  assign new_new_n3806__ = po041 & ~new_new_n3805__;
  assign new_new_n3807__ = pi065 & ~new_new_n3497__;
  assign new_new_n3808__ = pi040 & ~new_new_n3807__;
  assign new_new_n3809__ = ~new_new_n3806__ & new_new_n3808__;
  assign new_new_n3810__ = ~new_new_n3802__ & ~new_new_n3804__;
  assign new_new_n3811__ = ~new_new_n3809__ & new_new_n3810__;
  assign new_new_n3812__ = pi041 & ~new_new_n3811__;
  assign new_new_n3813__ = ~new_new_n3497__ & ~new_new_n3805__;
  assign new_new_n3814__ = pi040 & ~new_new_n3509__;
  assign new_new_n3815__ = pi064 & ~new_new_n3814__;
  assign new_new_n3816__ = ~new_new_n3813__ & ~new_new_n3815__;
  assign new_new_n3817__ = ~pi065 & po040;
  assign new_new_n3818__ = ~po041 & ~new_new_n3817__;
  assign new_new_n3819__ = pi064 & ~new_new_n3785__;
  assign new_new_n3820__ = ~new_new_n3800__ & new_new_n3819__;
  assign new_new_n3821__ = ~new_new_n3818__ & new_new_n3820__;
  assign new_new_n3822__ = ~new_new_n3816__ & ~new_new_n3821__;
  assign new_new_n3823__ = ~pi041 & ~new_new_n3822__;
  assign new_new_n3824__ = ~new_new_n3812__ & ~new_new_n3823__;
  assign new_new_n3825__ = ~new_new_n3798__ & new_new_n3824__;
  assign new_new_n3826__ = ~new_new_n3797__ & ~new_new_n3825__;
  assign new_new_n3827__ = ~new_new_n3784__ & ~new_new_n3826__;
  assign new_new_n3828__ = ~new_new_n3783__ & ~new_new_n3827__;
  assign new_new_n3829__ = ~new_new_n3777__ & ~new_new_n3828__;
  assign new_new_n3830__ = ~new_new_n3776__ & ~new_new_n3829__;
  assign new_new_n3831__ = ~new_new_n3768__ & new_new_n3830__;
  assign new_new_n3832__ = ~new_new_n3767__ & ~new_new_n3831__;
  assign new_new_n3833__ = ~new_new_n3759__ & ~new_new_n3832__;
  assign new_new_n3834__ = ~new_new_n3758__ & ~new_new_n3833__;
  assign new_new_n3835__ = ~new_new_n3750__ & ~new_new_n3834__;
  assign new_new_n3836__ = ~new_new_n3749__ & ~new_new_n3835__;
  assign new_new_n3837__ = ~new_new_n3741__ & ~new_new_n3836__;
  assign new_new_n3838__ = ~new_new_n3740__ & ~new_new_n3837__;
  assign new_new_n3839__ = ~new_new_n3732__ & ~new_new_n3838__;
  assign new_new_n3840__ = ~new_new_n3731__ & ~new_new_n3839__;
  assign new_new_n3841__ = ~new_new_n3723__ & ~new_new_n3840__;
  assign new_new_n3842__ = ~new_new_n3722__ & ~new_new_n3841__;
  assign new_new_n3843__ = ~new_new_n3714__ & new_new_n3842__;
  assign new_new_n3844__ = ~new_new_n3713__ & ~new_new_n3843__;
  assign new_new_n3845__ = ~new_new_n3705__ & new_new_n3844__;
  assign new_new_n3846__ = ~new_new_n3704__ & ~new_new_n3845__;
  assign new_new_n3847__ = ~new_new_n3696__ & ~new_new_n3846__;
  assign new_new_n3848__ = ~new_new_n3695__ & ~new_new_n3847__;
  assign new_new_n3849__ = ~new_new_n3687__ & new_new_n3848__;
  assign new_new_n3850__ = ~new_new_n3686__ & ~new_new_n3849__;
  assign new_new_n3851__ = ~new_new_n3678__ & ~new_new_n3850__;
  assign new_new_n3852__ = ~new_new_n3677__ & ~new_new_n3851__;
  assign new_new_n3853__ = ~new_new_n3669__ & ~new_new_n3852__;
  assign new_new_n3854__ = ~new_new_n3668__ & ~new_new_n3853__;
  assign new_new_n3855__ = ~new_new_n3662__ & new_new_n3854__;
  assign new_new_n3856__ = ~new_new_n3661__ & ~new_new_n3855__;
  assign new_new_n3857__ = ~new_new_n3653__ & ~new_new_n3856__;
  assign new_new_n3858__ = ~new_new_n3652__ & ~new_new_n3857__;
  assign new_new_n3859__ = ~new_new_n3644__ & ~new_new_n3858__;
  assign new_new_n3860__ = ~new_new_n3643__ & ~new_new_n3859__;
  assign new_new_n3861__ = ~new_new_n3635__ & new_new_n3860__;
  assign new_new_n3862__ = ~new_new_n3634__ & ~new_new_n3861__;
  assign new_new_n3863__ = ~new_new_n3626__ & ~new_new_n3862__;
  assign new_new_n3864__ = ~new_new_n3625__ & ~new_new_n3863__;
  assign new_new_n3865__ = ~new_new_n3624__ & ~new_new_n3864__;
  assign new_new_n3866__ = ~new_new_n3623__ & ~new_new_n3865__;
  assign new_new_n3867__ = pi087 & ~new_new_n3866__;
  assign new_new_n3868__ = ~new_new_n3615__ & ~new_new_n3867__;
  assign new_new_n3869__ = ~pi087 & new_new_n3866__;
  assign new_new_n3870__ = pi086 & new_new_n3599__;
  assign new_new_n3871__ = ~pi086 & ~new_new_n3599__;
  assign new_new_n3872__ = ~new_new_n3870__ & ~new_new_n3871__;
  assign new_new_n3873__ = new_new_n3577__ & ~new_new_n3872__;
  assign new_new_n3874__ = ~new_new_n3584__ & ~new_new_n3873__;
  assign new_new_n3875__ = new_new_n3334__ & new_new_n3602__;
  assign new_new_n3876__ = new_new_n3584__ & new_new_n3875__;
  assign new_new_n3877__ = ~new_new_n3872__ & new_new_n3876__;
  assign new_new_n3878__ = ~new_new_n3874__ & ~new_new_n3877__;
  assign new_new_n3879__ = ~new_new_n3869__ & new_new_n3878__;
  assign new_new_n3880__ = new_new_n3868__ & ~new_new_n3879__;
  assign new_new_n3881__ = ~new_new_n3614__ & ~new_new_n3880__;
  assign new_new_n3882__ = new_new_n257__ & new_new_n294__;
  assign po039 = ~new_new_n3881__ & new_new_n3882__;
  assign new_new_n3884__ = pi085 & ~new_new_n3862__;
  assign new_new_n3885__ = ~pi085 & new_new_n3862__;
  assign new_new_n3886__ = ~new_new_n3884__ & ~new_new_n3885__;
  assign new_new_n3887__ = po039 & new_new_n3886__;
  assign new_new_n3888__ = new_new_n3610__ & new_new_n3887__;
  assign new_new_n3889__ = ~new_new_n3610__ & ~new_new_n3887__;
  assign new_new_n3890__ = ~new_new_n3888__ & ~new_new_n3889__;
  assign new_new_n3891__ = pi086 & ~new_new_n3890__;
  assign new_new_n3892__ = ~pi086 & new_new_n3890__;
  assign new_new_n3893__ = ~new_new_n3891__ & ~new_new_n3892__;
  assign new_new_n3894__ = ~new_new_n3634__ & ~new_new_n3635__;
  assign new_new_n3895__ = ~new_new_n3860__ & po039;
  assign new_new_n3896__ = ~pi084 & ~po039;
  assign new_new_n3897__ = ~new_new_n3895__ & ~new_new_n3896__;
  assign new_new_n3898__ = new_new_n3894__ & ~new_new_n3897__;
  assign new_new_n3899__ = ~new_new_n3894__ & new_new_n3897__;
  assign new_new_n3900__ = ~new_new_n3898__ & ~new_new_n3899__;
  assign new_new_n3901__ = pi085 & ~new_new_n3900__;
  assign new_new_n3902__ = ~pi085 & new_new_n3900__;
  assign new_new_n3903__ = ~pi083 & ~new_new_n3858__;
  assign new_new_n3904__ = pi083 & new_new_n3858__;
  assign new_new_n3905__ = ~new_new_n3903__ & ~new_new_n3904__;
  assign new_new_n3906__ = po039 & new_new_n3905__;
  assign new_new_n3907__ = new_new_n3642__ & new_new_n3906__;
  assign new_new_n3908__ = ~new_new_n3642__ & ~new_new_n3906__;
  assign new_new_n3909__ = ~new_new_n3907__ & ~new_new_n3908__;
  assign new_new_n3910__ = pi084 & new_new_n3909__;
  assign new_new_n3911__ = ~pi084 & ~new_new_n3909__;
  assign new_new_n3912__ = ~new_new_n3652__ & ~new_new_n3653__;
  assign new_new_n3913__ = ~new_new_n3856__ & po039;
  assign new_new_n3914__ = ~pi082 & ~po039;
  assign new_new_n3915__ = ~new_new_n3913__ & ~new_new_n3914__;
  assign new_new_n3916__ = new_new_n3912__ & ~new_new_n3915__;
  assign new_new_n3917__ = ~new_new_n3912__ & new_new_n3915__;
  assign new_new_n3918__ = ~new_new_n3916__ & ~new_new_n3917__;
  assign new_new_n3919__ = pi083 & ~new_new_n3918__;
  assign new_new_n3920__ = ~pi083 & new_new_n3918__;
  assign new_new_n3921__ = ~new_new_n3661__ & ~new_new_n3662__;
  assign new_new_n3922__ = ~new_new_n3854__ & po039;
  assign new_new_n3923__ = pi081 & ~po039;
  assign new_new_n3924__ = ~new_new_n3922__ & ~new_new_n3923__;
  assign new_new_n3925__ = new_new_n3921__ & ~new_new_n3924__;
  assign new_new_n3926__ = ~new_new_n3921__ & new_new_n3924__;
  assign new_new_n3927__ = ~new_new_n3925__ & ~new_new_n3926__;
  assign new_new_n3928__ = pi082 & new_new_n3927__;
  assign new_new_n3929__ = ~pi082 & ~new_new_n3927__;
  assign new_new_n3930__ = ~new_new_n3668__ & ~new_new_n3669__;
  assign new_new_n3931__ = ~new_new_n3852__ & po039;
  assign new_new_n3932__ = pi080 & ~po039;
  assign new_new_n3933__ = ~new_new_n3931__ & ~new_new_n3932__;
  assign new_new_n3934__ = new_new_n3930__ & new_new_n3933__;
  assign new_new_n3935__ = ~new_new_n3930__ & ~new_new_n3933__;
  assign new_new_n3936__ = ~new_new_n3934__ & ~new_new_n3935__;
  assign new_new_n3937__ = pi081 & ~new_new_n3936__;
  assign new_new_n3938__ = ~pi081 & new_new_n3936__;
  assign new_new_n3939__ = pi079 & ~new_new_n3850__;
  assign new_new_n3940__ = ~pi079 & new_new_n3850__;
  assign new_new_n3941__ = ~new_new_n3939__ & ~new_new_n3940__;
  assign new_new_n3942__ = po039 & new_new_n3941__;
  assign new_new_n3943__ = new_new_n3676__ & new_new_n3942__;
  assign new_new_n3944__ = ~new_new_n3676__ & ~new_new_n3942__;
  assign new_new_n3945__ = ~new_new_n3943__ & ~new_new_n3944__;
  assign new_new_n3946__ = pi080 & ~new_new_n3945__;
  assign new_new_n3947__ = ~pi080 & new_new_n3945__;
  assign new_new_n3948__ = new_new_n3848__ & po039;
  assign new_new_n3949__ = pi078 & ~po039;
  assign new_new_n3950__ = ~new_new_n3948__ & ~new_new_n3949__;
  assign new_new_n3951__ = ~new_new_n3686__ & ~new_new_n3687__;
  assign new_new_n3952__ = ~new_new_n3950__ & ~new_new_n3951__;
  assign new_new_n3953__ = new_new_n3950__ & new_new_n3951__;
  assign new_new_n3954__ = ~new_new_n3952__ & ~new_new_n3953__;
  assign new_new_n3955__ = ~pi079 & new_new_n3954__;
  assign new_new_n3956__ = pi079 & ~new_new_n3954__;
  assign new_new_n3957__ = ~pi077 & ~new_new_n3846__;
  assign new_new_n3958__ = pi077 & new_new_n3846__;
  assign new_new_n3959__ = ~new_new_n3957__ & ~new_new_n3958__;
  assign new_new_n3960__ = po039 & new_new_n3959__;
  assign new_new_n3961__ = new_new_n3694__ & new_new_n3960__;
  assign new_new_n3962__ = ~new_new_n3694__ & ~new_new_n3960__;
  assign new_new_n3963__ = ~new_new_n3961__ & ~new_new_n3962__;
  assign new_new_n3964__ = ~pi078 & ~new_new_n3963__;
  assign new_new_n3965__ = pi078 & new_new_n3963__;
  assign new_new_n3966__ = ~new_new_n3704__ & ~new_new_n3705__;
  assign new_new_n3967__ = new_new_n3844__ & po039;
  assign new_new_n3968__ = ~pi076 & ~po039;
  assign new_new_n3969__ = ~new_new_n3967__ & ~new_new_n3968__;
  assign new_new_n3970__ = ~new_new_n3966__ & ~new_new_n3969__;
  assign new_new_n3971__ = new_new_n3966__ & new_new_n3969__;
  assign new_new_n3972__ = ~new_new_n3970__ & ~new_new_n3971__;
  assign new_new_n3973__ = ~pi077 & ~new_new_n3972__;
  assign new_new_n3974__ = pi077 & new_new_n3972__;
  assign new_new_n3975__ = new_new_n3842__ & po039;
  assign new_new_n3976__ = pi075 & ~po039;
  assign new_new_n3977__ = ~new_new_n3975__ & ~new_new_n3976__;
  assign new_new_n3978__ = ~new_new_n3713__ & ~new_new_n3714__;
  assign new_new_n3979__ = ~new_new_n3977__ & ~new_new_n3978__;
  assign new_new_n3980__ = new_new_n3977__ & new_new_n3978__;
  assign new_new_n3981__ = ~new_new_n3979__ & ~new_new_n3980__;
  assign new_new_n3982__ = pi076 & ~new_new_n3981__;
  assign new_new_n3983__ = ~pi076 & new_new_n3981__;
  assign new_new_n3984__ = ~new_new_n3722__ & ~new_new_n3723__;
  assign new_new_n3985__ = ~new_new_n3840__ & po039;
  assign new_new_n3986__ = ~pi074 & ~po039;
  assign new_new_n3987__ = ~new_new_n3985__ & ~new_new_n3986__;
  assign new_new_n3988__ = new_new_n3984__ & ~new_new_n3987__;
  assign new_new_n3989__ = ~new_new_n3984__ & new_new_n3987__;
  assign new_new_n3990__ = ~new_new_n3988__ & ~new_new_n3989__;
  assign new_new_n3991__ = pi075 & ~new_new_n3990__;
  assign new_new_n3992__ = ~pi075 & new_new_n3990__;
  assign new_new_n3993__ = ~pi073 & ~new_new_n3838__;
  assign new_new_n3994__ = pi073 & new_new_n3838__;
  assign new_new_n3995__ = ~new_new_n3993__ & ~new_new_n3994__;
  assign new_new_n3996__ = po039 & new_new_n3995__;
  assign new_new_n3997__ = new_new_n3730__ & new_new_n3996__;
  assign new_new_n3998__ = ~new_new_n3730__ & ~new_new_n3996__;
  assign new_new_n3999__ = ~new_new_n3997__ & ~new_new_n3998__;
  assign new_new_n4000__ = ~pi074 & ~new_new_n3999__;
  assign new_new_n4001__ = pi074 & new_new_n3999__;
  assign new_new_n4002__ = ~new_new_n3740__ & ~new_new_n3741__;
  assign new_new_n4003__ = ~new_new_n3836__ & po039;
  assign new_new_n4004__ = ~pi072 & ~po039;
  assign new_new_n4005__ = ~new_new_n4003__ & ~new_new_n4004__;
  assign new_new_n4006__ = new_new_n4002__ & ~new_new_n4005__;
  assign new_new_n4007__ = ~new_new_n4002__ & new_new_n4005__;
  assign new_new_n4008__ = ~new_new_n4006__ & ~new_new_n4007__;
  assign new_new_n4009__ = pi073 & ~new_new_n4008__;
  assign new_new_n4010__ = ~pi073 & new_new_n4008__;
  assign new_new_n4011__ = ~new_new_n3749__ & ~new_new_n3750__;
  assign new_new_n4012__ = ~new_new_n3834__ & po039;
  assign new_new_n4013__ = ~pi071 & ~po039;
  assign new_new_n4014__ = ~new_new_n4012__ & ~new_new_n4013__;
  assign new_new_n4015__ = new_new_n4011__ & ~new_new_n4014__;
  assign new_new_n4016__ = ~new_new_n4011__ & new_new_n4014__;
  assign new_new_n4017__ = ~new_new_n4015__ & ~new_new_n4016__;
  assign new_new_n4018__ = ~pi072 & new_new_n4017__;
  assign new_new_n4019__ = pi072 & ~new_new_n4017__;
  assign new_new_n4020__ = ~new_new_n3758__ & ~new_new_n3759__;
  assign new_new_n4021__ = ~new_new_n3832__ & po039;
  assign new_new_n4022__ = ~pi070 & ~po039;
  assign new_new_n4023__ = ~new_new_n4021__ & ~new_new_n4022__;
  assign new_new_n4024__ = new_new_n4020__ & ~new_new_n4023__;
  assign new_new_n4025__ = ~new_new_n4020__ & new_new_n4023__;
  assign new_new_n4026__ = ~new_new_n4024__ & ~new_new_n4025__;
  assign new_new_n4027__ = ~pi071 & new_new_n4026__;
  assign new_new_n4028__ = pi071 & ~new_new_n4026__;
  assign new_new_n4029__ = ~new_new_n3767__ & ~new_new_n3768__;
  assign new_new_n4030__ = new_new_n3830__ & po039;
  assign new_new_n4031__ = ~pi069 & ~po039;
  assign new_new_n4032__ = ~new_new_n4030__ & ~new_new_n4031__;
  assign new_new_n4033__ = ~new_new_n4029__ & ~new_new_n4032__;
  assign new_new_n4034__ = new_new_n4029__ & new_new_n4032__;
  assign new_new_n4035__ = ~new_new_n4033__ & ~new_new_n4034__;
  assign new_new_n4036__ = ~pi070 & ~new_new_n4035__;
  assign new_new_n4037__ = pi070 & new_new_n4035__;
  assign new_new_n4038__ = pi068 & ~new_new_n3828__;
  assign new_new_n4039__ = ~pi068 & new_new_n3828__;
  assign new_new_n4040__ = ~new_new_n4038__ & ~new_new_n4039__;
  assign new_new_n4041__ = po039 & new_new_n4040__;
  assign new_new_n4042__ = ~new_new_n3775__ & ~new_new_n4041__;
  assign new_new_n4043__ = new_new_n3775__ & new_new_n4041__;
  assign new_new_n4044__ = ~new_new_n4042__ & ~new_new_n4043__;
  assign new_new_n4045__ = ~pi069 & new_new_n4044__;
  assign new_new_n4046__ = pi069 & ~new_new_n4044__;
  assign new_new_n4047__ = ~new_new_n3783__ & ~new_new_n3784__;
  assign new_new_n4048__ = ~new_new_n3826__ & po039;
  assign new_new_n4049__ = pi067 & ~po039;
  assign new_new_n4050__ = ~new_new_n4048__ & ~new_new_n4049__;
  assign new_new_n4051__ = new_new_n4047__ & ~new_new_n4050__;
  assign new_new_n4052__ = ~new_new_n4047__ & new_new_n4050__;
  assign new_new_n4053__ = ~new_new_n4051__ & ~new_new_n4052__;
  assign new_new_n4054__ = ~pi068 & ~new_new_n4053__;
  assign new_new_n4055__ = pi068 & new_new_n4053__;
  assign new_new_n4056__ = ~new_new_n3797__ & ~new_new_n3798__;
  assign new_new_n4057__ = po039 & new_new_n4056__;
  assign new_new_n4058__ = new_new_n3824__ & ~new_new_n4057__;
  assign new_new_n4059__ = ~new_new_n3824__ & new_new_n4057__;
  assign new_new_n4060__ = ~new_new_n4058__ & ~new_new_n4059__;
  assign new_new_n4061__ = pi067 & ~new_new_n4060__;
  assign new_new_n4062__ = ~pi067 & new_new_n4060__;
  assign new_new_n4063__ = pi039 & po039;
  assign new_new_n4064__ = pi038 & ~pi065;
  assign new_new_n4065__ = new_new_n4063__ & ~new_new_n4064__;
  assign new_new_n4066__ = ~pi039 & ~po039;
  assign new_new_n4067__ = ~pi065 & ~new_new_n4066__;
  assign new_new_n4068__ = ~pi038 & ~new_new_n4067__;
  assign new_new_n4069__ = ~new_new_n4065__ & ~new_new_n4068__;
  assign new_new_n4070__ = pi064 & ~new_new_n4069__;
  assign new_new_n4071__ = pi064 & po039;
  assign new_new_n4072__ = ~pi039 & pi065;
  assign new_new_n4073__ = ~new_new_n4071__ & new_new_n4072__;
  assign new_new_n4074__ = ~new_new_n4070__ & ~new_new_n4073__;
  assign new_new_n4075__ = pi066 & ~new_new_n4074__;
  assign new_new_n4076__ = ~pi066 & new_new_n4074__;
  assign new_new_n4077__ = new_new_n426__ & ~po040;
  assign new_new_n4078__ = new_new_n3817__ & po039;
  assign new_new_n4079__ = ~new_new_n4077__ & ~new_new_n4078__;
  assign new_new_n4080__ = ~pi039 & ~new_new_n4079__;
  assign new_new_n4081__ = ~new_new_n332__ & po039;
  assign new_new_n4082__ = ~new_new_n3793__ & ~new_new_n4081__;
  assign new_new_n4083__ = pi065 & po039;
  assign new_new_n4084__ = po040 & ~new_new_n4083__;
  assign new_new_n4085__ = pi065 & ~new_new_n3793__;
  assign new_new_n4086__ = pi039 & ~new_new_n4085__;
  assign new_new_n4087__ = ~new_new_n4084__ & new_new_n4086__;
  assign new_new_n4088__ = ~new_new_n4080__ & ~new_new_n4082__;
  assign new_new_n4089__ = ~new_new_n4087__ & new_new_n4088__;
  assign new_new_n4090__ = pi040 & ~new_new_n4089__;
  assign new_new_n4091__ = ~new_new_n3793__ & ~new_new_n4083__;
  assign new_new_n4092__ = pi039 & ~new_new_n3805__;
  assign new_new_n4093__ = pi064 & ~new_new_n4092__;
  assign new_new_n4094__ = ~new_new_n4091__ & ~new_new_n4093__;
  assign new_new_n4095__ = ~pi065 & po039;
  assign new_new_n4096__ = ~po040 & ~new_new_n4095__;
  assign new_new_n4097__ = pi064 & ~new_new_n4063__;
  assign new_new_n4098__ = ~new_new_n4078__ & new_new_n4097__;
  assign new_new_n4099__ = ~new_new_n4096__ & new_new_n4098__;
  assign new_new_n4100__ = ~new_new_n4094__ & ~new_new_n4099__;
  assign new_new_n4101__ = ~pi040 & ~new_new_n4100__;
  assign new_new_n4102__ = ~new_new_n4090__ & ~new_new_n4101__;
  assign new_new_n4103__ = ~new_new_n4076__ & new_new_n4102__;
  assign new_new_n4104__ = ~new_new_n4075__ & ~new_new_n4103__;
  assign new_new_n4105__ = ~new_new_n4062__ & ~new_new_n4104__;
  assign new_new_n4106__ = ~new_new_n4061__ & ~new_new_n4105__;
  assign new_new_n4107__ = ~new_new_n4055__ & new_new_n4106__;
  assign new_new_n4108__ = ~new_new_n4054__ & ~new_new_n4107__;
  assign new_new_n4109__ = ~new_new_n4046__ & ~new_new_n4108__;
  assign new_new_n4110__ = ~new_new_n4045__ & ~new_new_n4109__;
  assign new_new_n4111__ = ~new_new_n4037__ & ~new_new_n4110__;
  assign new_new_n4112__ = ~new_new_n4036__ & ~new_new_n4111__;
  assign new_new_n4113__ = ~new_new_n4028__ & ~new_new_n4112__;
  assign new_new_n4114__ = ~new_new_n4027__ & ~new_new_n4113__;
  assign new_new_n4115__ = ~new_new_n4019__ & ~new_new_n4114__;
  assign new_new_n4116__ = ~new_new_n4018__ & ~new_new_n4115__;
  assign new_new_n4117__ = ~new_new_n4010__ & new_new_n4116__;
  assign new_new_n4118__ = ~new_new_n4009__ & ~new_new_n4117__;
  assign new_new_n4119__ = ~new_new_n4001__ & new_new_n4118__;
  assign new_new_n4120__ = ~new_new_n4000__ & ~new_new_n4119__;
  assign new_new_n4121__ = ~new_new_n3992__ & new_new_n4120__;
  assign new_new_n4122__ = ~new_new_n3991__ & ~new_new_n4121__;
  assign new_new_n4123__ = ~new_new_n3983__ & ~new_new_n4122__;
  assign new_new_n4124__ = ~new_new_n3982__ & ~new_new_n4123__;
  assign new_new_n4125__ = ~new_new_n3974__ & new_new_n4124__;
  assign new_new_n4126__ = ~new_new_n3973__ & ~new_new_n4125__;
  assign new_new_n4127__ = ~new_new_n3965__ & ~new_new_n4126__;
  assign new_new_n4128__ = ~new_new_n3964__ & ~new_new_n4127__;
  assign new_new_n4129__ = ~new_new_n3956__ & ~new_new_n4128__;
  assign new_new_n4130__ = ~new_new_n3955__ & ~new_new_n4129__;
  assign new_new_n4131__ = ~new_new_n3947__ & new_new_n4130__;
  assign new_new_n4132__ = ~new_new_n3946__ & ~new_new_n4131__;
  assign new_new_n4133__ = ~new_new_n3938__ & ~new_new_n4132__;
  assign new_new_n4134__ = ~new_new_n3937__ & ~new_new_n4133__;
  assign new_new_n4135__ = ~new_new_n3929__ & ~new_new_n4134__;
  assign new_new_n4136__ = ~new_new_n3928__ & ~new_new_n4135__;
  assign new_new_n4137__ = ~new_new_n3920__ & ~new_new_n4136__;
  assign new_new_n4138__ = ~new_new_n3919__ & ~new_new_n4137__;
  assign new_new_n4139__ = ~new_new_n3911__ & ~new_new_n4138__;
  assign new_new_n4140__ = ~new_new_n3910__ & ~new_new_n4139__;
  assign new_new_n4141__ = ~new_new_n3902__ & ~new_new_n4140__;
  assign new_new_n4142__ = ~new_new_n3901__ & ~new_new_n4141__;
  assign new_new_n4143__ = new_new_n3613__ & ~po039;
  assign new_new_n4144__ = ~new_new_n376__ & ~new_new_n4143__;
  assign new_new_n4145__ = ~pi089 & ~new_new_n4144__;
  assign new_new_n4146__ = ~new_new_n3869__ & new_new_n3882__;
  assign new_new_n4147__ = new_new_n3868__ & new_new_n4146__;
  assign new_new_n4148__ = ~new_new_n3878__ & ~new_new_n4147__;
  assign new_new_n4149__ = new_new_n3334__ & new_new_n3613__;
  assign new_new_n4150__ = ~new_new_n3867__ & new_new_n4149__;
  assign new_new_n4151__ = new_new_n3879__ & new_new_n4150__;
  assign new_new_n4152__ = ~new_new_n4148__ & ~new_new_n4151__;
  assign new_new_n4153__ = ~new_new_n3623__ & ~new_new_n3624__;
  assign new_new_n4154__ = ~new_new_n3864__ & po039;
  assign new_new_n4155__ = pi086 & ~po039;
  assign new_new_n4156__ = ~new_new_n4154__ & ~new_new_n4155__;
  assign new_new_n4157__ = new_new_n4153__ & new_new_n4156__;
  assign new_new_n4158__ = ~new_new_n4153__ & ~new_new_n4156__;
  assign new_new_n4159__ = ~new_new_n4157__ & ~new_new_n4158__;
  assign new_new_n4160__ = pi087 & ~new_new_n4159__;
  assign new_new_n4161__ = ~pi087 & new_new_n4159__;
  assign new_new_n4162__ = ~new_new_n3892__ & ~new_new_n4142__;
  assign new_new_n4163__ = ~new_new_n3891__ & ~new_new_n4162__;
  assign new_new_n4164__ = ~new_new_n4161__ & ~new_new_n4163__;
  assign new_new_n4165__ = ~new_new_n4160__ & ~new_new_n4164__;
  assign new_new_n4166__ = ~pi088 & new_new_n4165__;
  assign new_new_n4167__ = new_new_n4152__ & ~new_new_n4166__;
  assign new_new_n4168__ = pi088 & ~new_new_n4165__;
  assign new_new_n4169__ = pi089 & new_new_n4144__;
  assign new_new_n4170__ = ~new_new_n4168__ & ~new_new_n4169__;
  assign new_new_n4171__ = ~new_new_n4167__ & new_new_n4170__;
  assign new_new_n4172__ = ~new_new_n4145__ & ~new_new_n4171__;
  assign new_new_n4173__ = ~pi090 & ~new_new_n4172__;
  assign po038 = new_new_n3333__ & new_new_n4173__;
  assign new_new_n4175__ = ~new_new_n4142__ & po038;
  assign new_new_n4176__ = pi086 & ~po038;
  assign new_new_n4177__ = ~new_new_n4175__ & ~new_new_n4176__;
  assign new_new_n4178__ = new_new_n3893__ & ~new_new_n4177__;
  assign new_new_n4179__ = ~new_new_n3893__ & new_new_n4177__;
  assign new_new_n4180__ = ~new_new_n4178__ & ~new_new_n4179__;
  assign new_new_n4181__ = ~new_new_n4166__ & ~new_new_n4168__;
  assign new_new_n4182__ = po038 & new_new_n4181__;
  assign new_new_n4183__ = new_new_n4152__ & ~new_new_n4182__;
  assign new_new_n4184__ = ~new_new_n4152__ & new_new_n4182__;
  assign new_new_n4185__ = ~new_new_n4183__ & ~new_new_n4184__;
  assign new_new_n4186__ = ~pi089 & new_new_n4185__;
  assign new_new_n4187__ = pi089 & ~new_new_n4185__;
  assign new_new_n4188__ = ~pi087 & ~new_new_n4180__;
  assign new_new_n4189__ = pi087 & new_new_n4180__;
  assign new_new_n4190__ = ~new_new_n3901__ & ~new_new_n3902__;
  assign new_new_n4191__ = ~new_new_n4140__ & po038;
  assign new_new_n4192__ = pi085 & ~po038;
  assign new_new_n4193__ = ~new_new_n4191__ & ~new_new_n4192__;
  assign new_new_n4194__ = new_new_n4190__ & ~new_new_n4193__;
  assign new_new_n4195__ = ~new_new_n4190__ & new_new_n4193__;
  assign new_new_n4196__ = ~new_new_n4194__ & ~new_new_n4195__;
  assign new_new_n4197__ = ~pi086 & ~new_new_n4196__;
  assign new_new_n4198__ = pi086 & new_new_n4196__;
  assign new_new_n4199__ = ~new_new_n4138__ & po038;
  assign new_new_n4200__ = pi084 & ~po038;
  assign new_new_n4201__ = ~new_new_n4199__ & ~new_new_n4200__;
  assign new_new_n4202__ = ~new_new_n3910__ & ~new_new_n3911__;
  assign new_new_n4203__ = ~new_new_n4201__ & new_new_n4202__;
  assign new_new_n4204__ = new_new_n4201__ & ~new_new_n4202__;
  assign new_new_n4205__ = ~new_new_n4203__ & ~new_new_n4204__;
  assign new_new_n4206__ = ~pi085 & ~new_new_n4205__;
  assign new_new_n4207__ = pi085 & new_new_n4205__;
  assign new_new_n4208__ = ~new_new_n3919__ & ~new_new_n3920__;
  assign new_new_n4209__ = ~new_new_n4136__ & po038;
  assign new_new_n4210__ = pi083 & ~po038;
  assign new_new_n4211__ = ~new_new_n4209__ & ~new_new_n4210__;
  assign new_new_n4212__ = new_new_n4208__ & new_new_n4211__;
  assign new_new_n4213__ = ~new_new_n4208__ & ~new_new_n4211__;
  assign new_new_n4214__ = ~new_new_n4212__ & ~new_new_n4213__;
  assign new_new_n4215__ = ~pi084 & new_new_n4214__;
  assign new_new_n4216__ = pi084 & ~new_new_n4214__;
  assign new_new_n4217__ = new_new_n4134__ & po038;
  assign new_new_n4218__ = ~pi082 & ~po038;
  assign new_new_n4219__ = ~new_new_n4217__ & ~new_new_n4218__;
  assign new_new_n4220__ = ~new_new_n3928__ & ~new_new_n3929__;
  assign new_new_n4221__ = ~new_new_n4219__ & ~new_new_n4220__;
  assign new_new_n4222__ = new_new_n4219__ & new_new_n4220__;
  assign new_new_n4223__ = ~new_new_n4221__ & ~new_new_n4222__;
  assign new_new_n4224__ = ~pi083 & ~new_new_n4223__;
  assign new_new_n4225__ = pi083 & new_new_n4223__;
  assign new_new_n4226__ = ~new_new_n3937__ & ~new_new_n3938__;
  assign new_new_n4227__ = ~new_new_n4132__ & po038;
  assign new_new_n4228__ = pi081 & ~po038;
  assign new_new_n4229__ = ~new_new_n4227__ & ~new_new_n4228__;
  assign new_new_n4230__ = new_new_n4226__ & new_new_n4229__;
  assign new_new_n4231__ = ~new_new_n4226__ & ~new_new_n4229__;
  assign new_new_n4232__ = ~new_new_n4230__ & ~new_new_n4231__;
  assign new_new_n4233__ = pi082 & ~new_new_n4232__;
  assign new_new_n4234__ = ~pi082 & new_new_n4232__;
  assign new_new_n4235__ = new_new_n4130__ & po038;
  assign new_new_n4236__ = pi080 & ~po038;
  assign new_new_n4237__ = ~new_new_n4235__ & ~new_new_n4236__;
  assign new_new_n4238__ = ~new_new_n3946__ & ~new_new_n3947__;
  assign new_new_n4239__ = ~new_new_n4237__ & ~new_new_n4238__;
  assign new_new_n4240__ = new_new_n4237__ & new_new_n4238__;
  assign new_new_n4241__ = ~new_new_n4239__ & ~new_new_n4240__;
  assign new_new_n4242__ = ~pi081 & new_new_n4241__;
  assign new_new_n4243__ = pi081 & ~new_new_n4241__;
  assign new_new_n4244__ = ~new_new_n3955__ & ~new_new_n3956__;
  assign new_new_n4245__ = ~new_new_n4128__ & po038;
  assign new_new_n4246__ = ~pi079 & ~po038;
  assign new_new_n4247__ = ~new_new_n4245__ & ~new_new_n4246__;
  assign new_new_n4248__ = new_new_n4244__ & new_new_n4247__;
  assign new_new_n4249__ = ~new_new_n4244__ & ~new_new_n4247__;
  assign new_new_n4250__ = ~new_new_n4248__ & ~new_new_n4249__;
  assign new_new_n4251__ = ~pi080 & ~new_new_n4250__;
  assign new_new_n4252__ = pi080 & new_new_n4250__;
  assign new_new_n4253__ = ~pi078 & ~new_new_n4126__;
  assign new_new_n4254__ = pi078 & new_new_n4126__;
  assign new_new_n4255__ = ~new_new_n4253__ & ~new_new_n4254__;
  assign new_new_n4256__ = po038 & new_new_n4255__;
  assign new_new_n4257__ = new_new_n3963__ & new_new_n4256__;
  assign new_new_n4258__ = ~new_new_n3963__ & ~new_new_n4256__;
  assign new_new_n4259__ = ~new_new_n4257__ & ~new_new_n4258__;
  assign new_new_n4260__ = ~pi079 & ~new_new_n4259__;
  assign new_new_n4261__ = pi079 & new_new_n4259__;
  assign new_new_n4262__ = ~new_new_n3973__ & ~new_new_n3974__;
  assign new_new_n4263__ = new_new_n4124__ & po038;
  assign new_new_n4264__ = ~pi077 & ~po038;
  assign new_new_n4265__ = ~new_new_n4263__ & ~new_new_n4264__;
  assign new_new_n4266__ = ~new_new_n4262__ & ~new_new_n4265__;
  assign new_new_n4267__ = new_new_n4262__ & new_new_n4265__;
  assign new_new_n4268__ = ~new_new_n4266__ & ~new_new_n4267__;
  assign new_new_n4269__ = ~pi078 & ~new_new_n4268__;
  assign new_new_n4270__ = pi078 & new_new_n4268__;
  assign new_new_n4271__ = ~new_new_n3982__ & ~new_new_n3983__;
  assign new_new_n4272__ = ~new_new_n4122__ & po038;
  assign new_new_n4273__ = pi076 & ~po038;
  assign new_new_n4274__ = ~new_new_n4272__ & ~new_new_n4273__;
  assign new_new_n4275__ = new_new_n4271__ & ~new_new_n4274__;
  assign new_new_n4276__ = ~new_new_n4271__ & new_new_n4274__;
  assign new_new_n4277__ = ~new_new_n4275__ & ~new_new_n4276__;
  assign new_new_n4278__ = ~pi077 & ~new_new_n4277__;
  assign new_new_n4279__ = pi077 & new_new_n4277__;
  assign new_new_n4280__ = ~new_new_n3991__ & ~new_new_n3992__;
  assign new_new_n4281__ = ~new_new_n4120__ & po038;
  assign new_new_n4282__ = ~pi075 & ~po038;
  assign new_new_n4283__ = ~new_new_n4281__ & ~new_new_n4282__;
  assign new_new_n4284__ = new_new_n4280__ & ~new_new_n4283__;
  assign new_new_n4285__ = ~new_new_n4280__ & new_new_n4283__;
  assign new_new_n4286__ = ~new_new_n4284__ & ~new_new_n4285__;
  assign new_new_n4287__ = ~pi076 & new_new_n4286__;
  assign new_new_n4288__ = pi076 & ~new_new_n4286__;
  assign new_new_n4289__ = ~new_new_n4000__ & ~new_new_n4001__;
  assign new_new_n4290__ = new_new_n4118__ & po038;
  assign new_new_n4291__ = ~pi074 & ~po038;
  assign new_new_n4292__ = ~new_new_n4290__ & ~new_new_n4291__;
  assign new_new_n4293__ = ~new_new_n4289__ & ~new_new_n4292__;
  assign new_new_n4294__ = new_new_n4289__ & new_new_n4292__;
  assign new_new_n4295__ = ~new_new_n4293__ & ~new_new_n4294__;
  assign new_new_n4296__ = ~pi075 & ~new_new_n4295__;
  assign new_new_n4297__ = pi075 & new_new_n4295__;
  assign new_new_n4298__ = new_new_n4116__ & po038;
  assign new_new_n4299__ = pi073 & ~po038;
  assign new_new_n4300__ = ~new_new_n4298__ & ~new_new_n4299__;
  assign new_new_n4301__ = ~new_new_n4009__ & ~new_new_n4010__;
  assign new_new_n4302__ = ~new_new_n4300__ & ~new_new_n4301__;
  assign new_new_n4303__ = new_new_n4300__ & new_new_n4301__;
  assign new_new_n4304__ = ~new_new_n4302__ & ~new_new_n4303__;
  assign new_new_n4305__ = ~pi074 & new_new_n4304__;
  assign new_new_n4306__ = pi074 & ~new_new_n4304__;
  assign new_new_n4307__ = ~new_new_n4018__ & ~new_new_n4019__;
  assign new_new_n4308__ = ~new_new_n4114__ & po038;
  assign new_new_n4309__ = ~pi072 & ~po038;
  assign new_new_n4310__ = ~new_new_n4308__ & ~new_new_n4309__;
  assign new_new_n4311__ = new_new_n4307__ & new_new_n4310__;
  assign new_new_n4312__ = ~new_new_n4307__ & ~new_new_n4310__;
  assign new_new_n4313__ = ~new_new_n4311__ & ~new_new_n4312__;
  assign new_new_n4314__ = ~pi073 & ~new_new_n4313__;
  assign new_new_n4315__ = pi073 & new_new_n4313__;
  assign new_new_n4316__ = new_new_n4112__ & po038;
  assign new_new_n4317__ = pi071 & ~po038;
  assign new_new_n4318__ = ~new_new_n4316__ & ~new_new_n4317__;
  assign new_new_n4319__ = ~new_new_n4027__ & ~new_new_n4028__;
  assign new_new_n4320__ = ~new_new_n4318__ & ~new_new_n4319__;
  assign new_new_n4321__ = new_new_n4318__ & new_new_n4319__;
  assign new_new_n4322__ = ~new_new_n4320__ & ~new_new_n4321__;
  assign new_new_n4323__ = pi072 & ~new_new_n4322__;
  assign new_new_n4324__ = ~pi072 & new_new_n4322__;
  assign new_new_n4325__ = ~new_new_n4036__ & ~new_new_n4037__;
  assign new_new_n4326__ = ~new_new_n4110__ & po038;
  assign new_new_n4327__ = ~pi070 & ~po038;
  assign new_new_n4328__ = ~new_new_n4326__ & ~new_new_n4327__;
  assign new_new_n4329__ = new_new_n4325__ & ~new_new_n4328__;
  assign new_new_n4330__ = ~new_new_n4325__ & new_new_n4328__;
  assign new_new_n4331__ = ~new_new_n4329__ & ~new_new_n4330__;
  assign new_new_n4332__ = pi071 & ~new_new_n4331__;
  assign new_new_n4333__ = ~pi071 & new_new_n4331__;
  assign new_new_n4334__ = ~new_new_n4045__ & ~new_new_n4046__;
  assign new_new_n4335__ = ~new_new_n4108__ & po038;
  assign new_new_n4336__ = ~pi069 & ~po038;
  assign new_new_n4337__ = ~new_new_n4335__ & ~new_new_n4336__;
  assign new_new_n4338__ = new_new_n4334__ & ~new_new_n4337__;
  assign new_new_n4339__ = ~new_new_n4334__ & new_new_n4337__;
  assign new_new_n4340__ = ~new_new_n4338__ & ~new_new_n4339__;
  assign new_new_n4341__ = pi070 & ~new_new_n4340__;
  assign new_new_n4342__ = ~pi070 & new_new_n4340__;
  assign new_new_n4343__ = ~new_new_n4054__ & ~new_new_n4055__;
  assign new_new_n4344__ = new_new_n4106__ & po038;
  assign new_new_n4345__ = ~pi068 & ~po038;
  assign new_new_n4346__ = ~new_new_n4344__ & ~new_new_n4345__;
  assign new_new_n4347__ = ~new_new_n4343__ & ~new_new_n4346__;
  assign new_new_n4348__ = new_new_n4343__ & new_new_n4346__;
  assign new_new_n4349__ = ~new_new_n4347__ & ~new_new_n4348__;
  assign new_new_n4350__ = ~pi069 & ~new_new_n4349__;
  assign new_new_n4351__ = pi069 & new_new_n4349__;
  assign new_new_n4352__ = ~new_new_n4104__ & po038;
  assign new_new_n4353__ = pi067 & ~po038;
  assign new_new_n4354__ = ~new_new_n4352__ & ~new_new_n4353__;
  assign new_new_n4355__ = ~new_new_n4061__ & ~new_new_n4062__;
  assign new_new_n4356__ = ~new_new_n4354__ & new_new_n4355__;
  assign new_new_n4357__ = new_new_n4354__ & ~new_new_n4355__;
  assign new_new_n4358__ = ~new_new_n4356__ & ~new_new_n4357__;
  assign new_new_n4359__ = ~pi068 & ~new_new_n4358__;
  assign new_new_n4360__ = pi068 & new_new_n4358__;
  assign new_new_n4361__ = ~new_new_n4075__ & ~new_new_n4076__;
  assign new_new_n4362__ = po038 & new_new_n4361__;
  assign new_new_n4363__ = new_new_n4102__ & ~new_new_n4362__;
  assign new_new_n4364__ = ~new_new_n4102__ & new_new_n4362__;
  assign new_new_n4365__ = ~new_new_n4363__ & ~new_new_n4364__;
  assign new_new_n4366__ = ~pi067 & new_new_n4365__;
  assign new_new_n4367__ = pi067 & ~new_new_n4365__;
  assign new_new_n4368__ = ~pi038 & ~po038;
  assign new_new_n4369__ = ~pi065 & ~new_new_n4368__;
  assign new_new_n4370__ = ~pi037 & ~new_new_n4369__;
  assign new_new_n4371__ = pi037 & ~pi065;
  assign new_new_n4372__ = pi038 & ~new_new_n4371__;
  assign new_new_n4373__ = po038 & new_new_n4372__;
  assign new_new_n4374__ = ~new_new_n4370__ & ~new_new_n4373__;
  assign new_new_n4375__ = pi064 & ~new_new_n4374__;
  assign new_new_n4376__ = pi064 & po038;
  assign new_new_n4377__ = ~pi038 & pi065;
  assign new_new_n4378__ = ~new_new_n4376__ & new_new_n4377__;
  assign new_new_n4379__ = ~new_new_n4375__ & ~new_new_n4378__;
  assign new_new_n4380__ = ~pi066 & new_new_n4379__;
  assign new_new_n4381__ = pi066 & ~new_new_n4379__;
  assign new_new_n4382__ = ~pi065 & ~po039;
  assign new_new_n4383__ = new_new_n4083__ & new_new_n4376__;
  assign new_new_n4384__ = ~new_new_n4382__ & ~new_new_n4383__;
  assign new_new_n4385__ = pi038 & ~new_new_n4384__;
  assign new_new_n4386__ = ~new_new_n332__ & po038;
  assign new_new_n4387__ = ~new_new_n4071__ & ~new_new_n4386__;
  assign new_new_n4388__ = po039 & ~new_new_n4173__;
  assign new_new_n4389__ = ~new_new_n426__ & ~po039;
  assign new_new_n4390__ = ~pi038 & ~new_new_n4083__;
  assign new_new_n4391__ = ~new_new_n4389__ & new_new_n4390__;
  assign new_new_n4392__ = ~new_new_n4388__ & new_new_n4391__;
  assign new_new_n4393__ = ~new_new_n4387__ & ~new_new_n4392__;
  assign new_new_n4394__ = ~new_new_n4385__ & new_new_n4393__;
  assign new_new_n4395__ = pi039 & ~new_new_n4394__;
  assign new_new_n4396__ = po038 & new_new_n4382__;
  assign new_new_n4397__ = ~new_new_n4083__ & ~new_new_n4396__;
  assign new_new_n4398__ = ~pi038 & ~new_new_n4397__;
  assign new_new_n4399__ = ~new_new_n4388__ & ~new_new_n4398__;
  assign new_new_n4400__ = pi064 & ~new_new_n4399__;
  assign new_new_n4401__ = pi065 & po038;
  assign new_new_n4402__ = ~new_new_n4071__ & ~new_new_n4401__;
  assign new_new_n4403__ = pi038 & ~new_new_n4083__;
  assign new_new_n4404__ = pi064 & ~new_new_n4403__;
  assign new_new_n4405__ = ~new_new_n4402__ & ~new_new_n4404__;
  assign new_new_n4406__ = ~new_new_n4400__ & ~new_new_n4405__;
  assign new_new_n4407__ = ~pi039 & ~new_new_n4406__;
  assign new_new_n4408__ = ~new_new_n4395__ & ~new_new_n4407__;
  assign new_new_n4409__ = ~new_new_n4381__ & ~new_new_n4408__;
  assign new_new_n4410__ = ~new_new_n4380__ & ~new_new_n4409__;
  assign new_new_n4411__ = ~new_new_n4367__ & ~new_new_n4410__;
  assign new_new_n4412__ = ~new_new_n4366__ & ~new_new_n4411__;
  assign new_new_n4413__ = ~new_new_n4360__ & ~new_new_n4412__;
  assign new_new_n4414__ = ~new_new_n4359__ & ~new_new_n4413__;
  assign new_new_n4415__ = ~new_new_n4351__ & ~new_new_n4414__;
  assign new_new_n4416__ = ~new_new_n4350__ & ~new_new_n4415__;
  assign new_new_n4417__ = ~new_new_n4342__ & new_new_n4416__;
  assign new_new_n4418__ = ~new_new_n4341__ & ~new_new_n4417__;
  assign new_new_n4419__ = ~new_new_n4333__ & ~new_new_n4418__;
  assign new_new_n4420__ = ~new_new_n4332__ & ~new_new_n4419__;
  assign new_new_n4421__ = ~new_new_n4324__ & ~new_new_n4420__;
  assign new_new_n4422__ = ~new_new_n4323__ & ~new_new_n4421__;
  assign new_new_n4423__ = ~new_new_n4315__ & new_new_n4422__;
  assign new_new_n4424__ = ~new_new_n4314__ & ~new_new_n4423__;
  assign new_new_n4425__ = ~new_new_n4306__ & ~new_new_n4424__;
  assign new_new_n4426__ = ~new_new_n4305__ & ~new_new_n4425__;
  assign new_new_n4427__ = ~new_new_n4297__ & ~new_new_n4426__;
  assign new_new_n4428__ = ~new_new_n4296__ & ~new_new_n4427__;
  assign new_new_n4429__ = ~new_new_n4288__ & ~new_new_n4428__;
  assign new_new_n4430__ = ~new_new_n4287__ & ~new_new_n4429__;
  assign new_new_n4431__ = ~new_new_n4279__ & ~new_new_n4430__;
  assign new_new_n4432__ = ~new_new_n4278__ & ~new_new_n4431__;
  assign new_new_n4433__ = ~new_new_n4270__ & ~new_new_n4432__;
  assign new_new_n4434__ = ~new_new_n4269__ & ~new_new_n4433__;
  assign new_new_n4435__ = ~new_new_n4261__ & ~new_new_n4434__;
  assign new_new_n4436__ = ~new_new_n4260__ & ~new_new_n4435__;
  assign new_new_n4437__ = ~new_new_n4252__ & ~new_new_n4436__;
  assign new_new_n4438__ = ~new_new_n4251__ & ~new_new_n4437__;
  assign new_new_n4439__ = ~new_new_n4243__ & ~new_new_n4438__;
  assign new_new_n4440__ = ~new_new_n4242__ & ~new_new_n4439__;
  assign new_new_n4441__ = ~new_new_n4234__ & new_new_n4440__;
  assign new_new_n4442__ = ~new_new_n4233__ & ~new_new_n4441__;
  assign new_new_n4443__ = ~new_new_n4225__ & new_new_n4442__;
  assign new_new_n4444__ = ~new_new_n4224__ & ~new_new_n4443__;
  assign new_new_n4445__ = ~new_new_n4216__ & ~new_new_n4444__;
  assign new_new_n4446__ = ~new_new_n4215__ & ~new_new_n4445__;
  assign new_new_n4447__ = ~new_new_n4207__ & ~new_new_n4446__;
  assign new_new_n4448__ = ~new_new_n4206__ & ~new_new_n4447__;
  assign new_new_n4449__ = ~new_new_n4198__ & ~new_new_n4448__;
  assign new_new_n4450__ = ~new_new_n4197__ & ~new_new_n4449__;
  assign new_new_n4451__ = ~new_new_n4189__ & ~new_new_n4450__;
  assign new_new_n4452__ = ~new_new_n4188__ & ~new_new_n4451__;
  assign new_new_n4453__ = ~pi088 & ~new_new_n4452__;
  assign new_new_n4454__ = pi088 & new_new_n4452__;
  assign new_new_n4455__ = ~new_new_n4160__ & ~new_new_n4161__;
  assign new_new_n4456__ = ~new_new_n4163__ & po038;
  assign new_new_n4457__ = pi087 & ~po038;
  assign new_new_n4458__ = ~new_new_n4456__ & ~new_new_n4457__;
  assign new_new_n4459__ = new_new_n4455__ & new_new_n4458__;
  assign new_new_n4460__ = ~new_new_n4455__ & ~new_new_n4458__;
  assign new_new_n4461__ = ~new_new_n4459__ & ~new_new_n4460__;
  assign new_new_n4462__ = ~new_new_n4454__ & new_new_n4461__;
  assign new_new_n4463__ = ~new_new_n4453__ & ~new_new_n4462__;
  assign new_new_n4464__ = ~new_new_n4187__ & ~new_new_n4463__;
  assign new_new_n4465__ = ~new_new_n4186__ & ~new_new_n4464__;
  assign new_new_n4466__ = pi090 & new_new_n4465__;
  assign new_new_n4467__ = new_new_n3333__ & ~new_new_n4466__;
  assign new_new_n4468__ = ~pi090 & ~new_new_n4465__;
  assign new_new_n4469__ = new_new_n4143__ & ~new_new_n4173__;
  assign new_new_n4470__ = ~new_new_n376__ & ~new_new_n4469__;
  assign new_new_n4471__ = ~new_new_n4468__ & new_new_n4470__;
  assign po037 = new_new_n4467__ & ~new_new_n4471__;
  assign new_new_n4473__ = ~pi087 & ~new_new_n4450__;
  assign new_new_n4474__ = pi087 & new_new_n4450__;
  assign new_new_n4475__ = ~new_new_n4473__ & ~new_new_n4474__;
  assign new_new_n4476__ = po037 & new_new_n4475__;
  assign new_new_n4477__ = new_new_n4180__ & new_new_n4476__;
  assign new_new_n4478__ = ~new_new_n4180__ & ~new_new_n4476__;
  assign new_new_n4479__ = ~new_new_n4477__ & ~new_new_n4478__;
  assign new_new_n4480__ = ~pi088 & ~new_new_n4479__;
  assign new_new_n4481__ = pi088 & new_new_n4479__;
  assign new_new_n4482__ = ~new_new_n4197__ & ~new_new_n4198__;
  assign new_new_n4483__ = ~new_new_n4448__ & po037;
  assign new_new_n4484__ = ~pi086 & ~po037;
  assign new_new_n4485__ = ~new_new_n4483__ & ~new_new_n4484__;
  assign new_new_n4486__ = ~new_new_n4482__ & ~new_new_n4485__;
  assign new_new_n4487__ = new_new_n4482__ & new_new_n4485__;
  assign new_new_n4488__ = ~new_new_n4486__ & ~new_new_n4487__;
  assign new_new_n4489__ = ~pi087 & ~new_new_n4488__;
  assign new_new_n4490__ = pi087 & new_new_n4488__;
  assign new_new_n4491__ = ~pi085 & ~new_new_n4446__;
  assign new_new_n4492__ = pi085 & new_new_n4446__;
  assign new_new_n4493__ = ~new_new_n4491__ & ~new_new_n4492__;
  assign new_new_n4494__ = po037 & new_new_n4493__;
  assign new_new_n4495__ = new_new_n4205__ & new_new_n4494__;
  assign new_new_n4496__ = ~new_new_n4205__ & ~new_new_n4494__;
  assign new_new_n4497__ = ~new_new_n4495__ & ~new_new_n4496__;
  assign new_new_n4498__ = ~pi086 & ~new_new_n4497__;
  assign new_new_n4499__ = pi086 & new_new_n4497__;
  assign new_new_n4500__ = ~new_new_n4215__ & ~new_new_n4216__;
  assign new_new_n4501__ = ~new_new_n4444__ & po037;
  assign new_new_n4502__ = ~pi084 & ~po037;
  assign new_new_n4503__ = ~new_new_n4501__ & ~new_new_n4502__;
  assign new_new_n4504__ = new_new_n4500__ & ~new_new_n4503__;
  assign new_new_n4505__ = ~new_new_n4500__ & new_new_n4503__;
  assign new_new_n4506__ = ~new_new_n4504__ & ~new_new_n4505__;
  assign new_new_n4507__ = pi085 & ~new_new_n4506__;
  assign new_new_n4508__ = ~pi085 & new_new_n4506__;
  assign new_new_n4509__ = ~new_new_n4224__ & ~new_new_n4225__;
  assign new_new_n4510__ = ~new_new_n4442__ & po037;
  assign new_new_n4511__ = pi083 & ~po037;
  assign new_new_n4512__ = ~new_new_n4510__ & ~new_new_n4511__;
  assign new_new_n4513__ = new_new_n4509__ & ~new_new_n4512__;
  assign new_new_n4514__ = ~new_new_n4509__ & new_new_n4512__;
  assign new_new_n4515__ = ~new_new_n4513__ & ~new_new_n4514__;
  assign new_new_n4516__ = pi084 & new_new_n4515__;
  assign new_new_n4517__ = ~pi084 & ~new_new_n4515__;
  assign new_new_n4518__ = ~new_new_n4233__ & ~new_new_n4234__;
  assign new_new_n4519__ = ~new_new_n4440__ & po037;
  assign new_new_n4520__ = ~pi082 & ~po037;
  assign new_new_n4521__ = ~new_new_n4519__ & ~new_new_n4520__;
  assign new_new_n4522__ = new_new_n4518__ & ~new_new_n4521__;
  assign new_new_n4523__ = ~new_new_n4518__ & new_new_n4521__;
  assign new_new_n4524__ = ~new_new_n4522__ & ~new_new_n4523__;
  assign new_new_n4525__ = pi083 & ~new_new_n4524__;
  assign new_new_n4526__ = ~pi083 & new_new_n4524__;
  assign new_new_n4527__ = ~new_new_n4242__ & ~new_new_n4243__;
  assign new_new_n4528__ = ~new_new_n4438__ & po037;
  assign new_new_n4529__ = ~pi081 & ~po037;
  assign new_new_n4530__ = ~new_new_n4528__ & ~new_new_n4529__;
  assign new_new_n4531__ = new_new_n4527__ & new_new_n4530__;
  assign new_new_n4532__ = ~new_new_n4527__ & ~new_new_n4530__;
  assign new_new_n4533__ = ~new_new_n4531__ & ~new_new_n4532__;
  assign new_new_n4534__ = ~pi082 & ~new_new_n4533__;
  assign new_new_n4535__ = pi082 & new_new_n4533__;
  assign new_new_n4536__ = ~pi080 & ~new_new_n4436__;
  assign new_new_n4537__ = pi080 & new_new_n4436__;
  assign new_new_n4538__ = ~new_new_n4536__ & ~new_new_n4537__;
  assign new_new_n4539__ = po037 & new_new_n4538__;
  assign new_new_n4540__ = new_new_n4250__ & new_new_n4539__;
  assign new_new_n4541__ = ~new_new_n4250__ & ~new_new_n4539__;
  assign new_new_n4542__ = ~new_new_n4540__ & ~new_new_n4541__;
  assign new_new_n4543__ = ~pi081 & ~new_new_n4542__;
  assign new_new_n4544__ = pi081 & new_new_n4542__;
  assign new_new_n4545__ = ~pi079 & ~new_new_n4434__;
  assign new_new_n4546__ = pi079 & new_new_n4434__;
  assign new_new_n4547__ = ~new_new_n4545__ & ~new_new_n4546__;
  assign new_new_n4548__ = po037 & new_new_n4547__;
  assign new_new_n4549__ = ~new_new_n4259__ & new_new_n4548__;
  assign new_new_n4550__ = new_new_n4259__ & ~new_new_n4548__;
  assign new_new_n4551__ = ~new_new_n4549__ & ~new_new_n4550__;
  assign new_new_n4552__ = pi080 & ~new_new_n4551__;
  assign new_new_n4553__ = ~pi080 & new_new_n4551__;
  assign new_new_n4554__ = ~new_new_n4269__ & ~new_new_n4270__;
  assign new_new_n4555__ = ~new_new_n4432__ & po037;
  assign new_new_n4556__ = ~pi078 & ~po037;
  assign new_new_n4557__ = ~new_new_n4555__ & ~new_new_n4556__;
  assign new_new_n4558__ = new_new_n4554__ & ~new_new_n4557__;
  assign new_new_n4559__ = ~new_new_n4554__ & new_new_n4557__;
  assign new_new_n4560__ = ~new_new_n4558__ & ~new_new_n4559__;
  assign new_new_n4561__ = pi079 & ~new_new_n4560__;
  assign new_new_n4562__ = ~pi079 & new_new_n4560__;
  assign new_new_n4563__ = ~new_new_n4278__ & ~new_new_n4279__;
  assign new_new_n4564__ = ~new_new_n4430__ & po037;
  assign new_new_n4565__ = ~pi077 & ~po037;
  assign new_new_n4566__ = ~new_new_n4564__ & ~new_new_n4565__;
  assign new_new_n4567__ = ~new_new_n4563__ & ~new_new_n4566__;
  assign new_new_n4568__ = new_new_n4563__ & new_new_n4566__;
  assign new_new_n4569__ = ~new_new_n4567__ & ~new_new_n4568__;
  assign new_new_n4570__ = ~pi078 & ~new_new_n4569__;
  assign new_new_n4571__ = pi078 & new_new_n4569__;
  assign new_new_n4572__ = new_new_n4428__ & po037;
  assign new_new_n4573__ = pi076 & ~po037;
  assign new_new_n4574__ = ~new_new_n4572__ & ~new_new_n4573__;
  assign new_new_n4575__ = ~new_new_n4287__ & ~new_new_n4288__;
  assign new_new_n4576__ = ~new_new_n4574__ & ~new_new_n4575__;
  assign new_new_n4577__ = new_new_n4574__ & new_new_n4575__;
  assign new_new_n4578__ = ~new_new_n4576__ & ~new_new_n4577__;
  assign new_new_n4579__ = pi077 & ~new_new_n4578__;
  assign new_new_n4580__ = ~pi077 & new_new_n4578__;
  assign new_new_n4581__ = ~new_new_n4296__ & ~new_new_n4297__;
  assign new_new_n4582__ = ~new_new_n4426__ & po037;
  assign new_new_n4583__ = ~pi075 & ~po037;
  assign new_new_n4584__ = ~new_new_n4582__ & ~new_new_n4583__;
  assign new_new_n4585__ = new_new_n4581__ & ~new_new_n4584__;
  assign new_new_n4586__ = ~new_new_n4581__ & new_new_n4584__;
  assign new_new_n4587__ = ~new_new_n4585__ & ~new_new_n4586__;
  assign new_new_n4588__ = pi076 & ~new_new_n4587__;
  assign new_new_n4589__ = ~pi076 & new_new_n4587__;
  assign new_new_n4590__ = ~new_new_n4305__ & ~new_new_n4306__;
  assign new_new_n4591__ = ~new_new_n4424__ & po037;
  assign new_new_n4592__ = ~pi074 & ~po037;
  assign new_new_n4593__ = ~new_new_n4591__ & ~new_new_n4592__;
  assign new_new_n4594__ = new_new_n4590__ & ~new_new_n4593__;
  assign new_new_n4595__ = ~new_new_n4590__ & new_new_n4593__;
  assign new_new_n4596__ = ~new_new_n4594__ & ~new_new_n4595__;
  assign new_new_n4597__ = pi075 & ~new_new_n4596__;
  assign new_new_n4598__ = ~pi075 & new_new_n4596__;
  assign new_new_n4599__ = ~new_new_n4422__ & po037;
  assign new_new_n4600__ = pi073 & ~po037;
  assign new_new_n4601__ = ~new_new_n4599__ & ~new_new_n4600__;
  assign new_new_n4602__ = ~new_new_n4314__ & ~new_new_n4315__;
  assign new_new_n4603__ = ~new_new_n4601__ & new_new_n4602__;
  assign new_new_n4604__ = new_new_n4601__ & ~new_new_n4602__;
  assign new_new_n4605__ = ~new_new_n4603__ & ~new_new_n4604__;
  assign new_new_n4606__ = pi074 & new_new_n4605__;
  assign new_new_n4607__ = ~pi074 & ~new_new_n4605__;
  assign new_new_n4608__ = ~new_new_n4323__ & ~new_new_n4324__;
  assign new_new_n4609__ = ~new_new_n4420__ & po037;
  assign new_new_n4610__ = pi072 & ~po037;
  assign new_new_n4611__ = ~new_new_n4609__ & ~new_new_n4610__;
  assign new_new_n4612__ = new_new_n4608__ & ~new_new_n4611__;
  assign new_new_n4613__ = ~new_new_n4608__ & new_new_n4611__;
  assign new_new_n4614__ = ~new_new_n4612__ & ~new_new_n4613__;
  assign new_new_n4615__ = pi073 & new_new_n4614__;
  assign new_new_n4616__ = ~pi073 & ~new_new_n4614__;
  assign new_new_n4617__ = pi071 & ~new_new_n4418__;
  assign new_new_n4618__ = ~pi071 & new_new_n4418__;
  assign new_new_n4619__ = ~new_new_n4617__ & ~new_new_n4618__;
  assign new_new_n4620__ = po037 & new_new_n4619__;
  assign new_new_n4621__ = new_new_n4331__ & new_new_n4620__;
  assign new_new_n4622__ = ~new_new_n4331__ & ~new_new_n4620__;
  assign new_new_n4623__ = ~new_new_n4621__ & ~new_new_n4622__;
  assign new_new_n4624__ = pi072 & ~new_new_n4623__;
  assign new_new_n4625__ = ~pi072 & new_new_n4623__;
  assign new_new_n4626__ = ~new_new_n4341__ & ~new_new_n4342__;
  assign new_new_n4627__ = ~new_new_n4416__ & po037;
  assign new_new_n4628__ = ~pi070 & ~po037;
  assign new_new_n4629__ = ~new_new_n4627__ & ~new_new_n4628__;
  assign new_new_n4630__ = new_new_n4626__ & ~new_new_n4629__;
  assign new_new_n4631__ = ~new_new_n4626__ & new_new_n4629__;
  assign new_new_n4632__ = ~new_new_n4630__ & ~new_new_n4631__;
  assign new_new_n4633__ = pi071 & ~new_new_n4632__;
  assign new_new_n4634__ = ~pi071 & new_new_n4632__;
  assign new_new_n4635__ = ~new_new_n4350__ & ~new_new_n4351__;
  assign new_new_n4636__ = ~new_new_n4414__ & po037;
  assign new_new_n4637__ = ~pi069 & ~po037;
  assign new_new_n4638__ = ~new_new_n4636__ & ~new_new_n4637__;
  assign new_new_n4639__ = new_new_n4635__ & ~new_new_n4638__;
  assign new_new_n4640__ = ~new_new_n4635__ & new_new_n4638__;
  assign new_new_n4641__ = ~new_new_n4639__ & ~new_new_n4640__;
  assign new_new_n4642__ = ~pi070 & new_new_n4641__;
  assign new_new_n4643__ = pi070 & ~new_new_n4641__;
  assign new_new_n4644__ = ~new_new_n4359__ & ~new_new_n4360__;
  assign new_new_n4645__ = ~new_new_n4412__ & po037;
  assign new_new_n4646__ = ~pi068 & ~po037;
  assign new_new_n4647__ = ~new_new_n4645__ & ~new_new_n4646__;
  assign new_new_n4648__ = ~new_new_n4644__ & ~new_new_n4647__;
  assign new_new_n4649__ = new_new_n4644__ & new_new_n4647__;
  assign new_new_n4650__ = ~new_new_n4648__ & ~new_new_n4649__;
  assign new_new_n4651__ = ~pi069 & ~new_new_n4650__;
  assign new_new_n4652__ = pi069 & new_new_n4650__;
  assign new_new_n4653__ = ~new_new_n4366__ & ~new_new_n4367__;
  assign new_new_n4654__ = ~new_new_n4410__ & po037;
  assign new_new_n4655__ = ~pi067 & ~po037;
  assign new_new_n4656__ = ~new_new_n4654__ & ~new_new_n4655__;
  assign new_new_n4657__ = new_new_n4653__ & ~new_new_n4656__;
  assign new_new_n4658__ = ~new_new_n4653__ & new_new_n4656__;
  assign new_new_n4659__ = ~new_new_n4657__ & ~new_new_n4658__;
  assign new_new_n4660__ = pi068 & ~new_new_n4659__;
  assign new_new_n4661__ = ~pi068 & new_new_n4659__;
  assign new_new_n4662__ = ~new_new_n4380__ & ~new_new_n4381__;
  assign new_new_n4663__ = po037 & new_new_n4662__;
  assign new_new_n4664__ = new_new_n4408__ & ~new_new_n4663__;
  assign new_new_n4665__ = ~new_new_n4408__ & new_new_n4663__;
  assign new_new_n4666__ = ~new_new_n4664__ & ~new_new_n4665__;
  assign new_new_n4667__ = pi067 & ~new_new_n4666__;
  assign new_new_n4668__ = ~pi067 & new_new_n4666__;
  assign new_new_n4669__ = pi037 & po037;
  assign new_new_n4670__ = ~pi037 & ~po037;
  assign new_new_n4671__ = ~pi065 & ~new_new_n4669__;
  assign new_new_n4672__ = ~new_new_n4670__ & new_new_n4671__;
  assign new_new_n4673__ = ~pi036 & ~new_new_n4672__;
  assign new_new_n4674__ = pi065 & new_new_n4669__;
  assign new_new_n4675__ = ~new_new_n4673__ & ~new_new_n4674__;
  assign new_new_n4676__ = pi064 & ~new_new_n4675__;
  assign new_new_n4677__ = pi064 & po037;
  assign new_new_n4678__ = ~pi037 & pi065;
  assign new_new_n4679__ = ~new_new_n4677__ & new_new_n4678__;
  assign new_new_n4680__ = ~new_new_n4676__ & ~new_new_n4679__;
  assign new_new_n4681__ = pi066 & ~new_new_n4680__;
  assign new_new_n4682__ = ~pi066 & new_new_n4680__;
  assign new_new_n4683__ = pi065 & po037;
  assign new_new_n4684__ = ~pi064 & new_new_n4683__;
  assign new_new_n4685__ = ~new_new_n4376__ & ~new_new_n4683__;
  assign new_new_n4686__ = pi037 & ~new_new_n4401__;
  assign new_new_n4687__ = ~new_new_n4685__ & new_new_n4686__;
  assign new_new_n4688__ = ~pi065 & po037;
  assign new_new_n4689__ = po038 & new_new_n4688__;
  assign new_new_n4690__ = ~po038 & ~new_new_n4688__;
  assign new_new_n4691__ = pi064 & ~new_new_n4669__;
  assign new_new_n4692__ = ~new_new_n4689__ & new_new_n4691__;
  assign new_new_n4693__ = ~new_new_n4690__ & new_new_n4692__;
  assign new_new_n4694__ = ~new_new_n4684__ & ~new_new_n4687__;
  assign new_new_n4695__ = ~new_new_n4693__ & new_new_n4694__;
  assign new_new_n4696__ = ~pi038 & ~new_new_n4695__;
  assign new_new_n4697__ = pi038 & new_new_n4695__;
  assign new_new_n4698__ = ~new_new_n4696__ & ~new_new_n4697__;
  assign new_new_n4699__ = ~new_new_n4682__ & new_new_n4698__;
  assign new_new_n4700__ = ~new_new_n4681__ & ~new_new_n4699__;
  assign new_new_n4701__ = ~new_new_n4668__ & ~new_new_n4700__;
  assign new_new_n4702__ = ~new_new_n4667__ & ~new_new_n4701__;
  assign new_new_n4703__ = ~new_new_n4661__ & ~new_new_n4702__;
  assign new_new_n4704__ = ~new_new_n4660__ & ~new_new_n4703__;
  assign new_new_n4705__ = ~new_new_n4652__ & new_new_n4704__;
  assign new_new_n4706__ = ~new_new_n4651__ & ~new_new_n4705__;
  assign new_new_n4707__ = ~new_new_n4643__ & ~new_new_n4706__;
  assign new_new_n4708__ = ~new_new_n4642__ & ~new_new_n4707__;
  assign new_new_n4709__ = ~new_new_n4634__ & new_new_n4708__;
  assign new_new_n4710__ = ~new_new_n4633__ & ~new_new_n4709__;
  assign new_new_n4711__ = ~new_new_n4625__ & ~new_new_n4710__;
  assign new_new_n4712__ = ~new_new_n4624__ & ~new_new_n4711__;
  assign new_new_n4713__ = ~new_new_n4616__ & ~new_new_n4712__;
  assign new_new_n4714__ = ~new_new_n4615__ & ~new_new_n4713__;
  assign new_new_n4715__ = ~new_new_n4607__ & ~new_new_n4714__;
  assign new_new_n4716__ = ~new_new_n4606__ & ~new_new_n4715__;
  assign new_new_n4717__ = ~new_new_n4598__ & ~new_new_n4716__;
  assign new_new_n4718__ = ~new_new_n4597__ & ~new_new_n4717__;
  assign new_new_n4719__ = ~new_new_n4589__ & ~new_new_n4718__;
  assign new_new_n4720__ = ~new_new_n4588__ & ~new_new_n4719__;
  assign new_new_n4721__ = ~new_new_n4580__ & ~new_new_n4720__;
  assign new_new_n4722__ = ~new_new_n4579__ & ~new_new_n4721__;
  assign new_new_n4723__ = ~new_new_n4571__ & new_new_n4722__;
  assign new_new_n4724__ = ~new_new_n4570__ & ~new_new_n4723__;
  assign new_new_n4725__ = ~new_new_n4562__ & new_new_n4724__;
  assign new_new_n4726__ = ~new_new_n4561__ & ~new_new_n4725__;
  assign new_new_n4727__ = ~new_new_n4553__ & ~new_new_n4726__;
  assign new_new_n4728__ = ~new_new_n4552__ & ~new_new_n4727__;
  assign new_new_n4729__ = ~new_new_n4544__ & new_new_n4728__;
  assign new_new_n4730__ = ~new_new_n4543__ & ~new_new_n4729__;
  assign new_new_n4731__ = ~new_new_n4535__ & ~new_new_n4730__;
  assign new_new_n4732__ = ~new_new_n4534__ & ~new_new_n4731__;
  assign new_new_n4733__ = ~new_new_n4526__ & new_new_n4732__;
  assign new_new_n4734__ = ~new_new_n4525__ & ~new_new_n4733__;
  assign new_new_n4735__ = ~new_new_n4517__ & ~new_new_n4734__;
  assign new_new_n4736__ = ~new_new_n4516__ & ~new_new_n4735__;
  assign new_new_n4737__ = ~new_new_n4508__ & ~new_new_n4736__;
  assign new_new_n4738__ = ~new_new_n4507__ & ~new_new_n4737__;
  assign new_new_n4739__ = ~new_new_n4499__ & new_new_n4738__;
  assign new_new_n4740__ = ~new_new_n4498__ & ~new_new_n4739__;
  assign new_new_n4741__ = ~new_new_n4490__ & ~new_new_n4740__;
  assign new_new_n4742__ = ~new_new_n4489__ & ~new_new_n4741__;
  assign new_new_n4743__ = ~new_new_n4481__ & ~new_new_n4742__;
  assign new_new_n4744__ = ~new_new_n4480__ & ~new_new_n4743__;
  assign new_new_n4745__ = new_new_n4143__ & ~new_new_n4467__;
  assign new_new_n4746__ = ~new_new_n376__ & ~new_new_n4745__;
  assign new_new_n4747__ = ~pi091 & ~new_new_n4746__;
  assign new_new_n4748__ = ~new_new_n4453__ & ~new_new_n4454__;
  assign new_new_n4749__ = po037 & new_new_n4748__;
  assign new_new_n4750__ = ~new_new_n4461__ & ~new_new_n4749__;
  assign new_new_n4751__ = new_new_n4461__ & new_new_n4749__;
  assign new_new_n4752__ = ~new_new_n4750__ & ~new_new_n4751__;
  assign new_new_n4753__ = pi089 & ~new_new_n4752__;
  assign new_new_n4754__ = ~pi089 & new_new_n4752__;
  assign new_new_n4755__ = new_new_n4744__ & ~new_new_n4754__;
  assign new_new_n4756__ = ~new_new_n4753__ & ~new_new_n4755__;
  assign new_new_n4757__ = ~pi090 & new_new_n4756__;
  assign new_new_n4758__ = ~new_new_n4186__ & ~new_new_n4187__;
  assign new_new_n4759__ = ~new_new_n4463__ & po037;
  assign new_new_n4760__ = ~pi089 & ~po037;
  assign new_new_n4761__ = ~new_new_n4759__ & ~new_new_n4760__;
  assign new_new_n4762__ = new_new_n4758__ & ~new_new_n4761__;
  assign new_new_n4763__ = ~new_new_n4758__ & new_new_n4761__;
  assign new_new_n4764__ = ~new_new_n4762__ & ~new_new_n4763__;
  assign new_new_n4765__ = ~new_new_n4757__ & ~new_new_n4764__;
  assign new_new_n4766__ = pi091 & new_new_n4746__;
  assign new_new_n4767__ = pi090 & ~new_new_n4756__;
  assign new_new_n4768__ = ~new_new_n4766__ & ~new_new_n4767__;
  assign new_new_n4769__ = ~new_new_n4765__ & new_new_n4768__;
  assign new_new_n4770__ = ~new_new_n4747__ & ~new_new_n4769__;
  assign new_new_n4771__ = ~pi094 & new_new_n3332__;
  assign new_new_n4772__ = ~pi093 & new_new_n4771__;
  assign new_new_n4773__ = ~pi092 & new_new_n4772__;
  assign po036 = ~new_new_n4770__ & new_new_n4773__;
  assign new_new_n4775__ = new_new_n4744__ & po036;
  assign new_new_n4776__ = pi089 & ~po036;
  assign new_new_n4777__ = ~new_new_n4775__ & ~new_new_n4776__;
  assign new_new_n4778__ = ~new_new_n4753__ & ~new_new_n4754__;
  assign new_new_n4779__ = ~new_new_n4777__ & ~new_new_n4778__;
  assign new_new_n4780__ = new_new_n4777__ & new_new_n4778__;
  assign new_new_n4781__ = ~new_new_n4779__ & ~new_new_n4780__;
  assign new_new_n4782__ = pi090 & ~new_new_n4781__;
  assign new_new_n4783__ = ~pi090 & new_new_n4781__;
  assign new_new_n4784__ = ~new_new_n4782__ & ~new_new_n4783__;
  assign new_new_n4785__ = ~new_new_n4480__ & ~new_new_n4481__;
  assign new_new_n4786__ = ~new_new_n4742__ & po036;
  assign new_new_n4787__ = ~pi088 & ~po036;
  assign new_new_n4788__ = ~new_new_n4786__ & ~new_new_n4787__;
  assign new_new_n4789__ = new_new_n4785__ & ~new_new_n4788__;
  assign new_new_n4790__ = ~new_new_n4785__ & new_new_n4788__;
  assign new_new_n4791__ = ~new_new_n4789__ & ~new_new_n4790__;
  assign new_new_n4792__ = pi089 & ~new_new_n4791__;
  assign new_new_n4793__ = ~pi089 & new_new_n4791__;
  assign new_new_n4794__ = ~pi087 & ~new_new_n4740__;
  assign new_new_n4795__ = pi087 & new_new_n4740__;
  assign new_new_n4796__ = ~new_new_n4794__ & ~new_new_n4795__;
  assign new_new_n4797__ = po036 & new_new_n4796__;
  assign new_new_n4798__ = ~new_new_n4488__ & new_new_n4797__;
  assign new_new_n4799__ = new_new_n4488__ & ~new_new_n4797__;
  assign new_new_n4800__ = ~new_new_n4798__ & ~new_new_n4799__;
  assign new_new_n4801__ = ~pi088 & new_new_n4800__;
  assign new_new_n4802__ = pi088 & ~new_new_n4800__;
  assign new_new_n4803__ = ~new_new_n4738__ & po036;
  assign new_new_n4804__ = pi086 & ~po036;
  assign new_new_n4805__ = ~new_new_n4803__ & ~new_new_n4804__;
  assign new_new_n4806__ = ~new_new_n4498__ & ~new_new_n4499__;
  assign new_new_n4807__ = ~new_new_n4805__ & new_new_n4806__;
  assign new_new_n4808__ = new_new_n4805__ & ~new_new_n4806__;
  assign new_new_n4809__ = ~new_new_n4807__ & ~new_new_n4808__;
  assign new_new_n4810__ = ~pi087 & ~new_new_n4809__;
  assign new_new_n4811__ = pi087 & new_new_n4809__;
  assign new_new_n4812__ = ~new_new_n4507__ & ~new_new_n4508__;
  assign new_new_n4813__ = ~new_new_n4736__ & po036;
  assign new_new_n4814__ = pi085 & ~po036;
  assign new_new_n4815__ = ~new_new_n4813__ & ~new_new_n4814__;
  assign new_new_n4816__ = new_new_n4812__ & ~new_new_n4815__;
  assign new_new_n4817__ = ~new_new_n4812__ & new_new_n4815__;
  assign new_new_n4818__ = ~new_new_n4816__ & ~new_new_n4817__;
  assign new_new_n4819__ = ~pi086 & ~new_new_n4818__;
  assign new_new_n4820__ = pi086 & new_new_n4818__;
  assign new_new_n4821__ = ~new_new_n4734__ & po036;
  assign new_new_n4822__ = pi084 & ~po036;
  assign new_new_n4823__ = ~new_new_n4821__ & ~new_new_n4822__;
  assign new_new_n4824__ = ~new_new_n4516__ & ~new_new_n4517__;
  assign new_new_n4825__ = ~new_new_n4823__ & new_new_n4824__;
  assign new_new_n4826__ = new_new_n4823__ & ~new_new_n4824__;
  assign new_new_n4827__ = ~new_new_n4825__ & ~new_new_n4826__;
  assign new_new_n4828__ = ~pi085 & ~new_new_n4827__;
  assign new_new_n4829__ = pi085 & new_new_n4827__;
  assign new_new_n4830__ = ~new_new_n4525__ & ~new_new_n4526__;
  assign new_new_n4831__ = ~new_new_n4732__ & po036;
  assign new_new_n4832__ = ~pi083 & ~po036;
  assign new_new_n4833__ = ~new_new_n4831__ & ~new_new_n4832__;
  assign new_new_n4834__ = new_new_n4830__ & ~new_new_n4833__;
  assign new_new_n4835__ = ~new_new_n4830__ & new_new_n4833__;
  assign new_new_n4836__ = ~new_new_n4834__ & ~new_new_n4835__;
  assign new_new_n4837__ = ~pi084 & new_new_n4836__;
  assign new_new_n4838__ = pi084 & ~new_new_n4836__;
  assign new_new_n4839__ = ~pi082 & ~new_new_n4730__;
  assign new_new_n4840__ = pi082 & new_new_n4730__;
  assign new_new_n4841__ = ~new_new_n4839__ & ~new_new_n4840__;
  assign new_new_n4842__ = po036 & new_new_n4841__;
  assign new_new_n4843__ = new_new_n4533__ & new_new_n4842__;
  assign new_new_n4844__ = ~new_new_n4533__ & ~new_new_n4842__;
  assign new_new_n4845__ = ~new_new_n4843__ & ~new_new_n4844__;
  assign new_new_n4846__ = ~pi083 & ~new_new_n4845__;
  assign new_new_n4847__ = pi083 & new_new_n4845__;
  assign new_new_n4848__ = ~new_new_n4543__ & ~new_new_n4544__;
  assign new_new_n4849__ = new_new_n4728__ & po036;
  assign new_new_n4850__ = ~pi081 & ~po036;
  assign new_new_n4851__ = ~new_new_n4849__ & ~new_new_n4850__;
  assign new_new_n4852__ = ~new_new_n4848__ & ~new_new_n4851__;
  assign new_new_n4853__ = new_new_n4848__ & new_new_n4851__;
  assign new_new_n4854__ = ~new_new_n4852__ & ~new_new_n4853__;
  assign new_new_n4855__ = ~pi082 & ~new_new_n4854__;
  assign new_new_n4856__ = pi082 & new_new_n4854__;
  assign new_new_n4857__ = ~new_new_n4726__ & po036;
  assign new_new_n4858__ = pi080 & ~po036;
  assign new_new_n4859__ = ~new_new_n4857__ & ~new_new_n4858__;
  assign new_new_n4860__ = ~new_new_n4552__ & ~new_new_n4553__;
  assign new_new_n4861__ = ~new_new_n4859__ & new_new_n4860__;
  assign new_new_n4862__ = new_new_n4859__ & ~new_new_n4860__;
  assign new_new_n4863__ = ~new_new_n4861__ & ~new_new_n4862__;
  assign new_new_n4864__ = pi081 & new_new_n4863__;
  assign new_new_n4865__ = ~pi081 & ~new_new_n4863__;
  assign new_new_n4866__ = ~new_new_n4561__ & ~new_new_n4562__;
  assign new_new_n4867__ = ~new_new_n4724__ & po036;
  assign new_new_n4868__ = ~pi079 & ~po036;
  assign new_new_n4869__ = ~new_new_n4867__ & ~new_new_n4868__;
  assign new_new_n4870__ = new_new_n4866__ & ~new_new_n4869__;
  assign new_new_n4871__ = ~new_new_n4866__ & new_new_n4869__;
  assign new_new_n4872__ = ~new_new_n4870__ & ~new_new_n4871__;
  assign new_new_n4873__ = pi080 & ~new_new_n4872__;
  assign new_new_n4874__ = ~pi080 & new_new_n4872__;
  assign new_new_n4875__ = ~new_new_n4722__ & po036;
  assign new_new_n4876__ = pi078 & ~po036;
  assign new_new_n4877__ = ~new_new_n4875__ & ~new_new_n4876__;
  assign new_new_n4878__ = ~new_new_n4570__ & ~new_new_n4571__;
  assign new_new_n4879__ = ~new_new_n4877__ & new_new_n4878__;
  assign new_new_n4880__ = new_new_n4877__ & ~new_new_n4878__;
  assign new_new_n4881__ = ~new_new_n4879__ & ~new_new_n4880__;
  assign new_new_n4882__ = ~pi079 & ~new_new_n4881__;
  assign new_new_n4883__ = pi079 & new_new_n4881__;
  assign new_new_n4884__ = ~new_new_n4579__ & ~new_new_n4580__;
  assign new_new_n4885__ = ~new_new_n4720__ & po036;
  assign new_new_n4886__ = pi077 & ~po036;
  assign new_new_n4887__ = ~new_new_n4885__ & ~new_new_n4886__;
  assign new_new_n4888__ = new_new_n4884__ & new_new_n4887__;
  assign new_new_n4889__ = ~new_new_n4884__ & ~new_new_n4887__;
  assign new_new_n4890__ = ~new_new_n4888__ & ~new_new_n4889__;
  assign new_new_n4891__ = pi078 & ~new_new_n4890__;
  assign new_new_n4892__ = ~pi078 & new_new_n4890__;
  assign new_new_n4893__ = pi076 & ~new_new_n4718__;
  assign new_new_n4894__ = ~pi076 & new_new_n4718__;
  assign new_new_n4895__ = ~new_new_n4893__ & ~new_new_n4894__;
  assign new_new_n4896__ = po036 & new_new_n4895__;
  assign new_new_n4897__ = new_new_n4587__ & new_new_n4896__;
  assign new_new_n4898__ = ~new_new_n4587__ & ~new_new_n4896__;
  assign new_new_n4899__ = ~new_new_n4897__ & ~new_new_n4898__;
  assign new_new_n4900__ = pi077 & ~new_new_n4899__;
  assign new_new_n4901__ = ~pi077 & new_new_n4899__;
  assign new_new_n4902__ = pi075 & ~new_new_n4716__;
  assign new_new_n4903__ = ~pi075 & new_new_n4716__;
  assign new_new_n4904__ = ~new_new_n4902__ & ~new_new_n4903__;
  assign new_new_n4905__ = po036 & new_new_n4904__;
  assign new_new_n4906__ = new_new_n4596__ & new_new_n4905__;
  assign new_new_n4907__ = ~new_new_n4596__ & ~new_new_n4905__;
  assign new_new_n4908__ = ~new_new_n4906__ & ~new_new_n4907__;
  assign new_new_n4909__ = ~pi076 & new_new_n4908__;
  assign new_new_n4910__ = pi076 & ~new_new_n4908__;
  assign new_new_n4911__ = ~new_new_n4606__ & ~new_new_n4607__;
  assign new_new_n4912__ = ~new_new_n4714__ & po036;
  assign new_new_n4913__ = pi074 & ~po036;
  assign new_new_n4914__ = ~new_new_n4912__ & ~new_new_n4913__;
  assign new_new_n4915__ = new_new_n4911__ & ~new_new_n4914__;
  assign new_new_n4916__ = ~new_new_n4911__ & new_new_n4914__;
  assign new_new_n4917__ = ~new_new_n4915__ & ~new_new_n4916__;
  assign new_new_n4918__ = ~pi075 & ~new_new_n4917__;
  assign new_new_n4919__ = pi075 & new_new_n4917__;
  assign new_new_n4920__ = ~new_new_n4615__ & ~new_new_n4616__;
  assign new_new_n4921__ = ~new_new_n4712__ & po036;
  assign new_new_n4922__ = pi073 & ~po036;
  assign new_new_n4923__ = ~new_new_n4921__ & ~new_new_n4922__;
  assign new_new_n4924__ = new_new_n4920__ & ~new_new_n4923__;
  assign new_new_n4925__ = ~new_new_n4920__ & new_new_n4923__;
  assign new_new_n4926__ = ~new_new_n4924__ & ~new_new_n4925__;
  assign new_new_n4927__ = ~pi074 & ~new_new_n4926__;
  assign new_new_n4928__ = pi074 & new_new_n4926__;
  assign new_new_n4929__ = ~new_new_n4633__ & ~new_new_n4634__;
  assign new_new_n4930__ = ~new_new_n4708__ & po036;
  assign new_new_n4931__ = ~pi071 & ~po036;
  assign new_new_n4932__ = ~new_new_n4930__ & ~new_new_n4931__;
  assign new_new_n4933__ = new_new_n4929__ & ~new_new_n4932__;
  assign new_new_n4934__ = ~new_new_n4929__ & new_new_n4932__;
  assign new_new_n4935__ = ~new_new_n4933__ & ~new_new_n4934__;
  assign new_new_n4936__ = ~pi072 & new_new_n4935__;
  assign new_new_n4937__ = pi072 & ~new_new_n4935__;
  assign new_new_n4938__ = ~new_new_n4642__ & ~new_new_n4643__;
  assign new_new_n4939__ = ~new_new_n4706__ & po036;
  assign new_new_n4940__ = ~pi070 & ~po036;
  assign new_new_n4941__ = ~new_new_n4939__ & ~new_new_n4940__;
  assign new_new_n4942__ = new_new_n4938__ & ~new_new_n4941__;
  assign new_new_n4943__ = ~new_new_n4938__ & new_new_n4941__;
  assign new_new_n4944__ = ~new_new_n4942__ & ~new_new_n4943__;
  assign new_new_n4945__ = ~pi071 & new_new_n4944__;
  assign new_new_n4946__ = pi071 & ~new_new_n4944__;
  assign new_new_n4947__ = ~new_new_n4704__ & po036;
  assign new_new_n4948__ = pi069 & ~po036;
  assign new_new_n4949__ = ~new_new_n4947__ & ~new_new_n4948__;
  assign new_new_n4950__ = ~new_new_n4651__ & ~new_new_n4652__;
  assign new_new_n4951__ = ~new_new_n4949__ & new_new_n4950__;
  assign new_new_n4952__ = new_new_n4949__ & ~new_new_n4950__;
  assign new_new_n4953__ = ~new_new_n4951__ & ~new_new_n4952__;
  assign new_new_n4954__ = ~pi070 & ~new_new_n4953__;
  assign new_new_n4955__ = pi070 & new_new_n4953__;
  assign new_new_n4956__ = pi068 & ~new_new_n4702__;
  assign new_new_n4957__ = ~pi068 & new_new_n4702__;
  assign new_new_n4958__ = ~new_new_n4956__ & ~new_new_n4957__;
  assign new_new_n4959__ = po036 & new_new_n4958__;
  assign new_new_n4960__ = new_new_n4659__ & new_new_n4959__;
  assign new_new_n4961__ = ~new_new_n4659__ & ~new_new_n4959__;
  assign new_new_n4962__ = ~new_new_n4960__ & ~new_new_n4961__;
  assign new_new_n4963__ = ~pi069 & new_new_n4962__;
  assign new_new_n4964__ = pi069 & ~new_new_n4962__;
  assign new_new_n4965__ = ~new_new_n4681__ & ~new_new_n4682__;
  assign new_new_n4966__ = po036 & new_new_n4965__;
  assign new_new_n4967__ = ~new_new_n4698__ & ~new_new_n4966__;
  assign new_new_n4968__ = new_new_n4698__ & new_new_n4966__;
  assign new_new_n4969__ = ~new_new_n4967__ & ~new_new_n4968__;
  assign new_new_n4970__ = ~pi067 & ~new_new_n4969__;
  assign new_new_n4971__ = pi067 & new_new_n4969__;
  assign new_new_n4972__ = pi036 & po036;
  assign new_new_n4973__ = ~pi036 & ~po036;
  assign new_new_n4974__ = ~pi065 & ~new_new_n4972__;
  assign new_new_n4975__ = ~new_new_n4973__ & new_new_n4974__;
  assign new_new_n4976__ = ~pi035 & ~new_new_n4975__;
  assign new_new_n4977__ = pi065 & new_new_n4972__;
  assign new_new_n4978__ = ~new_new_n4976__ & ~new_new_n4977__;
  assign new_new_n4979__ = pi064 & ~new_new_n4978__;
  assign new_new_n4980__ = pi064 & po036;
  assign new_new_n4981__ = ~pi036 & pi065;
  assign new_new_n4982__ = ~new_new_n4980__ & new_new_n4981__;
  assign new_new_n4983__ = ~new_new_n4979__ & ~new_new_n4982__;
  assign new_new_n4984__ = pi066 & ~new_new_n4983__;
  assign new_new_n4985__ = new_new_n426__ & ~po037;
  assign new_new_n4986__ = new_new_n4688__ & po036;
  assign new_new_n4987__ = ~new_new_n4985__ & ~new_new_n4986__;
  assign new_new_n4988__ = ~pi036 & ~new_new_n4987__;
  assign new_new_n4989__ = ~new_new_n332__ & po036;
  assign new_new_n4990__ = ~new_new_n4677__ & ~new_new_n4989__;
  assign new_new_n4991__ = pi065 & po036;
  assign new_new_n4992__ = po037 & ~new_new_n4991__;
  assign new_new_n4993__ = pi065 & ~new_new_n4677__;
  assign new_new_n4994__ = pi036 & ~new_new_n4993__;
  assign new_new_n4995__ = ~new_new_n4992__ & new_new_n4994__;
  assign new_new_n4996__ = ~new_new_n4988__ & ~new_new_n4990__;
  assign new_new_n4997__ = ~new_new_n4995__ & new_new_n4996__;
  assign new_new_n4998__ = ~pi037 & ~new_new_n4997__;
  assign new_new_n4999__ = ~pi064 & ~new_new_n4991__;
  assign new_new_n5000__ = ~pi065 & po036;
  assign new_new_n5001__ = ~po037 & ~new_new_n5000__;
  assign new_new_n5002__ = ~new_new_n4972__ & ~new_new_n4986__;
  assign new_new_n5003__ = ~new_new_n5001__ & new_new_n5002__;
  assign new_new_n5004__ = pi064 & ~new_new_n5003__;
  assign new_new_n5005__ = ~new_new_n4999__ & ~new_new_n5004__;
  assign new_new_n5006__ = ~new_new_n4677__ & ~new_new_n4991__;
  assign new_new_n5007__ = pi036 & ~new_new_n4683__;
  assign new_new_n5008__ = ~new_new_n5006__ & new_new_n5007__;
  assign new_new_n5009__ = ~new_new_n5005__ & ~new_new_n5008__;
  assign new_new_n5010__ = pi037 & ~new_new_n5009__;
  assign new_new_n5011__ = ~new_new_n4998__ & ~new_new_n5010__;
  assign new_new_n5012__ = ~pi066 & new_new_n4983__;
  assign new_new_n5013__ = ~new_new_n5011__ & ~new_new_n5012__;
  assign new_new_n5014__ = ~new_new_n4984__ & ~new_new_n5013__;
  assign new_new_n5015__ = ~new_new_n4971__ & new_new_n5014__;
  assign new_new_n5016__ = ~new_new_n4970__ & ~new_new_n5015__;
  assign new_new_n5017__ = ~pi068 & ~new_new_n5016__;
  assign new_new_n5018__ = pi068 & new_new_n5016__;
  assign new_new_n5019__ = ~new_new_n4700__ & po036;
  assign new_new_n5020__ = pi067 & ~po036;
  assign new_new_n5021__ = ~new_new_n5019__ & ~new_new_n5020__;
  assign new_new_n5022__ = ~new_new_n4667__ & ~new_new_n4668__;
  assign new_new_n5023__ = ~new_new_n5021__ & new_new_n5022__;
  assign new_new_n5024__ = new_new_n5021__ & ~new_new_n5022__;
  assign new_new_n5025__ = ~new_new_n5023__ & ~new_new_n5024__;
  assign new_new_n5026__ = ~new_new_n5018__ & ~new_new_n5025__;
  assign new_new_n5027__ = ~new_new_n5017__ & ~new_new_n5026__;
  assign new_new_n5028__ = ~new_new_n4964__ & ~new_new_n5027__;
  assign new_new_n5029__ = ~new_new_n4963__ & ~new_new_n5028__;
  assign new_new_n5030__ = ~new_new_n4955__ & ~new_new_n5029__;
  assign new_new_n5031__ = ~new_new_n4954__ & ~new_new_n5030__;
  assign new_new_n5032__ = ~new_new_n4946__ & ~new_new_n5031__;
  assign new_new_n5033__ = ~new_new_n4945__ & ~new_new_n5032__;
  assign new_new_n5034__ = ~new_new_n4937__ & ~new_new_n5033__;
  assign new_new_n5035__ = ~new_new_n4936__ & ~new_new_n5034__;
  assign new_new_n5036__ = ~pi073 & ~new_new_n5035__;
  assign new_new_n5037__ = pi073 & new_new_n5035__;
  assign new_new_n5038__ = ~new_new_n4624__ & ~new_new_n4625__;
  assign new_new_n5039__ = ~new_new_n4710__ & po036;
  assign new_new_n5040__ = pi072 & ~po036;
  assign new_new_n5041__ = ~new_new_n5039__ & ~new_new_n5040__;
  assign new_new_n5042__ = new_new_n5038__ & ~new_new_n5041__;
  assign new_new_n5043__ = ~new_new_n5038__ & new_new_n5041__;
  assign new_new_n5044__ = ~new_new_n5042__ & ~new_new_n5043__;
  assign new_new_n5045__ = ~new_new_n5037__ & ~new_new_n5044__;
  assign new_new_n5046__ = ~new_new_n5036__ & ~new_new_n5045__;
  assign new_new_n5047__ = ~new_new_n4928__ & ~new_new_n5046__;
  assign new_new_n5048__ = ~new_new_n4927__ & ~new_new_n5047__;
  assign new_new_n5049__ = ~new_new_n4919__ & ~new_new_n5048__;
  assign new_new_n5050__ = ~new_new_n4918__ & ~new_new_n5049__;
  assign new_new_n5051__ = ~new_new_n4910__ & ~new_new_n5050__;
  assign new_new_n5052__ = ~new_new_n4909__ & ~new_new_n5051__;
  assign new_new_n5053__ = ~new_new_n4901__ & new_new_n5052__;
  assign new_new_n5054__ = ~new_new_n4900__ & ~new_new_n5053__;
  assign new_new_n5055__ = ~new_new_n4892__ & ~new_new_n5054__;
  assign new_new_n5056__ = ~new_new_n4891__ & ~new_new_n5055__;
  assign new_new_n5057__ = ~new_new_n4883__ & new_new_n5056__;
  assign new_new_n5058__ = ~new_new_n4882__ & ~new_new_n5057__;
  assign new_new_n5059__ = ~new_new_n4874__ & new_new_n5058__;
  assign new_new_n5060__ = ~new_new_n4873__ & ~new_new_n5059__;
  assign new_new_n5061__ = ~new_new_n4865__ & ~new_new_n5060__;
  assign new_new_n5062__ = ~new_new_n4864__ & ~new_new_n5061__;
  assign new_new_n5063__ = ~new_new_n4856__ & new_new_n5062__;
  assign new_new_n5064__ = ~new_new_n4855__ & ~new_new_n5063__;
  assign new_new_n5065__ = ~new_new_n4847__ & ~new_new_n5064__;
  assign new_new_n5066__ = ~new_new_n4846__ & ~new_new_n5065__;
  assign new_new_n5067__ = ~new_new_n4838__ & ~new_new_n5066__;
  assign new_new_n5068__ = ~new_new_n4837__ & ~new_new_n5067__;
  assign new_new_n5069__ = ~new_new_n4829__ & ~new_new_n5068__;
  assign new_new_n5070__ = ~new_new_n4828__ & ~new_new_n5069__;
  assign new_new_n5071__ = ~new_new_n4820__ & ~new_new_n5070__;
  assign new_new_n5072__ = ~new_new_n4819__ & ~new_new_n5071__;
  assign new_new_n5073__ = ~new_new_n4811__ & ~new_new_n5072__;
  assign new_new_n5074__ = ~new_new_n4810__ & ~new_new_n5073__;
  assign new_new_n5075__ = ~new_new_n4802__ & ~new_new_n5074__;
  assign new_new_n5076__ = ~new_new_n4801__ & ~new_new_n5075__;
  assign new_new_n5077__ = ~new_new_n4793__ & new_new_n5076__;
  assign new_new_n5078__ = ~new_new_n4792__ & ~new_new_n5077__;
  assign new_new_n5079__ = new_new_n4745__ & ~po036;
  assign new_new_n5080__ = ~new_new_n376__ & ~new_new_n5079__;
  assign new_new_n5081__ = ~pi092 & ~new_new_n5080__;
  assign new_new_n5082__ = ~new_new_n4783__ & ~new_new_n5078__;
  assign new_new_n5083__ = ~new_new_n4782__ & ~new_new_n5082__;
  assign new_new_n5084__ = ~pi091 & new_new_n5083__;
  assign new_new_n5085__ = ~new_new_n4757__ & new_new_n4773__;
  assign new_new_n5086__ = new_new_n4768__ & new_new_n5085__;
  assign new_new_n5087__ = new_new_n4764__ & ~new_new_n5086__;
  assign new_new_n5088__ = new_new_n4747__ & new_new_n4773__;
  assign new_new_n5089__ = ~new_new_n4767__ & new_new_n5088__;
  assign new_new_n5090__ = new_new_n4765__ & new_new_n5089__;
  assign new_new_n5091__ = ~new_new_n5087__ & ~new_new_n5090__;
  assign new_new_n5092__ = ~new_new_n5084__ & new_new_n5091__;
  assign new_new_n5093__ = pi092 & new_new_n5080__;
  assign new_new_n5094__ = pi091 & ~new_new_n5083__;
  assign new_new_n5095__ = ~new_new_n5093__ & ~new_new_n5094__;
  assign new_new_n5096__ = ~new_new_n5092__ & new_new_n5095__;
  assign new_new_n5097__ = ~new_new_n5081__ & ~new_new_n5096__;
  assign po035 = new_new_n4772__ & ~new_new_n5097__;
  assign new_new_n5099__ = ~new_new_n5078__ & po035;
  assign new_new_n5100__ = pi090 & ~po035;
  assign new_new_n5101__ = ~new_new_n5099__ & ~new_new_n5100__;
  assign new_new_n5102__ = new_new_n4784__ & ~new_new_n5101__;
  assign new_new_n5103__ = ~new_new_n4784__ & new_new_n5101__;
  assign new_new_n5104__ = ~new_new_n5102__ & ~new_new_n5103__;
  assign new_new_n5105__ = ~pi091 & ~new_new_n5104__;
  assign new_new_n5106__ = pi091 & new_new_n5104__;
  assign new_new_n5107__ = ~new_new_n4792__ & ~new_new_n4793__;
  assign new_new_n5108__ = ~new_new_n5076__ & po035;
  assign new_new_n5109__ = ~pi089 & ~po035;
  assign new_new_n5110__ = ~new_new_n5108__ & ~new_new_n5109__;
  assign new_new_n5111__ = new_new_n5107__ & ~new_new_n5110__;
  assign new_new_n5112__ = ~new_new_n5107__ & new_new_n5110__;
  assign new_new_n5113__ = ~new_new_n5111__ & ~new_new_n5112__;
  assign new_new_n5114__ = ~pi090 & new_new_n5113__;
  assign new_new_n5115__ = pi090 & ~new_new_n5113__;
  assign new_new_n5116__ = ~new_new_n4801__ & ~new_new_n4802__;
  assign new_new_n5117__ = ~new_new_n5074__ & po035;
  assign new_new_n5118__ = ~pi088 & ~po035;
  assign new_new_n5119__ = ~new_new_n5117__ & ~new_new_n5118__;
  assign new_new_n5120__ = new_new_n5116__ & ~new_new_n5119__;
  assign new_new_n5121__ = ~new_new_n5116__ & new_new_n5119__;
  assign new_new_n5122__ = ~new_new_n5120__ & ~new_new_n5121__;
  assign new_new_n5123__ = ~pi089 & new_new_n5122__;
  assign new_new_n5124__ = pi089 & ~new_new_n5122__;
  assign new_new_n5125__ = ~pi087 & ~new_new_n5072__;
  assign new_new_n5126__ = pi087 & new_new_n5072__;
  assign new_new_n5127__ = ~new_new_n5125__ & ~new_new_n5126__;
  assign new_new_n5128__ = po035 & new_new_n5127__;
  assign new_new_n5129__ = new_new_n4809__ & new_new_n5128__;
  assign new_new_n5130__ = ~new_new_n4809__ & ~new_new_n5128__;
  assign new_new_n5131__ = ~new_new_n5129__ & ~new_new_n5130__;
  assign new_new_n5132__ = ~pi088 & ~new_new_n5131__;
  assign new_new_n5133__ = pi088 & new_new_n5131__;
  assign new_new_n5134__ = ~new_new_n4819__ & ~new_new_n4820__;
  assign new_new_n5135__ = ~new_new_n5070__ & po035;
  assign new_new_n5136__ = ~pi086 & ~po035;
  assign new_new_n5137__ = ~new_new_n5135__ & ~new_new_n5136__;
  assign new_new_n5138__ = new_new_n5134__ & ~new_new_n5137__;
  assign new_new_n5139__ = ~new_new_n5134__ & new_new_n5137__;
  assign new_new_n5140__ = ~new_new_n5138__ & ~new_new_n5139__;
  assign new_new_n5141__ = pi087 & ~new_new_n5140__;
  assign new_new_n5142__ = ~pi087 & new_new_n5140__;
  assign new_new_n5143__ = ~new_new_n4828__ & ~new_new_n4829__;
  assign new_new_n5144__ = ~new_new_n5068__ & po035;
  assign new_new_n5145__ = ~pi085 & ~po035;
  assign new_new_n5146__ = ~new_new_n5144__ & ~new_new_n5145__;
  assign new_new_n5147__ = ~new_new_n5143__ & ~new_new_n5146__;
  assign new_new_n5148__ = new_new_n5143__ & new_new_n5146__;
  assign new_new_n5149__ = ~new_new_n5147__ & ~new_new_n5148__;
  assign new_new_n5150__ = ~pi086 & ~new_new_n5149__;
  assign new_new_n5151__ = pi086 & new_new_n5149__;
  assign new_new_n5152__ = new_new_n5066__ & po035;
  assign new_new_n5153__ = pi084 & ~po035;
  assign new_new_n5154__ = ~new_new_n5152__ & ~new_new_n5153__;
  assign new_new_n5155__ = ~new_new_n4837__ & ~new_new_n4838__;
  assign new_new_n5156__ = ~new_new_n5154__ & ~new_new_n5155__;
  assign new_new_n5157__ = new_new_n5154__ & new_new_n5155__;
  assign new_new_n5158__ = ~new_new_n5156__ & ~new_new_n5157__;
  assign new_new_n5159__ = pi085 & ~new_new_n5158__;
  assign new_new_n5160__ = ~pi085 & new_new_n5158__;
  assign new_new_n5161__ = ~new_new_n4846__ & ~new_new_n4847__;
  assign new_new_n5162__ = ~new_new_n5064__ & po035;
  assign new_new_n5163__ = ~pi083 & ~po035;
  assign new_new_n5164__ = ~new_new_n5162__ & ~new_new_n5163__;
  assign new_new_n5165__ = new_new_n5161__ & ~new_new_n5164__;
  assign new_new_n5166__ = ~new_new_n5161__ & new_new_n5164__;
  assign new_new_n5167__ = ~new_new_n5165__ & ~new_new_n5166__;
  assign new_new_n5168__ = ~pi084 & new_new_n5167__;
  assign new_new_n5169__ = pi084 & ~new_new_n5167__;
  assign new_new_n5170__ = new_new_n5062__ & po035;
  assign new_new_n5171__ = ~pi082 & ~po035;
  assign new_new_n5172__ = ~new_new_n5170__ & ~new_new_n5171__;
  assign new_new_n5173__ = ~new_new_n4855__ & ~new_new_n4856__;
  assign new_new_n5174__ = ~new_new_n5172__ & ~new_new_n5173__;
  assign new_new_n5175__ = new_new_n5172__ & new_new_n5173__;
  assign new_new_n5176__ = ~new_new_n5174__ & ~new_new_n5175__;
  assign new_new_n5177__ = ~pi083 & ~new_new_n5176__;
  assign new_new_n5178__ = pi083 & new_new_n5176__;
  assign new_new_n5179__ = ~new_new_n5060__ & po035;
  assign new_new_n5180__ = pi081 & ~po035;
  assign new_new_n5181__ = ~new_new_n5179__ & ~new_new_n5180__;
  assign new_new_n5182__ = ~new_new_n4864__ & ~new_new_n4865__;
  assign new_new_n5183__ = ~new_new_n5181__ & new_new_n5182__;
  assign new_new_n5184__ = new_new_n5181__ & ~new_new_n5182__;
  assign new_new_n5185__ = ~new_new_n5183__ & ~new_new_n5184__;
  assign new_new_n5186__ = ~pi082 & ~new_new_n5185__;
  assign new_new_n5187__ = pi082 & new_new_n5185__;
  assign new_new_n5188__ = ~new_new_n4873__ & ~new_new_n4874__;
  assign new_new_n5189__ = ~new_new_n5058__ & po035;
  assign new_new_n5190__ = ~pi080 & ~po035;
  assign new_new_n5191__ = ~new_new_n5189__ & ~new_new_n5190__;
  assign new_new_n5192__ = new_new_n5188__ & ~new_new_n5191__;
  assign new_new_n5193__ = ~new_new_n5188__ & new_new_n5191__;
  assign new_new_n5194__ = ~new_new_n5192__ & ~new_new_n5193__;
  assign new_new_n5195__ = ~pi081 & new_new_n5194__;
  assign new_new_n5196__ = pi081 & ~new_new_n5194__;
  assign new_new_n5197__ = ~new_new_n5056__ & po035;
  assign new_new_n5198__ = pi079 & ~po035;
  assign new_new_n5199__ = ~new_new_n5197__ & ~new_new_n5198__;
  assign new_new_n5200__ = ~new_new_n4882__ & ~new_new_n4883__;
  assign new_new_n5201__ = ~new_new_n5199__ & new_new_n5200__;
  assign new_new_n5202__ = new_new_n5199__ & ~new_new_n5200__;
  assign new_new_n5203__ = ~new_new_n5201__ & ~new_new_n5202__;
  assign new_new_n5204__ = ~pi080 & ~new_new_n5203__;
  assign new_new_n5205__ = pi080 & new_new_n5203__;
  assign new_new_n5206__ = pi078 & ~new_new_n5054__;
  assign new_new_n5207__ = ~pi078 & new_new_n5054__;
  assign new_new_n5208__ = ~new_new_n5206__ & ~new_new_n5207__;
  assign new_new_n5209__ = po035 & new_new_n5208__;
  assign new_new_n5210__ = new_new_n4890__ & new_new_n5209__;
  assign new_new_n5211__ = ~new_new_n4890__ & ~new_new_n5209__;
  assign new_new_n5212__ = ~new_new_n5210__ & ~new_new_n5211__;
  assign new_new_n5213__ = pi079 & ~new_new_n5212__;
  assign new_new_n5214__ = ~pi079 & new_new_n5212__;
  assign new_new_n5215__ = ~new_new_n4900__ & ~new_new_n4901__;
  assign new_new_n5216__ = ~new_new_n5052__ & po035;
  assign new_new_n5217__ = ~pi077 & ~po035;
  assign new_new_n5218__ = ~new_new_n5216__ & ~new_new_n5217__;
  assign new_new_n5219__ = new_new_n5215__ & ~new_new_n5218__;
  assign new_new_n5220__ = ~new_new_n5215__ & new_new_n5218__;
  assign new_new_n5221__ = ~new_new_n5219__ & ~new_new_n5220__;
  assign new_new_n5222__ = pi078 & ~new_new_n5221__;
  assign new_new_n5223__ = ~pi078 & new_new_n5221__;
  assign new_new_n5224__ = ~new_new_n4909__ & ~new_new_n4910__;
  assign new_new_n5225__ = ~new_new_n5050__ & po035;
  assign new_new_n5226__ = ~pi076 & ~po035;
  assign new_new_n5227__ = ~new_new_n5225__ & ~new_new_n5226__;
  assign new_new_n5228__ = new_new_n5224__ & ~new_new_n5227__;
  assign new_new_n5229__ = ~new_new_n5224__ & new_new_n5227__;
  assign new_new_n5230__ = ~new_new_n5228__ & ~new_new_n5229__;
  assign new_new_n5231__ = pi077 & ~new_new_n5230__;
  assign new_new_n5232__ = ~pi077 & new_new_n5230__;
  assign new_new_n5233__ = ~pi075 & ~new_new_n5048__;
  assign new_new_n5234__ = pi075 & new_new_n5048__;
  assign new_new_n5235__ = ~new_new_n5233__ & ~new_new_n5234__;
  assign new_new_n5236__ = po035 & new_new_n5235__;
  assign new_new_n5237__ = new_new_n4917__ & new_new_n5236__;
  assign new_new_n5238__ = ~new_new_n4917__ & ~new_new_n5236__;
  assign new_new_n5239__ = ~new_new_n5237__ & ~new_new_n5238__;
  assign new_new_n5240__ = ~pi076 & ~new_new_n5239__;
  assign new_new_n5241__ = pi076 & new_new_n5239__;
  assign new_new_n5242__ = ~pi074 & ~new_new_n5046__;
  assign new_new_n5243__ = pi074 & new_new_n5046__;
  assign new_new_n5244__ = ~new_new_n5242__ & ~new_new_n5243__;
  assign new_new_n5245__ = po035 & new_new_n5244__;
  assign new_new_n5246__ = new_new_n4926__ & new_new_n5245__;
  assign new_new_n5247__ = ~new_new_n4926__ & ~new_new_n5245__;
  assign new_new_n5248__ = ~new_new_n5246__ & ~new_new_n5247__;
  assign new_new_n5249__ = pi075 & new_new_n5248__;
  assign new_new_n5250__ = ~pi075 & ~new_new_n5248__;
  assign new_new_n5251__ = ~new_new_n5036__ & ~new_new_n5037__;
  assign new_new_n5252__ = po035 & new_new_n5251__;
  assign new_new_n5253__ = new_new_n5044__ & new_new_n5252__;
  assign new_new_n5254__ = ~new_new_n5044__ & ~new_new_n5252__;
  assign new_new_n5255__ = ~new_new_n5253__ & ~new_new_n5254__;
  assign new_new_n5256__ = pi074 & new_new_n5255__;
  assign new_new_n5257__ = ~pi074 & ~new_new_n5255__;
  assign new_new_n5258__ = ~new_new_n4936__ & ~new_new_n4937__;
  assign new_new_n5259__ = ~new_new_n5033__ & po035;
  assign new_new_n5260__ = ~pi072 & ~po035;
  assign new_new_n5261__ = ~new_new_n5259__ & ~new_new_n5260__;
  assign new_new_n5262__ = new_new_n5258__ & ~new_new_n5261__;
  assign new_new_n5263__ = ~new_new_n5258__ & new_new_n5261__;
  assign new_new_n5264__ = ~new_new_n5262__ & ~new_new_n5263__;
  assign new_new_n5265__ = pi073 & ~new_new_n5264__;
  assign new_new_n5266__ = ~pi073 & new_new_n5264__;
  assign new_new_n5267__ = ~new_new_n4945__ & ~new_new_n4946__;
  assign new_new_n5268__ = ~new_new_n5031__ & po035;
  assign new_new_n5269__ = ~pi071 & ~po035;
  assign new_new_n5270__ = ~new_new_n5268__ & ~new_new_n5269__;
  assign new_new_n5271__ = new_new_n5267__ & ~new_new_n5270__;
  assign new_new_n5272__ = ~new_new_n5267__ & new_new_n5270__;
  assign new_new_n5273__ = ~new_new_n5271__ & ~new_new_n5272__;
  assign new_new_n5274__ = pi072 & ~new_new_n5273__;
  assign new_new_n5275__ = ~pi072 & new_new_n5273__;
  assign new_new_n5276__ = ~pi070 & ~new_new_n5029__;
  assign new_new_n5277__ = pi070 & new_new_n5029__;
  assign new_new_n5278__ = ~new_new_n5276__ & ~new_new_n5277__;
  assign new_new_n5279__ = po035 & new_new_n5278__;
  assign new_new_n5280__ = new_new_n4953__ & new_new_n5279__;
  assign new_new_n5281__ = ~new_new_n4953__ & ~new_new_n5279__;
  assign new_new_n5282__ = ~new_new_n5280__ & ~new_new_n5281__;
  assign new_new_n5283__ = ~pi071 & ~new_new_n5282__;
  assign new_new_n5284__ = pi071 & new_new_n5282__;
  assign new_new_n5285__ = ~new_new_n4963__ & ~new_new_n4964__;
  assign new_new_n5286__ = ~new_new_n5027__ & po035;
  assign new_new_n5287__ = ~pi069 & ~po035;
  assign new_new_n5288__ = ~new_new_n5286__ & ~new_new_n5287__;
  assign new_new_n5289__ = new_new_n5285__ & ~new_new_n5288__;
  assign new_new_n5290__ = ~new_new_n5285__ & new_new_n5288__;
  assign new_new_n5291__ = ~new_new_n5289__ & ~new_new_n5290__;
  assign new_new_n5292__ = pi070 & ~new_new_n5291__;
  assign new_new_n5293__ = ~pi070 & new_new_n5291__;
  assign new_new_n5294__ = ~new_new_n5017__ & ~new_new_n5018__;
  assign new_new_n5295__ = po035 & new_new_n5294__;
  assign new_new_n5296__ = ~new_new_n5025__ & ~new_new_n5295__;
  assign new_new_n5297__ = new_new_n5025__ & new_new_n5295__;
  assign new_new_n5298__ = ~new_new_n5296__ & ~new_new_n5297__;
  assign new_new_n5299__ = ~pi069 & ~new_new_n5298__;
  assign new_new_n5300__ = pi069 & new_new_n5298__;
  assign new_new_n5301__ = ~new_new_n4970__ & ~new_new_n4971__;
  assign new_new_n5302__ = ~new_new_n5014__ & po035;
  assign new_new_n5303__ = pi067 & ~po035;
  assign new_new_n5304__ = ~new_new_n5302__ & ~new_new_n5303__;
  assign new_new_n5305__ = new_new_n5301__ & ~new_new_n5304__;
  assign new_new_n5306__ = ~new_new_n5301__ & new_new_n5304__;
  assign new_new_n5307__ = ~new_new_n5305__ & ~new_new_n5306__;
  assign new_new_n5308__ = ~pi068 & ~new_new_n5307__;
  assign new_new_n5309__ = pi068 & new_new_n5307__;
  assign new_new_n5310__ = ~new_new_n4984__ & po035;
  assign new_new_n5311__ = ~new_new_n5012__ & new_new_n5310__;
  assign new_new_n5312__ = new_new_n5011__ & ~new_new_n5311__;
  assign new_new_n5313__ = new_new_n5013__ & new_new_n5310__;
  assign new_new_n5314__ = ~new_new_n5312__ & ~new_new_n5313__;
  assign new_new_n5315__ = ~pi067 & ~new_new_n5314__;
  assign new_new_n5316__ = pi067 & new_new_n5314__;
  assign new_new_n5317__ = pi035 & po035;
  assign new_new_n5318__ = ~pi035 & ~po035;
  assign new_new_n5319__ = ~new_new_n5317__ & ~new_new_n5318__;
  assign new_new_n5320__ = ~pi034 & ~new_new_n5319__;
  assign new_new_n5321__ = ~pi034 & pi065;
  assign new_new_n5322__ = pi065 & new_new_n5317__;
  assign new_new_n5323__ = ~new_new_n5321__ & ~new_new_n5322__;
  assign new_new_n5324__ = ~new_new_n5320__ & new_new_n5323__;
  assign new_new_n5325__ = pi064 & ~new_new_n5324__;
  assign new_new_n5326__ = pi064 & po035;
  assign new_new_n5327__ = ~pi035 & pi065;
  assign new_new_n5328__ = ~new_new_n5326__ & new_new_n5327__;
  assign new_new_n5329__ = ~new_new_n5325__ & ~new_new_n5328__;
  assign new_new_n5330__ = ~pi066 & new_new_n5329__;
  assign new_new_n5331__ = pi066 & ~new_new_n5329__;
  assign new_new_n5332__ = new_new_n426__ & ~po036;
  assign new_new_n5333__ = new_new_n5000__ & po035;
  assign new_new_n5334__ = ~new_new_n5332__ & ~new_new_n5333__;
  assign new_new_n5335__ = ~pi035 & ~new_new_n5334__;
  assign new_new_n5336__ = ~new_new_n332__ & po035;
  assign new_new_n5337__ = ~new_new_n4980__ & ~new_new_n5336__;
  assign new_new_n5338__ = pi065 & po035;
  assign new_new_n5339__ = po036 & ~new_new_n5338__;
  assign new_new_n5340__ = pi065 & ~new_new_n4980__;
  assign new_new_n5341__ = pi035 & ~new_new_n5340__;
  assign new_new_n5342__ = ~new_new_n5339__ & new_new_n5341__;
  assign new_new_n5343__ = ~new_new_n5335__ & ~new_new_n5337__;
  assign new_new_n5344__ = ~new_new_n5342__ & new_new_n5343__;
  assign new_new_n5345__ = pi036 & ~new_new_n5344__;
  assign new_new_n5346__ = ~new_new_n4980__ & ~new_new_n5338__;
  assign new_new_n5347__ = pi035 & ~new_new_n4991__;
  assign new_new_n5348__ = pi064 & ~new_new_n5347__;
  assign new_new_n5349__ = ~new_new_n5346__ & ~new_new_n5348__;
  assign new_new_n5350__ = ~pi065 & po035;
  assign new_new_n5351__ = ~po036 & ~new_new_n5350__;
  assign new_new_n5352__ = pi064 & ~new_new_n5317__;
  assign new_new_n5353__ = ~new_new_n5333__ & new_new_n5352__;
  assign new_new_n5354__ = ~new_new_n5351__ & new_new_n5353__;
  assign new_new_n5355__ = ~new_new_n5349__ & ~new_new_n5354__;
  assign new_new_n5356__ = ~pi036 & ~new_new_n5355__;
  assign new_new_n5357__ = ~new_new_n5345__ & ~new_new_n5356__;
  assign new_new_n5358__ = ~new_new_n5331__ & ~new_new_n5357__;
  assign new_new_n5359__ = ~new_new_n5330__ & ~new_new_n5358__;
  assign new_new_n5360__ = ~new_new_n5316__ & ~new_new_n5359__;
  assign new_new_n5361__ = ~new_new_n5315__ & ~new_new_n5360__;
  assign new_new_n5362__ = ~new_new_n5309__ & ~new_new_n5361__;
  assign new_new_n5363__ = ~new_new_n5308__ & ~new_new_n5362__;
  assign new_new_n5364__ = ~new_new_n5300__ & ~new_new_n5363__;
  assign new_new_n5365__ = ~new_new_n5299__ & ~new_new_n5364__;
  assign new_new_n5366__ = ~new_new_n5293__ & new_new_n5365__;
  assign new_new_n5367__ = ~new_new_n5292__ & ~new_new_n5366__;
  assign new_new_n5368__ = ~new_new_n5284__ & new_new_n5367__;
  assign new_new_n5369__ = ~new_new_n5283__ & ~new_new_n5368__;
  assign new_new_n5370__ = ~new_new_n5275__ & new_new_n5369__;
  assign new_new_n5371__ = ~new_new_n5274__ & ~new_new_n5370__;
  assign new_new_n5372__ = ~new_new_n5266__ & ~new_new_n5371__;
  assign new_new_n5373__ = ~new_new_n5265__ & ~new_new_n5372__;
  assign new_new_n5374__ = ~new_new_n5257__ & ~new_new_n5373__;
  assign new_new_n5375__ = ~new_new_n5256__ & ~new_new_n5374__;
  assign new_new_n5376__ = ~new_new_n5250__ & ~new_new_n5375__;
  assign new_new_n5377__ = ~new_new_n5249__ & ~new_new_n5376__;
  assign new_new_n5378__ = ~new_new_n5241__ & new_new_n5377__;
  assign new_new_n5379__ = ~new_new_n5240__ & ~new_new_n5378__;
  assign new_new_n5380__ = ~new_new_n5232__ & new_new_n5379__;
  assign new_new_n5381__ = ~new_new_n5231__ & ~new_new_n5380__;
  assign new_new_n5382__ = ~new_new_n5223__ & ~new_new_n5381__;
  assign new_new_n5383__ = ~new_new_n5222__ & ~new_new_n5382__;
  assign new_new_n5384__ = ~new_new_n5214__ & ~new_new_n5383__;
  assign new_new_n5385__ = ~new_new_n5213__ & ~new_new_n5384__;
  assign new_new_n5386__ = ~new_new_n5205__ & new_new_n5385__;
  assign new_new_n5387__ = ~new_new_n5204__ & ~new_new_n5386__;
  assign new_new_n5388__ = ~new_new_n5196__ & ~new_new_n5387__;
  assign new_new_n5389__ = ~new_new_n5195__ & ~new_new_n5388__;
  assign new_new_n5390__ = ~new_new_n5187__ & ~new_new_n5389__;
  assign new_new_n5391__ = ~new_new_n5186__ & ~new_new_n5390__;
  assign new_new_n5392__ = ~new_new_n5178__ & ~new_new_n5391__;
  assign new_new_n5393__ = ~new_new_n5177__ & ~new_new_n5392__;
  assign new_new_n5394__ = ~new_new_n5169__ & ~new_new_n5393__;
  assign new_new_n5395__ = ~new_new_n5168__ & ~new_new_n5394__;
  assign new_new_n5396__ = ~new_new_n5160__ & new_new_n5395__;
  assign new_new_n5397__ = ~new_new_n5159__ & ~new_new_n5396__;
  assign new_new_n5398__ = ~new_new_n5151__ & new_new_n5397__;
  assign new_new_n5399__ = ~new_new_n5150__ & ~new_new_n5398__;
  assign new_new_n5400__ = ~new_new_n5142__ & new_new_n5399__;
  assign new_new_n5401__ = ~new_new_n5141__ & ~new_new_n5400__;
  assign new_new_n5402__ = ~new_new_n5133__ & new_new_n5401__;
  assign new_new_n5403__ = ~new_new_n5132__ & ~new_new_n5402__;
  assign new_new_n5404__ = ~new_new_n5124__ & ~new_new_n5403__;
  assign new_new_n5405__ = ~new_new_n5123__ & ~new_new_n5404__;
  assign new_new_n5406__ = ~new_new_n5115__ & ~new_new_n5405__;
  assign new_new_n5407__ = ~new_new_n5114__ & ~new_new_n5406__;
  assign new_new_n5408__ = ~new_new_n5106__ & ~new_new_n5407__;
  assign new_new_n5409__ = ~new_new_n5105__ & ~new_new_n5408__;
  assign new_new_n5410__ = ~pi092 & ~new_new_n5409__;
  assign new_new_n5411__ = pi092 & new_new_n5409__;
  assign new_new_n5412__ = ~new_new_n5410__ & ~new_new_n5411__;
  assign new_new_n5413__ = ~new_new_n376__ & po035;
  assign new_new_n5414__ = ~new_new_n5080__ & ~new_new_n5413__;
  assign new_new_n5415__ = pi093 & ~new_new_n5414__;
  assign new_new_n5416__ = new_new_n4771__ & ~new_new_n5415__;
  assign new_new_n5417__ = new_new_n5412__ & new_new_n5416__;
  assign new_new_n5418__ = new_new_n4772__ & ~new_new_n5084__;
  assign new_new_n5419__ = new_new_n5095__ & new_new_n5418__;
  assign new_new_n5420__ = ~new_new_n5091__ & ~new_new_n5419__;
  assign new_new_n5421__ = new_new_n5081__ & new_new_n5091__;
  assign new_new_n5422__ = ~new_new_n5094__ & new_new_n5421__;
  assign new_new_n5423__ = new_new_n5418__ & new_new_n5422__;
  assign new_new_n5424__ = ~new_new_n5420__ & ~new_new_n5423__;
  assign new_new_n5425__ = ~new_new_n5417__ & ~new_new_n5424__;
  assign new_new_n5426__ = ~pi093 & new_new_n5414__;
  assign new_new_n5427__ = new_new_n4771__ & new_new_n5426__;
  assign new_new_n5428__ = new_new_n5424__ & new_new_n5427__;
  assign new_new_n5429__ = new_new_n5412__ & new_new_n5428__;
  assign new_new_n5430__ = ~new_new_n5425__ & ~new_new_n5429__;
  assign new_new_n5431__ = ~pi093 & ~new_new_n5430__;
  assign new_new_n5432__ = pi093 & new_new_n5430__;
  assign new_new_n5433__ = ~new_new_n5431__ & ~new_new_n5432__;
  assign new_new_n5434__ = ~new_new_n5410__ & new_new_n5424__;
  assign new_new_n5435__ = new_new_n5416__ & ~new_new_n5426__;
  assign new_new_n5436__ = ~new_new_n5411__ & new_new_n5435__;
  assign new_new_n5437__ = ~new_new_n5434__ & new_new_n5436__;
  assign po034 = new_new_n5427__ | new_new_n5437__;
  assign new_new_n5439__ = ~pi091 & ~new_new_n5407__;
  assign new_new_n5440__ = pi091 & new_new_n5407__;
  assign new_new_n5441__ = ~new_new_n5439__ & ~new_new_n5440__;
  assign new_new_n5442__ = po034 & new_new_n5441__;
  assign new_new_n5443__ = new_new_n5104__ & new_new_n5442__;
  assign new_new_n5444__ = ~new_new_n5104__ & ~new_new_n5442__;
  assign new_new_n5445__ = ~new_new_n5443__ & ~new_new_n5444__;
  assign new_new_n5446__ = pi092 & new_new_n5445__;
  assign new_new_n5447__ = ~pi092 & ~new_new_n5445__;
  assign new_new_n5448__ = ~new_new_n5114__ & ~new_new_n5115__;
  assign new_new_n5449__ = ~pi090 & ~po034;
  assign new_new_n5450__ = ~new_new_n5405__ & po034;
  assign new_new_n5451__ = ~new_new_n5449__ & ~new_new_n5450__;
  assign new_new_n5452__ = new_new_n5448__ & ~new_new_n5451__;
  assign new_new_n5453__ = ~new_new_n5448__ & new_new_n5451__;
  assign new_new_n5454__ = ~new_new_n5452__ & ~new_new_n5453__;
  assign new_new_n5455__ = pi091 & ~new_new_n5454__;
  assign new_new_n5456__ = ~new_new_n5123__ & ~new_new_n5124__;
  assign new_new_n5457__ = ~pi089 & ~po034;
  assign new_new_n5458__ = ~new_new_n5403__ & po034;
  assign new_new_n5459__ = ~new_new_n5457__ & ~new_new_n5458__;
  assign new_new_n5460__ = new_new_n5456__ & ~new_new_n5459__;
  assign new_new_n5461__ = ~new_new_n5456__ & new_new_n5459__;
  assign new_new_n5462__ = ~new_new_n5460__ & ~new_new_n5461__;
  assign new_new_n5463__ = pi090 & ~new_new_n5462__;
  assign new_new_n5464__ = ~pi090 & new_new_n5462__;
  assign new_new_n5465__ = ~new_new_n5132__ & ~new_new_n5133__;
  assign new_new_n5466__ = ~pi088 & ~po034;
  assign new_new_n5467__ = new_new_n5401__ & po034;
  assign new_new_n5468__ = ~new_new_n5466__ & ~new_new_n5467__;
  assign new_new_n5469__ = new_new_n5465__ & ~new_new_n5468__;
  assign new_new_n5470__ = ~new_new_n5465__ & new_new_n5468__;
  assign new_new_n5471__ = ~new_new_n5469__ & ~new_new_n5470__;
  assign new_new_n5472__ = pi089 & ~new_new_n5471__;
  assign new_new_n5473__ = ~pi089 & new_new_n5471__;
  assign new_new_n5474__ = new_new_n5399__ & po034;
  assign new_new_n5475__ = pi087 & ~po034;
  assign new_new_n5476__ = ~new_new_n5474__ & ~new_new_n5475__;
  assign new_new_n5477__ = ~new_new_n5141__ & ~new_new_n5142__;
  assign new_new_n5478__ = ~new_new_n5476__ & ~new_new_n5477__;
  assign new_new_n5479__ = new_new_n5476__ & new_new_n5477__;
  assign new_new_n5480__ = ~new_new_n5478__ & ~new_new_n5479__;
  assign new_new_n5481__ = pi088 & ~new_new_n5480__;
  assign new_new_n5482__ = ~pi088 & new_new_n5480__;
  assign new_new_n5483__ = ~new_new_n5150__ & ~new_new_n5151__;
  assign new_new_n5484__ = new_new_n5397__ & po034;
  assign new_new_n5485__ = ~pi086 & ~po034;
  assign new_new_n5486__ = ~new_new_n5484__ & ~new_new_n5485__;
  assign new_new_n5487__ = ~new_new_n5483__ & ~new_new_n5486__;
  assign new_new_n5488__ = new_new_n5483__ & new_new_n5486__;
  assign new_new_n5489__ = ~new_new_n5487__ & ~new_new_n5488__;
  assign new_new_n5490__ = pi087 & new_new_n5489__;
  assign new_new_n5491__ = ~pi087 & ~new_new_n5489__;
  assign new_new_n5492__ = ~new_new_n5159__ & ~new_new_n5160__;
  assign new_new_n5493__ = ~new_new_n5395__ & po034;
  assign new_new_n5494__ = ~pi085 & ~po034;
  assign new_new_n5495__ = ~new_new_n5493__ & ~new_new_n5494__;
  assign new_new_n5496__ = new_new_n5492__ & new_new_n5495__;
  assign new_new_n5497__ = ~new_new_n5492__ & ~new_new_n5495__;
  assign new_new_n5498__ = ~new_new_n5496__ & ~new_new_n5497__;
  assign new_new_n5499__ = pi086 & new_new_n5498__;
  assign new_new_n5500__ = ~pi086 & ~new_new_n5498__;
  assign new_new_n5501__ = new_new_n5393__ & po034;
  assign new_new_n5502__ = pi084 & ~po034;
  assign new_new_n5503__ = ~new_new_n5501__ & ~new_new_n5502__;
  assign new_new_n5504__ = ~new_new_n5168__ & ~new_new_n5169__;
  assign new_new_n5505__ = ~new_new_n5503__ & ~new_new_n5504__;
  assign new_new_n5506__ = new_new_n5503__ & new_new_n5504__;
  assign new_new_n5507__ = ~new_new_n5505__ & ~new_new_n5506__;
  assign new_new_n5508__ = pi085 & ~new_new_n5507__;
  assign new_new_n5509__ = ~pi085 & new_new_n5507__;
  assign new_new_n5510__ = ~pi083 & ~new_new_n5391__;
  assign new_new_n5511__ = pi083 & new_new_n5391__;
  assign new_new_n5512__ = ~new_new_n5510__ & ~new_new_n5511__;
  assign new_new_n5513__ = po034 & new_new_n5512__;
  assign new_new_n5514__ = new_new_n5176__ & new_new_n5513__;
  assign new_new_n5515__ = ~new_new_n5176__ & ~new_new_n5513__;
  assign new_new_n5516__ = ~new_new_n5514__ & ~new_new_n5515__;
  assign new_new_n5517__ = ~pi084 & ~new_new_n5516__;
  assign new_new_n5518__ = pi084 & new_new_n5516__;
  assign new_new_n5519__ = ~new_new_n5186__ & ~new_new_n5187__;
  assign new_new_n5520__ = ~new_new_n5389__ & po034;
  assign new_new_n5521__ = ~pi082 & ~po034;
  assign new_new_n5522__ = ~new_new_n5520__ & ~new_new_n5521__;
  assign new_new_n5523__ = ~new_new_n5519__ & ~new_new_n5522__;
  assign new_new_n5524__ = new_new_n5519__ & new_new_n5522__;
  assign new_new_n5525__ = ~new_new_n5523__ & ~new_new_n5524__;
  assign new_new_n5526__ = ~pi083 & ~new_new_n5525__;
  assign new_new_n5527__ = pi083 & new_new_n5525__;
  assign new_new_n5528__ = new_new_n5387__ & po034;
  assign new_new_n5529__ = pi081 & ~po034;
  assign new_new_n5530__ = ~new_new_n5528__ & ~new_new_n5529__;
  assign new_new_n5531__ = ~new_new_n5195__ & ~new_new_n5196__;
  assign new_new_n5532__ = ~new_new_n5530__ & ~new_new_n5531__;
  assign new_new_n5533__ = new_new_n5530__ & new_new_n5531__;
  assign new_new_n5534__ = ~new_new_n5532__ & ~new_new_n5533__;
  assign new_new_n5535__ = ~pi082 & new_new_n5534__;
  assign new_new_n5536__ = pi082 & ~new_new_n5534__;
  assign new_new_n5537__ = new_new_n5385__ & po034;
  assign new_new_n5538__ = ~pi080 & ~po034;
  assign new_new_n5539__ = ~new_new_n5537__ & ~new_new_n5538__;
  assign new_new_n5540__ = ~new_new_n5204__ & ~new_new_n5205__;
  assign new_new_n5541__ = ~new_new_n5539__ & ~new_new_n5540__;
  assign new_new_n5542__ = new_new_n5539__ & new_new_n5540__;
  assign new_new_n5543__ = ~new_new_n5541__ & ~new_new_n5542__;
  assign new_new_n5544__ = ~pi081 & ~new_new_n5543__;
  assign new_new_n5545__ = pi081 & new_new_n5543__;
  assign new_new_n5546__ = ~new_new_n5213__ & ~new_new_n5214__;
  assign new_new_n5547__ = new_new_n5383__ & po034;
  assign new_new_n5548__ = ~pi079 & ~po034;
  assign new_new_n5549__ = ~new_new_n5547__ & ~new_new_n5548__;
  assign new_new_n5550__ = new_new_n5546__ & new_new_n5549__;
  assign new_new_n5551__ = ~new_new_n5546__ & ~new_new_n5549__;
  assign new_new_n5552__ = ~new_new_n5550__ & ~new_new_n5551__;
  assign new_new_n5553__ = ~pi080 & ~new_new_n5552__;
  assign new_new_n5554__ = pi080 & new_new_n5552__;
  assign new_new_n5555__ = pi078 & ~new_new_n5381__;
  assign new_new_n5556__ = ~pi078 & new_new_n5381__;
  assign new_new_n5557__ = ~new_new_n5555__ & ~new_new_n5556__;
  assign new_new_n5558__ = po034 & new_new_n5557__;
  assign new_new_n5559__ = new_new_n5221__ & new_new_n5558__;
  assign new_new_n5560__ = ~new_new_n5221__ & ~new_new_n5558__;
  assign new_new_n5561__ = ~new_new_n5559__ & ~new_new_n5560__;
  assign new_new_n5562__ = pi079 & ~new_new_n5561__;
  assign new_new_n5563__ = ~pi079 & new_new_n5561__;
  assign new_new_n5564__ = ~new_new_n5231__ & ~new_new_n5232__;
  assign new_new_n5565__ = ~pi077 & ~po034;
  assign new_new_n5566__ = ~new_new_n5379__ & po034;
  assign new_new_n5567__ = ~new_new_n5565__ & ~new_new_n5566__;
  assign new_new_n5568__ = new_new_n5564__ & ~new_new_n5567__;
  assign new_new_n5569__ = ~new_new_n5564__ & new_new_n5567__;
  assign new_new_n5570__ = ~new_new_n5568__ & ~new_new_n5569__;
  assign new_new_n5571__ = pi078 & ~new_new_n5570__;
  assign new_new_n5572__ = ~pi078 & new_new_n5570__;
  assign new_new_n5573__ = ~new_new_n5240__ & ~new_new_n5241__;
  assign new_new_n5574__ = new_new_n5377__ & po034;
  assign new_new_n5575__ = ~pi076 & ~po034;
  assign new_new_n5576__ = ~new_new_n5574__ & ~new_new_n5575__;
  assign new_new_n5577__ = ~new_new_n5573__ & ~new_new_n5576__;
  assign new_new_n5578__ = new_new_n5573__ & new_new_n5576__;
  assign new_new_n5579__ = ~new_new_n5577__ & ~new_new_n5578__;
  assign new_new_n5580__ = ~pi077 & ~new_new_n5579__;
  assign new_new_n5581__ = pi077 & new_new_n5579__;
  assign new_new_n5582__ = ~new_new_n5249__ & ~new_new_n5250__;
  assign new_new_n5583__ = new_new_n5375__ & po034;
  assign new_new_n5584__ = ~pi075 & ~po034;
  assign new_new_n5585__ = ~new_new_n5583__ & ~new_new_n5584__;
  assign new_new_n5586__ = ~new_new_n5582__ & ~new_new_n5585__;
  assign new_new_n5587__ = new_new_n5582__ & new_new_n5585__;
  assign new_new_n5588__ = ~new_new_n5586__ & ~new_new_n5587__;
  assign new_new_n5589__ = pi076 & new_new_n5588__;
  assign new_new_n5590__ = ~pi076 & ~new_new_n5588__;
  assign new_new_n5591__ = ~new_new_n5256__ & ~new_new_n5257__;
  assign new_new_n5592__ = new_new_n5373__ & po034;
  assign new_new_n5593__ = ~pi074 & ~po034;
  assign new_new_n5594__ = ~new_new_n5592__ & ~new_new_n5593__;
  assign new_new_n5595__ = new_new_n5591__ & ~new_new_n5594__;
  assign new_new_n5596__ = ~new_new_n5591__ & new_new_n5594__;
  assign new_new_n5597__ = ~new_new_n5595__ & ~new_new_n5596__;
  assign new_new_n5598__ = pi075 & ~new_new_n5597__;
  assign new_new_n5599__ = ~pi075 & new_new_n5597__;
  assign new_new_n5600__ = pi073 & ~new_new_n5371__;
  assign new_new_n5601__ = ~pi073 & new_new_n5371__;
  assign new_new_n5602__ = ~new_new_n5600__ & ~new_new_n5601__;
  assign new_new_n5603__ = po034 & new_new_n5602__;
  assign new_new_n5604__ = ~new_new_n5264__ & ~new_new_n5603__;
  assign new_new_n5605__ = new_new_n5264__ & new_new_n5603__;
  assign new_new_n5606__ = ~new_new_n5604__ & ~new_new_n5605__;
  assign new_new_n5607__ = pi074 & ~new_new_n5606__;
  assign new_new_n5608__ = ~pi074 & new_new_n5606__;
  assign new_new_n5609__ = ~new_new_n5274__ & ~new_new_n5275__;
  assign new_new_n5610__ = ~pi072 & ~po034;
  assign new_new_n5611__ = ~new_new_n5369__ & po034;
  assign new_new_n5612__ = ~new_new_n5610__ & ~new_new_n5611__;
  assign new_new_n5613__ = new_new_n5609__ & ~new_new_n5612__;
  assign new_new_n5614__ = ~new_new_n5609__ & new_new_n5612__;
  assign new_new_n5615__ = ~new_new_n5613__ & ~new_new_n5614__;
  assign new_new_n5616__ = ~pi073 & new_new_n5615__;
  assign new_new_n5617__ = pi073 & ~new_new_n5615__;
  assign new_new_n5618__ = ~new_new_n5283__ & ~new_new_n5284__;
  assign new_new_n5619__ = new_new_n5367__ & po034;
  assign new_new_n5620__ = ~pi071 & ~po034;
  assign new_new_n5621__ = ~new_new_n5619__ & ~new_new_n5620__;
  assign new_new_n5622__ = ~new_new_n5618__ & ~new_new_n5621__;
  assign new_new_n5623__ = new_new_n5618__ & new_new_n5621__;
  assign new_new_n5624__ = ~new_new_n5622__ & ~new_new_n5623__;
  assign new_new_n5625__ = ~pi072 & ~new_new_n5624__;
  assign new_new_n5626__ = pi072 & new_new_n5624__;
  assign new_new_n5627__ = ~new_new_n5292__ & ~new_new_n5293__;
  assign new_new_n5628__ = ~pi070 & ~po034;
  assign new_new_n5629__ = ~new_new_n5365__ & po034;
  assign new_new_n5630__ = ~new_new_n5628__ & ~new_new_n5629__;
  assign new_new_n5631__ = new_new_n5627__ & ~new_new_n5630__;
  assign new_new_n5632__ = ~new_new_n5627__ & new_new_n5630__;
  assign new_new_n5633__ = ~new_new_n5631__ & ~new_new_n5632__;
  assign new_new_n5634__ = pi071 & ~new_new_n5633__;
  assign new_new_n5635__ = ~pi071 & new_new_n5633__;
  assign new_new_n5636__ = ~new_new_n5299__ & ~new_new_n5300__;
  assign new_new_n5637__ = ~new_new_n5363__ & po034;
  assign new_new_n5638__ = ~pi069 & ~po034;
  assign new_new_n5639__ = ~new_new_n5637__ & ~new_new_n5638__;
  assign new_new_n5640__ = ~new_new_n5636__ & ~new_new_n5639__;
  assign new_new_n5641__ = new_new_n5636__ & new_new_n5639__;
  assign new_new_n5642__ = ~new_new_n5640__ & ~new_new_n5641__;
  assign new_new_n5643__ = pi070 & new_new_n5642__;
  assign new_new_n5644__ = ~pi070 & ~new_new_n5642__;
  assign new_new_n5645__ = ~pi068 & ~new_new_n5361__;
  assign new_new_n5646__ = pi068 & new_new_n5361__;
  assign new_new_n5647__ = ~new_new_n5645__ & ~new_new_n5646__;
  assign new_new_n5648__ = po034 & new_new_n5647__;
  assign new_new_n5649__ = ~new_new_n5307__ & ~new_new_n5648__;
  assign new_new_n5650__ = new_new_n5307__ & new_new_n5648__;
  assign new_new_n5651__ = ~new_new_n5649__ & ~new_new_n5650__;
  assign new_new_n5652__ = pi069 & new_new_n5651__;
  assign new_new_n5653__ = ~pi069 & ~new_new_n5651__;
  assign new_new_n5654__ = ~new_new_n5315__ & ~new_new_n5316__;
  assign new_new_n5655__ = ~pi067 & ~po034;
  assign new_new_n5656__ = ~new_new_n5359__ & po034;
  assign new_new_n5657__ = ~new_new_n5655__ & ~new_new_n5656__;
  assign new_new_n5658__ = new_new_n5654__ & ~new_new_n5657__;
  assign new_new_n5659__ = ~new_new_n5654__ & new_new_n5657__;
  assign new_new_n5660__ = ~new_new_n5658__ & ~new_new_n5659__;
  assign new_new_n5661__ = pi068 & ~new_new_n5660__;
  assign new_new_n5662__ = ~pi068 & new_new_n5660__;
  assign new_new_n5663__ = ~new_new_n5330__ & ~new_new_n5331__;
  assign new_new_n5664__ = po034 & new_new_n5663__;
  assign new_new_n5665__ = new_new_n5357__ & ~new_new_n5664__;
  assign new_new_n5666__ = ~new_new_n5357__ & new_new_n5664__;
  assign new_new_n5667__ = ~new_new_n5665__ & ~new_new_n5666__;
  assign new_new_n5668__ = pi067 & ~new_new_n5667__;
  assign new_new_n5669__ = ~pi067 & new_new_n5667__;
  assign new_new_n5670__ = pi034 & po034;
  assign new_new_n5671__ = pi033 & ~pi065;
  assign new_new_n5672__ = new_new_n5670__ & ~new_new_n5671__;
  assign new_new_n5673__ = ~pi034 & ~po034;
  assign new_new_n5674__ = ~pi065 & ~new_new_n5673__;
  assign new_new_n5675__ = ~pi033 & ~new_new_n5674__;
  assign new_new_n5676__ = ~new_new_n5672__ & ~new_new_n5675__;
  assign new_new_n5677__ = pi064 & ~new_new_n5676__;
  assign new_new_n5678__ = pi064 & po034;
  assign new_new_n5679__ = new_new_n5321__ & ~new_new_n5678__;
  assign new_new_n5680__ = ~new_new_n5677__ & ~new_new_n5679__;
  assign new_new_n5681__ = pi066 & ~new_new_n5680__;
  assign new_new_n5682__ = pi065 & po034;
  assign new_new_n5683__ = ~new_new_n5326__ & ~new_new_n5682__;
  assign new_new_n5684__ = ~new_new_n5678__ & new_new_n5683__;
  assign new_new_n5685__ = new_new_n426__ & ~po035;
  assign new_new_n5686__ = new_new_n5350__ & po034;
  assign new_new_n5687__ = ~new_new_n5685__ & ~new_new_n5686__;
  assign new_new_n5688__ = ~pi034 & ~new_new_n5687__;
  assign new_new_n5689__ = po035 & ~new_new_n5682__;
  assign new_new_n5690__ = pi065 & ~new_new_n5326__;
  assign new_new_n5691__ = pi034 & ~new_new_n5690__;
  assign new_new_n5692__ = ~new_new_n5689__ & new_new_n5691__;
  assign new_new_n5693__ = ~new_new_n5684__ & ~new_new_n5688__;
  assign new_new_n5694__ = ~new_new_n5692__ & new_new_n5693__;
  assign new_new_n5695__ = ~pi035 & ~new_new_n5694__;
  assign new_new_n5696__ = pi034 & ~new_new_n5338__;
  assign new_new_n5697__ = pi064 & ~new_new_n5696__;
  assign new_new_n5698__ = ~new_new_n5683__ & ~new_new_n5697__;
  assign new_new_n5699__ = ~pi065 & po034;
  assign new_new_n5700__ = ~po035 & ~new_new_n5699__;
  assign new_new_n5701__ = pi064 & ~new_new_n5670__;
  assign new_new_n5702__ = ~new_new_n5686__ & new_new_n5701__;
  assign new_new_n5703__ = ~new_new_n5700__ & new_new_n5702__;
  assign new_new_n5704__ = ~new_new_n5698__ & ~new_new_n5703__;
  assign new_new_n5705__ = pi035 & ~new_new_n5704__;
  assign new_new_n5706__ = ~new_new_n5695__ & ~new_new_n5705__;
  assign new_new_n5707__ = ~pi066 & new_new_n5680__;
  assign new_new_n5708__ = ~new_new_n5706__ & ~new_new_n5707__;
  assign new_new_n5709__ = ~new_new_n5681__ & ~new_new_n5708__;
  assign new_new_n5710__ = ~new_new_n5669__ & ~new_new_n5709__;
  assign new_new_n5711__ = ~new_new_n5668__ & ~new_new_n5710__;
  assign new_new_n5712__ = ~new_new_n5662__ & ~new_new_n5711__;
  assign new_new_n5713__ = ~new_new_n5661__ & ~new_new_n5712__;
  assign new_new_n5714__ = ~new_new_n5653__ & ~new_new_n5713__;
  assign new_new_n5715__ = ~new_new_n5652__ & ~new_new_n5714__;
  assign new_new_n5716__ = ~new_new_n5644__ & ~new_new_n5715__;
  assign new_new_n5717__ = ~new_new_n5643__ & ~new_new_n5716__;
  assign new_new_n5718__ = ~new_new_n5635__ & ~new_new_n5717__;
  assign new_new_n5719__ = ~new_new_n5634__ & ~new_new_n5718__;
  assign new_new_n5720__ = ~new_new_n5626__ & new_new_n5719__;
  assign new_new_n5721__ = ~new_new_n5625__ & ~new_new_n5720__;
  assign new_new_n5722__ = ~new_new_n5617__ & ~new_new_n5721__;
  assign new_new_n5723__ = ~new_new_n5616__ & ~new_new_n5722__;
  assign new_new_n5724__ = ~new_new_n5608__ & new_new_n5723__;
  assign new_new_n5725__ = ~new_new_n5607__ & ~new_new_n5724__;
  assign new_new_n5726__ = ~new_new_n5599__ & ~new_new_n5725__;
  assign new_new_n5727__ = ~new_new_n5598__ & ~new_new_n5726__;
  assign new_new_n5728__ = ~new_new_n5590__ & ~new_new_n5727__;
  assign new_new_n5729__ = ~new_new_n5589__ & ~new_new_n5728__;
  assign new_new_n5730__ = ~new_new_n5581__ & new_new_n5729__;
  assign new_new_n5731__ = ~new_new_n5580__ & ~new_new_n5730__;
  assign new_new_n5732__ = ~new_new_n5572__ & new_new_n5731__;
  assign new_new_n5733__ = ~new_new_n5571__ & ~new_new_n5732__;
  assign new_new_n5734__ = ~new_new_n5563__ & ~new_new_n5733__;
  assign new_new_n5735__ = ~new_new_n5562__ & ~new_new_n5734__;
  assign new_new_n5736__ = ~new_new_n5554__ & new_new_n5735__;
  assign new_new_n5737__ = ~new_new_n5553__ & ~new_new_n5736__;
  assign new_new_n5738__ = ~new_new_n5545__ & ~new_new_n5737__;
  assign new_new_n5739__ = ~new_new_n5544__ & ~new_new_n5738__;
  assign new_new_n5740__ = ~new_new_n5536__ & ~new_new_n5739__;
  assign new_new_n5741__ = ~new_new_n5535__ & ~new_new_n5740__;
  assign new_new_n5742__ = ~new_new_n5527__ & ~new_new_n5741__;
  assign new_new_n5743__ = ~new_new_n5526__ & ~new_new_n5742__;
  assign new_new_n5744__ = ~new_new_n5518__ & ~new_new_n5743__;
  assign new_new_n5745__ = ~new_new_n5517__ & ~new_new_n5744__;
  assign new_new_n5746__ = ~new_new_n5509__ & new_new_n5745__;
  assign new_new_n5747__ = ~new_new_n5508__ & ~new_new_n5746__;
  assign new_new_n5748__ = ~new_new_n5500__ & ~new_new_n5747__;
  assign new_new_n5749__ = ~new_new_n5499__ & ~new_new_n5748__;
  assign new_new_n5750__ = ~new_new_n5491__ & ~new_new_n5749__;
  assign new_new_n5751__ = ~new_new_n5490__ & ~new_new_n5750__;
  assign new_new_n5752__ = ~new_new_n5482__ & ~new_new_n5751__;
  assign new_new_n5753__ = ~new_new_n5481__ & ~new_new_n5752__;
  assign new_new_n5754__ = ~new_new_n5473__ & ~new_new_n5753__;
  assign new_new_n5755__ = ~new_new_n5472__ & ~new_new_n5754__;
  assign new_new_n5756__ = ~new_new_n5464__ & ~new_new_n5755__;
  assign new_new_n5757__ = ~new_new_n5463__ & ~new_new_n5756__;
  assign new_new_n5758__ = ~pi091 & new_new_n5454__;
  assign new_new_n5759__ = ~new_new_n5757__ & ~new_new_n5758__;
  assign new_new_n5760__ = ~new_new_n5455__ & ~new_new_n5759__;
  assign new_new_n5761__ = ~new_new_n5447__ & ~new_new_n5760__;
  assign new_new_n5762__ = ~new_new_n5446__ & ~new_new_n5761__;
  assign new_new_n5763__ = new_new_n5414__ & ~po034;
  assign new_new_n5764__ = ~pi094 & new_new_n5763__;
  assign new_new_n5765__ = ~new_new_n5431__ & ~new_new_n5762__;
  assign new_new_n5766__ = pi094 & ~new_new_n5763__;
  assign new_new_n5767__ = ~new_new_n5432__ & ~new_new_n5766__;
  assign new_new_n5768__ = ~new_new_n5765__ & new_new_n5767__;
  assign new_new_n5769__ = ~new_new_n5764__ & ~new_new_n5768__;
  assign po033 = new_new_n3332__ & ~new_new_n5769__;
  assign new_new_n5771__ = new_new_n5762__ & po033;
  assign new_new_n5772__ = ~pi093 & ~po033;
  assign new_new_n5773__ = ~new_new_n5771__ & ~new_new_n5772__;
  assign new_new_n5774__ = ~new_new_n5433__ & ~new_new_n5773__;
  assign new_new_n5775__ = new_new_n5433__ & new_new_n5773__;
  assign new_new_n5776__ = ~new_new_n5774__ & ~new_new_n5775__;
  assign new_new_n5777__ = new_new_n5763__ & ~po033;
  assign new_new_n5778__ = ~new_new_n376__ & ~new_new_n5777__;
  assign new_new_n5779__ = pi095 & new_new_n5778__;
  assign new_new_n5780__ = new_new_n5760__ & po033;
  assign new_new_n5781__ = ~pi092 & ~po033;
  assign new_new_n5782__ = ~new_new_n5780__ & ~new_new_n5781__;
  assign new_new_n5783__ = ~new_new_n5446__ & ~new_new_n5447__;
  assign new_new_n5784__ = ~new_new_n5782__ & ~new_new_n5783__;
  assign new_new_n5785__ = new_new_n5782__ & new_new_n5783__;
  assign new_new_n5786__ = ~new_new_n5784__ & ~new_new_n5785__;
  assign new_new_n5787__ = ~pi093 & ~new_new_n5786__;
  assign new_new_n5788__ = pi093 & new_new_n5786__;
  assign new_new_n5789__ = ~new_new_n5455__ & ~new_new_n5758__;
  assign new_new_n5790__ = pi091 & ~po033;
  assign new_new_n5791__ = ~new_new_n5757__ & po033;
  assign new_new_n5792__ = ~new_new_n5790__ & ~new_new_n5791__;
  assign new_new_n5793__ = new_new_n5789__ & new_new_n5792__;
  assign new_new_n5794__ = ~new_new_n5789__ & ~new_new_n5792__;
  assign new_new_n5795__ = ~new_new_n5793__ & ~new_new_n5794__;
  assign new_new_n5796__ = ~pi092 & new_new_n5795__;
  assign new_new_n5797__ = pi092 & ~new_new_n5795__;
  assign new_new_n5798__ = ~new_new_n5755__ & po033;
  assign new_new_n5799__ = pi090 & ~po033;
  assign new_new_n5800__ = ~new_new_n5798__ & ~new_new_n5799__;
  assign new_new_n5801__ = ~new_new_n5463__ & ~new_new_n5464__;
  assign new_new_n5802__ = ~new_new_n5800__ & new_new_n5801__;
  assign new_new_n5803__ = new_new_n5800__ & ~new_new_n5801__;
  assign new_new_n5804__ = ~new_new_n5802__ & ~new_new_n5803__;
  assign new_new_n5805__ = ~pi091 & ~new_new_n5804__;
  assign new_new_n5806__ = pi091 & new_new_n5804__;
  assign new_new_n5807__ = pi089 & ~new_new_n5753__;
  assign new_new_n5808__ = ~pi089 & new_new_n5753__;
  assign new_new_n5809__ = ~new_new_n5807__ & ~new_new_n5808__;
  assign new_new_n5810__ = po033 & new_new_n5809__;
  assign new_new_n5811__ = new_new_n5471__ & new_new_n5810__;
  assign new_new_n5812__ = ~new_new_n5471__ & ~new_new_n5810__;
  assign new_new_n5813__ = ~new_new_n5811__ & ~new_new_n5812__;
  assign new_new_n5814__ = pi090 & ~new_new_n5813__;
  assign new_new_n5815__ = ~pi090 & new_new_n5813__;
  assign new_new_n5816__ = ~new_new_n5481__ & ~new_new_n5482__;
  assign new_new_n5817__ = ~new_new_n5751__ & po033;
  assign new_new_n5818__ = pi088 & ~po033;
  assign new_new_n5819__ = ~new_new_n5817__ & ~new_new_n5818__;
  assign new_new_n5820__ = new_new_n5816__ & ~new_new_n5819__;
  assign new_new_n5821__ = ~new_new_n5816__ & new_new_n5819__;
  assign new_new_n5822__ = ~new_new_n5820__ & ~new_new_n5821__;
  assign new_new_n5823__ = ~pi089 & ~new_new_n5822__;
  assign new_new_n5824__ = pi089 & new_new_n5822__;
  assign new_new_n5825__ = ~new_new_n5749__ & po033;
  assign new_new_n5826__ = pi087 & ~po033;
  assign new_new_n5827__ = ~new_new_n5825__ & ~new_new_n5826__;
  assign new_new_n5828__ = ~new_new_n5490__ & ~new_new_n5491__;
  assign new_new_n5829__ = ~new_new_n5827__ & new_new_n5828__;
  assign new_new_n5830__ = new_new_n5827__ & ~new_new_n5828__;
  assign new_new_n5831__ = ~new_new_n5829__ & ~new_new_n5830__;
  assign new_new_n5832__ = ~pi088 & ~new_new_n5831__;
  assign new_new_n5833__ = pi088 & new_new_n5831__;
  assign new_new_n5834__ = ~new_new_n5499__ & ~new_new_n5500__;
  assign new_new_n5835__ = ~new_new_n5747__ & po033;
  assign new_new_n5836__ = pi086 & ~po033;
  assign new_new_n5837__ = ~new_new_n5835__ & ~new_new_n5836__;
  assign new_new_n5838__ = new_new_n5834__ & ~new_new_n5837__;
  assign new_new_n5839__ = ~new_new_n5834__ & new_new_n5837__;
  assign new_new_n5840__ = ~new_new_n5838__ & ~new_new_n5839__;
  assign new_new_n5841__ = ~pi087 & ~new_new_n5840__;
  assign new_new_n5842__ = pi087 & new_new_n5840__;
  assign new_new_n5843__ = ~new_new_n5508__ & ~new_new_n5509__;
  assign new_new_n5844__ = ~new_new_n5745__ & po033;
  assign new_new_n5845__ = ~pi085 & ~po033;
  assign new_new_n5846__ = ~new_new_n5844__ & ~new_new_n5845__;
  assign new_new_n5847__ = new_new_n5843__ & ~new_new_n5846__;
  assign new_new_n5848__ = ~new_new_n5843__ & new_new_n5846__;
  assign new_new_n5849__ = ~new_new_n5847__ & ~new_new_n5848__;
  assign new_new_n5850__ = pi086 & ~new_new_n5849__;
  assign new_new_n5851__ = ~pi086 & new_new_n5849__;
  assign new_new_n5852__ = ~new_new_n5517__ & ~new_new_n5518__;
  assign new_new_n5853__ = ~new_new_n5743__ & po033;
  assign new_new_n5854__ = ~pi084 & ~po033;
  assign new_new_n5855__ = ~new_new_n5853__ & ~new_new_n5854__;
  assign new_new_n5856__ = new_new_n5852__ & ~new_new_n5855__;
  assign new_new_n5857__ = ~new_new_n5852__ & new_new_n5855__;
  assign new_new_n5858__ = ~new_new_n5856__ & ~new_new_n5857__;
  assign new_new_n5859__ = pi085 & ~new_new_n5858__;
  assign new_new_n5860__ = ~pi085 & new_new_n5858__;
  assign new_new_n5861__ = ~pi083 & ~new_new_n5741__;
  assign new_new_n5862__ = pi083 & new_new_n5741__;
  assign new_new_n5863__ = ~new_new_n5861__ & ~new_new_n5862__;
  assign new_new_n5864__ = po033 & new_new_n5863__;
  assign new_new_n5865__ = ~new_new_n5525__ & new_new_n5864__;
  assign new_new_n5866__ = new_new_n5525__ & ~new_new_n5864__;
  assign new_new_n5867__ = ~new_new_n5865__ & ~new_new_n5866__;
  assign new_new_n5868__ = pi084 & ~new_new_n5867__;
  assign new_new_n5869__ = ~pi084 & new_new_n5867__;
  assign new_new_n5870__ = ~new_new_n5535__ & ~new_new_n5536__;
  assign new_new_n5871__ = ~new_new_n5739__ & po033;
  assign new_new_n5872__ = ~pi082 & ~po033;
  assign new_new_n5873__ = ~new_new_n5871__ & ~new_new_n5872__;
  assign new_new_n5874__ = new_new_n5870__ & ~new_new_n5873__;
  assign new_new_n5875__ = ~new_new_n5870__ & new_new_n5873__;
  assign new_new_n5876__ = ~new_new_n5874__ & ~new_new_n5875__;
  assign new_new_n5877__ = pi083 & ~new_new_n5876__;
  assign new_new_n5878__ = ~pi083 & new_new_n5876__;
  assign new_new_n5879__ = ~pi081 & ~new_new_n5737__;
  assign new_new_n5880__ = pi081 & new_new_n5737__;
  assign new_new_n5881__ = ~new_new_n5879__ & ~new_new_n5880__;
  assign new_new_n5882__ = po033 & new_new_n5881__;
  assign new_new_n5883__ = new_new_n5543__ & ~new_new_n5882__;
  assign new_new_n5884__ = ~new_new_n5543__ & new_new_n5882__;
  assign new_new_n5885__ = ~new_new_n5883__ & ~new_new_n5884__;
  assign new_new_n5886__ = pi082 & ~new_new_n5885__;
  assign new_new_n5887__ = ~pi082 & new_new_n5885__;
  assign new_new_n5888__ = ~new_new_n5553__ & ~new_new_n5554__;
  assign new_new_n5889__ = ~new_new_n5735__ & po033;
  assign new_new_n5890__ = pi080 & ~po033;
  assign new_new_n5891__ = ~new_new_n5889__ & ~new_new_n5890__;
  assign new_new_n5892__ = new_new_n5888__ & ~new_new_n5891__;
  assign new_new_n5893__ = ~new_new_n5888__ & new_new_n5891__;
  assign new_new_n5894__ = ~new_new_n5892__ & ~new_new_n5893__;
  assign new_new_n5895__ = ~pi081 & ~new_new_n5894__;
  assign new_new_n5896__ = pi081 & new_new_n5894__;
  assign new_new_n5897__ = pi079 & ~new_new_n5733__;
  assign new_new_n5898__ = ~pi079 & new_new_n5733__;
  assign new_new_n5899__ = ~new_new_n5897__ & ~new_new_n5898__;
  assign new_new_n5900__ = po033 & new_new_n5899__;
  assign new_new_n5901__ = ~new_new_n5561__ & ~new_new_n5900__;
  assign new_new_n5902__ = new_new_n5561__ & new_new_n5900__;
  assign new_new_n5903__ = ~new_new_n5901__ & ~new_new_n5902__;
  assign new_new_n5904__ = pi080 & ~new_new_n5903__;
  assign new_new_n5905__ = ~pi080 & new_new_n5903__;
  assign new_new_n5906__ = ~new_new_n5571__ & ~new_new_n5572__;
  assign new_new_n5907__ = ~new_new_n5731__ & po033;
  assign new_new_n5908__ = ~pi078 & ~po033;
  assign new_new_n5909__ = ~new_new_n5907__ & ~new_new_n5908__;
  assign new_new_n5910__ = new_new_n5906__ & ~new_new_n5909__;
  assign new_new_n5911__ = ~new_new_n5906__ & new_new_n5909__;
  assign new_new_n5912__ = ~new_new_n5910__ & ~new_new_n5911__;
  assign new_new_n5913__ = pi079 & ~new_new_n5912__;
  assign new_new_n5914__ = ~pi079 & new_new_n5912__;
  assign new_new_n5915__ = ~new_new_n5729__ & po033;
  assign new_new_n5916__ = pi077 & ~po033;
  assign new_new_n5917__ = ~new_new_n5915__ & ~new_new_n5916__;
  assign new_new_n5918__ = ~new_new_n5580__ & ~new_new_n5581__;
  assign new_new_n5919__ = ~new_new_n5917__ & new_new_n5918__;
  assign new_new_n5920__ = new_new_n5917__ & ~new_new_n5918__;
  assign new_new_n5921__ = ~new_new_n5919__ & ~new_new_n5920__;
  assign new_new_n5922__ = pi078 & new_new_n5921__;
  assign new_new_n5923__ = ~pi078 & ~new_new_n5921__;
  assign new_new_n5924__ = ~new_new_n5727__ & po033;
  assign new_new_n5925__ = pi076 & ~po033;
  assign new_new_n5926__ = ~new_new_n5924__ & ~new_new_n5925__;
  assign new_new_n5927__ = ~new_new_n5589__ & ~new_new_n5590__;
  assign new_new_n5928__ = ~new_new_n5926__ & new_new_n5927__;
  assign new_new_n5929__ = new_new_n5926__ & ~new_new_n5927__;
  assign new_new_n5930__ = ~new_new_n5928__ & ~new_new_n5929__;
  assign new_new_n5931__ = pi077 & new_new_n5930__;
  assign new_new_n5932__ = ~pi077 & ~new_new_n5930__;
  assign new_new_n5933__ = ~new_new_n5598__ & ~new_new_n5599__;
  assign new_new_n5934__ = ~new_new_n5725__ & po033;
  assign new_new_n5935__ = pi075 & ~po033;
  assign new_new_n5936__ = ~new_new_n5934__ & ~new_new_n5935__;
  assign new_new_n5937__ = new_new_n5933__ & new_new_n5936__;
  assign new_new_n5938__ = ~new_new_n5933__ & ~new_new_n5936__;
  assign new_new_n5939__ = ~new_new_n5937__ & ~new_new_n5938__;
  assign new_new_n5940__ = pi076 & ~new_new_n5939__;
  assign new_new_n5941__ = ~pi076 & new_new_n5939__;
  assign new_new_n5942__ = new_new_n5723__ & po033;
  assign new_new_n5943__ = pi074 & ~po033;
  assign new_new_n5944__ = ~new_new_n5942__ & ~new_new_n5943__;
  assign new_new_n5945__ = ~new_new_n5607__ & ~new_new_n5608__;
  assign new_new_n5946__ = ~new_new_n5944__ & ~new_new_n5945__;
  assign new_new_n5947__ = new_new_n5944__ & new_new_n5945__;
  assign new_new_n5948__ = ~new_new_n5946__ & ~new_new_n5947__;
  assign new_new_n5949__ = pi075 & ~new_new_n5948__;
  assign new_new_n5950__ = ~pi075 & new_new_n5948__;
  assign new_new_n5951__ = ~new_new_n5616__ & ~new_new_n5617__;
  assign new_new_n5952__ = ~new_new_n5721__ & po033;
  assign new_new_n5953__ = ~pi073 & ~po033;
  assign new_new_n5954__ = ~new_new_n5952__ & ~new_new_n5953__;
  assign new_new_n5955__ = new_new_n5951__ & ~new_new_n5954__;
  assign new_new_n5956__ = ~new_new_n5951__ & new_new_n5954__;
  assign new_new_n5957__ = ~new_new_n5955__ & ~new_new_n5956__;
  assign new_new_n5958__ = ~pi074 & new_new_n5957__;
  assign new_new_n5959__ = pi074 & ~new_new_n5957__;
  assign new_new_n5960__ = ~new_new_n5719__ & po033;
  assign new_new_n5961__ = pi072 & ~po033;
  assign new_new_n5962__ = ~new_new_n5960__ & ~new_new_n5961__;
  assign new_new_n5963__ = ~new_new_n5625__ & ~new_new_n5626__;
  assign new_new_n5964__ = ~new_new_n5962__ & new_new_n5963__;
  assign new_new_n5965__ = new_new_n5962__ & ~new_new_n5963__;
  assign new_new_n5966__ = ~new_new_n5964__ & ~new_new_n5965__;
  assign new_new_n5967__ = ~pi073 & ~new_new_n5966__;
  assign new_new_n5968__ = pi073 & new_new_n5966__;
  assign new_new_n5969__ = pi071 & ~new_new_n5717__;
  assign new_new_n5970__ = ~pi071 & new_new_n5717__;
  assign new_new_n5971__ = ~new_new_n5969__ & ~new_new_n5970__;
  assign new_new_n5972__ = po033 & new_new_n5971__;
  assign new_new_n5973__ = new_new_n5633__ & new_new_n5972__;
  assign new_new_n5974__ = ~new_new_n5633__ & ~new_new_n5972__;
  assign new_new_n5975__ = ~new_new_n5973__ & ~new_new_n5974__;
  assign new_new_n5976__ = ~pi072 & new_new_n5975__;
  assign new_new_n5977__ = pi072 & ~new_new_n5975__;
  assign new_new_n5978__ = ~new_new_n5715__ & po033;
  assign new_new_n5979__ = pi070 & ~po033;
  assign new_new_n5980__ = ~new_new_n5978__ & ~new_new_n5979__;
  assign new_new_n5981__ = ~new_new_n5643__ & ~new_new_n5644__;
  assign new_new_n5982__ = ~new_new_n5980__ & new_new_n5981__;
  assign new_new_n5983__ = new_new_n5980__ & ~new_new_n5981__;
  assign new_new_n5984__ = ~new_new_n5982__ & ~new_new_n5983__;
  assign new_new_n5985__ = ~pi071 & ~new_new_n5984__;
  assign new_new_n5986__ = pi071 & new_new_n5984__;
  assign new_new_n5987__ = ~new_new_n5652__ & ~new_new_n5653__;
  assign new_new_n5988__ = new_new_n5713__ & po033;
  assign new_new_n5989__ = ~pi069 & ~po033;
  assign new_new_n5990__ = ~new_new_n5988__ & ~new_new_n5989__;
  assign new_new_n5991__ = ~new_new_n5987__ & ~new_new_n5990__;
  assign new_new_n5992__ = new_new_n5987__ & new_new_n5990__;
  assign new_new_n5993__ = ~new_new_n5991__ & ~new_new_n5992__;
  assign new_new_n5994__ = ~pi070 & ~new_new_n5993__;
  assign new_new_n5995__ = pi070 & new_new_n5993__;
  assign new_new_n5996__ = ~new_new_n5661__ & ~new_new_n5662__;
  assign new_new_n5997__ = ~new_new_n5711__ & po033;
  assign new_new_n5998__ = pi068 & ~po033;
  assign new_new_n5999__ = ~new_new_n5997__ & ~new_new_n5998__;
  assign new_new_n6000__ = new_new_n5996__ & new_new_n5999__;
  assign new_new_n6001__ = ~new_new_n5996__ & ~new_new_n5999__;
  assign new_new_n6002__ = ~new_new_n6000__ & ~new_new_n6001__;
  assign new_new_n6003__ = pi069 & ~new_new_n6002__;
  assign new_new_n6004__ = ~pi069 & new_new_n6002__;
  assign new_new_n6005__ = pi067 & ~new_new_n5709__;
  assign new_new_n6006__ = ~pi067 & new_new_n5709__;
  assign new_new_n6007__ = ~new_new_n6005__ & ~new_new_n6006__;
  assign new_new_n6008__ = po033 & new_new_n6007__;
  assign new_new_n6009__ = new_new_n5667__ & new_new_n6008__;
  assign new_new_n6010__ = ~new_new_n5667__ & ~new_new_n6008__;
  assign new_new_n6011__ = ~new_new_n6009__ & ~new_new_n6010__;
  assign new_new_n6012__ = pi068 & ~new_new_n6011__;
  assign new_new_n6013__ = ~pi068 & new_new_n6011__;
  assign new_new_n6014__ = ~new_new_n5681__ & ~new_new_n5707__;
  assign new_new_n6015__ = po033 & new_new_n6014__;
  assign new_new_n6016__ = new_new_n5706__ & ~new_new_n6015__;
  assign new_new_n6017__ = ~new_new_n5706__ & new_new_n6015__;
  assign new_new_n6018__ = ~new_new_n6016__ & ~new_new_n6017__;
  assign new_new_n6019__ = ~pi067 & ~new_new_n6018__;
  assign new_new_n6020__ = pi067 & new_new_n6018__;
  assign new_new_n6021__ = pi033 & po033;
  assign new_new_n6022__ = ~pi033 & ~po033;
  assign new_new_n6023__ = ~pi065 & ~new_new_n6021__;
  assign new_new_n6024__ = ~new_new_n6022__ & new_new_n6023__;
  assign new_new_n6025__ = ~pi032 & ~new_new_n6024__;
  assign new_new_n6026__ = pi065 & new_new_n6021__;
  assign new_new_n6027__ = ~new_new_n6025__ & ~new_new_n6026__;
  assign new_new_n6028__ = pi064 & ~new_new_n6027__;
  assign new_new_n6029__ = pi064 & po033;
  assign new_new_n6030__ = ~pi033 & pi065;
  assign new_new_n6031__ = ~new_new_n6029__ & new_new_n6030__;
  assign new_new_n6032__ = ~new_new_n6028__ & ~new_new_n6031__;
  assign new_new_n6033__ = pi066 & ~new_new_n6032__;
  assign new_new_n6034__ = ~pi066 & new_new_n6032__;
  assign new_new_n6035__ = pi065 & po033;
  assign new_new_n6036__ = ~pi064 & ~new_new_n6035__;
  assign new_new_n6037__ = ~pi065 & po033;
  assign new_new_n6038__ = ~po034 & ~new_new_n6037__;
  assign new_new_n6039__ = new_new_n5699__ & po033;
  assign new_new_n6040__ = ~new_new_n6021__ & ~new_new_n6039__;
  assign new_new_n6041__ = ~new_new_n6038__ & new_new_n6040__;
  assign new_new_n6042__ = pi064 & ~new_new_n6041__;
  assign new_new_n6043__ = ~new_new_n6036__ & ~new_new_n6042__;
  assign new_new_n6044__ = ~new_new_n5678__ & ~new_new_n6035__;
  assign new_new_n6045__ = pi033 & ~new_new_n5682__;
  assign new_new_n6046__ = ~new_new_n6044__ & new_new_n6045__;
  assign new_new_n6047__ = ~new_new_n6043__ & ~new_new_n6046__;
  assign new_new_n6048__ = pi034 & ~new_new_n6047__;
  assign new_new_n6049__ = pi065 & ~new_new_n5678__;
  assign new_new_n6050__ = po034 & ~new_new_n6035__;
  assign new_new_n6051__ = pi033 & ~new_new_n6049__;
  assign new_new_n6052__ = ~new_new_n6050__ & new_new_n6051__;
  assign new_new_n6053__ = new_new_n426__ & ~po034;
  assign new_new_n6054__ = ~new_new_n6039__ & ~new_new_n6053__;
  assign new_new_n6055__ = ~pi033 & ~new_new_n6054__;
  assign new_new_n6056__ = ~po034 & ~po033;
  assign new_new_n6057__ = ~new_new_n6036__ & ~new_new_n6056__;
  assign new_new_n6058__ = ~new_new_n6052__ & new_new_n6057__;
  assign new_new_n6059__ = ~new_new_n6055__ & new_new_n6058__;
  assign new_new_n6060__ = ~pi034 & ~new_new_n6059__;
  assign new_new_n6061__ = ~new_new_n6048__ & ~new_new_n6060__;
  assign new_new_n6062__ = ~new_new_n6034__ & ~new_new_n6061__;
  assign new_new_n6063__ = ~new_new_n6033__ & ~new_new_n6062__;
  assign new_new_n6064__ = ~new_new_n6020__ & new_new_n6063__;
  assign new_new_n6065__ = ~new_new_n6019__ & ~new_new_n6064__;
  assign new_new_n6066__ = ~new_new_n6013__ & new_new_n6065__;
  assign new_new_n6067__ = ~new_new_n6012__ & ~new_new_n6066__;
  assign new_new_n6068__ = ~new_new_n6004__ & ~new_new_n6067__;
  assign new_new_n6069__ = ~new_new_n6003__ & ~new_new_n6068__;
  assign new_new_n6070__ = ~new_new_n5995__ & new_new_n6069__;
  assign new_new_n6071__ = ~new_new_n5994__ & ~new_new_n6070__;
  assign new_new_n6072__ = ~new_new_n5986__ & ~new_new_n6071__;
  assign new_new_n6073__ = ~new_new_n5985__ & ~new_new_n6072__;
  assign new_new_n6074__ = ~new_new_n5977__ & ~new_new_n6073__;
  assign new_new_n6075__ = ~new_new_n5976__ & ~new_new_n6074__;
  assign new_new_n6076__ = ~new_new_n5968__ & ~new_new_n6075__;
  assign new_new_n6077__ = ~new_new_n5967__ & ~new_new_n6076__;
  assign new_new_n6078__ = ~new_new_n5959__ & ~new_new_n6077__;
  assign new_new_n6079__ = ~new_new_n5958__ & ~new_new_n6078__;
  assign new_new_n6080__ = ~new_new_n5950__ & new_new_n6079__;
  assign new_new_n6081__ = ~new_new_n5949__ & ~new_new_n6080__;
  assign new_new_n6082__ = ~new_new_n5941__ & ~new_new_n6081__;
  assign new_new_n6083__ = ~new_new_n5940__ & ~new_new_n6082__;
  assign new_new_n6084__ = ~new_new_n5932__ & ~new_new_n6083__;
  assign new_new_n6085__ = ~new_new_n5931__ & ~new_new_n6084__;
  assign new_new_n6086__ = ~new_new_n5923__ & ~new_new_n6085__;
  assign new_new_n6087__ = ~new_new_n5922__ & ~new_new_n6086__;
  assign new_new_n6088__ = ~new_new_n5914__ & ~new_new_n6087__;
  assign new_new_n6089__ = ~new_new_n5913__ & ~new_new_n6088__;
  assign new_new_n6090__ = ~new_new_n5905__ & ~new_new_n6089__;
  assign new_new_n6091__ = ~new_new_n5904__ & ~new_new_n6090__;
  assign new_new_n6092__ = ~new_new_n5896__ & new_new_n6091__;
  assign new_new_n6093__ = ~new_new_n5895__ & ~new_new_n6092__;
  assign new_new_n6094__ = ~new_new_n5887__ & new_new_n6093__;
  assign new_new_n6095__ = ~new_new_n5886__ & ~new_new_n6094__;
  assign new_new_n6096__ = ~new_new_n5878__ & ~new_new_n6095__;
  assign new_new_n6097__ = ~new_new_n5877__ & ~new_new_n6096__;
  assign new_new_n6098__ = ~new_new_n5869__ & ~new_new_n6097__;
  assign new_new_n6099__ = ~new_new_n5868__ & ~new_new_n6098__;
  assign new_new_n6100__ = ~new_new_n5860__ & ~new_new_n6099__;
  assign new_new_n6101__ = ~new_new_n5859__ & ~new_new_n6100__;
  assign new_new_n6102__ = ~new_new_n5851__ & ~new_new_n6101__;
  assign new_new_n6103__ = ~new_new_n5850__ & ~new_new_n6102__;
  assign new_new_n6104__ = ~new_new_n5842__ & new_new_n6103__;
  assign new_new_n6105__ = ~new_new_n5841__ & ~new_new_n6104__;
  assign new_new_n6106__ = ~new_new_n5833__ & ~new_new_n6105__;
  assign new_new_n6107__ = ~new_new_n5832__ & ~new_new_n6106__;
  assign new_new_n6108__ = ~new_new_n5824__ & ~new_new_n6107__;
  assign new_new_n6109__ = ~new_new_n5823__ & ~new_new_n6108__;
  assign new_new_n6110__ = ~new_new_n5815__ & new_new_n6109__;
  assign new_new_n6111__ = ~new_new_n5814__ & ~new_new_n6110__;
  assign new_new_n6112__ = ~new_new_n5806__ & new_new_n6111__;
  assign new_new_n6113__ = ~new_new_n5805__ & ~new_new_n6112__;
  assign new_new_n6114__ = ~new_new_n5797__ & ~new_new_n6113__;
  assign new_new_n6115__ = ~new_new_n5796__ & ~new_new_n6114__;
  assign new_new_n6116__ = ~new_new_n5788__ & ~new_new_n6115__;
  assign new_new_n6117__ = ~new_new_n5787__ & ~new_new_n6116__;
  assign new_new_n6118__ = pi094 & new_new_n6117__;
  assign new_new_n6119__ = ~new_new_n5779__ & ~new_new_n6118__;
  assign new_new_n6120__ = ~pi094 & ~new_new_n6117__;
  assign new_new_n6121__ = new_new_n289__ & ~new_new_n6120__;
  assign new_new_n6122__ = new_new_n6119__ & new_new_n6121__;
  assign new_new_n6123__ = ~new_new_n5776__ & ~new_new_n6122__;
  assign new_new_n6124__ = new_new_n5776__ & ~new_new_n6120__;
  assign new_new_n6125__ = ~pi095 & ~new_new_n5778__;
  assign new_new_n6126__ = new_new_n289__ & new_new_n6125__;
  assign new_new_n6127__ = ~new_new_n6118__ & new_new_n6126__;
  assign new_new_n6128__ = new_new_n6124__ & new_new_n6127__;
  assign new_new_n6129__ = ~new_new_n6123__ & ~new_new_n6128__;
  assign new_new_n6130__ = ~pi095 & ~new_new_n6129__;
  assign new_new_n6131__ = pi095 & new_new_n6129__;
  assign new_new_n6132__ = ~new_new_n6130__ & ~new_new_n6131__;
  assign new_new_n6133__ = ~new_new_n5787__ & ~new_new_n5788__;
  assign new_new_n6134__ = new_new_n6119__ & ~new_new_n6124__;
  assign new_new_n6135__ = ~new_new_n6125__ & ~new_new_n6134__;
  assign po032 = new_new_n289__ & ~new_new_n6135__;
  assign new_new_n6137__ = ~new_new_n6115__ & po032;
  assign new_new_n6138__ = ~pi093 & ~po032;
  assign new_new_n6139__ = ~new_new_n6137__ & ~new_new_n6138__;
  assign new_new_n6140__ = new_new_n6133__ & ~new_new_n6139__;
  assign new_new_n6141__ = ~new_new_n6133__ & new_new_n6139__;
  assign new_new_n6142__ = ~new_new_n6140__ & ~new_new_n6141__;
  assign new_new_n6143__ = pi094 & ~new_new_n6142__;
  assign new_new_n6144__ = ~pi094 & new_new_n6142__;
  assign new_new_n6145__ = ~new_new_n5796__ & ~new_new_n5797__;
  assign new_new_n6146__ = ~new_new_n6113__ & po032;
  assign new_new_n6147__ = ~pi092 & ~po032;
  assign new_new_n6148__ = ~new_new_n6146__ & ~new_new_n6147__;
  assign new_new_n6149__ = new_new_n6145__ & ~new_new_n6148__;
  assign new_new_n6150__ = ~new_new_n6145__ & new_new_n6148__;
  assign new_new_n6151__ = ~new_new_n6149__ & ~new_new_n6150__;
  assign new_new_n6152__ = pi093 & ~new_new_n6151__;
  assign new_new_n6153__ = ~pi093 & new_new_n6151__;
  assign new_new_n6154__ = ~new_new_n5805__ & ~new_new_n5806__;
  assign new_new_n6155__ = ~new_new_n6111__ & po032;
  assign new_new_n6156__ = pi091 & ~po032;
  assign new_new_n6157__ = ~new_new_n6155__ & ~new_new_n6156__;
  assign new_new_n6158__ = new_new_n6154__ & ~new_new_n6157__;
  assign new_new_n6159__ = ~new_new_n6154__ & new_new_n6157__;
  assign new_new_n6160__ = ~new_new_n6158__ & ~new_new_n6159__;
  assign new_new_n6161__ = pi092 & new_new_n6160__;
  assign new_new_n6162__ = ~pi092 & ~new_new_n6160__;
  assign new_new_n6163__ = ~new_new_n5814__ & ~new_new_n5815__;
  assign new_new_n6164__ = ~new_new_n6109__ & po032;
  assign new_new_n6165__ = ~pi090 & ~po032;
  assign new_new_n6166__ = ~new_new_n6164__ & ~new_new_n6165__;
  assign new_new_n6167__ = new_new_n6163__ & ~new_new_n6166__;
  assign new_new_n6168__ = ~new_new_n6163__ & new_new_n6166__;
  assign new_new_n6169__ = ~new_new_n6167__ & ~new_new_n6168__;
  assign new_new_n6170__ = pi091 & ~new_new_n6169__;
  assign new_new_n6171__ = ~pi091 & new_new_n6169__;
  assign new_new_n6172__ = ~new_new_n5832__ & ~new_new_n5833__;
  assign new_new_n6173__ = ~new_new_n6105__ & po032;
  assign new_new_n6174__ = ~pi088 & ~po032;
  assign new_new_n6175__ = ~new_new_n6173__ & ~new_new_n6174__;
  assign new_new_n6176__ = new_new_n6172__ & ~new_new_n6175__;
  assign new_new_n6177__ = ~new_new_n6172__ & new_new_n6175__;
  assign new_new_n6178__ = ~new_new_n6176__ & ~new_new_n6177__;
  assign new_new_n6179__ = pi089 & ~new_new_n6178__;
  assign new_new_n6180__ = ~pi089 & new_new_n6178__;
  assign new_new_n6181__ = ~new_new_n6103__ & po032;
  assign new_new_n6182__ = pi087 & ~po032;
  assign new_new_n6183__ = ~new_new_n6181__ & ~new_new_n6182__;
  assign new_new_n6184__ = ~new_new_n5841__ & ~new_new_n5842__;
  assign new_new_n6185__ = ~new_new_n6183__ & new_new_n6184__;
  assign new_new_n6186__ = new_new_n6183__ & ~new_new_n6184__;
  assign new_new_n6187__ = ~new_new_n6185__ & ~new_new_n6186__;
  assign new_new_n6188__ = ~pi088 & ~new_new_n6187__;
  assign new_new_n6189__ = pi088 & new_new_n6187__;
  assign new_new_n6190__ = ~new_new_n5850__ & ~new_new_n5851__;
  assign new_new_n6191__ = ~new_new_n6101__ & po032;
  assign new_new_n6192__ = pi086 & ~po032;
  assign new_new_n6193__ = ~new_new_n6191__ & ~new_new_n6192__;
  assign new_new_n6194__ = new_new_n6190__ & new_new_n6193__;
  assign new_new_n6195__ = ~new_new_n6190__ & ~new_new_n6193__;
  assign new_new_n6196__ = ~new_new_n6194__ & ~new_new_n6195__;
  assign new_new_n6197__ = pi087 & ~new_new_n6196__;
  assign new_new_n6198__ = ~pi087 & new_new_n6196__;
  assign new_new_n6199__ = pi085 & ~new_new_n6099__;
  assign new_new_n6200__ = ~pi085 & new_new_n6099__;
  assign new_new_n6201__ = ~new_new_n6199__ & ~new_new_n6200__;
  assign new_new_n6202__ = po032 & new_new_n6201__;
  assign new_new_n6203__ = ~new_new_n5858__ & ~new_new_n6202__;
  assign new_new_n6204__ = new_new_n5858__ & new_new_n6202__;
  assign new_new_n6205__ = ~new_new_n6203__ & ~new_new_n6204__;
  assign new_new_n6206__ = pi086 & ~new_new_n6205__;
  assign new_new_n6207__ = ~pi086 & new_new_n6205__;
  assign new_new_n6208__ = ~new_new_n6097__ & po032;
  assign new_new_n6209__ = pi084 & ~po032;
  assign new_new_n6210__ = ~new_new_n6208__ & ~new_new_n6209__;
  assign new_new_n6211__ = ~new_new_n5868__ & ~new_new_n5869__;
  assign new_new_n6212__ = ~new_new_n6210__ & new_new_n6211__;
  assign new_new_n6213__ = new_new_n6210__ & ~new_new_n6211__;
  assign new_new_n6214__ = ~new_new_n6212__ & ~new_new_n6213__;
  assign new_new_n6215__ = pi085 & new_new_n6214__;
  assign new_new_n6216__ = ~pi085 & ~new_new_n6214__;
  assign new_new_n6217__ = ~new_new_n5877__ & ~new_new_n5878__;
  assign new_new_n6218__ = ~new_new_n6095__ & po032;
  assign new_new_n6219__ = pi083 & ~po032;
  assign new_new_n6220__ = ~new_new_n6218__ & ~new_new_n6219__;
  assign new_new_n6221__ = new_new_n6217__ & new_new_n6220__;
  assign new_new_n6222__ = ~new_new_n6217__ & ~new_new_n6220__;
  assign new_new_n6223__ = ~new_new_n6221__ & ~new_new_n6222__;
  assign new_new_n6224__ = pi084 & ~new_new_n6223__;
  assign new_new_n6225__ = ~pi084 & new_new_n6223__;
  assign new_new_n6226__ = new_new_n6093__ & po032;
  assign new_new_n6227__ = pi082 & ~po032;
  assign new_new_n6228__ = ~new_new_n6226__ & ~new_new_n6227__;
  assign new_new_n6229__ = ~new_new_n5886__ & ~new_new_n5887__;
  assign new_new_n6230__ = ~new_new_n6228__ & ~new_new_n6229__;
  assign new_new_n6231__ = new_new_n6228__ & new_new_n6229__;
  assign new_new_n6232__ = ~new_new_n6230__ & ~new_new_n6231__;
  assign new_new_n6233__ = pi083 & ~new_new_n6232__;
  assign new_new_n6234__ = ~pi083 & new_new_n6232__;
  assign new_new_n6235__ = ~new_new_n5895__ & ~new_new_n5896__;
  assign new_new_n6236__ = ~new_new_n6091__ & po032;
  assign new_new_n6237__ = pi081 & ~po032;
  assign new_new_n6238__ = ~new_new_n6236__ & ~new_new_n6237__;
  assign new_new_n6239__ = new_new_n6235__ & ~new_new_n6238__;
  assign new_new_n6240__ = ~new_new_n6235__ & new_new_n6238__;
  assign new_new_n6241__ = ~new_new_n6239__ & ~new_new_n6240__;
  assign new_new_n6242__ = pi082 & new_new_n6241__;
  assign new_new_n6243__ = ~pi082 & ~new_new_n6241__;
  assign new_new_n6244__ = ~new_new_n6089__ & po032;
  assign new_new_n6245__ = pi080 & ~po032;
  assign new_new_n6246__ = ~new_new_n6244__ & ~new_new_n6245__;
  assign new_new_n6247__ = ~new_new_n5904__ & ~new_new_n5905__;
  assign new_new_n6248__ = ~new_new_n6246__ & new_new_n6247__;
  assign new_new_n6249__ = new_new_n6246__ & ~new_new_n6247__;
  assign new_new_n6250__ = ~new_new_n6248__ & ~new_new_n6249__;
  assign new_new_n6251__ = pi081 & new_new_n6250__;
  assign new_new_n6252__ = ~pi081 & ~new_new_n6250__;
  assign new_new_n6253__ = pi079 & ~new_new_n6087__;
  assign new_new_n6254__ = ~pi079 & new_new_n6087__;
  assign new_new_n6255__ = ~new_new_n6253__ & ~new_new_n6254__;
  assign new_new_n6256__ = po032 & new_new_n6255__;
  assign new_new_n6257__ = new_new_n5912__ & new_new_n6256__;
  assign new_new_n6258__ = ~new_new_n5912__ & ~new_new_n6256__;
  assign new_new_n6259__ = ~new_new_n6257__ & ~new_new_n6258__;
  assign new_new_n6260__ = pi080 & ~new_new_n6259__;
  assign new_new_n6261__ = ~pi080 & new_new_n6259__;
  assign new_new_n6262__ = ~new_new_n5922__ & ~new_new_n5923__;
  assign new_new_n6263__ = ~new_new_n6085__ & po032;
  assign new_new_n6264__ = pi078 & ~po032;
  assign new_new_n6265__ = ~new_new_n6263__ & ~new_new_n6264__;
  assign new_new_n6266__ = new_new_n6262__ & ~new_new_n6265__;
  assign new_new_n6267__ = ~new_new_n6262__ & new_new_n6265__;
  assign new_new_n6268__ = ~new_new_n6266__ & ~new_new_n6267__;
  assign new_new_n6269__ = pi079 & new_new_n6268__;
  assign new_new_n6270__ = ~pi079 & ~new_new_n6268__;
  assign new_new_n6271__ = ~new_new_n6083__ & po032;
  assign new_new_n6272__ = pi077 & ~po032;
  assign new_new_n6273__ = ~new_new_n6271__ & ~new_new_n6272__;
  assign new_new_n6274__ = ~new_new_n5931__ & ~new_new_n5932__;
  assign new_new_n6275__ = ~new_new_n6273__ & new_new_n6274__;
  assign new_new_n6276__ = new_new_n6273__ & ~new_new_n6274__;
  assign new_new_n6277__ = ~new_new_n6275__ & ~new_new_n6276__;
  assign new_new_n6278__ = pi078 & new_new_n6277__;
  assign new_new_n6279__ = ~pi078 & ~new_new_n6277__;
  assign new_new_n6280__ = ~new_new_n5940__ & ~new_new_n5941__;
  assign new_new_n6281__ = ~new_new_n6081__ & po032;
  assign new_new_n6282__ = pi076 & ~po032;
  assign new_new_n6283__ = ~new_new_n6281__ & ~new_new_n6282__;
  assign new_new_n6284__ = new_new_n6280__ & new_new_n6283__;
  assign new_new_n6285__ = ~new_new_n6280__ & ~new_new_n6283__;
  assign new_new_n6286__ = ~new_new_n6284__ & ~new_new_n6285__;
  assign new_new_n6287__ = pi077 & ~new_new_n6286__;
  assign new_new_n6288__ = ~pi077 & new_new_n6286__;
  assign new_new_n6289__ = new_new_n6079__ & po032;
  assign new_new_n6290__ = pi075 & ~po032;
  assign new_new_n6291__ = ~new_new_n6289__ & ~new_new_n6290__;
  assign new_new_n6292__ = ~new_new_n5949__ & ~new_new_n5950__;
  assign new_new_n6293__ = ~new_new_n6291__ & ~new_new_n6292__;
  assign new_new_n6294__ = new_new_n6291__ & new_new_n6292__;
  assign new_new_n6295__ = ~new_new_n6293__ & ~new_new_n6294__;
  assign new_new_n6296__ = pi076 & ~new_new_n6295__;
  assign new_new_n6297__ = ~pi076 & new_new_n6295__;
  assign new_new_n6298__ = ~new_new_n5958__ & ~new_new_n5959__;
  assign new_new_n6299__ = ~new_new_n6077__ & po032;
  assign new_new_n6300__ = ~pi074 & ~po032;
  assign new_new_n6301__ = ~new_new_n6299__ & ~new_new_n6300__;
  assign new_new_n6302__ = new_new_n6298__ & ~new_new_n6301__;
  assign new_new_n6303__ = ~new_new_n6298__ & new_new_n6301__;
  assign new_new_n6304__ = ~new_new_n6302__ & ~new_new_n6303__;
  assign new_new_n6305__ = pi075 & ~new_new_n6304__;
  assign new_new_n6306__ = ~pi075 & new_new_n6304__;
  assign new_new_n6307__ = ~pi073 & ~new_new_n6075__;
  assign new_new_n6308__ = pi073 & new_new_n6075__;
  assign new_new_n6309__ = ~new_new_n6307__ & ~new_new_n6308__;
  assign new_new_n6310__ = po032 & new_new_n6309__;
  assign new_new_n6311__ = new_new_n5966__ & new_new_n6310__;
  assign new_new_n6312__ = ~new_new_n5966__ & ~new_new_n6310__;
  assign new_new_n6313__ = ~new_new_n6311__ & ~new_new_n6312__;
  assign new_new_n6314__ = ~pi074 & ~new_new_n6313__;
  assign new_new_n6315__ = pi074 & new_new_n6313__;
  assign new_new_n6316__ = ~new_new_n5976__ & ~new_new_n5977__;
  assign new_new_n6317__ = ~new_new_n6073__ & po032;
  assign new_new_n6318__ = ~pi072 & ~po032;
  assign new_new_n6319__ = ~new_new_n6317__ & ~new_new_n6318__;
  assign new_new_n6320__ = new_new_n6316__ & new_new_n6319__;
  assign new_new_n6321__ = ~new_new_n6316__ & ~new_new_n6319__;
  assign new_new_n6322__ = ~new_new_n6320__ & ~new_new_n6321__;
  assign new_new_n6323__ = ~pi073 & ~new_new_n6322__;
  assign new_new_n6324__ = pi073 & new_new_n6322__;
  assign new_new_n6325__ = ~new_new_n5985__ & ~new_new_n5986__;
  assign new_new_n6326__ = ~new_new_n6071__ & po032;
  assign new_new_n6327__ = ~pi071 & ~po032;
  assign new_new_n6328__ = ~new_new_n6326__ & ~new_new_n6327__;
  assign new_new_n6329__ = new_new_n6325__ & ~new_new_n6328__;
  assign new_new_n6330__ = ~new_new_n6325__ & new_new_n6328__;
  assign new_new_n6331__ = ~new_new_n6329__ & ~new_new_n6330__;
  assign new_new_n6332__ = ~pi072 & new_new_n6331__;
  assign new_new_n6333__ = pi072 & ~new_new_n6331__;
  assign new_new_n6334__ = new_new_n6069__ & po032;
  assign new_new_n6335__ = ~pi070 & ~po032;
  assign new_new_n6336__ = ~new_new_n6334__ & ~new_new_n6335__;
  assign new_new_n6337__ = ~new_new_n5994__ & ~new_new_n5995__;
  assign new_new_n6338__ = ~new_new_n6336__ & ~new_new_n6337__;
  assign new_new_n6339__ = new_new_n6336__ & new_new_n6337__;
  assign new_new_n6340__ = ~new_new_n6338__ & ~new_new_n6339__;
  assign new_new_n6341__ = ~pi071 & ~new_new_n6340__;
  assign new_new_n6342__ = pi071 & new_new_n6340__;
  assign new_new_n6343__ = ~new_new_n6003__ & ~new_new_n6004__;
  assign new_new_n6344__ = ~new_new_n6067__ & po032;
  assign new_new_n6345__ = pi069 & ~po032;
  assign new_new_n6346__ = ~new_new_n6344__ & ~new_new_n6345__;
  assign new_new_n6347__ = new_new_n6343__ & new_new_n6346__;
  assign new_new_n6348__ = ~new_new_n6343__ & ~new_new_n6346__;
  assign new_new_n6349__ = ~new_new_n6347__ & ~new_new_n6348__;
  assign new_new_n6350__ = ~pi070 & new_new_n6349__;
  assign new_new_n6351__ = pi070 & ~new_new_n6349__;
  assign new_new_n6352__ = new_new_n6065__ & po032;
  assign new_new_n6353__ = pi068 & ~po032;
  assign new_new_n6354__ = ~new_new_n6352__ & ~new_new_n6353__;
  assign new_new_n6355__ = ~new_new_n6012__ & ~new_new_n6013__;
  assign new_new_n6356__ = ~new_new_n6354__ & ~new_new_n6355__;
  assign new_new_n6357__ = new_new_n6354__ & new_new_n6355__;
  assign new_new_n6358__ = ~new_new_n6356__ & ~new_new_n6357__;
  assign new_new_n6359__ = ~pi069 & new_new_n6358__;
  assign new_new_n6360__ = pi069 & ~new_new_n6358__;
  assign new_new_n6361__ = ~new_new_n6019__ & ~new_new_n6020__;
  assign new_new_n6362__ = new_new_n6063__ & po032;
  assign new_new_n6363__ = ~pi067 & ~po032;
  assign new_new_n6364__ = ~new_new_n6362__ & ~new_new_n6363__;
  assign new_new_n6365__ = ~new_new_n6361__ & ~new_new_n6364__;
  assign new_new_n6366__ = new_new_n6361__ & new_new_n6364__;
  assign new_new_n6367__ = ~new_new_n6365__ & ~new_new_n6366__;
  assign new_new_n6368__ = ~pi068 & ~new_new_n6367__;
  assign new_new_n6369__ = pi068 & new_new_n6367__;
  assign new_new_n6370__ = ~new_new_n6033__ & ~new_new_n6034__;
  assign new_new_n6371__ = po032 & new_new_n6370__;
  assign new_new_n6372__ = new_new_n6061__ & ~new_new_n6371__;
  assign new_new_n6373__ = ~new_new_n6061__ & new_new_n6371__;
  assign new_new_n6374__ = ~new_new_n6372__ & ~new_new_n6373__;
  assign new_new_n6375__ = pi067 & new_new_n6374__;
  assign new_new_n6376__ = ~pi067 & ~new_new_n6374__;
  assign new_new_n6377__ = pi032 & po032;
  assign new_new_n6378__ = pi031 & ~pi065;
  assign new_new_n6379__ = new_new_n6377__ & ~new_new_n6378__;
  assign new_new_n6380__ = ~pi032 & ~po032;
  assign new_new_n6381__ = ~pi065 & ~new_new_n6380__;
  assign new_new_n6382__ = ~pi031 & ~new_new_n6381__;
  assign new_new_n6383__ = ~new_new_n6379__ & ~new_new_n6382__;
  assign new_new_n6384__ = pi064 & ~new_new_n6383__;
  assign new_new_n6385__ = pi064 & po032;
  assign new_new_n6386__ = ~pi032 & pi065;
  assign new_new_n6387__ = ~new_new_n6385__ & new_new_n6386__;
  assign new_new_n6388__ = ~new_new_n6384__ & ~new_new_n6387__;
  assign new_new_n6389__ = pi066 & ~new_new_n6388__;
  assign new_new_n6390__ = ~pi066 & new_new_n6388__;
  assign new_new_n6391__ = new_new_n426__ & ~po033;
  assign new_new_n6392__ = new_new_n6037__ & po032;
  assign new_new_n6393__ = ~new_new_n6391__ & ~new_new_n6392__;
  assign new_new_n6394__ = ~pi032 & ~new_new_n6393__;
  assign new_new_n6395__ = ~new_new_n332__ & po032;
  assign new_new_n6396__ = ~new_new_n6029__ & ~new_new_n6395__;
  assign new_new_n6397__ = pi065 & po032;
  assign new_new_n6398__ = po033 & ~new_new_n6397__;
  assign new_new_n6399__ = pi065 & ~new_new_n6029__;
  assign new_new_n6400__ = pi032 & ~new_new_n6399__;
  assign new_new_n6401__ = ~new_new_n6398__ & new_new_n6400__;
  assign new_new_n6402__ = ~new_new_n6394__ & ~new_new_n6396__;
  assign new_new_n6403__ = ~new_new_n6401__ & new_new_n6402__;
  assign new_new_n6404__ = pi033 & ~new_new_n6403__;
  assign new_new_n6405__ = ~new_new_n6029__ & ~new_new_n6397__;
  assign new_new_n6406__ = pi032 & ~new_new_n6035__;
  assign new_new_n6407__ = pi064 & ~new_new_n6406__;
  assign new_new_n6408__ = ~new_new_n6405__ & ~new_new_n6407__;
  assign new_new_n6409__ = ~pi065 & po032;
  assign new_new_n6410__ = ~po033 & ~new_new_n6409__;
  assign new_new_n6411__ = pi064 & ~new_new_n6377__;
  assign new_new_n6412__ = ~new_new_n6392__ & new_new_n6411__;
  assign new_new_n6413__ = ~new_new_n6410__ & new_new_n6412__;
  assign new_new_n6414__ = ~new_new_n6408__ & ~new_new_n6413__;
  assign new_new_n6415__ = ~pi033 & ~new_new_n6414__;
  assign new_new_n6416__ = ~new_new_n6404__ & ~new_new_n6415__;
  assign new_new_n6417__ = ~new_new_n6390__ & new_new_n6416__;
  assign new_new_n6418__ = ~new_new_n6389__ & ~new_new_n6417__;
  assign new_new_n6419__ = ~new_new_n6376__ & ~new_new_n6418__;
  assign new_new_n6420__ = ~new_new_n6375__ & ~new_new_n6419__;
  assign new_new_n6421__ = ~new_new_n6369__ & new_new_n6420__;
  assign new_new_n6422__ = ~new_new_n6368__ & ~new_new_n6421__;
  assign new_new_n6423__ = ~new_new_n6360__ & ~new_new_n6422__;
  assign new_new_n6424__ = ~new_new_n6359__ & ~new_new_n6423__;
  assign new_new_n6425__ = ~new_new_n6351__ & ~new_new_n6424__;
  assign new_new_n6426__ = ~new_new_n6350__ & ~new_new_n6425__;
  assign new_new_n6427__ = ~new_new_n6342__ & ~new_new_n6426__;
  assign new_new_n6428__ = ~new_new_n6341__ & ~new_new_n6427__;
  assign new_new_n6429__ = ~new_new_n6333__ & ~new_new_n6428__;
  assign new_new_n6430__ = ~new_new_n6332__ & ~new_new_n6429__;
  assign new_new_n6431__ = ~new_new_n6324__ & ~new_new_n6430__;
  assign new_new_n6432__ = ~new_new_n6323__ & ~new_new_n6431__;
  assign new_new_n6433__ = ~new_new_n6315__ & ~new_new_n6432__;
  assign new_new_n6434__ = ~new_new_n6314__ & ~new_new_n6433__;
  assign new_new_n6435__ = ~new_new_n6306__ & new_new_n6434__;
  assign new_new_n6436__ = ~new_new_n6305__ & ~new_new_n6435__;
  assign new_new_n6437__ = ~new_new_n6297__ & ~new_new_n6436__;
  assign new_new_n6438__ = ~new_new_n6296__ & ~new_new_n6437__;
  assign new_new_n6439__ = ~new_new_n6288__ & ~new_new_n6438__;
  assign new_new_n6440__ = ~new_new_n6287__ & ~new_new_n6439__;
  assign new_new_n6441__ = ~new_new_n6279__ & ~new_new_n6440__;
  assign new_new_n6442__ = ~new_new_n6278__ & ~new_new_n6441__;
  assign new_new_n6443__ = ~new_new_n6270__ & ~new_new_n6442__;
  assign new_new_n6444__ = ~new_new_n6269__ & ~new_new_n6443__;
  assign new_new_n6445__ = ~new_new_n6261__ & ~new_new_n6444__;
  assign new_new_n6446__ = ~new_new_n6260__ & ~new_new_n6445__;
  assign new_new_n6447__ = ~new_new_n6252__ & ~new_new_n6446__;
  assign new_new_n6448__ = ~new_new_n6251__ & ~new_new_n6447__;
  assign new_new_n6449__ = ~new_new_n6243__ & ~new_new_n6448__;
  assign new_new_n6450__ = ~new_new_n6242__ & ~new_new_n6449__;
  assign new_new_n6451__ = ~new_new_n6234__ & ~new_new_n6450__;
  assign new_new_n6452__ = ~new_new_n6233__ & ~new_new_n6451__;
  assign new_new_n6453__ = ~new_new_n6225__ & ~new_new_n6452__;
  assign new_new_n6454__ = ~new_new_n6224__ & ~new_new_n6453__;
  assign new_new_n6455__ = ~new_new_n6216__ & ~new_new_n6454__;
  assign new_new_n6456__ = ~new_new_n6215__ & ~new_new_n6455__;
  assign new_new_n6457__ = ~new_new_n6207__ & ~new_new_n6456__;
  assign new_new_n6458__ = ~new_new_n6206__ & ~new_new_n6457__;
  assign new_new_n6459__ = ~new_new_n6198__ & ~new_new_n6458__;
  assign new_new_n6460__ = ~new_new_n6197__ & ~new_new_n6459__;
  assign new_new_n6461__ = ~new_new_n6189__ & new_new_n6460__;
  assign new_new_n6462__ = ~new_new_n6188__ & ~new_new_n6461__;
  assign new_new_n6463__ = ~new_new_n6180__ & new_new_n6462__;
  assign new_new_n6464__ = ~new_new_n6179__ & ~new_new_n6463__;
  assign new_new_n6465__ = pi090 & ~new_new_n6464__;
  assign new_new_n6466__ = ~pi090 & new_new_n6464__;
  assign new_new_n6467__ = ~pi089 & ~new_new_n6107__;
  assign new_new_n6468__ = pi089 & new_new_n6107__;
  assign new_new_n6469__ = ~new_new_n6467__ & ~new_new_n6468__;
  assign new_new_n6470__ = po032 & new_new_n6469__;
  assign new_new_n6471__ = new_new_n5822__ & new_new_n6470__;
  assign new_new_n6472__ = ~new_new_n5822__ & ~new_new_n6470__;
  assign new_new_n6473__ = ~new_new_n6471__ & ~new_new_n6472__;
  assign new_new_n6474__ = ~new_new_n6466__ & new_new_n6473__;
  assign new_new_n6475__ = ~new_new_n6465__ & ~new_new_n6474__;
  assign new_new_n6476__ = ~new_new_n6171__ & ~new_new_n6475__;
  assign new_new_n6477__ = ~new_new_n6170__ & ~new_new_n6476__;
  assign new_new_n6478__ = ~new_new_n6162__ & ~new_new_n6477__;
  assign new_new_n6479__ = ~new_new_n6161__ & ~new_new_n6478__;
  assign new_new_n6480__ = ~new_new_n6153__ & ~new_new_n6479__;
  assign new_new_n6481__ = ~new_new_n6152__ & ~new_new_n6480__;
  assign new_new_n6482__ = ~new_new_n6144__ & ~new_new_n6481__;
  assign new_new_n6483__ = ~new_new_n6143__ & ~new_new_n6482__;
  assign new_new_n6484__ = ~new_new_n6130__ & ~new_new_n6483__;
  assign new_new_n6485__ = ~new_new_n6131__ & ~new_new_n6484__;
  assign new_new_n6486__ = ~pi096 & new_new_n6485__;
  assign new_new_n6487__ = ~new_new_n376__ & po032;
  assign new_new_n6488__ = ~new_new_n5778__ & ~new_new_n6487__;
  assign new_new_n6489__ = ~new_new_n6486__ & ~new_new_n6488__;
  assign new_new_n6490__ = pi096 & ~new_new_n6485__;
  assign new_new_n6491__ = new_new_n259__ & new_new_n287__;
  assign new_new_n6492__ = ~new_new_n6490__ & new_new_n6491__;
  assign po031 = ~new_new_n6489__ & new_new_n6492__;
  assign new_new_n6494__ = new_new_n6483__ & po031;
  assign new_new_n6495__ = ~pi095 & ~po031;
  assign new_new_n6496__ = ~new_new_n6494__ & ~new_new_n6495__;
  assign new_new_n6497__ = ~new_new_n6132__ & ~new_new_n6496__;
  assign new_new_n6498__ = new_new_n6132__ & new_new_n6496__;
  assign new_new_n6499__ = ~new_new_n6497__ & ~new_new_n6498__;
  assign new_new_n6500__ = ~new_new_n6143__ & ~new_new_n6144__;
  assign new_new_n6501__ = pi094 & ~po031;
  assign new_new_n6502__ = ~new_new_n6481__ & po031;
  assign new_new_n6503__ = ~new_new_n6501__ & ~new_new_n6502__;
  assign new_new_n6504__ = new_new_n6500__ & new_new_n6503__;
  assign new_new_n6505__ = ~new_new_n6500__ & ~new_new_n6503__;
  assign new_new_n6506__ = ~new_new_n6504__ & ~new_new_n6505__;
  assign new_new_n6507__ = pi095 & ~new_new_n6506__;
  assign new_new_n6508__ = ~pi095 & new_new_n6506__;
  assign new_new_n6509__ = ~new_new_n6152__ & ~new_new_n6153__;
  assign new_new_n6510__ = ~new_new_n6479__ & po031;
  assign new_new_n6511__ = pi093 & ~po031;
  assign new_new_n6512__ = ~new_new_n6510__ & ~new_new_n6511__;
  assign new_new_n6513__ = new_new_n6509__ & new_new_n6512__;
  assign new_new_n6514__ = ~new_new_n6509__ & ~new_new_n6512__;
  assign new_new_n6515__ = ~new_new_n6513__ & ~new_new_n6514__;
  assign new_new_n6516__ = pi094 & ~new_new_n6515__;
  assign new_new_n6517__ = ~pi094 & new_new_n6515__;
  assign new_new_n6518__ = new_new_n6477__ & po031;
  assign new_new_n6519__ = ~pi092 & ~po031;
  assign new_new_n6520__ = ~new_new_n6518__ & ~new_new_n6519__;
  assign new_new_n6521__ = ~new_new_n6161__ & ~new_new_n6162__;
  assign new_new_n6522__ = ~new_new_n6520__ & ~new_new_n6521__;
  assign new_new_n6523__ = new_new_n6520__ & new_new_n6521__;
  assign new_new_n6524__ = ~new_new_n6522__ & ~new_new_n6523__;
  assign new_new_n6525__ = ~pi093 & ~new_new_n6524__;
  assign new_new_n6526__ = pi093 & new_new_n6524__;
  assign new_new_n6527__ = pi091 & ~new_new_n6475__;
  assign new_new_n6528__ = ~pi091 & new_new_n6475__;
  assign new_new_n6529__ = ~new_new_n6527__ & ~new_new_n6528__;
  assign new_new_n6530__ = po031 & new_new_n6529__;
  assign new_new_n6531__ = new_new_n6169__ & new_new_n6530__;
  assign new_new_n6532__ = ~new_new_n6169__ & ~new_new_n6530__;
  assign new_new_n6533__ = ~new_new_n6531__ & ~new_new_n6532__;
  assign new_new_n6534__ = pi092 & ~new_new_n6533__;
  assign new_new_n6535__ = ~pi092 & new_new_n6533__;
  assign new_new_n6536__ = ~new_new_n6465__ & ~new_new_n6466__;
  assign new_new_n6537__ = po031 & new_new_n6536__;
  assign new_new_n6538__ = new_new_n6473__ & new_new_n6537__;
  assign new_new_n6539__ = ~new_new_n6473__ & ~new_new_n6537__;
  assign new_new_n6540__ = ~new_new_n6538__ & ~new_new_n6539__;
  assign new_new_n6541__ = ~pi091 & ~new_new_n6540__;
  assign new_new_n6542__ = pi091 & new_new_n6540__;
  assign new_new_n6543__ = ~new_new_n6179__ & ~new_new_n6180__;
  assign new_new_n6544__ = ~new_new_n6462__ & po031;
  assign new_new_n6545__ = ~pi089 & ~po031;
  assign new_new_n6546__ = ~new_new_n6544__ & ~new_new_n6545__;
  assign new_new_n6547__ = new_new_n6543__ & ~new_new_n6546__;
  assign new_new_n6548__ = ~new_new_n6543__ & new_new_n6546__;
  assign new_new_n6549__ = ~new_new_n6547__ & ~new_new_n6548__;
  assign new_new_n6550__ = pi090 & ~new_new_n6549__;
  assign new_new_n6551__ = ~pi090 & new_new_n6549__;
  assign new_new_n6552__ = ~new_new_n6460__ & po031;
  assign new_new_n6553__ = pi088 & ~po031;
  assign new_new_n6554__ = ~new_new_n6552__ & ~new_new_n6553__;
  assign new_new_n6555__ = ~new_new_n6188__ & ~new_new_n6189__;
  assign new_new_n6556__ = ~new_new_n6554__ & new_new_n6555__;
  assign new_new_n6557__ = new_new_n6554__ & ~new_new_n6555__;
  assign new_new_n6558__ = ~new_new_n6556__ & ~new_new_n6557__;
  assign new_new_n6559__ = pi089 & new_new_n6558__;
  assign new_new_n6560__ = ~pi089 & ~new_new_n6558__;
  assign new_new_n6561__ = pi087 & ~new_new_n6458__;
  assign new_new_n6562__ = ~pi087 & new_new_n6458__;
  assign new_new_n6563__ = ~new_new_n6561__ & ~new_new_n6562__;
  assign new_new_n6564__ = po031 & new_new_n6563__;
  assign new_new_n6565__ = new_new_n6196__ & new_new_n6564__;
  assign new_new_n6566__ = ~new_new_n6196__ & ~new_new_n6564__;
  assign new_new_n6567__ = ~new_new_n6565__ & ~new_new_n6566__;
  assign new_new_n6568__ = pi088 & ~new_new_n6567__;
  assign new_new_n6569__ = ~pi088 & new_new_n6567__;
  assign new_new_n6570__ = ~new_new_n6456__ & po031;
  assign new_new_n6571__ = pi086 & ~po031;
  assign new_new_n6572__ = ~new_new_n6570__ & ~new_new_n6571__;
  assign new_new_n6573__ = ~new_new_n6206__ & ~new_new_n6207__;
  assign new_new_n6574__ = ~new_new_n6572__ & new_new_n6573__;
  assign new_new_n6575__ = new_new_n6572__ & ~new_new_n6573__;
  assign new_new_n6576__ = ~new_new_n6574__ & ~new_new_n6575__;
  assign new_new_n6577__ = ~pi087 & ~new_new_n6576__;
  assign new_new_n6578__ = pi087 & new_new_n6576__;
  assign new_new_n6579__ = ~new_new_n6454__ & po031;
  assign new_new_n6580__ = pi085 & ~po031;
  assign new_new_n6581__ = ~new_new_n6579__ & ~new_new_n6580__;
  assign new_new_n6582__ = ~new_new_n6215__ & ~new_new_n6216__;
  assign new_new_n6583__ = ~new_new_n6581__ & new_new_n6582__;
  assign new_new_n6584__ = new_new_n6581__ & ~new_new_n6582__;
  assign new_new_n6585__ = ~new_new_n6583__ & ~new_new_n6584__;
  assign new_new_n6586__ = ~pi086 & ~new_new_n6585__;
  assign new_new_n6587__ = pi086 & new_new_n6585__;
  assign new_new_n6588__ = pi084 & ~new_new_n6452__;
  assign new_new_n6589__ = ~pi084 & new_new_n6452__;
  assign new_new_n6590__ = ~new_new_n6588__ & ~new_new_n6589__;
  assign new_new_n6591__ = po031 & new_new_n6590__;
  assign new_new_n6592__ = ~new_new_n6223__ & ~new_new_n6591__;
  assign new_new_n6593__ = new_new_n6223__ & new_new_n6591__;
  assign new_new_n6594__ = ~new_new_n6592__ & ~new_new_n6593__;
  assign new_new_n6595__ = ~pi085 & new_new_n6594__;
  assign new_new_n6596__ = pi085 & ~new_new_n6594__;
  assign new_new_n6597__ = ~new_new_n6233__ & ~new_new_n6234__;
  assign new_new_n6598__ = ~new_new_n6450__ & po031;
  assign new_new_n6599__ = pi083 & ~po031;
  assign new_new_n6600__ = ~new_new_n6598__ & ~new_new_n6599__;
  assign new_new_n6601__ = new_new_n6597__ & new_new_n6600__;
  assign new_new_n6602__ = ~new_new_n6597__ & ~new_new_n6600__;
  assign new_new_n6603__ = ~new_new_n6601__ & ~new_new_n6602__;
  assign new_new_n6604__ = ~pi084 & new_new_n6603__;
  assign new_new_n6605__ = pi084 & ~new_new_n6603__;
  assign new_new_n6606__ = new_new_n6448__ & po031;
  assign new_new_n6607__ = ~pi082 & ~po031;
  assign new_new_n6608__ = ~new_new_n6606__ & ~new_new_n6607__;
  assign new_new_n6609__ = ~new_new_n6242__ & ~new_new_n6243__;
  assign new_new_n6610__ = ~new_new_n6608__ & ~new_new_n6609__;
  assign new_new_n6611__ = new_new_n6608__ & new_new_n6609__;
  assign new_new_n6612__ = ~new_new_n6610__ & ~new_new_n6611__;
  assign new_new_n6613__ = ~pi083 & ~new_new_n6612__;
  assign new_new_n6614__ = pi083 & new_new_n6612__;
  assign new_new_n6615__ = new_new_n6446__ & po031;
  assign new_new_n6616__ = ~pi081 & ~po031;
  assign new_new_n6617__ = ~new_new_n6615__ & ~new_new_n6616__;
  assign new_new_n6618__ = ~new_new_n6251__ & ~new_new_n6252__;
  assign new_new_n6619__ = ~new_new_n6617__ & ~new_new_n6618__;
  assign new_new_n6620__ = new_new_n6617__ & new_new_n6618__;
  assign new_new_n6621__ = ~new_new_n6619__ & ~new_new_n6620__;
  assign new_new_n6622__ = ~pi082 & ~new_new_n6621__;
  assign new_new_n6623__ = pi082 & new_new_n6621__;
  assign new_new_n6624__ = ~new_new_n6260__ & ~new_new_n6261__;
  assign new_new_n6625__ = ~new_new_n6444__ & po031;
  assign new_new_n6626__ = pi080 & ~po031;
  assign new_new_n6627__ = ~new_new_n6625__ & ~new_new_n6626__;
  assign new_new_n6628__ = new_new_n6624__ & new_new_n6627__;
  assign new_new_n6629__ = ~new_new_n6624__ & ~new_new_n6627__;
  assign new_new_n6630__ = ~new_new_n6628__ & ~new_new_n6629__;
  assign new_new_n6631__ = pi081 & ~new_new_n6630__;
  assign new_new_n6632__ = ~pi081 & new_new_n6630__;
  assign new_new_n6633__ = new_new_n6442__ & po031;
  assign new_new_n6634__ = ~pi079 & ~po031;
  assign new_new_n6635__ = ~new_new_n6633__ & ~new_new_n6634__;
  assign new_new_n6636__ = ~new_new_n6269__ & ~new_new_n6270__;
  assign new_new_n6637__ = ~new_new_n6635__ & ~new_new_n6636__;
  assign new_new_n6638__ = new_new_n6635__ & new_new_n6636__;
  assign new_new_n6639__ = ~new_new_n6637__ & ~new_new_n6638__;
  assign new_new_n6640__ = pi080 & new_new_n6639__;
  assign new_new_n6641__ = ~pi080 & ~new_new_n6639__;
  assign new_new_n6642__ = new_new_n6440__ & po031;
  assign new_new_n6643__ = ~pi078 & ~po031;
  assign new_new_n6644__ = ~new_new_n6642__ & ~new_new_n6643__;
  assign new_new_n6645__ = ~new_new_n6278__ & ~new_new_n6279__;
  assign new_new_n6646__ = ~new_new_n6644__ & ~new_new_n6645__;
  assign new_new_n6647__ = new_new_n6644__ & new_new_n6645__;
  assign new_new_n6648__ = ~new_new_n6646__ & ~new_new_n6647__;
  assign new_new_n6649__ = pi079 & new_new_n6648__;
  assign new_new_n6650__ = ~pi079 & ~new_new_n6648__;
  assign new_new_n6651__ = ~new_new_n6287__ & ~new_new_n6288__;
  assign new_new_n6652__ = ~new_new_n6438__ & po031;
  assign new_new_n6653__ = pi077 & ~po031;
  assign new_new_n6654__ = ~new_new_n6652__ & ~new_new_n6653__;
  assign new_new_n6655__ = new_new_n6651__ & new_new_n6654__;
  assign new_new_n6656__ = ~new_new_n6651__ & ~new_new_n6654__;
  assign new_new_n6657__ = ~new_new_n6655__ & ~new_new_n6656__;
  assign new_new_n6658__ = pi078 & ~new_new_n6657__;
  assign new_new_n6659__ = ~pi078 & new_new_n6657__;
  assign new_new_n6660__ = pi076 & ~new_new_n6436__;
  assign new_new_n6661__ = ~pi076 & new_new_n6436__;
  assign new_new_n6662__ = ~new_new_n6660__ & ~new_new_n6661__;
  assign new_new_n6663__ = po031 & new_new_n6662__;
  assign new_new_n6664__ = ~new_new_n6295__ & ~new_new_n6663__;
  assign new_new_n6665__ = new_new_n6295__ & new_new_n6663__;
  assign new_new_n6666__ = ~new_new_n6664__ & ~new_new_n6665__;
  assign new_new_n6667__ = pi077 & ~new_new_n6666__;
  assign new_new_n6668__ = ~pi077 & new_new_n6666__;
  assign new_new_n6669__ = new_new_n6434__ & po031;
  assign new_new_n6670__ = pi075 & ~po031;
  assign new_new_n6671__ = ~new_new_n6669__ & ~new_new_n6670__;
  assign new_new_n6672__ = ~new_new_n6305__ & ~new_new_n6306__;
  assign new_new_n6673__ = ~new_new_n6671__ & ~new_new_n6672__;
  assign new_new_n6674__ = new_new_n6671__ & new_new_n6672__;
  assign new_new_n6675__ = ~new_new_n6673__ & ~new_new_n6674__;
  assign new_new_n6676__ = pi076 & ~new_new_n6675__;
  assign new_new_n6677__ = ~pi076 & new_new_n6675__;
  assign new_new_n6678__ = ~new_new_n6314__ & ~new_new_n6315__;
  assign new_new_n6679__ = ~new_new_n6432__ & po031;
  assign new_new_n6680__ = ~pi074 & ~po031;
  assign new_new_n6681__ = ~new_new_n6679__ & ~new_new_n6680__;
  assign new_new_n6682__ = ~new_new_n6678__ & ~new_new_n6681__;
  assign new_new_n6683__ = new_new_n6678__ & new_new_n6681__;
  assign new_new_n6684__ = ~new_new_n6682__ & ~new_new_n6683__;
  assign new_new_n6685__ = ~pi075 & ~new_new_n6684__;
  assign new_new_n6686__ = pi075 & new_new_n6684__;
  assign new_new_n6687__ = ~new_new_n6323__ & ~new_new_n6324__;
  assign new_new_n6688__ = ~new_new_n6430__ & po031;
  assign new_new_n6689__ = ~pi073 & ~po031;
  assign new_new_n6690__ = ~new_new_n6688__ & ~new_new_n6689__;
  assign new_new_n6691__ = ~new_new_n6687__ & ~new_new_n6690__;
  assign new_new_n6692__ = new_new_n6687__ & new_new_n6690__;
  assign new_new_n6693__ = ~new_new_n6691__ & ~new_new_n6692__;
  assign new_new_n6694__ = ~pi074 & ~new_new_n6693__;
  assign new_new_n6695__ = pi074 & new_new_n6693__;
  assign new_new_n6696__ = new_new_n6428__ & po031;
  assign new_new_n6697__ = pi072 & ~po031;
  assign new_new_n6698__ = ~new_new_n6696__ & ~new_new_n6697__;
  assign new_new_n6699__ = ~new_new_n6332__ & ~new_new_n6333__;
  assign new_new_n6700__ = ~new_new_n6698__ & ~new_new_n6699__;
  assign new_new_n6701__ = new_new_n6698__ & new_new_n6699__;
  assign new_new_n6702__ = ~new_new_n6700__ & ~new_new_n6701__;
  assign new_new_n6703__ = pi073 & ~new_new_n6702__;
  assign new_new_n6704__ = ~pi073 & new_new_n6702__;
  assign new_new_n6705__ = ~new_new_n6341__ & ~new_new_n6342__;
  assign new_new_n6706__ = ~new_new_n6426__ & po031;
  assign new_new_n6707__ = ~pi071 & ~po031;
  assign new_new_n6708__ = ~new_new_n6706__ & ~new_new_n6707__;
  assign new_new_n6709__ = new_new_n6705__ & ~new_new_n6708__;
  assign new_new_n6710__ = ~new_new_n6705__ & new_new_n6708__;
  assign new_new_n6711__ = ~new_new_n6709__ & ~new_new_n6710__;
  assign new_new_n6712__ = pi072 & ~new_new_n6711__;
  assign new_new_n6713__ = ~pi072 & new_new_n6711__;
  assign new_new_n6714__ = ~new_new_n6350__ & ~new_new_n6351__;
  assign new_new_n6715__ = ~new_new_n6424__ & po031;
  assign new_new_n6716__ = ~pi070 & ~po031;
  assign new_new_n6717__ = ~new_new_n6715__ & ~new_new_n6716__;
  assign new_new_n6718__ = new_new_n6714__ & ~new_new_n6717__;
  assign new_new_n6719__ = ~new_new_n6714__ & new_new_n6717__;
  assign new_new_n6720__ = ~new_new_n6718__ & ~new_new_n6719__;
  assign new_new_n6721__ = pi071 & ~new_new_n6720__;
  assign new_new_n6722__ = ~pi071 & new_new_n6720__;
  assign new_new_n6723__ = ~new_new_n6359__ & ~new_new_n6360__;
  assign new_new_n6724__ = ~new_new_n6422__ & po031;
  assign new_new_n6725__ = ~pi069 & ~po031;
  assign new_new_n6726__ = ~new_new_n6724__ & ~new_new_n6725__;
  assign new_new_n6727__ = new_new_n6723__ & ~new_new_n6726__;
  assign new_new_n6728__ = ~new_new_n6723__ & new_new_n6726__;
  assign new_new_n6729__ = ~new_new_n6727__ & ~new_new_n6728__;
  assign new_new_n6730__ = pi070 & ~new_new_n6729__;
  assign new_new_n6731__ = ~pi070 & new_new_n6729__;
  assign new_new_n6732__ = new_new_n6420__ & po031;
  assign new_new_n6733__ = ~pi068 & ~po031;
  assign new_new_n6734__ = ~new_new_n6732__ & ~new_new_n6733__;
  assign new_new_n6735__ = ~new_new_n6368__ & ~new_new_n6369__;
  assign new_new_n6736__ = ~new_new_n6734__ & ~new_new_n6735__;
  assign new_new_n6737__ = new_new_n6734__ & new_new_n6735__;
  assign new_new_n6738__ = ~new_new_n6736__ & ~new_new_n6737__;
  assign new_new_n6739__ = ~pi069 & ~new_new_n6738__;
  assign new_new_n6740__ = pi069 & new_new_n6738__;
  assign new_new_n6741__ = ~new_new_n6375__ & ~new_new_n6376__;
  assign new_new_n6742__ = ~new_new_n6418__ & po031;
  assign new_new_n6743__ = pi067 & ~po031;
  assign new_new_n6744__ = ~new_new_n6742__ & ~new_new_n6743__;
  assign new_new_n6745__ = new_new_n6741__ & ~new_new_n6744__;
  assign new_new_n6746__ = ~new_new_n6741__ & new_new_n6744__;
  assign new_new_n6747__ = ~new_new_n6745__ & ~new_new_n6746__;
  assign new_new_n6748__ = pi068 & new_new_n6747__;
  assign new_new_n6749__ = ~pi068 & ~new_new_n6747__;
  assign new_new_n6750__ = ~new_new_n6389__ & ~new_new_n6390__;
  assign new_new_n6751__ = po031 & new_new_n6750__;
  assign new_new_n6752__ = ~new_new_n6416__ & new_new_n6751__;
  assign new_new_n6753__ = new_new_n6416__ & ~new_new_n6751__;
  assign new_new_n6754__ = ~new_new_n6752__ & ~new_new_n6753__;
  assign new_new_n6755__ = pi067 & ~new_new_n6754__;
  assign new_new_n6756__ = ~pi067 & new_new_n6754__;
  assign new_new_n6757__ = pi031 & po031;
  assign new_new_n6758__ = pi030 & ~pi065;
  assign new_new_n6759__ = new_new_n6757__ & ~new_new_n6758__;
  assign new_new_n6760__ = ~pi031 & ~po031;
  assign new_new_n6761__ = ~pi065 & ~new_new_n6760__;
  assign new_new_n6762__ = ~pi030 & ~new_new_n6761__;
  assign new_new_n6763__ = ~new_new_n6759__ & ~new_new_n6762__;
  assign new_new_n6764__ = pi064 & ~new_new_n6763__;
  assign new_new_n6765__ = pi064 & po031;
  assign new_new_n6766__ = ~pi031 & pi065;
  assign new_new_n6767__ = ~new_new_n6765__ & new_new_n6766__;
  assign new_new_n6768__ = ~new_new_n6764__ & ~new_new_n6767__;
  assign new_new_n6769__ = pi066 & ~new_new_n6768__;
  assign new_new_n6770__ = ~pi066 & new_new_n6768__;
  assign new_new_n6771__ = new_new_n426__ & ~po032;
  assign new_new_n6772__ = new_new_n6409__ & po031;
  assign new_new_n6773__ = ~new_new_n6771__ & ~new_new_n6772__;
  assign new_new_n6774__ = ~pi031 & ~new_new_n6773__;
  assign new_new_n6775__ = ~new_new_n332__ & po031;
  assign new_new_n6776__ = ~new_new_n6385__ & ~new_new_n6775__;
  assign new_new_n6777__ = pi065 & po031;
  assign new_new_n6778__ = po032 & ~new_new_n6777__;
  assign new_new_n6779__ = pi065 & ~new_new_n6385__;
  assign new_new_n6780__ = pi031 & ~new_new_n6779__;
  assign new_new_n6781__ = ~new_new_n6778__ & new_new_n6780__;
  assign new_new_n6782__ = ~new_new_n6774__ & ~new_new_n6776__;
  assign new_new_n6783__ = ~new_new_n6781__ & new_new_n6782__;
  assign new_new_n6784__ = pi032 & ~new_new_n6783__;
  assign new_new_n6785__ = ~new_new_n6385__ & ~new_new_n6777__;
  assign new_new_n6786__ = pi031 & ~new_new_n6397__;
  assign new_new_n6787__ = pi064 & ~new_new_n6786__;
  assign new_new_n6788__ = ~new_new_n6785__ & ~new_new_n6787__;
  assign new_new_n6789__ = ~pi065 & po031;
  assign new_new_n6790__ = ~po032 & ~new_new_n6789__;
  assign new_new_n6791__ = pi064 & ~new_new_n6757__;
  assign new_new_n6792__ = ~new_new_n6772__ & new_new_n6791__;
  assign new_new_n6793__ = ~new_new_n6790__ & new_new_n6792__;
  assign new_new_n6794__ = ~new_new_n6788__ & ~new_new_n6793__;
  assign new_new_n6795__ = ~pi032 & ~new_new_n6794__;
  assign new_new_n6796__ = ~new_new_n6784__ & ~new_new_n6795__;
  assign new_new_n6797__ = ~new_new_n6770__ & new_new_n6796__;
  assign new_new_n6798__ = ~new_new_n6769__ & ~new_new_n6797__;
  assign new_new_n6799__ = ~new_new_n6756__ & ~new_new_n6798__;
  assign new_new_n6800__ = ~new_new_n6755__ & ~new_new_n6799__;
  assign new_new_n6801__ = ~new_new_n6749__ & ~new_new_n6800__;
  assign new_new_n6802__ = ~new_new_n6748__ & ~new_new_n6801__;
  assign new_new_n6803__ = ~new_new_n6740__ & new_new_n6802__;
  assign new_new_n6804__ = ~new_new_n6739__ & ~new_new_n6803__;
  assign new_new_n6805__ = ~new_new_n6731__ & new_new_n6804__;
  assign new_new_n6806__ = ~new_new_n6730__ & ~new_new_n6805__;
  assign new_new_n6807__ = ~new_new_n6722__ & ~new_new_n6806__;
  assign new_new_n6808__ = ~new_new_n6721__ & ~new_new_n6807__;
  assign new_new_n6809__ = ~new_new_n6713__ & ~new_new_n6808__;
  assign new_new_n6810__ = ~new_new_n6712__ & ~new_new_n6809__;
  assign new_new_n6811__ = ~new_new_n6704__ & ~new_new_n6810__;
  assign new_new_n6812__ = ~new_new_n6703__ & ~new_new_n6811__;
  assign new_new_n6813__ = ~new_new_n6695__ & new_new_n6812__;
  assign new_new_n6814__ = ~new_new_n6694__ & ~new_new_n6813__;
  assign new_new_n6815__ = ~new_new_n6686__ & ~new_new_n6814__;
  assign new_new_n6816__ = ~new_new_n6685__ & ~new_new_n6815__;
  assign new_new_n6817__ = ~new_new_n6677__ & new_new_n6816__;
  assign new_new_n6818__ = ~new_new_n6676__ & ~new_new_n6817__;
  assign new_new_n6819__ = ~new_new_n6668__ & ~new_new_n6818__;
  assign new_new_n6820__ = ~new_new_n6667__ & ~new_new_n6819__;
  assign new_new_n6821__ = ~new_new_n6659__ & ~new_new_n6820__;
  assign new_new_n6822__ = ~new_new_n6658__ & ~new_new_n6821__;
  assign new_new_n6823__ = ~new_new_n6650__ & ~new_new_n6822__;
  assign new_new_n6824__ = ~new_new_n6649__ & ~new_new_n6823__;
  assign new_new_n6825__ = ~new_new_n6641__ & ~new_new_n6824__;
  assign new_new_n6826__ = ~new_new_n6640__ & ~new_new_n6825__;
  assign new_new_n6827__ = ~new_new_n6632__ & ~new_new_n6826__;
  assign new_new_n6828__ = ~new_new_n6631__ & ~new_new_n6827__;
  assign new_new_n6829__ = ~new_new_n6623__ & new_new_n6828__;
  assign new_new_n6830__ = ~new_new_n6622__ & ~new_new_n6829__;
  assign new_new_n6831__ = ~new_new_n6614__ & ~new_new_n6830__;
  assign new_new_n6832__ = ~new_new_n6613__ & ~new_new_n6831__;
  assign new_new_n6833__ = ~new_new_n6605__ & ~new_new_n6832__;
  assign new_new_n6834__ = ~new_new_n6604__ & ~new_new_n6833__;
  assign new_new_n6835__ = ~new_new_n6596__ & ~new_new_n6834__;
  assign new_new_n6836__ = ~new_new_n6595__ & ~new_new_n6835__;
  assign new_new_n6837__ = ~new_new_n6587__ & ~new_new_n6836__;
  assign new_new_n6838__ = ~new_new_n6586__ & ~new_new_n6837__;
  assign new_new_n6839__ = ~new_new_n6578__ & ~new_new_n6838__;
  assign new_new_n6840__ = ~new_new_n6577__ & ~new_new_n6839__;
  assign new_new_n6841__ = ~new_new_n6569__ & new_new_n6840__;
  assign new_new_n6842__ = ~new_new_n6568__ & ~new_new_n6841__;
  assign new_new_n6843__ = ~new_new_n6560__ & ~new_new_n6842__;
  assign new_new_n6844__ = ~new_new_n6559__ & ~new_new_n6843__;
  assign new_new_n6845__ = ~new_new_n6551__ & ~new_new_n6844__;
  assign new_new_n6846__ = ~new_new_n6550__ & ~new_new_n6845__;
  assign new_new_n6847__ = ~new_new_n6542__ & new_new_n6846__;
  assign new_new_n6848__ = ~new_new_n6541__ & ~new_new_n6847__;
  assign new_new_n6849__ = ~new_new_n6535__ & new_new_n6848__;
  assign new_new_n6850__ = ~new_new_n6534__ & ~new_new_n6849__;
  assign new_new_n6851__ = ~new_new_n6526__ & new_new_n6850__;
  assign new_new_n6852__ = ~new_new_n6525__ & ~new_new_n6851__;
  assign new_new_n6853__ = ~new_new_n6517__ & new_new_n6852__;
  assign new_new_n6854__ = ~new_new_n6516__ & ~new_new_n6853__;
  assign new_new_n6855__ = ~new_new_n6508__ & ~new_new_n6854__;
  assign new_new_n6856__ = ~new_new_n6507__ & ~new_new_n6855__;
  assign new_new_n6857__ = ~pi096 & new_new_n6856__;
  assign new_new_n6858__ = pi096 & ~new_new_n6856__;
  assign new_new_n6859__ = new_new_n6488__ & ~new_new_n6492__;
  assign new_new_n6860__ = ~new_new_n376__ & ~new_new_n6859__;
  assign new_new_n6861__ = pi097 & new_new_n6860__;
  assign new_new_n6862__ = ~new_new_n6499__ & ~new_new_n6858__;
  assign new_new_n6863__ = ~pi097 & ~new_new_n6860__;
  assign new_new_n6864__ = ~new_new_n6857__ & ~new_new_n6863__;
  assign new_new_n6865__ = ~new_new_n6862__ & new_new_n6864__;
  assign new_new_n6866__ = ~pi098 & new_new_n287__;
  assign new_new_n6867__ = ~new_new_n6861__ & new_new_n6866__;
  assign po030 = ~new_new_n6865__ & new_new_n6867__;
  assign new_new_n6869__ = ~new_new_n6857__ & ~new_new_n6858__;
  assign new_new_n6870__ = po030 & new_new_n6869__;
  assign new_new_n6871__ = ~new_new_n6499__ & ~new_new_n6870__;
  assign new_new_n6872__ = new_new_n6499__ & new_new_n6870__;
  assign new_new_n6873__ = ~new_new_n6871__ & ~new_new_n6872__;
  assign new_new_n6874__ = ~pi097 & ~new_new_n6873__;
  assign new_new_n6875__ = pi097 & new_new_n6873__;
  assign new_new_n6876__ = ~new_new_n6507__ & ~new_new_n6508__;
  assign new_new_n6877__ = ~new_new_n6854__ & po030;
  assign new_new_n6878__ = pi095 & ~po030;
  assign new_new_n6879__ = ~new_new_n6877__ & ~new_new_n6878__;
  assign new_new_n6880__ = new_new_n6876__ & ~new_new_n6879__;
  assign new_new_n6881__ = ~new_new_n6876__ & new_new_n6879__;
  assign new_new_n6882__ = ~new_new_n6880__ & ~new_new_n6881__;
  assign new_new_n6883__ = ~pi096 & ~new_new_n6882__;
  assign new_new_n6884__ = pi096 & new_new_n6882__;
  assign new_new_n6885__ = ~new_new_n6516__ & ~new_new_n6517__;
  assign new_new_n6886__ = ~new_new_n6852__ & po030;
  assign new_new_n6887__ = ~pi094 & ~po030;
  assign new_new_n6888__ = ~new_new_n6886__ & ~new_new_n6887__;
  assign new_new_n6889__ = new_new_n6885__ & ~new_new_n6888__;
  assign new_new_n6890__ = ~new_new_n6885__ & new_new_n6888__;
  assign new_new_n6891__ = ~new_new_n6889__ & ~new_new_n6890__;
  assign new_new_n6892__ = ~pi095 & new_new_n6891__;
  assign new_new_n6893__ = pi095 & ~new_new_n6891__;
  assign new_new_n6894__ = ~new_new_n6525__ & ~new_new_n6526__;
  assign new_new_n6895__ = ~new_new_n6850__ & po030;
  assign new_new_n6896__ = pi093 & ~po030;
  assign new_new_n6897__ = ~new_new_n6895__ & ~new_new_n6896__;
  assign new_new_n6898__ = new_new_n6894__ & ~new_new_n6897__;
  assign new_new_n6899__ = ~new_new_n6894__ & new_new_n6897__;
  assign new_new_n6900__ = ~new_new_n6898__ & ~new_new_n6899__;
  assign new_new_n6901__ = ~pi094 & ~new_new_n6900__;
  assign new_new_n6902__ = pi094 & new_new_n6900__;
  assign new_new_n6903__ = ~new_new_n6534__ & ~new_new_n6535__;
  assign new_new_n6904__ = ~new_new_n6848__ & po030;
  assign new_new_n6905__ = ~pi092 & ~po030;
  assign new_new_n6906__ = ~new_new_n6904__ & ~new_new_n6905__;
  assign new_new_n6907__ = new_new_n6903__ & ~new_new_n6906__;
  assign new_new_n6908__ = ~new_new_n6903__ & new_new_n6906__;
  assign new_new_n6909__ = ~new_new_n6907__ & ~new_new_n6908__;
  assign new_new_n6910__ = pi093 & ~new_new_n6909__;
  assign new_new_n6911__ = ~pi093 & new_new_n6909__;
  assign new_new_n6912__ = ~new_new_n6846__ & po030;
  assign new_new_n6913__ = pi091 & ~po030;
  assign new_new_n6914__ = ~new_new_n6912__ & ~new_new_n6913__;
  assign new_new_n6915__ = ~new_new_n6541__ & ~new_new_n6542__;
  assign new_new_n6916__ = ~new_new_n6914__ & new_new_n6915__;
  assign new_new_n6917__ = new_new_n6914__ & ~new_new_n6915__;
  assign new_new_n6918__ = ~new_new_n6916__ & ~new_new_n6917__;
  assign new_new_n6919__ = ~pi092 & ~new_new_n6918__;
  assign new_new_n6920__ = pi092 & new_new_n6918__;
  assign new_new_n6921__ = ~new_new_n6550__ & ~new_new_n6551__;
  assign new_new_n6922__ = ~new_new_n6844__ & po030;
  assign new_new_n6923__ = pi090 & ~po030;
  assign new_new_n6924__ = ~new_new_n6922__ & ~new_new_n6923__;
  assign new_new_n6925__ = new_new_n6921__ & new_new_n6924__;
  assign new_new_n6926__ = ~new_new_n6921__ & ~new_new_n6924__;
  assign new_new_n6927__ = ~new_new_n6925__ & ~new_new_n6926__;
  assign new_new_n6928__ = pi091 & ~new_new_n6927__;
  assign new_new_n6929__ = ~pi091 & new_new_n6927__;
  assign new_new_n6930__ = new_new_n6842__ & po030;
  assign new_new_n6931__ = ~pi089 & ~po030;
  assign new_new_n6932__ = ~new_new_n6930__ & ~new_new_n6931__;
  assign new_new_n6933__ = ~new_new_n6559__ & ~new_new_n6560__;
  assign new_new_n6934__ = ~new_new_n6932__ & ~new_new_n6933__;
  assign new_new_n6935__ = new_new_n6932__ & new_new_n6933__;
  assign new_new_n6936__ = ~new_new_n6934__ & ~new_new_n6935__;
  assign new_new_n6937__ = pi090 & new_new_n6936__;
  assign new_new_n6938__ = ~pi090 & ~new_new_n6936__;
  assign new_new_n6939__ = new_new_n6840__ & po030;
  assign new_new_n6940__ = pi088 & ~po030;
  assign new_new_n6941__ = ~new_new_n6939__ & ~new_new_n6940__;
  assign new_new_n6942__ = ~new_new_n6568__ & ~new_new_n6569__;
  assign new_new_n6943__ = ~new_new_n6941__ & ~new_new_n6942__;
  assign new_new_n6944__ = new_new_n6941__ & new_new_n6942__;
  assign new_new_n6945__ = ~new_new_n6943__ & ~new_new_n6944__;
  assign new_new_n6946__ = pi089 & ~new_new_n6945__;
  assign new_new_n6947__ = ~pi089 & new_new_n6945__;
  assign new_new_n6948__ = ~pi087 & ~new_new_n6838__;
  assign new_new_n6949__ = pi087 & new_new_n6838__;
  assign new_new_n6950__ = ~new_new_n6948__ & ~new_new_n6949__;
  assign new_new_n6951__ = po030 & new_new_n6950__;
  assign new_new_n6952__ = new_new_n6576__ & new_new_n6951__;
  assign new_new_n6953__ = ~new_new_n6576__ & ~new_new_n6951__;
  assign new_new_n6954__ = ~new_new_n6952__ & ~new_new_n6953__;
  assign new_new_n6955__ = pi088 & new_new_n6954__;
  assign new_new_n6956__ = ~pi088 & ~new_new_n6954__;
  assign new_new_n6957__ = ~pi086 & ~new_new_n6836__;
  assign new_new_n6958__ = pi086 & new_new_n6836__;
  assign new_new_n6959__ = ~new_new_n6957__ & ~new_new_n6958__;
  assign new_new_n6960__ = po030 & new_new_n6959__;
  assign new_new_n6961__ = new_new_n6585__ & new_new_n6960__;
  assign new_new_n6962__ = ~new_new_n6585__ & ~new_new_n6960__;
  assign new_new_n6963__ = ~new_new_n6961__ & ~new_new_n6962__;
  assign new_new_n6964__ = pi087 & new_new_n6963__;
  assign new_new_n6965__ = ~pi087 & ~new_new_n6963__;
  assign new_new_n6966__ = ~new_new_n6595__ & ~new_new_n6596__;
  assign new_new_n6967__ = ~new_new_n6834__ & po030;
  assign new_new_n6968__ = ~pi085 & ~po030;
  assign new_new_n6969__ = ~new_new_n6967__ & ~new_new_n6968__;
  assign new_new_n6970__ = new_new_n6966__ & new_new_n6969__;
  assign new_new_n6971__ = ~new_new_n6966__ & ~new_new_n6969__;
  assign new_new_n6972__ = ~new_new_n6970__ & ~new_new_n6971__;
  assign new_new_n6973__ = pi086 & new_new_n6972__;
  assign new_new_n6974__ = ~pi086 & ~new_new_n6972__;
  assign new_new_n6975__ = new_new_n6832__ & po030;
  assign new_new_n6976__ = pi084 & ~po030;
  assign new_new_n6977__ = ~new_new_n6975__ & ~new_new_n6976__;
  assign new_new_n6978__ = ~new_new_n6604__ & ~new_new_n6605__;
  assign new_new_n6979__ = ~new_new_n6977__ & ~new_new_n6978__;
  assign new_new_n6980__ = new_new_n6977__ & new_new_n6978__;
  assign new_new_n6981__ = ~new_new_n6979__ & ~new_new_n6980__;
  assign new_new_n6982__ = pi085 & ~new_new_n6981__;
  assign new_new_n6983__ = ~pi085 & new_new_n6981__;
  assign new_new_n6984__ = ~pi083 & ~new_new_n6830__;
  assign new_new_n6985__ = pi083 & new_new_n6830__;
  assign new_new_n6986__ = ~new_new_n6984__ & ~new_new_n6985__;
  assign new_new_n6987__ = po030 & new_new_n6986__;
  assign new_new_n6988__ = ~new_new_n6612__ & new_new_n6987__;
  assign new_new_n6989__ = new_new_n6612__ & ~new_new_n6987__;
  assign new_new_n6990__ = ~new_new_n6988__ & ~new_new_n6989__;
  assign new_new_n6991__ = pi084 & ~new_new_n6990__;
  assign new_new_n6992__ = ~pi084 & new_new_n6990__;
  assign new_new_n6993__ = ~new_new_n6622__ & ~new_new_n6623__;
  assign new_new_n6994__ = ~new_new_n6828__ & po030;
  assign new_new_n6995__ = pi082 & ~po030;
  assign new_new_n6996__ = ~new_new_n6994__ & ~new_new_n6995__;
  assign new_new_n6997__ = new_new_n6993__ & ~new_new_n6996__;
  assign new_new_n6998__ = ~new_new_n6993__ & new_new_n6996__;
  assign new_new_n6999__ = ~new_new_n6997__ & ~new_new_n6998__;
  assign new_new_n7000__ = ~pi083 & ~new_new_n6999__;
  assign new_new_n7001__ = pi083 & new_new_n6999__;
  assign new_new_n7002__ = ~new_new_n6631__ & ~new_new_n6632__;
  assign new_new_n7003__ = ~new_new_n6826__ & po030;
  assign new_new_n7004__ = pi081 & ~po030;
  assign new_new_n7005__ = ~new_new_n7003__ & ~new_new_n7004__;
  assign new_new_n7006__ = new_new_n7002__ & ~new_new_n7005__;
  assign new_new_n7007__ = ~new_new_n7002__ & new_new_n7005__;
  assign new_new_n7008__ = ~new_new_n7006__ & ~new_new_n7007__;
  assign new_new_n7009__ = ~pi082 & ~new_new_n7008__;
  assign new_new_n7010__ = pi082 & new_new_n7008__;
  assign new_new_n7011__ = ~new_new_n6824__ & po030;
  assign new_new_n7012__ = pi080 & ~po030;
  assign new_new_n7013__ = ~new_new_n7011__ & ~new_new_n7012__;
  assign new_new_n7014__ = ~new_new_n6640__ & ~new_new_n6641__;
  assign new_new_n7015__ = ~new_new_n7013__ & new_new_n7014__;
  assign new_new_n7016__ = new_new_n7013__ & ~new_new_n7014__;
  assign new_new_n7017__ = ~new_new_n7015__ & ~new_new_n7016__;
  assign new_new_n7018__ = ~pi081 & ~new_new_n7017__;
  assign new_new_n7019__ = pi081 & new_new_n7017__;
  assign new_new_n7020__ = ~new_new_n6822__ & po030;
  assign new_new_n7021__ = pi079 & ~po030;
  assign new_new_n7022__ = ~new_new_n7020__ & ~new_new_n7021__;
  assign new_new_n7023__ = ~new_new_n6649__ & ~new_new_n6650__;
  assign new_new_n7024__ = ~new_new_n7022__ & new_new_n7023__;
  assign new_new_n7025__ = new_new_n7022__ & ~new_new_n7023__;
  assign new_new_n7026__ = ~new_new_n7024__ & ~new_new_n7025__;
  assign new_new_n7027__ = pi080 & new_new_n7026__;
  assign new_new_n7028__ = ~pi080 & ~new_new_n7026__;
  assign new_new_n7029__ = pi078 & ~new_new_n6820__;
  assign new_new_n7030__ = ~pi078 & new_new_n6820__;
  assign new_new_n7031__ = ~new_new_n7029__ & ~new_new_n7030__;
  assign new_new_n7032__ = po030 & new_new_n7031__;
  assign new_new_n7033__ = new_new_n6657__ & new_new_n7032__;
  assign new_new_n7034__ = ~new_new_n6657__ & ~new_new_n7032__;
  assign new_new_n7035__ = ~new_new_n7033__ & ~new_new_n7034__;
  assign new_new_n7036__ = pi079 & ~new_new_n7035__;
  assign new_new_n7037__ = ~pi079 & new_new_n7035__;
  assign new_new_n7038__ = ~new_new_n6818__ & po030;
  assign new_new_n7039__ = pi077 & ~po030;
  assign new_new_n7040__ = ~new_new_n7038__ & ~new_new_n7039__;
  assign new_new_n7041__ = ~new_new_n6667__ & ~new_new_n6668__;
  assign new_new_n7042__ = ~new_new_n7040__ & new_new_n7041__;
  assign new_new_n7043__ = new_new_n7040__ & ~new_new_n7041__;
  assign new_new_n7044__ = ~new_new_n7042__ & ~new_new_n7043__;
  assign new_new_n7045__ = ~pi078 & ~new_new_n7044__;
  assign new_new_n7046__ = pi078 & new_new_n7044__;
  assign new_new_n7047__ = ~new_new_n6676__ & ~new_new_n6677__;
  assign new_new_n7048__ = ~new_new_n6816__ & po030;
  assign new_new_n7049__ = ~pi076 & ~po030;
  assign new_new_n7050__ = ~new_new_n7048__ & ~new_new_n7049__;
  assign new_new_n7051__ = new_new_n7047__ & ~new_new_n7050__;
  assign new_new_n7052__ = ~new_new_n7047__ & new_new_n7050__;
  assign new_new_n7053__ = ~new_new_n7051__ & ~new_new_n7052__;
  assign new_new_n7054__ = pi077 & ~new_new_n7053__;
  assign new_new_n7055__ = ~pi077 & new_new_n7053__;
  assign new_new_n7056__ = ~pi075 & ~new_new_n6814__;
  assign new_new_n7057__ = pi075 & new_new_n6814__;
  assign new_new_n7058__ = ~new_new_n7056__ & ~new_new_n7057__;
  assign new_new_n7059__ = po030 & new_new_n7058__;
  assign new_new_n7060__ = new_new_n6684__ & ~new_new_n7059__;
  assign new_new_n7061__ = ~new_new_n6684__ & new_new_n7059__;
  assign new_new_n7062__ = ~new_new_n7060__ & ~new_new_n7061__;
  assign new_new_n7063__ = pi076 & ~new_new_n7062__;
  assign new_new_n7064__ = ~pi076 & new_new_n7062__;
  assign new_new_n7065__ = ~new_new_n6812__ & po030;
  assign new_new_n7066__ = pi074 & ~po030;
  assign new_new_n7067__ = ~new_new_n7065__ & ~new_new_n7066__;
  assign new_new_n7068__ = ~new_new_n6694__ & ~new_new_n6695__;
  assign new_new_n7069__ = ~new_new_n7067__ & new_new_n7068__;
  assign new_new_n7070__ = new_new_n7067__ & ~new_new_n7068__;
  assign new_new_n7071__ = ~new_new_n7069__ & ~new_new_n7070__;
  assign new_new_n7072__ = pi075 & new_new_n7071__;
  assign new_new_n7073__ = ~pi075 & ~new_new_n7071__;
  assign new_new_n7074__ = pi073 & ~new_new_n6810__;
  assign new_new_n7075__ = ~pi073 & new_new_n6810__;
  assign new_new_n7076__ = ~new_new_n7074__ & ~new_new_n7075__;
  assign new_new_n7077__ = po030 & new_new_n7076__;
  assign new_new_n7078__ = new_new_n6702__ & new_new_n7077__;
  assign new_new_n7079__ = ~new_new_n6702__ & ~new_new_n7077__;
  assign new_new_n7080__ = ~new_new_n7078__ & ~new_new_n7079__;
  assign new_new_n7081__ = pi074 & ~new_new_n7080__;
  assign new_new_n7082__ = ~pi074 & new_new_n7080__;
  assign new_new_n7083__ = pi072 & ~new_new_n6808__;
  assign new_new_n7084__ = ~pi072 & new_new_n6808__;
  assign new_new_n7085__ = ~new_new_n7083__ & ~new_new_n7084__;
  assign new_new_n7086__ = po030 & new_new_n7085__;
  assign new_new_n7087__ = new_new_n6711__ & new_new_n7086__;
  assign new_new_n7088__ = ~new_new_n6711__ & ~new_new_n7086__;
  assign new_new_n7089__ = ~new_new_n7087__ & ~new_new_n7088__;
  assign new_new_n7090__ = pi073 & ~new_new_n7089__;
  assign new_new_n7091__ = ~pi073 & new_new_n7089__;
  assign new_new_n7092__ = ~new_new_n6721__ & ~new_new_n6722__;
  assign new_new_n7093__ = ~new_new_n6806__ & po030;
  assign new_new_n7094__ = pi071 & ~po030;
  assign new_new_n7095__ = ~new_new_n7093__ & ~new_new_n7094__;
  assign new_new_n7096__ = new_new_n7092__ & ~new_new_n7095__;
  assign new_new_n7097__ = ~new_new_n7092__ & new_new_n7095__;
  assign new_new_n7098__ = ~new_new_n7096__ & ~new_new_n7097__;
  assign new_new_n7099__ = pi072 & new_new_n7098__;
  assign new_new_n7100__ = ~pi072 & ~new_new_n7098__;
  assign new_new_n7101__ = ~new_new_n6730__ & ~new_new_n6731__;
  assign new_new_n7102__ = ~new_new_n6804__ & po030;
  assign new_new_n7103__ = ~pi070 & ~po030;
  assign new_new_n7104__ = ~new_new_n7102__ & ~new_new_n7103__;
  assign new_new_n7105__ = new_new_n7101__ & ~new_new_n7104__;
  assign new_new_n7106__ = ~new_new_n7101__ & new_new_n7104__;
  assign new_new_n7107__ = ~new_new_n7105__ & ~new_new_n7106__;
  assign new_new_n7108__ = pi071 & ~new_new_n7107__;
  assign new_new_n7109__ = ~pi071 & new_new_n7107__;
  assign new_new_n7110__ = ~new_new_n6739__ & ~new_new_n6740__;
  assign new_new_n7111__ = new_new_n6802__ & po030;
  assign new_new_n7112__ = ~pi069 & ~po030;
  assign new_new_n7113__ = ~new_new_n7111__ & ~new_new_n7112__;
  assign new_new_n7114__ = ~new_new_n7110__ & ~new_new_n7113__;
  assign new_new_n7115__ = new_new_n7110__ & new_new_n7113__;
  assign new_new_n7116__ = ~new_new_n7114__ & ~new_new_n7115__;
  assign new_new_n7117__ = ~pi070 & ~new_new_n7116__;
  assign new_new_n7118__ = pi070 & new_new_n7116__;
  assign new_new_n7119__ = new_new_n6800__ & po030;
  assign new_new_n7120__ = ~pi068 & ~po030;
  assign new_new_n7121__ = ~new_new_n7119__ & ~new_new_n7120__;
  assign new_new_n7122__ = ~new_new_n6748__ & ~new_new_n6749__;
  assign new_new_n7123__ = ~new_new_n7121__ & ~new_new_n7122__;
  assign new_new_n7124__ = new_new_n7121__ & new_new_n7122__;
  assign new_new_n7125__ = ~new_new_n7123__ & ~new_new_n7124__;
  assign new_new_n7126__ = pi069 & new_new_n7125__;
  assign new_new_n7127__ = ~pi069 & ~new_new_n7125__;
  assign new_new_n7128__ = ~new_new_n6769__ & ~new_new_n6770__;
  assign new_new_n7129__ = po030 & new_new_n7128__;
  assign new_new_n7130__ = new_new_n6796__ & ~new_new_n7129__;
  assign new_new_n7131__ = ~new_new_n6796__ & new_new_n7129__;
  assign new_new_n7132__ = ~new_new_n7130__ & ~new_new_n7131__;
  assign new_new_n7133__ = pi067 & ~new_new_n7132__;
  assign new_new_n7134__ = ~pi067 & new_new_n7132__;
  assign new_new_n7135__ = pi030 & po030;
  assign new_new_n7136__ = pi029 & ~pi065;
  assign new_new_n7137__ = new_new_n7135__ & ~new_new_n7136__;
  assign new_new_n7138__ = ~pi030 & ~po030;
  assign new_new_n7139__ = ~pi065 & ~new_new_n7138__;
  assign new_new_n7140__ = ~pi029 & ~new_new_n7139__;
  assign new_new_n7141__ = ~new_new_n7137__ & ~new_new_n7140__;
  assign new_new_n7142__ = pi064 & ~new_new_n7141__;
  assign new_new_n7143__ = pi064 & po030;
  assign new_new_n7144__ = ~pi030 & pi065;
  assign new_new_n7145__ = ~new_new_n7143__ & new_new_n7144__;
  assign new_new_n7146__ = ~new_new_n7142__ & ~new_new_n7145__;
  assign new_new_n7147__ = pi066 & ~new_new_n7146__;
  assign new_new_n7148__ = new_new_n426__ & ~po031;
  assign new_new_n7149__ = new_new_n6789__ & po030;
  assign new_new_n7150__ = ~new_new_n7148__ & ~new_new_n7149__;
  assign new_new_n7151__ = ~pi030 & ~new_new_n7150__;
  assign new_new_n7152__ = ~new_new_n332__ & po030;
  assign new_new_n7153__ = ~new_new_n6765__ & ~new_new_n7152__;
  assign new_new_n7154__ = pi065 & po030;
  assign new_new_n7155__ = po031 & ~new_new_n7154__;
  assign new_new_n7156__ = pi065 & ~new_new_n6765__;
  assign new_new_n7157__ = pi030 & ~new_new_n7156__;
  assign new_new_n7158__ = ~new_new_n7155__ & new_new_n7157__;
  assign new_new_n7159__ = ~new_new_n7151__ & ~new_new_n7153__;
  assign new_new_n7160__ = ~new_new_n7158__ & new_new_n7159__;
  assign new_new_n7161__ = ~pi031 & ~new_new_n7160__;
  assign new_new_n7162__ = ~new_new_n6765__ & ~new_new_n7154__;
  assign new_new_n7163__ = pi030 & ~new_new_n6777__;
  assign new_new_n7164__ = pi064 & ~new_new_n7163__;
  assign new_new_n7165__ = ~new_new_n7162__ & ~new_new_n7164__;
  assign new_new_n7166__ = ~pi065 & po030;
  assign new_new_n7167__ = ~po031 & ~new_new_n7166__;
  assign new_new_n7168__ = pi064 & ~new_new_n7135__;
  assign new_new_n7169__ = ~new_new_n7149__ & new_new_n7168__;
  assign new_new_n7170__ = ~new_new_n7167__ & new_new_n7169__;
  assign new_new_n7171__ = ~new_new_n7165__ & ~new_new_n7170__;
  assign new_new_n7172__ = pi031 & ~new_new_n7171__;
  assign new_new_n7173__ = ~new_new_n7161__ & ~new_new_n7172__;
  assign new_new_n7174__ = ~pi066 & new_new_n7146__;
  assign new_new_n7175__ = ~new_new_n7173__ & ~new_new_n7174__;
  assign new_new_n7176__ = ~new_new_n7147__ & ~new_new_n7175__;
  assign new_new_n7177__ = ~new_new_n7134__ & ~new_new_n7176__;
  assign new_new_n7178__ = ~new_new_n7133__ & ~new_new_n7177__;
  assign new_new_n7179__ = pi068 & ~new_new_n7178__;
  assign new_new_n7180__ = ~pi068 & new_new_n7178__;
  assign new_new_n7181__ = ~new_new_n6755__ & ~new_new_n6756__;
  assign new_new_n7182__ = ~new_new_n6798__ & po030;
  assign new_new_n7183__ = pi067 & ~po030;
  assign new_new_n7184__ = ~new_new_n7182__ & ~new_new_n7183__;
  assign new_new_n7185__ = new_new_n7181__ & ~new_new_n7184__;
  assign new_new_n7186__ = ~new_new_n7181__ & new_new_n7184__;
  assign new_new_n7187__ = ~new_new_n7185__ & ~new_new_n7186__;
  assign new_new_n7188__ = ~new_new_n7180__ & new_new_n7187__;
  assign new_new_n7189__ = ~new_new_n7179__ & ~new_new_n7188__;
  assign new_new_n7190__ = ~new_new_n7127__ & ~new_new_n7189__;
  assign new_new_n7191__ = ~new_new_n7126__ & ~new_new_n7190__;
  assign new_new_n7192__ = ~new_new_n7118__ & new_new_n7191__;
  assign new_new_n7193__ = ~new_new_n7117__ & ~new_new_n7192__;
  assign new_new_n7194__ = ~new_new_n7109__ & new_new_n7193__;
  assign new_new_n7195__ = ~new_new_n7108__ & ~new_new_n7194__;
  assign new_new_n7196__ = ~new_new_n7100__ & ~new_new_n7195__;
  assign new_new_n7197__ = ~new_new_n7099__ & ~new_new_n7196__;
  assign new_new_n7198__ = ~new_new_n7091__ & ~new_new_n7197__;
  assign new_new_n7199__ = ~new_new_n7090__ & ~new_new_n7198__;
  assign new_new_n7200__ = ~new_new_n7082__ & ~new_new_n7199__;
  assign new_new_n7201__ = ~new_new_n7081__ & ~new_new_n7200__;
  assign new_new_n7202__ = ~new_new_n7073__ & ~new_new_n7201__;
  assign new_new_n7203__ = ~new_new_n7072__ & ~new_new_n7202__;
  assign new_new_n7204__ = ~new_new_n7064__ & ~new_new_n7203__;
  assign new_new_n7205__ = ~new_new_n7063__ & ~new_new_n7204__;
  assign new_new_n7206__ = ~new_new_n7055__ & ~new_new_n7205__;
  assign new_new_n7207__ = ~new_new_n7054__ & ~new_new_n7206__;
  assign new_new_n7208__ = ~new_new_n7046__ & new_new_n7207__;
  assign new_new_n7209__ = ~new_new_n7045__ & ~new_new_n7208__;
  assign new_new_n7210__ = ~new_new_n7037__ & new_new_n7209__;
  assign new_new_n7211__ = ~new_new_n7036__ & ~new_new_n7210__;
  assign new_new_n7212__ = ~new_new_n7028__ & ~new_new_n7211__;
  assign new_new_n7213__ = ~new_new_n7027__ & ~new_new_n7212__;
  assign new_new_n7214__ = ~new_new_n7019__ & new_new_n7213__;
  assign new_new_n7215__ = ~new_new_n7018__ & ~new_new_n7214__;
  assign new_new_n7216__ = ~new_new_n7010__ & ~new_new_n7215__;
  assign new_new_n7217__ = ~new_new_n7009__ & ~new_new_n7216__;
  assign new_new_n7218__ = ~new_new_n7001__ & ~new_new_n7217__;
  assign new_new_n7219__ = ~new_new_n7000__ & ~new_new_n7218__;
  assign new_new_n7220__ = ~new_new_n6992__ & new_new_n7219__;
  assign new_new_n7221__ = ~new_new_n6991__ & ~new_new_n7220__;
  assign new_new_n7222__ = ~new_new_n6983__ & ~new_new_n7221__;
  assign new_new_n7223__ = ~new_new_n6982__ & ~new_new_n7222__;
  assign new_new_n7224__ = ~new_new_n6974__ & ~new_new_n7223__;
  assign new_new_n7225__ = ~new_new_n6973__ & ~new_new_n7224__;
  assign new_new_n7226__ = ~new_new_n6965__ & ~new_new_n7225__;
  assign new_new_n7227__ = ~new_new_n6964__ & ~new_new_n7226__;
  assign new_new_n7228__ = ~new_new_n6956__ & ~new_new_n7227__;
  assign new_new_n7229__ = ~new_new_n6955__ & ~new_new_n7228__;
  assign new_new_n7230__ = ~new_new_n6947__ & ~new_new_n7229__;
  assign new_new_n7231__ = ~new_new_n6946__ & ~new_new_n7230__;
  assign new_new_n7232__ = ~new_new_n6938__ & ~new_new_n7231__;
  assign new_new_n7233__ = ~new_new_n6937__ & ~new_new_n7232__;
  assign new_new_n7234__ = ~new_new_n6929__ & ~new_new_n7233__;
  assign new_new_n7235__ = ~new_new_n6928__ & ~new_new_n7234__;
  assign new_new_n7236__ = ~new_new_n6920__ & new_new_n7235__;
  assign new_new_n7237__ = ~new_new_n6919__ & ~new_new_n7236__;
  assign new_new_n7238__ = ~new_new_n6911__ & new_new_n7237__;
  assign new_new_n7239__ = ~new_new_n6910__ & ~new_new_n7238__;
  assign new_new_n7240__ = ~new_new_n6902__ & new_new_n7239__;
  assign new_new_n7241__ = ~new_new_n6901__ & ~new_new_n7240__;
  assign new_new_n7242__ = ~new_new_n6893__ & ~new_new_n7241__;
  assign new_new_n7243__ = ~new_new_n6892__ & ~new_new_n7242__;
  assign new_new_n7244__ = ~new_new_n6884__ & ~new_new_n7243__;
  assign new_new_n7245__ = ~new_new_n6883__ & ~new_new_n7244__;
  assign new_new_n7246__ = ~new_new_n6875__ & ~new_new_n7245__;
  assign new_new_n7247__ = ~new_new_n6874__ & ~new_new_n7246__;
  assign new_new_n7248__ = pi098 & new_new_n7247__;
  assign new_new_n7249__ = new_new_n287__ & ~new_new_n7248__;
  assign new_new_n7250__ = new_new_n6859__ & new_new_n6865__;
  assign new_new_n7251__ = pi098 & ~new_new_n6859__;
  assign new_new_n7252__ = ~new_new_n7247__ & ~new_new_n7251__;
  assign new_new_n7253__ = ~new_new_n376__ & ~new_new_n7250__;
  assign new_new_n7254__ = ~new_new_n7252__ & new_new_n7253__;
  assign po029 = new_new_n7249__ & ~new_new_n7254__;
  assign new_new_n7256__ = ~pi097 & ~new_new_n7245__;
  assign new_new_n7257__ = pi097 & new_new_n7245__;
  assign new_new_n7258__ = ~new_new_n7256__ & ~new_new_n7257__;
  assign new_new_n7259__ = po029 & new_new_n7258__;
  assign new_new_n7260__ = ~new_new_n6873__ & ~new_new_n7259__;
  assign new_new_n7261__ = new_new_n6873__ & new_new_n7259__;
  assign new_new_n7262__ = ~new_new_n7260__ & ~new_new_n7261__;
  assign new_new_n7263__ = ~pi098 & ~new_new_n7262__;
  assign new_new_n7264__ = pi098 & new_new_n7262__;
  assign new_new_n7265__ = ~pi096 & ~new_new_n7243__;
  assign new_new_n7266__ = pi096 & new_new_n7243__;
  assign new_new_n7267__ = ~new_new_n7265__ & ~new_new_n7266__;
  assign new_new_n7268__ = po029 & new_new_n7267__;
  assign new_new_n7269__ = new_new_n6882__ & new_new_n7268__;
  assign new_new_n7270__ = ~new_new_n6882__ & ~new_new_n7268__;
  assign new_new_n7271__ = ~new_new_n7269__ & ~new_new_n7270__;
  assign new_new_n7272__ = ~pi097 & ~new_new_n7271__;
  assign new_new_n7273__ = pi097 & new_new_n7271__;
  assign new_new_n7274__ = ~new_new_n6892__ & ~new_new_n6893__;
  assign new_new_n7275__ = ~new_new_n7241__ & po029;
  assign new_new_n7276__ = ~pi095 & ~po029;
  assign new_new_n7277__ = ~new_new_n7275__ & ~new_new_n7276__;
  assign new_new_n7278__ = new_new_n7274__ & ~new_new_n7277__;
  assign new_new_n7279__ = ~new_new_n7274__ & new_new_n7277__;
  assign new_new_n7280__ = ~new_new_n7278__ & ~new_new_n7279__;
  assign new_new_n7281__ = ~pi096 & new_new_n7280__;
  assign new_new_n7282__ = pi096 & ~new_new_n7280__;
  assign new_new_n7283__ = ~new_new_n6901__ & ~new_new_n6902__;
  assign new_new_n7284__ = pi094 & ~po029;
  assign new_new_n7285__ = ~new_new_n7239__ & po029;
  assign new_new_n7286__ = ~new_new_n7284__ & ~new_new_n7285__;
  assign new_new_n7287__ = new_new_n7283__ & ~new_new_n7286__;
  assign new_new_n7288__ = ~new_new_n7283__ & new_new_n7286__;
  assign new_new_n7289__ = ~new_new_n7287__ & ~new_new_n7288__;
  assign new_new_n7290__ = ~pi095 & ~new_new_n7289__;
  assign new_new_n7291__ = pi095 & new_new_n7289__;
  assign new_new_n7292__ = ~new_new_n6910__ & ~new_new_n6911__;
  assign new_new_n7293__ = ~new_new_n7237__ & po029;
  assign new_new_n7294__ = ~pi093 & ~po029;
  assign new_new_n7295__ = ~new_new_n7293__ & ~new_new_n7294__;
  assign new_new_n7296__ = new_new_n7292__ & ~new_new_n7295__;
  assign new_new_n7297__ = ~new_new_n7292__ & new_new_n7295__;
  assign new_new_n7298__ = ~new_new_n7296__ & ~new_new_n7297__;
  assign new_new_n7299__ = pi094 & ~new_new_n7298__;
  assign new_new_n7300__ = ~pi094 & new_new_n7298__;
  assign new_new_n7301__ = ~new_new_n7235__ & po029;
  assign new_new_n7302__ = pi092 & ~po029;
  assign new_new_n7303__ = ~new_new_n7301__ & ~new_new_n7302__;
  assign new_new_n7304__ = ~new_new_n6919__ & ~new_new_n6920__;
  assign new_new_n7305__ = ~new_new_n7303__ & new_new_n7304__;
  assign new_new_n7306__ = new_new_n7303__ & ~new_new_n7304__;
  assign new_new_n7307__ = ~new_new_n7305__ & ~new_new_n7306__;
  assign new_new_n7308__ = ~pi093 & ~new_new_n7307__;
  assign new_new_n7309__ = pi093 & new_new_n7307__;
  assign new_new_n7310__ = ~new_new_n6928__ & ~new_new_n6929__;
  assign new_new_n7311__ = pi091 & ~po029;
  assign new_new_n7312__ = ~new_new_n7233__ & po029;
  assign new_new_n7313__ = ~new_new_n7311__ & ~new_new_n7312__;
  assign new_new_n7314__ = new_new_n7310__ & new_new_n7313__;
  assign new_new_n7315__ = ~new_new_n7310__ & ~new_new_n7313__;
  assign new_new_n7316__ = ~new_new_n7314__ & ~new_new_n7315__;
  assign new_new_n7317__ = pi092 & ~new_new_n7316__;
  assign new_new_n7318__ = ~pi092 & new_new_n7316__;
  assign new_new_n7319__ = new_new_n7231__ & po029;
  assign new_new_n7320__ = ~pi090 & ~po029;
  assign new_new_n7321__ = ~new_new_n7319__ & ~new_new_n7320__;
  assign new_new_n7322__ = ~new_new_n6937__ & ~new_new_n6938__;
  assign new_new_n7323__ = ~new_new_n7321__ & ~new_new_n7322__;
  assign new_new_n7324__ = new_new_n7321__ & new_new_n7322__;
  assign new_new_n7325__ = ~new_new_n7323__ & ~new_new_n7324__;
  assign new_new_n7326__ = pi091 & new_new_n7325__;
  assign new_new_n7327__ = ~pi091 & ~new_new_n7325__;
  assign new_new_n7328__ = ~new_new_n6946__ & ~new_new_n6947__;
  assign new_new_n7329__ = pi089 & ~po029;
  assign new_new_n7330__ = ~new_new_n7229__ & po029;
  assign new_new_n7331__ = ~new_new_n7329__ & ~new_new_n7330__;
  assign new_new_n7332__ = new_new_n7328__ & new_new_n7331__;
  assign new_new_n7333__ = ~new_new_n7328__ & ~new_new_n7331__;
  assign new_new_n7334__ = ~new_new_n7332__ & ~new_new_n7333__;
  assign new_new_n7335__ = pi090 & ~new_new_n7334__;
  assign new_new_n7336__ = ~pi090 & new_new_n7334__;
  assign new_new_n7337__ = new_new_n7227__ & po029;
  assign new_new_n7338__ = ~pi088 & ~po029;
  assign new_new_n7339__ = ~new_new_n7337__ & ~new_new_n7338__;
  assign new_new_n7340__ = ~new_new_n6955__ & ~new_new_n6956__;
  assign new_new_n7341__ = ~new_new_n7339__ & ~new_new_n7340__;
  assign new_new_n7342__ = new_new_n7339__ & new_new_n7340__;
  assign new_new_n7343__ = ~new_new_n7341__ & ~new_new_n7342__;
  assign new_new_n7344__ = pi089 & new_new_n7343__;
  assign new_new_n7345__ = ~pi089 & ~new_new_n7343__;
  assign new_new_n7346__ = new_new_n7225__ & po029;
  assign new_new_n7347__ = ~pi087 & ~po029;
  assign new_new_n7348__ = ~new_new_n7346__ & ~new_new_n7347__;
  assign new_new_n7349__ = ~new_new_n6964__ & ~new_new_n6965__;
  assign new_new_n7350__ = ~new_new_n7348__ & ~new_new_n7349__;
  assign new_new_n7351__ = new_new_n7348__ & new_new_n7349__;
  assign new_new_n7352__ = ~new_new_n7350__ & ~new_new_n7351__;
  assign new_new_n7353__ = pi088 & new_new_n7352__;
  assign new_new_n7354__ = ~pi088 & ~new_new_n7352__;
  assign new_new_n7355__ = new_new_n7223__ & po029;
  assign new_new_n7356__ = ~pi086 & ~po029;
  assign new_new_n7357__ = ~new_new_n7355__ & ~new_new_n7356__;
  assign new_new_n7358__ = ~new_new_n6973__ & ~new_new_n6974__;
  assign new_new_n7359__ = ~new_new_n7357__ & ~new_new_n7358__;
  assign new_new_n7360__ = new_new_n7357__ & new_new_n7358__;
  assign new_new_n7361__ = ~new_new_n7359__ & ~new_new_n7360__;
  assign new_new_n7362__ = pi087 & new_new_n7361__;
  assign new_new_n7363__ = ~pi087 & ~new_new_n7361__;
  assign new_new_n7364__ = ~new_new_n6982__ & ~new_new_n6983__;
  assign new_new_n7365__ = pi085 & ~po029;
  assign new_new_n7366__ = ~new_new_n7221__ & po029;
  assign new_new_n7367__ = ~new_new_n7365__ & ~new_new_n7366__;
  assign new_new_n7368__ = new_new_n7364__ & new_new_n7367__;
  assign new_new_n7369__ = ~new_new_n7364__ & ~new_new_n7367__;
  assign new_new_n7370__ = ~new_new_n7368__ & ~new_new_n7369__;
  assign new_new_n7371__ = pi086 & ~new_new_n7370__;
  assign new_new_n7372__ = ~pi086 & new_new_n7370__;
  assign new_new_n7373__ = new_new_n7219__ & po029;
  assign new_new_n7374__ = pi084 & ~po029;
  assign new_new_n7375__ = ~new_new_n7373__ & ~new_new_n7374__;
  assign new_new_n7376__ = ~new_new_n6991__ & ~new_new_n6992__;
  assign new_new_n7377__ = ~new_new_n7375__ & ~new_new_n7376__;
  assign new_new_n7378__ = new_new_n7375__ & new_new_n7376__;
  assign new_new_n7379__ = ~new_new_n7377__ & ~new_new_n7378__;
  assign new_new_n7380__ = pi085 & ~new_new_n7379__;
  assign new_new_n7381__ = ~pi085 & new_new_n7379__;
  assign new_new_n7382__ = ~pi083 & ~new_new_n7217__;
  assign new_new_n7383__ = pi083 & new_new_n7217__;
  assign new_new_n7384__ = ~new_new_n7382__ & ~new_new_n7383__;
  assign new_new_n7385__ = po029 & new_new_n7384__;
  assign new_new_n7386__ = new_new_n6999__ & new_new_n7385__;
  assign new_new_n7387__ = ~new_new_n6999__ & ~new_new_n7385__;
  assign new_new_n7388__ = ~new_new_n7386__ & ~new_new_n7387__;
  assign new_new_n7389__ = pi084 & new_new_n7388__;
  assign new_new_n7390__ = ~pi084 & ~new_new_n7388__;
  assign new_new_n7391__ = ~pi082 & ~new_new_n7215__;
  assign new_new_n7392__ = pi082 & new_new_n7215__;
  assign new_new_n7393__ = ~new_new_n7391__ & ~new_new_n7392__;
  assign new_new_n7394__ = po029 & new_new_n7393__;
  assign new_new_n7395__ = new_new_n7008__ & new_new_n7394__;
  assign new_new_n7396__ = ~new_new_n7008__ & ~new_new_n7394__;
  assign new_new_n7397__ = ~new_new_n7395__ & ~new_new_n7396__;
  assign new_new_n7398__ = pi083 & new_new_n7397__;
  assign new_new_n7399__ = ~pi083 & ~new_new_n7397__;
  assign new_new_n7400__ = ~new_new_n7018__ & ~new_new_n7019__;
  assign new_new_n7401__ = new_new_n7213__ & po029;
  assign new_new_n7402__ = ~pi081 & ~po029;
  assign new_new_n7403__ = ~new_new_n7401__ & ~new_new_n7402__;
  assign new_new_n7404__ = ~new_new_n7400__ & ~new_new_n7403__;
  assign new_new_n7405__ = new_new_n7400__ & new_new_n7403__;
  assign new_new_n7406__ = ~new_new_n7404__ & ~new_new_n7405__;
  assign new_new_n7407__ = pi082 & new_new_n7406__;
  assign new_new_n7408__ = ~pi082 & ~new_new_n7406__;
  assign new_new_n7409__ = new_new_n7211__ & po029;
  assign new_new_n7410__ = ~pi080 & ~po029;
  assign new_new_n7411__ = ~new_new_n7409__ & ~new_new_n7410__;
  assign new_new_n7412__ = ~new_new_n7027__ & ~new_new_n7028__;
  assign new_new_n7413__ = ~new_new_n7411__ & ~new_new_n7412__;
  assign new_new_n7414__ = new_new_n7411__ & new_new_n7412__;
  assign new_new_n7415__ = ~new_new_n7413__ & ~new_new_n7414__;
  assign new_new_n7416__ = pi081 & new_new_n7415__;
  assign new_new_n7417__ = ~pi081 & ~new_new_n7415__;
  assign new_new_n7418__ = new_new_n7209__ & po029;
  assign new_new_n7419__ = pi079 & ~po029;
  assign new_new_n7420__ = ~new_new_n7418__ & ~new_new_n7419__;
  assign new_new_n7421__ = ~new_new_n7036__ & ~new_new_n7037__;
  assign new_new_n7422__ = ~new_new_n7420__ & ~new_new_n7421__;
  assign new_new_n7423__ = new_new_n7420__ & new_new_n7421__;
  assign new_new_n7424__ = ~new_new_n7422__ & ~new_new_n7423__;
  assign new_new_n7425__ = pi080 & ~new_new_n7424__;
  assign new_new_n7426__ = ~pi080 & new_new_n7424__;
  assign new_new_n7427__ = ~new_new_n7207__ & po029;
  assign new_new_n7428__ = pi078 & ~po029;
  assign new_new_n7429__ = ~new_new_n7427__ & ~new_new_n7428__;
  assign new_new_n7430__ = ~new_new_n7045__ & ~new_new_n7046__;
  assign new_new_n7431__ = new_new_n7429__ & new_new_n7430__;
  assign new_new_n7432__ = ~new_new_n7429__ & ~new_new_n7430__;
  assign new_new_n7433__ = ~new_new_n7431__ & ~new_new_n7432__;
  assign new_new_n7434__ = pi079 & ~new_new_n7433__;
  assign new_new_n7435__ = ~pi079 & new_new_n7433__;
  assign new_new_n7436__ = ~new_new_n7054__ & ~new_new_n7055__;
  assign new_new_n7437__ = pi077 & ~po029;
  assign new_new_n7438__ = ~new_new_n7205__ & po029;
  assign new_new_n7439__ = ~new_new_n7437__ & ~new_new_n7438__;
  assign new_new_n7440__ = new_new_n7436__ & new_new_n7439__;
  assign new_new_n7441__ = ~new_new_n7436__ & ~new_new_n7439__;
  assign new_new_n7442__ = ~new_new_n7440__ & ~new_new_n7441__;
  assign new_new_n7443__ = pi078 & ~new_new_n7442__;
  assign new_new_n7444__ = ~pi078 & new_new_n7442__;
  assign new_new_n7445__ = pi076 & ~new_new_n7203__;
  assign new_new_n7446__ = ~pi076 & new_new_n7203__;
  assign new_new_n7447__ = ~new_new_n7445__ & ~new_new_n7446__;
  assign new_new_n7448__ = po029 & new_new_n7447__;
  assign new_new_n7449__ = new_new_n7062__ & new_new_n7448__;
  assign new_new_n7450__ = ~new_new_n7062__ & ~new_new_n7448__;
  assign new_new_n7451__ = ~new_new_n7449__ & ~new_new_n7450__;
  assign new_new_n7452__ = pi077 & ~new_new_n7451__;
  assign new_new_n7453__ = ~pi077 & new_new_n7451__;
  assign new_new_n7454__ = new_new_n7201__ & po029;
  assign new_new_n7455__ = ~pi075 & ~po029;
  assign new_new_n7456__ = ~new_new_n7454__ & ~new_new_n7455__;
  assign new_new_n7457__ = ~new_new_n7072__ & ~new_new_n7073__;
  assign new_new_n7458__ = ~new_new_n7456__ & ~new_new_n7457__;
  assign new_new_n7459__ = new_new_n7456__ & new_new_n7457__;
  assign new_new_n7460__ = ~new_new_n7458__ & ~new_new_n7459__;
  assign new_new_n7461__ = ~pi076 & ~new_new_n7460__;
  assign new_new_n7462__ = pi076 & new_new_n7460__;
  assign new_new_n7463__ = ~new_new_n7081__ & ~new_new_n7082__;
  assign new_new_n7464__ = pi074 & ~po029;
  assign new_new_n7465__ = ~new_new_n7199__ & po029;
  assign new_new_n7466__ = ~new_new_n7464__ & ~new_new_n7465__;
  assign new_new_n7467__ = new_new_n7463__ & new_new_n7466__;
  assign new_new_n7468__ = ~new_new_n7463__ & ~new_new_n7466__;
  assign new_new_n7469__ = ~new_new_n7467__ & ~new_new_n7468__;
  assign new_new_n7470__ = ~pi075 & new_new_n7469__;
  assign new_new_n7471__ = pi075 & ~new_new_n7469__;
  assign new_new_n7472__ = ~new_new_n7090__ & ~new_new_n7091__;
  assign new_new_n7473__ = pi073 & ~po029;
  assign new_new_n7474__ = ~new_new_n7197__ & po029;
  assign new_new_n7475__ = ~new_new_n7473__ & ~new_new_n7474__;
  assign new_new_n7476__ = new_new_n7472__ & new_new_n7475__;
  assign new_new_n7477__ = ~new_new_n7472__ & ~new_new_n7475__;
  assign new_new_n7478__ = ~new_new_n7476__ & ~new_new_n7477__;
  assign new_new_n7479__ = ~pi074 & new_new_n7478__;
  assign new_new_n7480__ = pi074 & ~new_new_n7478__;
  assign new_new_n7481__ = new_new_n7195__ & po029;
  assign new_new_n7482__ = ~pi072 & ~po029;
  assign new_new_n7483__ = ~new_new_n7481__ & ~new_new_n7482__;
  assign new_new_n7484__ = ~new_new_n7099__ & ~new_new_n7100__;
  assign new_new_n7485__ = ~new_new_n7483__ & ~new_new_n7484__;
  assign new_new_n7486__ = new_new_n7483__ & new_new_n7484__;
  assign new_new_n7487__ = ~new_new_n7485__ & ~new_new_n7486__;
  assign new_new_n7488__ = ~pi073 & ~new_new_n7487__;
  assign new_new_n7489__ = pi073 & new_new_n7487__;
  assign new_new_n7490__ = new_new_n7193__ & po029;
  assign new_new_n7491__ = pi071 & ~po029;
  assign new_new_n7492__ = ~new_new_n7490__ & ~new_new_n7491__;
  assign new_new_n7493__ = ~new_new_n7108__ & ~new_new_n7109__;
  assign new_new_n7494__ = ~new_new_n7492__ & ~new_new_n7493__;
  assign new_new_n7495__ = new_new_n7492__ & new_new_n7493__;
  assign new_new_n7496__ = ~new_new_n7494__ & ~new_new_n7495__;
  assign new_new_n7497__ = pi072 & ~new_new_n7496__;
  assign new_new_n7498__ = ~pi072 & new_new_n7496__;
  assign new_new_n7499__ = new_new_n7191__ & po029;
  assign new_new_n7500__ = ~pi070 & ~po029;
  assign new_new_n7501__ = ~new_new_n7499__ & ~new_new_n7500__;
  assign new_new_n7502__ = ~new_new_n7117__ & ~new_new_n7118__;
  assign new_new_n7503__ = ~new_new_n7501__ & ~new_new_n7502__;
  assign new_new_n7504__ = new_new_n7501__ & new_new_n7502__;
  assign new_new_n7505__ = ~new_new_n7503__ & ~new_new_n7504__;
  assign new_new_n7506__ = ~pi071 & ~new_new_n7505__;
  assign new_new_n7507__ = pi071 & new_new_n7505__;
  assign new_new_n7508__ = ~new_new_n7126__ & ~new_new_n7127__;
  assign new_new_n7509__ = new_new_n7189__ & po029;
  assign new_new_n7510__ = ~pi069 & ~po029;
  assign new_new_n7511__ = ~new_new_n7509__ & ~new_new_n7510__;
  assign new_new_n7512__ = ~new_new_n7508__ & ~new_new_n7511__;
  assign new_new_n7513__ = new_new_n7508__ & new_new_n7511__;
  assign new_new_n7514__ = ~new_new_n7512__ & ~new_new_n7513__;
  assign new_new_n7515__ = ~pi070 & ~new_new_n7514__;
  assign new_new_n7516__ = pi070 & new_new_n7514__;
  assign new_new_n7517__ = ~new_new_n7179__ & ~new_new_n7180__;
  assign new_new_n7518__ = po029 & new_new_n7517__;
  assign new_new_n7519__ = new_new_n7187__ & new_new_n7518__;
  assign new_new_n7520__ = ~new_new_n7187__ & ~new_new_n7518__;
  assign new_new_n7521__ = ~new_new_n7519__ & ~new_new_n7520__;
  assign new_new_n7522__ = pi069 & new_new_n7521__;
  assign new_new_n7523__ = ~pi069 & ~new_new_n7521__;
  assign new_new_n7524__ = ~pi067 & ~new_new_n7176__;
  assign new_new_n7525__ = pi067 & new_new_n7176__;
  assign new_new_n7526__ = ~new_new_n7524__ & ~new_new_n7525__;
  assign new_new_n7527__ = po029 & ~new_new_n7526__;
  assign new_new_n7528__ = new_new_n7132__ & new_new_n7527__;
  assign new_new_n7529__ = ~new_new_n7132__ & ~new_new_n7527__;
  assign new_new_n7530__ = ~new_new_n7528__ & ~new_new_n7529__;
  assign new_new_n7531__ = pi068 & ~new_new_n7530__;
  assign new_new_n7532__ = ~pi068 & new_new_n7530__;
  assign new_new_n7533__ = pi029 & po029;
  assign new_new_n7534__ = pi028 & ~pi065;
  assign new_new_n7535__ = new_new_n7533__ & ~new_new_n7534__;
  assign new_new_n7536__ = ~pi029 & ~po029;
  assign new_new_n7537__ = ~pi065 & ~new_new_n7536__;
  assign new_new_n7538__ = ~pi028 & ~new_new_n7537__;
  assign new_new_n7539__ = ~new_new_n7535__ & ~new_new_n7538__;
  assign new_new_n7540__ = pi064 & ~new_new_n7539__;
  assign new_new_n7541__ = pi064 & po029;
  assign new_new_n7542__ = ~pi029 & pi065;
  assign new_new_n7543__ = ~new_new_n7541__ & new_new_n7542__;
  assign new_new_n7544__ = ~new_new_n7540__ & ~new_new_n7543__;
  assign new_new_n7545__ = pi066 & ~new_new_n7544__;
  assign new_new_n7546__ = ~pi066 & new_new_n7544__;
  assign new_new_n7547__ = new_new_n426__ & ~po030;
  assign new_new_n7548__ = new_new_n7166__ & po029;
  assign new_new_n7549__ = ~new_new_n7547__ & ~new_new_n7548__;
  assign new_new_n7550__ = ~pi029 & ~new_new_n7549__;
  assign new_new_n7551__ = ~new_new_n332__ & po029;
  assign new_new_n7552__ = ~new_new_n7143__ & ~new_new_n7551__;
  assign new_new_n7553__ = pi065 & po029;
  assign new_new_n7554__ = po030 & ~new_new_n7553__;
  assign new_new_n7555__ = pi065 & ~new_new_n7143__;
  assign new_new_n7556__ = pi029 & ~new_new_n7555__;
  assign new_new_n7557__ = ~new_new_n7554__ & new_new_n7556__;
  assign new_new_n7558__ = ~new_new_n7550__ & ~new_new_n7552__;
  assign new_new_n7559__ = ~new_new_n7557__ & new_new_n7558__;
  assign new_new_n7560__ = pi030 & ~new_new_n7559__;
  assign new_new_n7561__ = ~new_new_n7143__ & ~new_new_n7553__;
  assign new_new_n7562__ = pi029 & ~new_new_n7154__;
  assign new_new_n7563__ = pi064 & ~new_new_n7562__;
  assign new_new_n7564__ = ~new_new_n7561__ & ~new_new_n7563__;
  assign new_new_n7565__ = ~pi065 & po029;
  assign new_new_n7566__ = ~po030 & ~new_new_n7565__;
  assign new_new_n7567__ = pi064 & ~new_new_n7533__;
  assign new_new_n7568__ = ~new_new_n7548__ & new_new_n7567__;
  assign new_new_n7569__ = ~new_new_n7566__ & new_new_n7568__;
  assign new_new_n7570__ = ~new_new_n7564__ & ~new_new_n7569__;
  assign new_new_n7571__ = ~pi030 & ~new_new_n7570__;
  assign new_new_n7572__ = ~new_new_n7560__ & ~new_new_n7571__;
  assign new_new_n7573__ = ~new_new_n7546__ & new_new_n7572__;
  assign new_new_n7574__ = ~new_new_n7545__ & ~new_new_n7573__;
  assign new_new_n7575__ = pi067 & ~new_new_n7574__;
  assign new_new_n7576__ = ~new_new_n7147__ & po029;
  assign new_new_n7577__ = ~new_new_n7174__ & new_new_n7576__;
  assign new_new_n7578__ = new_new_n7173__ & ~new_new_n7577__;
  assign new_new_n7579__ = new_new_n7175__ & new_new_n7576__;
  assign new_new_n7580__ = ~new_new_n7578__ & ~new_new_n7579__;
  assign new_new_n7581__ = ~new_new_n7575__ & ~new_new_n7580__;
  assign new_new_n7582__ = ~pi067 & new_new_n7574__;
  assign new_new_n7583__ = ~new_new_n7581__ & ~new_new_n7582__;
  assign new_new_n7584__ = ~new_new_n7532__ & new_new_n7583__;
  assign new_new_n7585__ = ~new_new_n7531__ & ~new_new_n7584__;
  assign new_new_n7586__ = ~new_new_n7523__ & ~new_new_n7585__;
  assign new_new_n7587__ = ~new_new_n7522__ & ~new_new_n7586__;
  assign new_new_n7588__ = ~new_new_n7516__ & new_new_n7587__;
  assign new_new_n7589__ = ~new_new_n7515__ & ~new_new_n7588__;
  assign new_new_n7590__ = ~new_new_n7507__ & ~new_new_n7589__;
  assign new_new_n7591__ = ~new_new_n7506__ & ~new_new_n7590__;
  assign new_new_n7592__ = ~new_new_n7498__ & new_new_n7591__;
  assign new_new_n7593__ = ~new_new_n7497__ & ~new_new_n7592__;
  assign new_new_n7594__ = ~new_new_n7489__ & new_new_n7593__;
  assign new_new_n7595__ = ~new_new_n7488__ & ~new_new_n7594__;
  assign new_new_n7596__ = ~new_new_n7480__ & ~new_new_n7595__;
  assign new_new_n7597__ = ~new_new_n7479__ & ~new_new_n7596__;
  assign new_new_n7598__ = ~new_new_n7471__ & ~new_new_n7597__;
  assign new_new_n7599__ = ~new_new_n7470__ & ~new_new_n7598__;
  assign new_new_n7600__ = ~new_new_n7462__ & ~new_new_n7599__;
  assign new_new_n7601__ = ~new_new_n7461__ & ~new_new_n7600__;
  assign new_new_n7602__ = ~new_new_n7453__ & new_new_n7601__;
  assign new_new_n7603__ = ~new_new_n7452__ & ~new_new_n7602__;
  assign new_new_n7604__ = ~new_new_n7444__ & ~new_new_n7603__;
  assign new_new_n7605__ = ~new_new_n7443__ & ~new_new_n7604__;
  assign new_new_n7606__ = ~new_new_n7435__ & ~new_new_n7605__;
  assign new_new_n7607__ = ~new_new_n7434__ & ~new_new_n7606__;
  assign new_new_n7608__ = ~new_new_n7426__ & ~new_new_n7607__;
  assign new_new_n7609__ = ~new_new_n7425__ & ~new_new_n7608__;
  assign new_new_n7610__ = ~new_new_n7417__ & ~new_new_n7609__;
  assign new_new_n7611__ = ~new_new_n7416__ & ~new_new_n7610__;
  assign new_new_n7612__ = ~new_new_n7408__ & ~new_new_n7611__;
  assign new_new_n7613__ = ~new_new_n7407__ & ~new_new_n7612__;
  assign new_new_n7614__ = ~new_new_n7399__ & ~new_new_n7613__;
  assign new_new_n7615__ = ~new_new_n7398__ & ~new_new_n7614__;
  assign new_new_n7616__ = ~new_new_n7390__ & ~new_new_n7615__;
  assign new_new_n7617__ = ~new_new_n7389__ & ~new_new_n7616__;
  assign new_new_n7618__ = ~new_new_n7381__ & ~new_new_n7617__;
  assign new_new_n7619__ = ~new_new_n7380__ & ~new_new_n7618__;
  assign new_new_n7620__ = ~new_new_n7372__ & ~new_new_n7619__;
  assign new_new_n7621__ = ~new_new_n7371__ & ~new_new_n7620__;
  assign new_new_n7622__ = ~new_new_n7363__ & ~new_new_n7621__;
  assign new_new_n7623__ = ~new_new_n7362__ & ~new_new_n7622__;
  assign new_new_n7624__ = ~new_new_n7354__ & ~new_new_n7623__;
  assign new_new_n7625__ = ~new_new_n7353__ & ~new_new_n7624__;
  assign new_new_n7626__ = ~new_new_n7345__ & ~new_new_n7625__;
  assign new_new_n7627__ = ~new_new_n7344__ & ~new_new_n7626__;
  assign new_new_n7628__ = ~new_new_n7336__ & ~new_new_n7627__;
  assign new_new_n7629__ = ~new_new_n7335__ & ~new_new_n7628__;
  assign new_new_n7630__ = ~new_new_n7327__ & ~new_new_n7629__;
  assign new_new_n7631__ = ~new_new_n7326__ & ~new_new_n7630__;
  assign new_new_n7632__ = ~new_new_n7318__ & ~new_new_n7631__;
  assign new_new_n7633__ = ~new_new_n7317__ & ~new_new_n7632__;
  assign new_new_n7634__ = ~new_new_n7309__ & new_new_n7633__;
  assign new_new_n7635__ = ~new_new_n7308__ & ~new_new_n7634__;
  assign new_new_n7636__ = ~new_new_n7300__ & new_new_n7635__;
  assign new_new_n7637__ = ~new_new_n7299__ & ~new_new_n7636__;
  assign new_new_n7638__ = ~new_new_n7291__ & new_new_n7637__;
  assign new_new_n7639__ = ~new_new_n7290__ & ~new_new_n7638__;
  assign new_new_n7640__ = ~new_new_n7282__ & ~new_new_n7639__;
  assign new_new_n7641__ = ~new_new_n7281__ & ~new_new_n7640__;
  assign new_new_n7642__ = ~new_new_n7273__ & ~new_new_n7641__;
  assign new_new_n7643__ = ~new_new_n7272__ & ~new_new_n7642__;
  assign new_new_n7644__ = ~new_new_n7264__ & ~new_new_n7643__;
  assign new_new_n7645__ = ~new_new_n7263__ & ~new_new_n7644__;
  assign new_new_n7646__ = pi099 & new_new_n7645__;
  assign new_new_n7647__ = ~pi101 & new_new_n284__;
  assign new_new_n7648__ = ~pi100 & new_new_n7647__;
  assign new_new_n7649__ = ~new_new_n7646__ & new_new_n7648__;
  assign new_new_n7650__ = ~new_new_n376__ & new_new_n7249__;
  assign new_new_n7651__ = ~new_new_n6860__ & ~new_new_n7650__;
  assign new_new_n7652__ = ~new_new_n7649__ & new_new_n7651__;
  assign new_new_n7653__ = ~new_new_n7263__ & ~new_new_n7264__;
  assign new_new_n7654__ = ~pi099 & ~new_new_n7645__;
  assign new_new_n7655__ = ~new_new_n7651__ & ~new_new_n7654__;
  assign po028 = new_new_n7649__ & ~new_new_n7655__;
  assign new_new_n7657__ = ~new_new_n7643__ & po028;
  assign new_new_n7658__ = ~pi098 & ~po028;
  assign new_new_n7659__ = ~new_new_n7657__ & ~new_new_n7658__;
  assign new_new_n7660__ = new_new_n7653__ & ~new_new_n7659__;
  assign new_new_n7661__ = ~new_new_n7653__ & new_new_n7659__;
  assign new_new_n7662__ = ~new_new_n7660__ & ~new_new_n7661__;
  assign new_new_n7663__ = ~new_new_n7281__ & ~new_new_n7282__;
  assign new_new_n7664__ = ~new_new_n7639__ & po028;
  assign new_new_n7665__ = ~pi096 & ~po028;
  assign new_new_n7666__ = ~new_new_n7664__ & ~new_new_n7665__;
  assign new_new_n7667__ = new_new_n7663__ & ~new_new_n7666__;
  assign new_new_n7668__ = ~new_new_n7663__ & new_new_n7666__;
  assign new_new_n7669__ = ~new_new_n7667__ & ~new_new_n7668__;
  assign new_new_n7670__ = pi097 & ~new_new_n7669__;
  assign new_new_n7671__ = ~pi097 & new_new_n7669__;
  assign new_new_n7672__ = ~new_new_n7637__ & po028;
  assign new_new_n7673__ = pi095 & ~po028;
  assign new_new_n7674__ = ~new_new_n7672__ & ~new_new_n7673__;
  assign new_new_n7675__ = ~new_new_n7290__ & ~new_new_n7291__;
  assign new_new_n7676__ = ~new_new_n7674__ & new_new_n7675__;
  assign new_new_n7677__ = new_new_n7674__ & ~new_new_n7675__;
  assign new_new_n7678__ = ~new_new_n7676__ & ~new_new_n7677__;
  assign new_new_n7679__ = pi096 & new_new_n7678__;
  assign new_new_n7680__ = ~pi096 & ~new_new_n7678__;
  assign new_new_n7681__ = ~new_new_n7299__ & ~new_new_n7300__;
  assign new_new_n7682__ = ~new_new_n7635__ & po028;
  assign new_new_n7683__ = ~pi094 & ~po028;
  assign new_new_n7684__ = ~new_new_n7682__ & ~new_new_n7683__;
  assign new_new_n7685__ = new_new_n7681__ & ~new_new_n7684__;
  assign new_new_n7686__ = ~new_new_n7681__ & new_new_n7684__;
  assign new_new_n7687__ = ~new_new_n7685__ & ~new_new_n7686__;
  assign new_new_n7688__ = pi095 & ~new_new_n7687__;
  assign new_new_n7689__ = ~pi095 & new_new_n7687__;
  assign new_new_n7690__ = ~new_new_n7633__ & po028;
  assign new_new_n7691__ = pi093 & ~po028;
  assign new_new_n7692__ = ~new_new_n7690__ & ~new_new_n7691__;
  assign new_new_n7693__ = ~new_new_n7308__ & ~new_new_n7309__;
  assign new_new_n7694__ = ~new_new_n7692__ & new_new_n7693__;
  assign new_new_n7695__ = new_new_n7692__ & ~new_new_n7693__;
  assign new_new_n7696__ = ~new_new_n7694__ & ~new_new_n7695__;
  assign new_new_n7697__ = ~pi094 & ~new_new_n7696__;
  assign new_new_n7698__ = pi094 & new_new_n7696__;
  assign new_new_n7699__ = ~new_new_n7317__ & ~new_new_n7318__;
  assign new_new_n7700__ = ~new_new_n7631__ & po028;
  assign new_new_n7701__ = pi092 & ~po028;
  assign new_new_n7702__ = ~new_new_n7700__ & ~new_new_n7701__;
  assign new_new_n7703__ = new_new_n7699__ & ~new_new_n7702__;
  assign new_new_n7704__ = ~new_new_n7699__ & new_new_n7702__;
  assign new_new_n7705__ = ~new_new_n7703__ & ~new_new_n7704__;
  assign new_new_n7706__ = ~pi093 & ~new_new_n7705__;
  assign new_new_n7707__ = pi093 & new_new_n7705__;
  assign new_new_n7708__ = ~new_new_n7629__ & po028;
  assign new_new_n7709__ = pi091 & ~po028;
  assign new_new_n7710__ = ~new_new_n7708__ & ~new_new_n7709__;
  assign new_new_n7711__ = ~new_new_n7326__ & ~new_new_n7327__;
  assign new_new_n7712__ = ~new_new_n7710__ & new_new_n7711__;
  assign new_new_n7713__ = new_new_n7710__ & ~new_new_n7711__;
  assign new_new_n7714__ = ~new_new_n7712__ & ~new_new_n7713__;
  assign new_new_n7715__ = ~pi092 & ~new_new_n7714__;
  assign new_new_n7716__ = pi092 & new_new_n7714__;
  assign new_new_n7717__ = pi090 & ~new_new_n7627__;
  assign new_new_n7718__ = ~pi090 & new_new_n7627__;
  assign new_new_n7719__ = ~new_new_n7717__ & ~new_new_n7718__;
  assign new_new_n7720__ = po028 & new_new_n7719__;
  assign new_new_n7721__ = new_new_n7334__ & new_new_n7720__;
  assign new_new_n7722__ = ~new_new_n7334__ & ~new_new_n7720__;
  assign new_new_n7723__ = ~new_new_n7721__ & ~new_new_n7722__;
  assign new_new_n7724__ = pi091 & ~new_new_n7723__;
  assign new_new_n7725__ = ~pi091 & new_new_n7723__;
  assign new_new_n7726__ = ~new_new_n7344__ & ~new_new_n7345__;
  assign new_new_n7727__ = ~new_new_n7625__ & po028;
  assign new_new_n7728__ = pi089 & ~po028;
  assign new_new_n7729__ = ~new_new_n7727__ & ~new_new_n7728__;
  assign new_new_n7730__ = new_new_n7726__ & ~new_new_n7729__;
  assign new_new_n7731__ = ~new_new_n7726__ & new_new_n7729__;
  assign new_new_n7732__ = ~new_new_n7730__ & ~new_new_n7731__;
  assign new_new_n7733__ = ~pi090 & ~new_new_n7732__;
  assign new_new_n7734__ = pi090 & new_new_n7732__;
  assign new_new_n7735__ = ~new_new_n7353__ & ~new_new_n7354__;
  assign new_new_n7736__ = ~new_new_n7623__ & po028;
  assign new_new_n7737__ = pi088 & ~po028;
  assign new_new_n7738__ = ~new_new_n7736__ & ~new_new_n7737__;
  assign new_new_n7739__ = new_new_n7735__ & ~new_new_n7738__;
  assign new_new_n7740__ = ~new_new_n7735__ & new_new_n7738__;
  assign new_new_n7741__ = ~new_new_n7739__ & ~new_new_n7740__;
  assign new_new_n7742__ = ~pi089 & ~new_new_n7741__;
  assign new_new_n7743__ = pi089 & new_new_n7741__;
  assign new_new_n7744__ = ~new_new_n7621__ & po028;
  assign new_new_n7745__ = pi087 & ~po028;
  assign new_new_n7746__ = ~new_new_n7744__ & ~new_new_n7745__;
  assign new_new_n7747__ = ~new_new_n7362__ & ~new_new_n7363__;
  assign new_new_n7748__ = ~new_new_n7746__ & new_new_n7747__;
  assign new_new_n7749__ = new_new_n7746__ & ~new_new_n7747__;
  assign new_new_n7750__ = ~new_new_n7748__ & ~new_new_n7749__;
  assign new_new_n7751__ = ~pi088 & ~new_new_n7750__;
  assign new_new_n7752__ = pi088 & new_new_n7750__;
  assign new_new_n7753__ = ~new_new_n7371__ & ~new_new_n7372__;
  assign new_new_n7754__ = ~new_new_n7619__ & po028;
  assign new_new_n7755__ = pi086 & ~po028;
  assign new_new_n7756__ = ~new_new_n7754__ & ~new_new_n7755__;
  assign new_new_n7757__ = new_new_n7753__ & new_new_n7756__;
  assign new_new_n7758__ = ~new_new_n7753__ & ~new_new_n7756__;
  assign new_new_n7759__ = ~new_new_n7757__ & ~new_new_n7758__;
  assign new_new_n7760__ = ~pi087 & new_new_n7759__;
  assign new_new_n7761__ = pi087 & ~new_new_n7759__;
  assign new_new_n7762__ = ~new_new_n7617__ & po028;
  assign new_new_n7763__ = pi085 & ~po028;
  assign new_new_n7764__ = ~new_new_n7762__ & ~new_new_n7763__;
  assign new_new_n7765__ = ~new_new_n7380__ & ~new_new_n7381__;
  assign new_new_n7766__ = ~new_new_n7764__ & new_new_n7765__;
  assign new_new_n7767__ = new_new_n7764__ & ~new_new_n7765__;
  assign new_new_n7768__ = ~new_new_n7766__ & ~new_new_n7767__;
  assign new_new_n7769__ = ~pi086 & ~new_new_n7768__;
  assign new_new_n7770__ = ~new_new_n7389__ & ~new_new_n7390__;
  assign new_new_n7771__ = ~new_new_n7615__ & po028;
  assign new_new_n7772__ = pi084 & ~po028;
  assign new_new_n7773__ = ~new_new_n7771__ & ~new_new_n7772__;
  assign new_new_n7774__ = new_new_n7770__ & ~new_new_n7773__;
  assign new_new_n7775__ = ~new_new_n7770__ & new_new_n7773__;
  assign new_new_n7776__ = ~new_new_n7774__ & ~new_new_n7775__;
  assign new_new_n7777__ = ~pi085 & ~new_new_n7776__;
  assign new_new_n7778__ = pi085 & new_new_n7776__;
  assign new_new_n7779__ = ~new_new_n7613__ & po028;
  assign new_new_n7780__ = pi083 & ~po028;
  assign new_new_n7781__ = ~new_new_n7779__ & ~new_new_n7780__;
  assign new_new_n7782__ = ~new_new_n7398__ & ~new_new_n7399__;
  assign new_new_n7783__ = ~new_new_n7781__ & new_new_n7782__;
  assign new_new_n7784__ = new_new_n7781__ & ~new_new_n7782__;
  assign new_new_n7785__ = ~new_new_n7783__ & ~new_new_n7784__;
  assign new_new_n7786__ = ~pi084 & ~new_new_n7785__;
  assign new_new_n7787__ = pi084 & new_new_n7785__;
  assign new_new_n7788__ = ~new_new_n7407__ & ~new_new_n7408__;
  assign new_new_n7789__ = new_new_n7611__ & po028;
  assign new_new_n7790__ = ~pi082 & ~po028;
  assign new_new_n7791__ = ~new_new_n7789__ & ~new_new_n7790__;
  assign new_new_n7792__ = ~new_new_n7788__ & ~new_new_n7791__;
  assign new_new_n7793__ = new_new_n7788__ & new_new_n7791__;
  assign new_new_n7794__ = ~new_new_n7792__ & ~new_new_n7793__;
  assign new_new_n7795__ = ~pi083 & ~new_new_n7794__;
  assign new_new_n7796__ = pi083 & new_new_n7794__;
  assign new_new_n7797__ = new_new_n7609__ & po028;
  assign new_new_n7798__ = ~pi081 & ~po028;
  assign new_new_n7799__ = ~new_new_n7797__ & ~new_new_n7798__;
  assign new_new_n7800__ = ~new_new_n7416__ & ~new_new_n7417__;
  assign new_new_n7801__ = ~new_new_n7799__ & ~new_new_n7800__;
  assign new_new_n7802__ = new_new_n7799__ & new_new_n7800__;
  assign new_new_n7803__ = ~new_new_n7801__ & ~new_new_n7802__;
  assign new_new_n7804__ = pi082 & new_new_n7803__;
  assign new_new_n7805__ = ~pi082 & ~new_new_n7803__;
  assign new_new_n7806__ = ~new_new_n7607__ & po028;
  assign new_new_n7807__ = pi080 & ~po028;
  assign new_new_n7808__ = ~new_new_n7806__ & ~new_new_n7807__;
  assign new_new_n7809__ = ~new_new_n7425__ & ~new_new_n7426__;
  assign new_new_n7810__ = ~new_new_n7808__ & new_new_n7809__;
  assign new_new_n7811__ = new_new_n7808__ & ~new_new_n7809__;
  assign new_new_n7812__ = ~new_new_n7810__ & ~new_new_n7811__;
  assign new_new_n7813__ = pi081 & new_new_n7812__;
  assign new_new_n7814__ = ~pi081 & ~new_new_n7812__;
  assign new_new_n7815__ = ~new_new_n7434__ & ~new_new_n7435__;
  assign new_new_n7816__ = pi079 & ~po028;
  assign new_new_n7817__ = ~new_new_n7605__ & po028;
  assign new_new_n7818__ = ~new_new_n7816__ & ~new_new_n7817__;
  assign new_new_n7819__ = new_new_n7815__ & new_new_n7818__;
  assign new_new_n7820__ = ~new_new_n7815__ & ~new_new_n7818__;
  assign new_new_n7821__ = ~new_new_n7819__ & ~new_new_n7820__;
  assign new_new_n7822__ = pi080 & ~new_new_n7821__;
  assign new_new_n7823__ = ~pi080 & new_new_n7821__;
  assign new_new_n7824__ = ~new_new_n7443__ & ~new_new_n7444__;
  assign new_new_n7825__ = ~new_new_n7603__ & po028;
  assign new_new_n7826__ = pi078 & ~po028;
  assign new_new_n7827__ = ~new_new_n7825__ & ~new_new_n7826__;
  assign new_new_n7828__ = new_new_n7824__ & new_new_n7827__;
  assign new_new_n7829__ = ~new_new_n7824__ & ~new_new_n7827__;
  assign new_new_n7830__ = ~new_new_n7828__ & ~new_new_n7829__;
  assign new_new_n7831__ = pi079 & ~new_new_n7830__;
  assign new_new_n7832__ = ~pi079 & new_new_n7830__;
  assign new_new_n7833__ = new_new_n7601__ & po028;
  assign new_new_n7834__ = pi077 & ~po028;
  assign new_new_n7835__ = ~new_new_n7833__ & ~new_new_n7834__;
  assign new_new_n7836__ = ~new_new_n7452__ & ~new_new_n7453__;
  assign new_new_n7837__ = ~new_new_n7835__ & ~new_new_n7836__;
  assign new_new_n7838__ = new_new_n7835__ & new_new_n7836__;
  assign new_new_n7839__ = ~new_new_n7837__ & ~new_new_n7838__;
  assign new_new_n7840__ = pi078 & ~new_new_n7839__;
  assign new_new_n7841__ = ~pi078 & new_new_n7839__;
  assign new_new_n7842__ = ~new_new_n7461__ & ~new_new_n7462__;
  assign new_new_n7843__ = ~new_new_n7599__ & po028;
  assign new_new_n7844__ = ~pi076 & ~po028;
  assign new_new_n7845__ = ~new_new_n7843__ & ~new_new_n7844__;
  assign new_new_n7846__ = new_new_n7842__ & ~new_new_n7845__;
  assign new_new_n7847__ = ~new_new_n7842__ & new_new_n7845__;
  assign new_new_n7848__ = ~new_new_n7846__ & ~new_new_n7847__;
  assign new_new_n7849__ = pi077 & ~new_new_n7848__;
  assign new_new_n7850__ = ~pi077 & new_new_n7848__;
  assign new_new_n7851__ = ~new_new_n7470__ & ~new_new_n7471__;
  assign new_new_n7852__ = ~new_new_n7597__ & po028;
  assign new_new_n7853__ = ~pi075 & ~po028;
  assign new_new_n7854__ = ~new_new_n7852__ & ~new_new_n7853__;
  assign new_new_n7855__ = new_new_n7851__ & ~new_new_n7854__;
  assign new_new_n7856__ = ~new_new_n7851__ & new_new_n7854__;
  assign new_new_n7857__ = ~new_new_n7855__ & ~new_new_n7856__;
  assign new_new_n7858__ = pi076 & ~new_new_n7857__;
  assign new_new_n7859__ = ~pi076 & new_new_n7857__;
  assign new_new_n7860__ = ~new_new_n7479__ & ~new_new_n7480__;
  assign new_new_n7861__ = ~new_new_n7595__ & po028;
  assign new_new_n7862__ = ~pi074 & ~po028;
  assign new_new_n7863__ = ~new_new_n7861__ & ~new_new_n7862__;
  assign new_new_n7864__ = new_new_n7860__ & ~new_new_n7863__;
  assign new_new_n7865__ = ~new_new_n7860__ & new_new_n7863__;
  assign new_new_n7866__ = ~new_new_n7864__ & ~new_new_n7865__;
  assign new_new_n7867__ = pi075 & ~new_new_n7866__;
  assign new_new_n7868__ = ~pi075 & new_new_n7866__;
  assign new_new_n7869__ = ~new_new_n7593__ & po028;
  assign new_new_n7870__ = pi073 & ~po028;
  assign new_new_n7871__ = ~new_new_n7869__ & ~new_new_n7870__;
  assign new_new_n7872__ = ~new_new_n7488__ & ~new_new_n7489__;
  assign new_new_n7873__ = ~new_new_n7871__ & new_new_n7872__;
  assign new_new_n7874__ = new_new_n7871__ & ~new_new_n7872__;
  assign new_new_n7875__ = ~new_new_n7873__ & ~new_new_n7874__;
  assign new_new_n7876__ = ~pi074 & ~new_new_n7875__;
  assign new_new_n7877__ = pi074 & new_new_n7875__;
  assign new_new_n7878__ = ~new_new_n7497__ & ~new_new_n7498__;
  assign new_new_n7879__ = ~new_new_n7591__ & po028;
  assign new_new_n7880__ = ~pi072 & ~po028;
  assign new_new_n7881__ = ~new_new_n7879__ & ~new_new_n7880__;
  assign new_new_n7882__ = new_new_n7878__ & new_new_n7881__;
  assign new_new_n7883__ = ~new_new_n7878__ & ~new_new_n7881__;
  assign new_new_n7884__ = ~new_new_n7882__ & ~new_new_n7883__;
  assign new_new_n7885__ = ~pi073 & ~new_new_n7884__;
  assign new_new_n7886__ = pi073 & new_new_n7884__;
  assign new_new_n7887__ = ~pi071 & ~new_new_n7589__;
  assign new_new_n7888__ = pi071 & new_new_n7589__;
  assign new_new_n7889__ = ~new_new_n7887__ & ~new_new_n7888__;
  assign new_new_n7890__ = po028 & new_new_n7889__;
  assign new_new_n7891__ = ~new_new_n7505__ & ~new_new_n7890__;
  assign new_new_n7892__ = new_new_n7505__ & new_new_n7890__;
  assign new_new_n7893__ = ~new_new_n7891__ & ~new_new_n7892__;
  assign new_new_n7894__ = ~pi072 & ~new_new_n7893__;
  assign new_new_n7895__ = pi072 & new_new_n7893__;
  assign new_new_n7896__ = new_new_n7587__ & po028;
  assign new_new_n7897__ = ~pi070 & ~po028;
  assign new_new_n7898__ = ~new_new_n7896__ & ~new_new_n7897__;
  assign new_new_n7899__ = ~new_new_n7515__ & ~new_new_n7516__;
  assign new_new_n7900__ = ~new_new_n7898__ & ~new_new_n7899__;
  assign new_new_n7901__ = new_new_n7898__ & new_new_n7899__;
  assign new_new_n7902__ = ~new_new_n7900__ & ~new_new_n7901__;
  assign new_new_n7903__ = ~pi071 & ~new_new_n7902__;
  assign new_new_n7904__ = pi071 & new_new_n7902__;
  assign new_new_n7905__ = ~new_new_n7531__ & ~new_new_n7532__;
  assign new_new_n7906__ = ~new_new_n7583__ & po028;
  assign new_new_n7907__ = ~pi068 & ~po028;
  assign new_new_n7908__ = ~new_new_n7906__ & ~new_new_n7907__;
  assign new_new_n7909__ = new_new_n7905__ & ~new_new_n7908__;
  assign new_new_n7910__ = ~new_new_n7905__ & new_new_n7908__;
  assign new_new_n7911__ = ~new_new_n7909__ & ~new_new_n7910__;
  assign new_new_n7912__ = ~pi069 & new_new_n7911__;
  assign new_new_n7913__ = ~new_new_n7575__ & ~new_new_n7582__;
  assign new_new_n7914__ = po028 & new_new_n7913__;
  assign new_new_n7915__ = new_new_n7580__ & ~new_new_n7914__;
  assign new_new_n7916__ = ~new_new_n7580__ & new_new_n7914__;
  assign new_new_n7917__ = ~new_new_n7915__ & ~new_new_n7916__;
  assign new_new_n7918__ = pi068 & ~new_new_n7917__;
  assign new_new_n7919__ = ~pi068 & new_new_n7917__;
  assign new_new_n7920__ = ~new_new_n7545__ & ~new_new_n7546__;
  assign new_new_n7921__ = po028 & new_new_n7920__;
  assign new_new_n7922__ = new_new_n7572__ & ~new_new_n7921__;
  assign new_new_n7923__ = ~new_new_n7572__ & new_new_n7921__;
  assign new_new_n7924__ = ~new_new_n7922__ & ~new_new_n7923__;
  assign new_new_n7925__ = pi067 & ~new_new_n7924__;
  assign new_new_n7926__ = ~pi067 & new_new_n7924__;
  assign new_new_n7927__ = pi028 & po028;
  assign new_new_n7928__ = pi027 & ~pi065;
  assign new_new_n7929__ = new_new_n7927__ & ~new_new_n7928__;
  assign new_new_n7930__ = ~pi028 & ~po028;
  assign new_new_n7931__ = ~pi065 & ~new_new_n7930__;
  assign new_new_n7932__ = ~pi027 & ~new_new_n7931__;
  assign new_new_n7933__ = ~new_new_n7929__ & ~new_new_n7932__;
  assign new_new_n7934__ = pi064 & ~new_new_n7933__;
  assign new_new_n7935__ = pi064 & po028;
  assign new_new_n7936__ = ~pi028 & pi065;
  assign new_new_n7937__ = ~new_new_n7935__ & new_new_n7936__;
  assign new_new_n7938__ = ~new_new_n7934__ & ~new_new_n7937__;
  assign new_new_n7939__ = pi066 & ~new_new_n7938__;
  assign new_new_n7940__ = new_new_n426__ & ~po029;
  assign new_new_n7941__ = new_new_n7565__ & po028;
  assign new_new_n7942__ = ~new_new_n7940__ & ~new_new_n7941__;
  assign new_new_n7943__ = ~pi028 & ~new_new_n7942__;
  assign new_new_n7944__ = ~new_new_n332__ & po028;
  assign new_new_n7945__ = ~new_new_n7541__ & ~new_new_n7944__;
  assign new_new_n7946__ = pi065 & po028;
  assign new_new_n7947__ = po029 & ~new_new_n7946__;
  assign new_new_n7948__ = pi065 & ~new_new_n7541__;
  assign new_new_n7949__ = pi028 & ~new_new_n7948__;
  assign new_new_n7950__ = ~new_new_n7947__ & new_new_n7949__;
  assign new_new_n7951__ = ~new_new_n7943__ & ~new_new_n7945__;
  assign new_new_n7952__ = ~new_new_n7950__ & new_new_n7951__;
  assign new_new_n7953__ = ~pi029 & ~new_new_n7952__;
  assign new_new_n7954__ = ~new_new_n7541__ & ~new_new_n7946__;
  assign new_new_n7955__ = pi028 & ~new_new_n7553__;
  assign new_new_n7956__ = pi064 & ~new_new_n7955__;
  assign new_new_n7957__ = ~new_new_n7954__ & ~new_new_n7956__;
  assign new_new_n7958__ = ~pi065 & po028;
  assign new_new_n7959__ = ~po029 & ~new_new_n7958__;
  assign new_new_n7960__ = pi064 & ~new_new_n7927__;
  assign new_new_n7961__ = ~new_new_n7941__ & new_new_n7960__;
  assign new_new_n7962__ = ~new_new_n7959__ & new_new_n7961__;
  assign new_new_n7963__ = ~new_new_n7957__ & ~new_new_n7962__;
  assign new_new_n7964__ = pi029 & ~new_new_n7963__;
  assign new_new_n7965__ = ~new_new_n7953__ & ~new_new_n7964__;
  assign new_new_n7966__ = ~pi066 & new_new_n7938__;
  assign new_new_n7967__ = ~new_new_n7965__ & ~new_new_n7966__;
  assign new_new_n7968__ = ~new_new_n7939__ & ~new_new_n7967__;
  assign new_new_n7969__ = ~new_new_n7926__ & ~new_new_n7968__;
  assign new_new_n7970__ = ~new_new_n7925__ & ~new_new_n7969__;
  assign new_new_n7971__ = ~new_new_n7919__ & ~new_new_n7970__;
  assign new_new_n7972__ = ~new_new_n7918__ & ~new_new_n7971__;
  assign new_new_n7973__ = ~new_new_n7912__ & ~new_new_n7972__;
  assign new_new_n7974__ = pi069 & ~new_new_n7911__;
  assign new_new_n7975__ = ~new_new_n7973__ & ~new_new_n7974__;
  assign new_new_n7976__ = pi070 & ~new_new_n7975__;
  assign new_new_n7977__ = ~pi070 & new_new_n7975__;
  assign new_new_n7978__ = ~new_new_n7522__ & ~new_new_n7523__;
  assign new_new_n7979__ = ~new_new_n7585__ & po028;
  assign new_new_n7980__ = pi069 & ~po028;
  assign new_new_n7981__ = ~new_new_n7979__ & ~new_new_n7980__;
  assign new_new_n7982__ = new_new_n7978__ & ~new_new_n7981__;
  assign new_new_n7983__ = ~new_new_n7978__ & new_new_n7981__;
  assign new_new_n7984__ = ~new_new_n7982__ & ~new_new_n7983__;
  assign new_new_n7985__ = ~new_new_n7977__ & new_new_n7984__;
  assign new_new_n7986__ = ~new_new_n7976__ & ~new_new_n7985__;
  assign new_new_n7987__ = ~new_new_n7904__ & new_new_n7986__;
  assign new_new_n7988__ = ~new_new_n7903__ & ~new_new_n7987__;
  assign new_new_n7989__ = ~new_new_n7895__ & ~new_new_n7988__;
  assign new_new_n7990__ = ~new_new_n7894__ & ~new_new_n7989__;
  assign new_new_n7991__ = ~new_new_n7886__ & ~new_new_n7990__;
  assign new_new_n7992__ = ~new_new_n7885__ & ~new_new_n7991__;
  assign new_new_n7993__ = ~new_new_n7877__ & ~new_new_n7992__;
  assign new_new_n7994__ = ~new_new_n7876__ & ~new_new_n7993__;
  assign new_new_n7995__ = ~new_new_n7868__ & new_new_n7994__;
  assign new_new_n7996__ = ~new_new_n7867__ & ~new_new_n7995__;
  assign new_new_n7997__ = ~new_new_n7859__ & ~new_new_n7996__;
  assign new_new_n7998__ = ~new_new_n7858__ & ~new_new_n7997__;
  assign new_new_n7999__ = ~new_new_n7850__ & ~new_new_n7998__;
  assign new_new_n8000__ = ~new_new_n7849__ & ~new_new_n7999__;
  assign new_new_n8001__ = ~new_new_n7841__ & ~new_new_n8000__;
  assign new_new_n8002__ = ~new_new_n7840__ & ~new_new_n8001__;
  assign new_new_n8003__ = ~new_new_n7832__ & ~new_new_n8002__;
  assign new_new_n8004__ = ~new_new_n7831__ & ~new_new_n8003__;
  assign new_new_n8005__ = ~new_new_n7823__ & ~new_new_n8004__;
  assign new_new_n8006__ = ~new_new_n7822__ & ~new_new_n8005__;
  assign new_new_n8007__ = ~new_new_n7814__ & ~new_new_n8006__;
  assign new_new_n8008__ = ~new_new_n7813__ & ~new_new_n8007__;
  assign new_new_n8009__ = ~new_new_n7805__ & ~new_new_n8008__;
  assign new_new_n8010__ = ~new_new_n7804__ & ~new_new_n8009__;
  assign new_new_n8011__ = ~new_new_n7796__ & new_new_n8010__;
  assign new_new_n8012__ = ~new_new_n7795__ & ~new_new_n8011__;
  assign new_new_n8013__ = ~new_new_n7787__ & ~new_new_n8012__;
  assign new_new_n8014__ = ~new_new_n7786__ & ~new_new_n8013__;
  assign new_new_n8015__ = ~new_new_n7778__ & ~new_new_n8014__;
  assign new_new_n8016__ = ~new_new_n7777__ & ~new_new_n8015__;
  assign new_new_n8017__ = pi086 & new_new_n7768__;
  assign new_new_n8018__ = ~new_new_n8016__ & ~new_new_n8017__;
  assign new_new_n8019__ = ~new_new_n7769__ & ~new_new_n8018__;
  assign new_new_n8020__ = ~new_new_n7761__ & ~new_new_n8019__;
  assign new_new_n8021__ = ~new_new_n7760__ & ~new_new_n8020__;
  assign new_new_n8022__ = ~new_new_n7752__ & ~new_new_n8021__;
  assign new_new_n8023__ = ~new_new_n7751__ & ~new_new_n8022__;
  assign new_new_n8024__ = ~new_new_n7743__ & ~new_new_n8023__;
  assign new_new_n8025__ = ~new_new_n7742__ & ~new_new_n8024__;
  assign new_new_n8026__ = ~new_new_n7734__ & ~new_new_n8025__;
  assign new_new_n8027__ = ~new_new_n7733__ & ~new_new_n8026__;
  assign new_new_n8028__ = ~new_new_n7725__ & new_new_n8027__;
  assign new_new_n8029__ = ~new_new_n7724__ & ~new_new_n8028__;
  assign new_new_n8030__ = ~new_new_n7716__ & new_new_n8029__;
  assign new_new_n8031__ = ~new_new_n7715__ & ~new_new_n8030__;
  assign new_new_n8032__ = ~new_new_n7707__ & ~new_new_n8031__;
  assign new_new_n8033__ = ~new_new_n7706__ & ~new_new_n8032__;
  assign new_new_n8034__ = ~new_new_n7698__ & ~new_new_n8033__;
  assign new_new_n8035__ = ~new_new_n7697__ & ~new_new_n8034__;
  assign new_new_n8036__ = ~new_new_n7689__ & new_new_n8035__;
  assign new_new_n8037__ = ~new_new_n7688__ & ~new_new_n8036__;
  assign new_new_n8038__ = ~new_new_n7680__ & ~new_new_n8037__;
  assign new_new_n8039__ = ~new_new_n7679__ & ~new_new_n8038__;
  assign new_new_n8040__ = ~new_new_n7671__ & ~new_new_n8039__;
  assign new_new_n8041__ = ~new_new_n7670__ & ~new_new_n8040__;
  assign new_new_n8042__ = pi098 & ~new_new_n8041__;
  assign new_new_n8043__ = ~pi098 & new_new_n8041__;
  assign new_new_n8044__ = ~pi097 & ~new_new_n7641__;
  assign new_new_n8045__ = pi097 & new_new_n7641__;
  assign new_new_n8046__ = ~new_new_n8044__ & ~new_new_n8045__;
  assign new_new_n8047__ = po028 & new_new_n8046__;
  assign new_new_n8048__ = new_new_n7271__ & new_new_n8047__;
  assign new_new_n8049__ = ~new_new_n7271__ & ~new_new_n8047__;
  assign new_new_n8050__ = ~new_new_n8048__ & ~new_new_n8049__;
  assign new_new_n8051__ = ~new_new_n8043__ & new_new_n8050__;
  assign new_new_n8052__ = ~new_new_n8042__ & ~new_new_n8051__;
  assign new_new_n8053__ = pi099 & ~new_new_n8052__;
  assign new_new_n8054__ = new_new_n7662__ & ~new_new_n8053__;
  assign new_new_n8055__ = ~pi099 & new_new_n8052__;
  assign new_new_n8056__ = ~new_new_n376__ & ~new_new_n7652__;
  assign new_new_n8057__ = ~pi100 & ~new_new_n8056__;
  assign new_new_n8058__ = ~new_new_n8055__ & ~new_new_n8057__;
  assign new_new_n8059__ = ~new_new_n8054__ & new_new_n8058__;
  assign new_new_n8060__ = pi100 & new_new_n8056__;
  assign new_new_n8061__ = new_new_n7647__ & ~new_new_n8060__;
  assign po027 = ~new_new_n8059__ & new_new_n8061__;
  assign new_new_n8063__ = new_new_n7652__ & ~po027;
  assign new_new_n8064__ = ~new_new_n376__ & ~new_new_n8063__;
  assign new_new_n8065__ = ~pi111 & new_new_n274__;
  assign new_new_n8066__ = ~pi110 & new_new_n8065__;
  assign new_new_n8067__ = new_new_n276__ & new_new_n280__;
  assign new_new_n8068__ = new_new_n8066__ & new_new_n8067__;
  assign new_new_n8069__ = ~pi104 & new_new_n8068__;
  assign new_new_n8070__ = ~pi103 & new_new_n8069__;
  assign new_new_n8071__ = ~new_new_n8053__ & ~new_new_n8055__;
  assign new_new_n8072__ = po027 & new_new_n8071__;
  assign new_new_n8073__ = ~new_new_n7662__ & ~new_new_n8072__;
  assign new_new_n8074__ = new_new_n7662__ & new_new_n8072__;
  assign new_new_n8075__ = ~new_new_n8073__ & ~new_new_n8074__;
  assign new_new_n8076__ = ~new_new_n8042__ & ~new_new_n8043__;
  assign new_new_n8077__ = po027 & new_new_n8076__;
  assign new_new_n8078__ = ~new_new_n8050__ & new_new_n8077__;
  assign new_new_n8079__ = new_new_n8050__ & ~new_new_n8077__;
  assign new_new_n8080__ = ~new_new_n8078__ & ~new_new_n8079__;
  assign new_new_n8081__ = pi099 & ~new_new_n8080__;
  assign new_new_n8082__ = ~pi099 & new_new_n8080__;
  assign new_new_n8083__ = ~new_new_n7670__ & ~new_new_n7671__;
  assign new_new_n8084__ = ~new_new_n8039__ & po027;
  assign new_new_n8085__ = pi097 & ~po027;
  assign new_new_n8086__ = ~new_new_n8084__ & ~new_new_n8085__;
  assign new_new_n8087__ = new_new_n8083__ & ~new_new_n8086__;
  assign new_new_n8088__ = ~new_new_n8083__ & new_new_n8086__;
  assign new_new_n8089__ = ~new_new_n8087__ & ~new_new_n8088__;
  assign new_new_n8090__ = ~pi098 & ~new_new_n8089__;
  assign new_new_n8091__ = pi098 & new_new_n8089__;
  assign new_new_n8092__ = ~new_new_n8037__ & po027;
  assign new_new_n8093__ = pi096 & ~po027;
  assign new_new_n8094__ = ~new_new_n8092__ & ~new_new_n8093__;
  assign new_new_n8095__ = ~new_new_n7679__ & ~new_new_n7680__;
  assign new_new_n8096__ = ~new_new_n8094__ & new_new_n8095__;
  assign new_new_n8097__ = new_new_n8094__ & ~new_new_n8095__;
  assign new_new_n8098__ = ~new_new_n8096__ & ~new_new_n8097__;
  assign new_new_n8099__ = ~pi097 & ~new_new_n8098__;
  assign new_new_n8100__ = pi097 & new_new_n8098__;
  assign new_new_n8101__ = ~new_new_n7688__ & ~new_new_n7689__;
  assign new_new_n8102__ = ~new_new_n8035__ & po027;
  assign new_new_n8103__ = ~pi095 & ~po027;
  assign new_new_n8104__ = ~new_new_n8102__ & ~new_new_n8103__;
  assign new_new_n8105__ = new_new_n8101__ & ~new_new_n8104__;
  assign new_new_n8106__ = ~new_new_n8101__ & new_new_n8104__;
  assign new_new_n8107__ = ~new_new_n8105__ & ~new_new_n8106__;
  assign new_new_n8108__ = ~pi096 & new_new_n8107__;
  assign new_new_n8109__ = pi096 & ~new_new_n8107__;
  assign new_new_n8110__ = ~pi094 & ~new_new_n8033__;
  assign new_new_n8111__ = pi094 & new_new_n8033__;
  assign new_new_n8112__ = ~new_new_n8110__ & ~new_new_n8111__;
  assign new_new_n8113__ = po027 & new_new_n8112__;
  assign new_new_n8114__ = new_new_n7696__ & new_new_n8113__;
  assign new_new_n8115__ = ~new_new_n7696__ & ~new_new_n8113__;
  assign new_new_n8116__ = ~new_new_n8114__ & ~new_new_n8115__;
  assign new_new_n8117__ = ~pi095 & ~new_new_n8116__;
  assign new_new_n8118__ = pi095 & new_new_n8116__;
  assign new_new_n8119__ = ~pi093 & ~new_new_n8031__;
  assign new_new_n8120__ = pi093 & new_new_n8031__;
  assign new_new_n8121__ = ~new_new_n8119__ & ~new_new_n8120__;
  assign new_new_n8122__ = po027 & new_new_n8121__;
  assign new_new_n8123__ = new_new_n7705__ & new_new_n8122__;
  assign new_new_n8124__ = ~new_new_n7705__ & ~new_new_n8122__;
  assign new_new_n8125__ = ~new_new_n8123__ & ~new_new_n8124__;
  assign new_new_n8126__ = ~pi094 & ~new_new_n8125__;
  assign new_new_n8127__ = pi094 & new_new_n8125__;
  assign new_new_n8128__ = ~new_new_n7715__ & ~new_new_n7716__;
  assign new_new_n8129__ = ~new_new_n8029__ & po027;
  assign new_new_n8130__ = pi092 & ~po027;
  assign new_new_n8131__ = ~new_new_n8129__ & ~new_new_n8130__;
  assign new_new_n8132__ = new_new_n8128__ & ~new_new_n8131__;
  assign new_new_n8133__ = ~new_new_n8128__ & new_new_n8131__;
  assign new_new_n8134__ = ~new_new_n8132__ & ~new_new_n8133__;
  assign new_new_n8135__ = ~pi093 & ~new_new_n8134__;
  assign new_new_n8136__ = pi093 & new_new_n8134__;
  assign new_new_n8137__ = ~new_new_n7724__ & ~new_new_n7725__;
  assign new_new_n8138__ = ~new_new_n8027__ & po027;
  assign new_new_n8139__ = ~pi091 & ~po027;
  assign new_new_n8140__ = ~new_new_n8138__ & ~new_new_n8139__;
  assign new_new_n8141__ = new_new_n8137__ & ~new_new_n8140__;
  assign new_new_n8142__ = ~new_new_n8137__ & new_new_n8140__;
  assign new_new_n8143__ = ~new_new_n8141__ & ~new_new_n8142__;
  assign new_new_n8144__ = pi092 & ~new_new_n8143__;
  assign new_new_n8145__ = ~pi092 & new_new_n8143__;
  assign new_new_n8146__ = ~pi090 & ~new_new_n8025__;
  assign new_new_n8147__ = pi090 & new_new_n8025__;
  assign new_new_n8148__ = ~new_new_n8146__ & ~new_new_n8147__;
  assign new_new_n8149__ = po027 & new_new_n8148__;
  assign new_new_n8150__ = new_new_n7732__ & new_new_n8149__;
  assign new_new_n8151__ = ~new_new_n7732__ & ~new_new_n8149__;
  assign new_new_n8152__ = ~new_new_n8150__ & ~new_new_n8151__;
  assign new_new_n8153__ = pi091 & new_new_n8152__;
  assign new_new_n8154__ = ~pi091 & ~new_new_n8152__;
  assign new_new_n8155__ = ~pi089 & ~new_new_n8023__;
  assign new_new_n8156__ = pi089 & new_new_n8023__;
  assign new_new_n8157__ = ~new_new_n8155__ & ~new_new_n8156__;
  assign new_new_n8158__ = po027 & new_new_n8157__;
  assign new_new_n8159__ = new_new_n7741__ & new_new_n8158__;
  assign new_new_n8160__ = ~new_new_n7741__ & ~new_new_n8158__;
  assign new_new_n8161__ = ~new_new_n8159__ & ~new_new_n8160__;
  assign new_new_n8162__ = pi090 & new_new_n8161__;
  assign new_new_n8163__ = ~pi090 & ~new_new_n8161__;
  assign new_new_n8164__ = ~new_new_n7751__ & ~new_new_n7752__;
  assign new_new_n8165__ = ~new_new_n8021__ & po027;
  assign new_new_n8166__ = ~pi088 & ~po027;
  assign new_new_n8167__ = ~new_new_n8165__ & ~new_new_n8166__;
  assign new_new_n8168__ = new_new_n8164__ & ~new_new_n8167__;
  assign new_new_n8169__ = ~new_new_n8164__ & new_new_n8167__;
  assign new_new_n8170__ = ~new_new_n8168__ & ~new_new_n8169__;
  assign new_new_n8171__ = pi089 & ~new_new_n8170__;
  assign new_new_n8172__ = ~pi089 & new_new_n8170__;
  assign new_new_n8173__ = ~new_new_n7760__ & ~new_new_n7761__;
  assign new_new_n8174__ = ~new_new_n8019__ & po027;
  assign new_new_n8175__ = ~pi087 & ~po027;
  assign new_new_n8176__ = ~new_new_n8174__ & ~new_new_n8175__;
  assign new_new_n8177__ = new_new_n8173__ & ~new_new_n8176__;
  assign new_new_n8178__ = ~new_new_n8173__ & new_new_n8176__;
  assign new_new_n8179__ = ~new_new_n8177__ & ~new_new_n8178__;
  assign new_new_n8180__ = pi088 & ~new_new_n8179__;
  assign new_new_n8181__ = ~pi088 & new_new_n8179__;
  assign new_new_n8182__ = ~new_new_n7769__ & ~new_new_n8017__;
  assign new_new_n8183__ = ~new_new_n8016__ & po027;
  assign new_new_n8184__ = ~pi086 & ~po027;
  assign new_new_n8185__ = ~new_new_n8183__ & ~new_new_n8184__;
  assign new_new_n8186__ = new_new_n8182__ & ~new_new_n8185__;
  assign new_new_n8187__ = ~new_new_n8182__ & new_new_n8185__;
  assign new_new_n8188__ = ~new_new_n8186__ & ~new_new_n8187__;
  assign new_new_n8189__ = pi087 & ~new_new_n8188__;
  assign new_new_n8190__ = ~pi087 & new_new_n8188__;
  assign new_new_n8191__ = ~pi085 & ~new_new_n8014__;
  assign new_new_n8192__ = pi085 & new_new_n8014__;
  assign new_new_n8193__ = ~new_new_n8191__ & ~new_new_n8192__;
  assign new_new_n8194__ = po027 & new_new_n8193__;
  assign new_new_n8195__ = new_new_n7776__ & new_new_n8194__;
  assign new_new_n8196__ = ~new_new_n7776__ & ~new_new_n8194__;
  assign new_new_n8197__ = ~new_new_n8195__ & ~new_new_n8196__;
  assign new_new_n8198__ = ~pi086 & ~new_new_n8197__;
  assign new_new_n8199__ = pi086 & new_new_n8197__;
  assign new_new_n8200__ = ~new_new_n7786__ & ~new_new_n7787__;
  assign new_new_n8201__ = ~new_new_n8012__ & po027;
  assign new_new_n8202__ = ~pi084 & ~po027;
  assign new_new_n8203__ = ~new_new_n8201__ & ~new_new_n8202__;
  assign new_new_n8204__ = ~new_new_n8200__ & ~new_new_n8203__;
  assign new_new_n8205__ = new_new_n8200__ & new_new_n8203__;
  assign new_new_n8206__ = ~new_new_n8204__ & ~new_new_n8205__;
  assign new_new_n8207__ = ~pi085 & ~new_new_n8206__;
  assign new_new_n8208__ = pi085 & new_new_n8206__;
  assign new_new_n8209__ = new_new_n8010__ & po027;
  assign new_new_n8210__ = ~pi083 & ~po027;
  assign new_new_n8211__ = ~new_new_n8209__ & ~new_new_n8210__;
  assign new_new_n8212__ = ~new_new_n7795__ & ~new_new_n7796__;
  assign new_new_n8213__ = ~new_new_n8211__ & ~new_new_n8212__;
  assign new_new_n8214__ = new_new_n8211__ & new_new_n8212__;
  assign new_new_n8215__ = ~new_new_n8213__ & ~new_new_n8214__;
  assign new_new_n8216__ = ~pi084 & ~new_new_n8215__;
  assign new_new_n8217__ = pi084 & new_new_n8215__;
  assign new_new_n8218__ = ~new_new_n8008__ & po027;
  assign new_new_n8219__ = pi082 & ~po027;
  assign new_new_n8220__ = ~new_new_n8218__ & ~new_new_n8219__;
  assign new_new_n8221__ = ~new_new_n7804__ & ~new_new_n7805__;
  assign new_new_n8222__ = ~new_new_n8220__ & new_new_n8221__;
  assign new_new_n8223__ = new_new_n8220__ & ~new_new_n8221__;
  assign new_new_n8224__ = ~new_new_n8222__ & ~new_new_n8223__;
  assign new_new_n8225__ = ~pi083 & ~new_new_n8224__;
  assign new_new_n8226__ = pi083 & new_new_n8224__;
  assign new_new_n8227__ = ~new_new_n8006__ & po027;
  assign new_new_n8228__ = pi081 & ~po027;
  assign new_new_n8229__ = ~new_new_n8227__ & ~new_new_n8228__;
  assign new_new_n8230__ = ~new_new_n7813__ & ~new_new_n7814__;
  assign new_new_n8231__ = ~new_new_n8229__ & new_new_n8230__;
  assign new_new_n8232__ = new_new_n8229__ & ~new_new_n8230__;
  assign new_new_n8233__ = ~new_new_n8231__ & ~new_new_n8232__;
  assign new_new_n8234__ = ~pi082 & ~new_new_n8233__;
  assign new_new_n8235__ = pi082 & new_new_n8233__;
  assign new_new_n8236__ = ~pi080 & ~new_new_n8004__;
  assign new_new_n8237__ = pi080 & new_new_n8004__;
  assign new_new_n8238__ = ~new_new_n8236__ & ~new_new_n8237__;
  assign new_new_n8239__ = po027 & ~new_new_n8238__;
  assign new_new_n8240__ = new_new_n7821__ & new_new_n8239__;
  assign new_new_n8241__ = ~new_new_n7821__ & ~new_new_n8239__;
  assign new_new_n8242__ = ~new_new_n8240__ & ~new_new_n8241__;
  assign new_new_n8243__ = pi081 & ~new_new_n8242__;
  assign new_new_n8244__ = ~pi081 & new_new_n8242__;
  assign new_new_n8245__ = ~pi079 & ~new_new_n8002__;
  assign new_new_n8246__ = pi079 & new_new_n8002__;
  assign new_new_n8247__ = ~new_new_n8245__ & ~new_new_n8246__;
  assign new_new_n8248__ = po027 & ~new_new_n8247__;
  assign new_new_n8249__ = new_new_n7830__ & new_new_n8248__;
  assign new_new_n8250__ = ~new_new_n7830__ & ~new_new_n8248__;
  assign new_new_n8251__ = ~new_new_n8249__ & ~new_new_n8250__;
  assign new_new_n8252__ = pi080 & ~new_new_n8251__;
  assign new_new_n8253__ = ~pi080 & new_new_n8251__;
  assign new_new_n8254__ = pi078 & ~new_new_n8000__;
  assign new_new_n8255__ = ~pi078 & new_new_n8000__;
  assign new_new_n8256__ = ~new_new_n8254__ & ~new_new_n8255__;
  assign new_new_n8257__ = po027 & new_new_n8256__;
  assign new_new_n8258__ = new_new_n7839__ & new_new_n8257__;
  assign new_new_n8259__ = ~new_new_n7839__ & ~new_new_n8257__;
  assign new_new_n8260__ = ~new_new_n8258__ & ~new_new_n8259__;
  assign new_new_n8261__ = pi079 & ~new_new_n8260__;
  assign new_new_n8262__ = ~pi079 & new_new_n8260__;
  assign new_new_n8263__ = pi077 & ~new_new_n7998__;
  assign new_new_n8264__ = ~pi077 & new_new_n7998__;
  assign new_new_n8265__ = ~new_new_n8263__ & ~new_new_n8264__;
  assign new_new_n8266__ = po027 & new_new_n8265__;
  assign new_new_n8267__ = new_new_n7848__ & new_new_n8266__;
  assign new_new_n8268__ = ~new_new_n7848__ & ~new_new_n8266__;
  assign new_new_n8269__ = ~new_new_n8267__ & ~new_new_n8268__;
  assign new_new_n8270__ = pi078 & ~new_new_n8269__;
  assign new_new_n8271__ = ~pi078 & new_new_n8269__;
  assign new_new_n8272__ = ~new_new_n7858__ & ~new_new_n7859__;
  assign new_new_n8273__ = ~new_new_n7996__ & po027;
  assign new_new_n8274__ = pi076 & ~po027;
  assign new_new_n8275__ = ~new_new_n8273__ & ~new_new_n8274__;
  assign new_new_n8276__ = new_new_n8272__ & ~new_new_n8275__;
  assign new_new_n8277__ = ~new_new_n8272__ & new_new_n8275__;
  assign new_new_n8278__ = ~new_new_n8276__ & ~new_new_n8277__;
  assign new_new_n8279__ = ~pi077 & ~new_new_n8278__;
  assign new_new_n8280__ = pi077 & new_new_n8278__;
  assign new_new_n8281__ = ~new_new_n7867__ & ~new_new_n7868__;
  assign new_new_n8282__ = ~new_new_n7994__ & po027;
  assign new_new_n8283__ = ~pi075 & ~po027;
  assign new_new_n8284__ = ~new_new_n8282__ & ~new_new_n8283__;
  assign new_new_n8285__ = new_new_n8281__ & ~new_new_n8284__;
  assign new_new_n8286__ = ~new_new_n8281__ & new_new_n8284__;
  assign new_new_n8287__ = ~new_new_n8285__ & ~new_new_n8286__;
  assign new_new_n8288__ = pi076 & ~new_new_n8287__;
  assign new_new_n8289__ = ~pi076 & new_new_n8287__;
  assign new_new_n8290__ = ~new_new_n7876__ & ~new_new_n7877__;
  assign new_new_n8291__ = ~new_new_n7992__ & po027;
  assign new_new_n8292__ = ~pi074 & ~po027;
  assign new_new_n8293__ = ~new_new_n8291__ & ~new_new_n8292__;
  assign new_new_n8294__ = new_new_n8290__ & ~new_new_n8293__;
  assign new_new_n8295__ = ~new_new_n8290__ & new_new_n8293__;
  assign new_new_n8296__ = ~new_new_n8294__ & ~new_new_n8295__;
  assign new_new_n8297__ = pi075 & ~new_new_n8296__;
  assign new_new_n8298__ = ~pi075 & new_new_n8296__;
  assign new_new_n8299__ = ~new_new_n7885__ & ~new_new_n7886__;
  assign new_new_n8300__ = ~new_new_n7990__ & po027;
  assign new_new_n8301__ = ~pi073 & ~po027;
  assign new_new_n8302__ = ~new_new_n8300__ & ~new_new_n8301__;
  assign new_new_n8303__ = ~new_new_n8299__ & ~new_new_n8302__;
  assign new_new_n8304__ = new_new_n8299__ & new_new_n8302__;
  assign new_new_n8305__ = ~new_new_n8303__ & ~new_new_n8304__;
  assign new_new_n8306__ = ~pi074 & ~new_new_n8305__;
  assign new_new_n8307__ = pi074 & new_new_n8305__;
  assign new_new_n8308__ = ~new_new_n7894__ & ~new_new_n7895__;
  assign new_new_n8309__ = ~new_new_n7988__ & po027;
  assign new_new_n8310__ = ~pi072 & ~po027;
  assign new_new_n8311__ = ~new_new_n8309__ & ~new_new_n8310__;
  assign new_new_n8312__ = ~new_new_n8308__ & ~new_new_n8311__;
  assign new_new_n8313__ = new_new_n8308__ & new_new_n8311__;
  assign new_new_n8314__ = ~new_new_n8312__ & ~new_new_n8313__;
  assign new_new_n8315__ = ~pi073 & ~new_new_n8314__;
  assign new_new_n8316__ = pi073 & new_new_n8314__;
  assign new_new_n8317__ = new_new_n7986__ & po027;
  assign new_new_n8318__ = ~pi071 & ~po027;
  assign new_new_n8319__ = ~new_new_n8317__ & ~new_new_n8318__;
  assign new_new_n8320__ = ~new_new_n7903__ & ~new_new_n7904__;
  assign new_new_n8321__ = ~new_new_n8319__ & ~new_new_n8320__;
  assign new_new_n8322__ = new_new_n8319__ & new_new_n8320__;
  assign new_new_n8323__ = ~new_new_n8321__ & ~new_new_n8322__;
  assign new_new_n8324__ = ~pi072 & ~new_new_n8323__;
  assign new_new_n8325__ = pi072 & new_new_n8323__;
  assign new_new_n8326__ = ~new_new_n7976__ & ~new_new_n7977__;
  assign new_new_n8327__ = po027 & new_new_n8326__;
  assign new_new_n8328__ = new_new_n7984__ & new_new_n8327__;
  assign new_new_n8329__ = ~new_new_n7984__ & ~new_new_n8327__;
  assign new_new_n8330__ = ~new_new_n8328__ & ~new_new_n8329__;
  assign new_new_n8331__ = pi071 & new_new_n8330__;
  assign new_new_n8332__ = ~pi071 & ~new_new_n8330__;
  assign new_new_n8333__ = pi068 & ~new_new_n7970__;
  assign new_new_n8334__ = ~pi068 & new_new_n7970__;
  assign new_new_n8335__ = ~new_new_n8333__ & ~new_new_n8334__;
  assign new_new_n8336__ = po027 & new_new_n8335__;
  assign new_new_n8337__ = ~new_new_n7917__ & ~new_new_n8336__;
  assign new_new_n8338__ = new_new_n7917__ & new_new_n8336__;
  assign new_new_n8339__ = ~new_new_n8337__ & ~new_new_n8338__;
  assign new_new_n8340__ = pi069 & ~new_new_n8339__;
  assign new_new_n8341__ = ~pi069 & new_new_n8339__;
  assign new_new_n8342__ = ~new_new_n7939__ & po027;
  assign new_new_n8343__ = ~new_new_n7966__ & new_new_n8342__;
  assign new_new_n8344__ = new_new_n7965__ & ~new_new_n8343__;
  assign new_new_n8345__ = new_new_n7967__ & new_new_n8342__;
  assign new_new_n8346__ = ~new_new_n8344__ & ~new_new_n8345__;
  assign new_new_n8347__ = ~pi067 & ~new_new_n8346__;
  assign new_new_n8348__ = pi067 & new_new_n8346__;
  assign new_new_n8349__ = pi027 & po027;
  assign new_new_n8350__ = ~pi027 & ~po027;
  assign new_new_n8351__ = ~pi065 & ~new_new_n8349__;
  assign new_new_n8352__ = ~new_new_n8350__ & new_new_n8351__;
  assign new_new_n8353__ = ~pi026 & ~new_new_n8352__;
  assign new_new_n8354__ = pi065 & new_new_n8349__;
  assign new_new_n8355__ = ~new_new_n8353__ & ~new_new_n8354__;
  assign new_new_n8356__ = pi064 & ~new_new_n8355__;
  assign new_new_n8357__ = pi064 & po027;
  assign new_new_n8358__ = ~pi027 & pi065;
  assign new_new_n8359__ = ~new_new_n8357__ & new_new_n8358__;
  assign new_new_n8360__ = ~new_new_n8356__ & ~new_new_n8359__;
  assign new_new_n8361__ = pi066 & ~new_new_n8360__;
  assign new_new_n8362__ = new_new_n426__ & ~po028;
  assign new_new_n8363__ = new_new_n7958__ & po027;
  assign new_new_n8364__ = ~new_new_n8362__ & ~new_new_n8363__;
  assign new_new_n8365__ = ~pi027 & ~new_new_n8364__;
  assign new_new_n8366__ = ~new_new_n332__ & po027;
  assign new_new_n8367__ = ~new_new_n7935__ & ~new_new_n8366__;
  assign new_new_n8368__ = pi065 & po027;
  assign new_new_n8369__ = po028 & ~new_new_n8368__;
  assign new_new_n8370__ = pi065 & ~new_new_n7935__;
  assign new_new_n8371__ = pi027 & ~new_new_n8370__;
  assign new_new_n8372__ = ~new_new_n8369__ & new_new_n8371__;
  assign new_new_n8373__ = ~new_new_n8365__ & ~new_new_n8367__;
  assign new_new_n8374__ = ~new_new_n8372__ & new_new_n8373__;
  assign new_new_n8375__ = ~pi028 & ~new_new_n8374__;
  assign new_new_n8376__ = ~pi064 & ~new_new_n8368__;
  assign new_new_n8377__ = ~pi065 & po027;
  assign new_new_n8378__ = ~po028 & ~new_new_n8377__;
  assign new_new_n8379__ = ~new_new_n8349__ & ~new_new_n8363__;
  assign new_new_n8380__ = ~new_new_n8378__ & new_new_n8379__;
  assign new_new_n8381__ = pi064 & ~new_new_n8380__;
  assign new_new_n8382__ = ~new_new_n8376__ & ~new_new_n8381__;
  assign new_new_n8383__ = ~new_new_n7935__ & ~new_new_n8368__;
  assign new_new_n8384__ = pi027 & ~new_new_n7946__;
  assign new_new_n8385__ = ~new_new_n8383__ & new_new_n8384__;
  assign new_new_n8386__ = ~new_new_n8382__ & ~new_new_n8385__;
  assign new_new_n8387__ = pi028 & ~new_new_n8386__;
  assign new_new_n8388__ = ~new_new_n8375__ & ~new_new_n8387__;
  assign new_new_n8389__ = ~pi066 & new_new_n8360__;
  assign new_new_n8390__ = ~new_new_n8388__ & ~new_new_n8389__;
  assign new_new_n8391__ = ~new_new_n8361__ & ~new_new_n8390__;
  assign new_new_n8392__ = ~new_new_n8348__ & new_new_n8391__;
  assign new_new_n8393__ = ~new_new_n8347__ & ~new_new_n8392__;
  assign new_new_n8394__ = ~pi068 & ~new_new_n8393__;
  assign new_new_n8395__ = pi068 & new_new_n8393__;
  assign new_new_n8396__ = ~pi067 & ~new_new_n7968__;
  assign new_new_n8397__ = pi067 & new_new_n7968__;
  assign new_new_n8398__ = ~new_new_n8396__ & ~new_new_n8397__;
  assign new_new_n8399__ = po027 & ~new_new_n8398__;
  assign new_new_n8400__ = new_new_n7924__ & new_new_n8399__;
  assign new_new_n8401__ = ~new_new_n7924__ & ~new_new_n8399__;
  assign new_new_n8402__ = ~new_new_n8400__ & ~new_new_n8401__;
  assign new_new_n8403__ = ~new_new_n8395__ & new_new_n8402__;
  assign new_new_n8404__ = ~new_new_n8394__ & ~new_new_n8403__;
  assign new_new_n8405__ = ~new_new_n8341__ & new_new_n8404__;
  assign new_new_n8406__ = ~new_new_n8340__ & ~new_new_n8405__;
  assign new_new_n8407__ = ~pi070 & new_new_n8406__;
  assign new_new_n8408__ = ~new_new_n7912__ & ~new_new_n7974__;
  assign new_new_n8409__ = ~new_new_n7972__ & po027;
  assign new_new_n8410__ = pi069 & ~po027;
  assign new_new_n8411__ = ~new_new_n8409__ & ~new_new_n8410__;
  assign new_new_n8412__ = new_new_n8408__ & new_new_n8411__;
  assign new_new_n8413__ = ~new_new_n8408__ & ~new_new_n8411__;
  assign new_new_n8414__ = ~new_new_n8412__ & ~new_new_n8413__;
  assign new_new_n8415__ = ~new_new_n8407__ & ~new_new_n8414__;
  assign new_new_n8416__ = pi070 & ~new_new_n8406__;
  assign new_new_n8417__ = ~new_new_n8415__ & ~new_new_n8416__;
  assign new_new_n8418__ = ~new_new_n8332__ & ~new_new_n8417__;
  assign new_new_n8419__ = ~new_new_n8331__ & ~new_new_n8418__;
  assign new_new_n8420__ = ~new_new_n8325__ & new_new_n8419__;
  assign new_new_n8421__ = ~new_new_n8324__ & ~new_new_n8420__;
  assign new_new_n8422__ = ~new_new_n8316__ & ~new_new_n8421__;
  assign new_new_n8423__ = ~new_new_n8315__ & ~new_new_n8422__;
  assign new_new_n8424__ = ~new_new_n8307__ & ~new_new_n8423__;
  assign new_new_n8425__ = ~new_new_n8306__ & ~new_new_n8424__;
  assign new_new_n8426__ = ~new_new_n8298__ & new_new_n8425__;
  assign new_new_n8427__ = ~new_new_n8297__ & ~new_new_n8426__;
  assign new_new_n8428__ = ~new_new_n8289__ & ~new_new_n8427__;
  assign new_new_n8429__ = ~new_new_n8288__ & ~new_new_n8428__;
  assign new_new_n8430__ = ~new_new_n8280__ & new_new_n8429__;
  assign new_new_n8431__ = ~new_new_n8279__ & ~new_new_n8430__;
  assign new_new_n8432__ = ~new_new_n8271__ & new_new_n8431__;
  assign new_new_n8433__ = ~new_new_n8270__ & ~new_new_n8432__;
  assign new_new_n8434__ = ~new_new_n8262__ & ~new_new_n8433__;
  assign new_new_n8435__ = ~new_new_n8261__ & ~new_new_n8434__;
  assign new_new_n8436__ = ~new_new_n8253__ & ~new_new_n8435__;
  assign new_new_n8437__ = ~new_new_n8252__ & ~new_new_n8436__;
  assign new_new_n8438__ = ~new_new_n8244__ & ~new_new_n8437__;
  assign new_new_n8439__ = ~new_new_n8243__ & ~new_new_n8438__;
  assign new_new_n8440__ = ~new_new_n8235__ & new_new_n8439__;
  assign new_new_n8441__ = ~new_new_n8234__ & ~new_new_n8440__;
  assign new_new_n8442__ = ~new_new_n8226__ & ~new_new_n8441__;
  assign new_new_n8443__ = ~new_new_n8225__ & ~new_new_n8442__;
  assign new_new_n8444__ = ~new_new_n8217__ & ~new_new_n8443__;
  assign new_new_n8445__ = ~new_new_n8216__ & ~new_new_n8444__;
  assign new_new_n8446__ = ~new_new_n8208__ & ~new_new_n8445__;
  assign new_new_n8447__ = ~new_new_n8207__ & ~new_new_n8446__;
  assign new_new_n8448__ = ~new_new_n8199__ & ~new_new_n8447__;
  assign new_new_n8449__ = ~new_new_n8198__ & ~new_new_n8448__;
  assign new_new_n8450__ = ~new_new_n8190__ & new_new_n8449__;
  assign new_new_n8451__ = ~new_new_n8189__ & ~new_new_n8450__;
  assign new_new_n8452__ = ~new_new_n8181__ & ~new_new_n8451__;
  assign new_new_n8453__ = ~new_new_n8180__ & ~new_new_n8452__;
  assign new_new_n8454__ = ~new_new_n8172__ & ~new_new_n8453__;
  assign new_new_n8455__ = ~new_new_n8171__ & ~new_new_n8454__;
  assign new_new_n8456__ = ~new_new_n8163__ & ~new_new_n8455__;
  assign new_new_n8457__ = ~new_new_n8162__ & ~new_new_n8456__;
  assign new_new_n8458__ = ~new_new_n8154__ & ~new_new_n8457__;
  assign new_new_n8459__ = ~new_new_n8153__ & ~new_new_n8458__;
  assign new_new_n8460__ = ~new_new_n8145__ & ~new_new_n8459__;
  assign new_new_n8461__ = ~new_new_n8144__ & ~new_new_n8460__;
  assign new_new_n8462__ = ~new_new_n8136__ & new_new_n8461__;
  assign new_new_n8463__ = ~new_new_n8135__ & ~new_new_n8462__;
  assign new_new_n8464__ = ~new_new_n8127__ & ~new_new_n8463__;
  assign new_new_n8465__ = ~new_new_n8126__ & ~new_new_n8464__;
  assign new_new_n8466__ = ~new_new_n8118__ & ~new_new_n8465__;
  assign new_new_n8467__ = ~new_new_n8117__ & ~new_new_n8466__;
  assign new_new_n8468__ = ~new_new_n8109__ & ~new_new_n8467__;
  assign new_new_n8469__ = ~new_new_n8108__ & ~new_new_n8468__;
  assign new_new_n8470__ = ~new_new_n8100__ & ~new_new_n8469__;
  assign new_new_n8471__ = ~new_new_n8099__ & ~new_new_n8470__;
  assign new_new_n8472__ = ~new_new_n8091__ & ~new_new_n8471__;
  assign new_new_n8473__ = ~new_new_n8090__ & ~new_new_n8472__;
  assign new_new_n8474__ = ~new_new_n8082__ & new_new_n8473__;
  assign new_new_n8475__ = ~new_new_n8081__ & ~new_new_n8474__;
  assign new_new_n8476__ = ~pi100 & new_new_n8475__;
  assign new_new_n8477__ = pi100 & ~new_new_n8475__;
  assign new_new_n8478__ = ~new_new_n8476__ & ~new_new_n8477__;
  assign new_new_n8479__ = pi101 & new_new_n8064__;
  assign new_new_n8480__ = new_new_n284__ & ~new_new_n8479__;
  assign new_new_n8481__ = new_new_n8478__ & new_new_n8480__;
  assign new_new_n8482__ = new_new_n8075__ & ~new_new_n8481__;
  assign new_new_n8483__ = pi101 & ~new_new_n8482__;
  assign new_new_n8484__ = ~pi101 & ~new_new_n8064__;
  assign new_new_n8485__ = new_new_n284__ & ~new_new_n8075__;
  assign new_new_n8486__ = new_new_n8484__ & new_new_n8485__;
  assign new_new_n8487__ = new_new_n8478__ & new_new_n8486__;
  assign new_new_n8488__ = ~new_new_n8482__ & ~new_new_n8487__;
  assign new_new_n8489__ = ~pi101 & ~new_new_n8488__;
  assign new_new_n8490__ = ~new_new_n8075__ & ~new_new_n8476__;
  assign new_new_n8491__ = ~new_new_n8477__ & ~new_new_n8479__;
  assign new_new_n8492__ = ~new_new_n8490__ & new_new_n8491__;
  assign new_new_n8493__ = ~new_new_n8484__ & ~new_new_n8492__;
  assign po026 = new_new_n284__ & ~new_new_n8493__;
  assign new_new_n8495__ = new_new_n8473__ & po026;
  assign new_new_n8496__ = pi099 & ~po026;
  assign new_new_n8497__ = ~new_new_n8495__ & ~new_new_n8496__;
  assign new_new_n8498__ = ~new_new_n8081__ & ~new_new_n8082__;
  assign new_new_n8499__ = ~new_new_n8497__ & ~new_new_n8498__;
  assign new_new_n8500__ = new_new_n8497__ & new_new_n8498__;
  assign new_new_n8501__ = ~new_new_n8499__ & ~new_new_n8500__;
  assign new_new_n8502__ = ~pi100 & new_new_n8501__;
  assign new_new_n8503__ = pi100 & ~new_new_n8501__;
  assign new_new_n8504__ = ~pi098 & ~new_new_n8471__;
  assign new_new_n8505__ = pi098 & new_new_n8471__;
  assign new_new_n8506__ = ~new_new_n8504__ & ~new_new_n8505__;
  assign new_new_n8507__ = po026 & new_new_n8506__;
  assign new_new_n8508__ = new_new_n8089__ & new_new_n8507__;
  assign new_new_n8509__ = ~new_new_n8089__ & ~new_new_n8507__;
  assign new_new_n8510__ = ~new_new_n8508__ & ~new_new_n8509__;
  assign new_new_n8511__ = ~pi099 & ~new_new_n8510__;
  assign new_new_n8512__ = pi099 & new_new_n8510__;
  assign new_new_n8513__ = ~pi097 & ~new_new_n8469__;
  assign new_new_n8514__ = pi097 & new_new_n8469__;
  assign new_new_n8515__ = ~new_new_n8513__ & ~new_new_n8514__;
  assign new_new_n8516__ = po026 & new_new_n8515__;
  assign new_new_n8517__ = new_new_n8098__ & new_new_n8516__;
  assign new_new_n8518__ = ~new_new_n8098__ & ~new_new_n8516__;
  assign new_new_n8519__ = ~new_new_n8517__ & ~new_new_n8518__;
  assign new_new_n8520__ = ~pi098 & ~new_new_n8519__;
  assign new_new_n8521__ = pi098 & new_new_n8519__;
  assign new_new_n8522__ = ~new_new_n8108__ & ~new_new_n8109__;
  assign new_new_n8523__ = ~new_new_n8467__ & po026;
  assign new_new_n8524__ = ~pi096 & ~po026;
  assign new_new_n8525__ = ~new_new_n8523__ & ~new_new_n8524__;
  assign new_new_n8526__ = new_new_n8522__ & ~new_new_n8525__;
  assign new_new_n8527__ = ~new_new_n8522__ & new_new_n8525__;
  assign new_new_n8528__ = ~new_new_n8526__ & ~new_new_n8527__;
  assign new_new_n8529__ = ~pi097 & new_new_n8528__;
  assign new_new_n8530__ = pi097 & ~new_new_n8528__;
  assign new_new_n8531__ = ~pi094 & ~new_new_n8463__;
  assign new_new_n8532__ = pi094 & new_new_n8463__;
  assign new_new_n8533__ = ~new_new_n8531__ & ~new_new_n8532__;
  assign new_new_n8534__ = po026 & new_new_n8533__;
  assign new_new_n8535__ = new_new_n8125__ & new_new_n8534__;
  assign new_new_n8536__ = ~new_new_n8125__ & ~new_new_n8534__;
  assign new_new_n8537__ = ~new_new_n8535__ & ~new_new_n8536__;
  assign new_new_n8538__ = ~pi095 & ~new_new_n8537__;
  assign new_new_n8539__ = pi095 & new_new_n8537__;
  assign new_new_n8540__ = ~new_new_n8135__ & ~new_new_n8136__;
  assign new_new_n8541__ = ~new_new_n8461__ & po026;
  assign new_new_n8542__ = pi093 & ~po026;
  assign new_new_n8543__ = ~new_new_n8541__ & ~new_new_n8542__;
  assign new_new_n8544__ = new_new_n8540__ & ~new_new_n8543__;
  assign new_new_n8545__ = ~new_new_n8540__ & new_new_n8543__;
  assign new_new_n8546__ = ~new_new_n8544__ & ~new_new_n8545__;
  assign new_new_n8547__ = ~pi094 & ~new_new_n8546__;
  assign new_new_n8548__ = pi094 & new_new_n8546__;
  assign new_new_n8549__ = ~new_new_n8144__ & ~new_new_n8145__;
  assign new_new_n8550__ = ~new_new_n8459__ & po026;
  assign new_new_n8551__ = pi092 & ~po026;
  assign new_new_n8552__ = ~new_new_n8550__ & ~new_new_n8551__;
  assign new_new_n8553__ = new_new_n8549__ & ~new_new_n8552__;
  assign new_new_n8554__ = ~new_new_n8549__ & new_new_n8552__;
  assign new_new_n8555__ = ~new_new_n8553__ & ~new_new_n8554__;
  assign new_new_n8556__ = ~pi093 & ~new_new_n8555__;
  assign new_new_n8557__ = pi093 & new_new_n8555__;
  assign new_new_n8558__ = ~new_new_n8457__ & po026;
  assign new_new_n8559__ = pi091 & ~po026;
  assign new_new_n8560__ = ~new_new_n8558__ & ~new_new_n8559__;
  assign new_new_n8561__ = ~new_new_n8153__ & ~new_new_n8154__;
  assign new_new_n8562__ = ~new_new_n8560__ & new_new_n8561__;
  assign new_new_n8563__ = new_new_n8560__ & ~new_new_n8561__;
  assign new_new_n8564__ = ~new_new_n8562__ & ~new_new_n8563__;
  assign new_new_n8565__ = ~pi092 & ~new_new_n8564__;
  assign new_new_n8566__ = pi092 & new_new_n8564__;
  assign new_new_n8567__ = ~new_new_n8162__ & ~new_new_n8163__;
  assign new_new_n8568__ = new_new_n8455__ & po026;
  assign new_new_n8569__ = ~pi090 & ~po026;
  assign new_new_n8570__ = ~new_new_n8568__ & ~new_new_n8569__;
  assign new_new_n8571__ = ~new_new_n8567__ & ~new_new_n8570__;
  assign new_new_n8572__ = new_new_n8567__ & new_new_n8570__;
  assign new_new_n8573__ = ~new_new_n8571__ & ~new_new_n8572__;
  assign new_new_n8574__ = ~pi091 & ~new_new_n8573__;
  assign new_new_n8575__ = pi091 & new_new_n8573__;
  assign new_new_n8576__ = pi089 & ~new_new_n8453__;
  assign new_new_n8577__ = ~pi089 & new_new_n8453__;
  assign new_new_n8578__ = ~new_new_n8576__ & ~new_new_n8577__;
  assign new_new_n8579__ = po026 & new_new_n8578__;
  assign new_new_n8580__ = new_new_n8170__ & new_new_n8579__;
  assign new_new_n8581__ = ~new_new_n8170__ & ~new_new_n8579__;
  assign new_new_n8582__ = ~new_new_n8580__ & ~new_new_n8581__;
  assign new_new_n8583__ = pi090 & ~new_new_n8582__;
  assign new_new_n8584__ = ~pi090 & new_new_n8582__;
  assign new_new_n8585__ = pi088 & ~new_new_n8451__;
  assign new_new_n8586__ = ~pi088 & new_new_n8451__;
  assign new_new_n8587__ = ~new_new_n8585__ & ~new_new_n8586__;
  assign new_new_n8588__ = po026 & new_new_n8587__;
  assign new_new_n8589__ = new_new_n8179__ & new_new_n8588__;
  assign new_new_n8590__ = ~new_new_n8179__ & ~new_new_n8588__;
  assign new_new_n8591__ = ~new_new_n8589__ & ~new_new_n8590__;
  assign new_new_n8592__ = pi089 & ~new_new_n8591__;
  assign new_new_n8593__ = ~pi089 & new_new_n8591__;
  assign new_new_n8594__ = ~new_new_n8189__ & ~new_new_n8190__;
  assign new_new_n8595__ = ~new_new_n8449__ & po026;
  assign new_new_n8596__ = ~pi087 & ~po026;
  assign new_new_n8597__ = ~new_new_n8595__ & ~new_new_n8596__;
  assign new_new_n8598__ = new_new_n8594__ & new_new_n8597__;
  assign new_new_n8599__ = ~new_new_n8594__ & ~new_new_n8597__;
  assign new_new_n8600__ = ~new_new_n8598__ & ~new_new_n8599__;
  assign new_new_n8601__ = ~pi088 & ~new_new_n8600__;
  assign new_new_n8602__ = pi088 & new_new_n8600__;
  assign new_new_n8603__ = ~pi086 & ~new_new_n8447__;
  assign new_new_n8604__ = pi086 & new_new_n8447__;
  assign new_new_n8605__ = ~new_new_n8603__ & ~new_new_n8604__;
  assign new_new_n8606__ = po026 & new_new_n8605__;
  assign new_new_n8607__ = new_new_n8197__ & new_new_n8606__;
  assign new_new_n8608__ = ~new_new_n8197__ & ~new_new_n8606__;
  assign new_new_n8609__ = ~new_new_n8607__ & ~new_new_n8608__;
  assign new_new_n8610__ = pi087 & new_new_n8609__;
  assign new_new_n8611__ = ~pi087 & ~new_new_n8609__;
  assign new_new_n8612__ = ~pi085 & ~new_new_n8445__;
  assign new_new_n8613__ = pi085 & new_new_n8445__;
  assign new_new_n8614__ = ~new_new_n8612__ & ~new_new_n8613__;
  assign new_new_n8615__ = po026 & new_new_n8614__;
  assign new_new_n8616__ = new_new_n8206__ & ~new_new_n8615__;
  assign new_new_n8617__ = ~new_new_n8206__ & new_new_n8615__;
  assign new_new_n8618__ = ~new_new_n8616__ & ~new_new_n8617__;
  assign new_new_n8619__ = pi086 & ~new_new_n8618__;
  assign new_new_n8620__ = ~pi086 & new_new_n8618__;
  assign new_new_n8621__ = ~new_new_n8216__ & ~new_new_n8217__;
  assign new_new_n8622__ = ~new_new_n8443__ & po026;
  assign new_new_n8623__ = ~pi084 & ~po026;
  assign new_new_n8624__ = ~new_new_n8622__ & ~new_new_n8623__;
  assign new_new_n8625__ = new_new_n8621__ & ~new_new_n8624__;
  assign new_new_n8626__ = ~new_new_n8621__ & new_new_n8624__;
  assign new_new_n8627__ = ~new_new_n8625__ & ~new_new_n8626__;
  assign new_new_n8628__ = pi085 & ~new_new_n8627__;
  assign new_new_n8629__ = ~pi083 & ~new_new_n8441__;
  assign new_new_n8630__ = pi083 & new_new_n8441__;
  assign new_new_n8631__ = ~new_new_n8629__ & ~new_new_n8630__;
  assign new_new_n8632__ = po026 & new_new_n8631__;
  assign new_new_n8633__ = new_new_n8224__ & new_new_n8632__;
  assign new_new_n8634__ = ~new_new_n8224__ & ~new_new_n8632__;
  assign new_new_n8635__ = ~new_new_n8633__ & ~new_new_n8634__;
  assign new_new_n8636__ = ~pi084 & ~new_new_n8635__;
  assign new_new_n8637__ = pi084 & new_new_n8635__;
  assign new_new_n8638__ = ~new_new_n8439__ & po026;
  assign new_new_n8639__ = pi082 & ~po026;
  assign new_new_n8640__ = ~new_new_n8638__ & ~new_new_n8639__;
  assign new_new_n8641__ = ~new_new_n8234__ & ~new_new_n8235__;
  assign new_new_n8642__ = ~new_new_n8640__ & new_new_n8641__;
  assign new_new_n8643__ = new_new_n8640__ & ~new_new_n8641__;
  assign new_new_n8644__ = ~new_new_n8642__ & ~new_new_n8643__;
  assign new_new_n8645__ = ~pi083 & ~new_new_n8644__;
  assign new_new_n8646__ = pi083 & new_new_n8644__;
  assign new_new_n8647__ = ~pi081 & ~new_new_n8437__;
  assign new_new_n8648__ = pi081 & new_new_n8437__;
  assign new_new_n8649__ = ~new_new_n8647__ & ~new_new_n8648__;
  assign new_new_n8650__ = po026 & ~new_new_n8649__;
  assign new_new_n8651__ = new_new_n8242__ & ~new_new_n8650__;
  assign new_new_n8652__ = ~new_new_n8242__ & new_new_n8650__;
  assign new_new_n8653__ = ~new_new_n8651__ & ~new_new_n8652__;
  assign new_new_n8654__ = ~pi082 & ~new_new_n8653__;
  assign new_new_n8655__ = pi082 & new_new_n8653__;
  assign new_new_n8656__ = pi080 & ~new_new_n8435__;
  assign new_new_n8657__ = ~pi080 & new_new_n8435__;
  assign new_new_n8658__ = ~new_new_n8656__ & ~new_new_n8657__;
  assign new_new_n8659__ = po026 & new_new_n8658__;
  assign new_new_n8660__ = ~new_new_n8251__ & new_new_n8659__;
  assign new_new_n8661__ = new_new_n8251__ & ~new_new_n8659__;
  assign new_new_n8662__ = ~new_new_n8660__ & ~new_new_n8661__;
  assign new_new_n8663__ = ~pi081 & ~new_new_n8662__;
  assign new_new_n8664__ = pi081 & new_new_n8662__;
  assign new_new_n8665__ = pi079 & ~new_new_n8433__;
  assign new_new_n8666__ = ~pi079 & new_new_n8433__;
  assign new_new_n8667__ = ~new_new_n8665__ & ~new_new_n8666__;
  assign new_new_n8668__ = po026 & new_new_n8667__;
  assign new_new_n8669__ = new_new_n8260__ & ~new_new_n8668__;
  assign new_new_n8670__ = ~new_new_n8260__ & new_new_n8668__;
  assign new_new_n8671__ = ~new_new_n8669__ & ~new_new_n8670__;
  assign new_new_n8672__ = ~pi080 & ~new_new_n8671__;
  assign new_new_n8673__ = pi080 & new_new_n8671__;
  assign new_new_n8674__ = ~new_new_n8270__ & ~new_new_n8271__;
  assign new_new_n8675__ = ~new_new_n8431__ & po026;
  assign new_new_n8676__ = ~pi078 & ~po026;
  assign new_new_n8677__ = ~new_new_n8675__ & ~new_new_n8676__;
  assign new_new_n8678__ = new_new_n8674__ & ~new_new_n8677__;
  assign new_new_n8679__ = ~new_new_n8674__ & new_new_n8677__;
  assign new_new_n8680__ = ~new_new_n8678__ & ~new_new_n8679__;
  assign new_new_n8681__ = ~pi079 & new_new_n8680__;
  assign new_new_n8682__ = pi079 & ~new_new_n8680__;
  assign new_new_n8683__ = ~new_new_n8429__ & po026;
  assign new_new_n8684__ = pi077 & ~po026;
  assign new_new_n8685__ = ~new_new_n8683__ & ~new_new_n8684__;
  assign new_new_n8686__ = ~new_new_n8279__ & ~new_new_n8280__;
  assign new_new_n8687__ = ~new_new_n8685__ & new_new_n8686__;
  assign new_new_n8688__ = new_new_n8685__ & ~new_new_n8686__;
  assign new_new_n8689__ = ~new_new_n8687__ & ~new_new_n8688__;
  assign new_new_n8690__ = ~pi078 & ~new_new_n8689__;
  assign new_new_n8691__ = pi078 & new_new_n8689__;
  assign new_new_n8692__ = ~new_new_n8288__ & ~new_new_n8289__;
  assign new_new_n8693__ = ~new_new_n8427__ & po026;
  assign new_new_n8694__ = pi076 & ~po026;
  assign new_new_n8695__ = ~new_new_n8693__ & ~new_new_n8694__;
  assign new_new_n8696__ = new_new_n8692__ & ~new_new_n8695__;
  assign new_new_n8697__ = ~new_new_n8692__ & new_new_n8695__;
  assign new_new_n8698__ = ~new_new_n8696__ & ~new_new_n8697__;
  assign new_new_n8699__ = ~pi077 & ~new_new_n8698__;
  assign new_new_n8700__ = pi077 & new_new_n8698__;
  assign new_new_n8701__ = ~new_new_n8297__ & ~new_new_n8298__;
  assign new_new_n8702__ = ~new_new_n8425__ & po026;
  assign new_new_n8703__ = ~pi075 & ~po026;
  assign new_new_n8704__ = ~new_new_n8702__ & ~new_new_n8703__;
  assign new_new_n8705__ = new_new_n8701__ & ~new_new_n8704__;
  assign new_new_n8706__ = ~new_new_n8701__ & new_new_n8704__;
  assign new_new_n8707__ = ~new_new_n8705__ & ~new_new_n8706__;
  assign new_new_n8708__ = pi076 & ~new_new_n8707__;
  assign new_new_n8709__ = ~pi076 & new_new_n8707__;
  assign new_new_n8710__ = ~pi074 & ~new_new_n8423__;
  assign new_new_n8711__ = pi074 & new_new_n8423__;
  assign new_new_n8712__ = ~new_new_n8710__ & ~new_new_n8711__;
  assign new_new_n8713__ = po026 & new_new_n8712__;
  assign new_new_n8714__ = ~new_new_n8305__ & new_new_n8713__;
  assign new_new_n8715__ = new_new_n8305__ & ~new_new_n8713__;
  assign new_new_n8716__ = ~new_new_n8714__ & ~new_new_n8715__;
  assign new_new_n8717__ = ~pi075 & new_new_n8716__;
  assign new_new_n8718__ = pi075 & ~new_new_n8716__;
  assign new_new_n8719__ = ~pi073 & ~new_new_n8421__;
  assign new_new_n8720__ = pi073 & new_new_n8421__;
  assign new_new_n8721__ = ~new_new_n8719__ & ~new_new_n8720__;
  assign new_new_n8722__ = po026 & new_new_n8721__;
  assign new_new_n8723__ = ~new_new_n8314__ & new_new_n8722__;
  assign new_new_n8724__ = new_new_n8314__ & ~new_new_n8722__;
  assign new_new_n8725__ = ~new_new_n8723__ & ~new_new_n8724__;
  assign new_new_n8726__ = ~pi074 & new_new_n8725__;
  assign new_new_n8727__ = pi074 & ~new_new_n8725__;
  assign new_new_n8728__ = ~new_new_n8324__ & ~new_new_n8325__;
  assign new_new_n8729__ = new_new_n8419__ & po026;
  assign new_new_n8730__ = ~pi072 & ~po026;
  assign new_new_n8731__ = ~new_new_n8729__ & ~new_new_n8730__;
  assign new_new_n8732__ = ~new_new_n8728__ & ~new_new_n8731__;
  assign new_new_n8733__ = new_new_n8728__ & new_new_n8731__;
  assign new_new_n8734__ = ~new_new_n8732__ & ~new_new_n8733__;
  assign new_new_n8735__ = ~pi073 & ~new_new_n8734__;
  assign new_new_n8736__ = pi073 & new_new_n8734__;
  assign new_new_n8737__ = new_new_n8417__ & po026;
  assign new_new_n8738__ = ~pi071 & ~po026;
  assign new_new_n8739__ = ~new_new_n8737__ & ~new_new_n8738__;
  assign new_new_n8740__ = ~new_new_n8331__ & ~new_new_n8332__;
  assign new_new_n8741__ = ~new_new_n8739__ & ~new_new_n8740__;
  assign new_new_n8742__ = new_new_n8739__ & new_new_n8740__;
  assign new_new_n8743__ = ~new_new_n8741__ & ~new_new_n8742__;
  assign new_new_n8744__ = ~pi072 & ~new_new_n8743__;
  assign new_new_n8745__ = pi072 & new_new_n8743__;
  assign new_new_n8746__ = ~new_new_n8407__ & ~new_new_n8416__;
  assign new_new_n8747__ = po026 & new_new_n8746__;
  assign new_new_n8748__ = new_new_n8414__ & new_new_n8747__;
  assign new_new_n8749__ = ~new_new_n8414__ & ~new_new_n8747__;
  assign new_new_n8750__ = ~new_new_n8748__ & ~new_new_n8749__;
  assign new_new_n8751__ = pi071 & ~new_new_n8750__;
  assign new_new_n8752__ = ~pi071 & new_new_n8750__;
  assign new_new_n8753__ = new_new_n8404__ & po026;
  assign new_new_n8754__ = pi069 & ~po026;
  assign new_new_n8755__ = ~new_new_n8753__ & ~new_new_n8754__;
  assign new_new_n8756__ = ~new_new_n8340__ & ~new_new_n8341__;
  assign new_new_n8757__ = ~new_new_n8755__ & ~new_new_n8756__;
  assign new_new_n8758__ = new_new_n8755__ & new_new_n8756__;
  assign new_new_n8759__ = ~new_new_n8757__ & ~new_new_n8758__;
  assign new_new_n8760__ = pi070 & ~new_new_n8759__;
  assign new_new_n8761__ = ~pi070 & new_new_n8759__;
  assign new_new_n8762__ = ~new_new_n8394__ & ~new_new_n8395__;
  assign new_new_n8763__ = po026 & new_new_n8762__;
  assign new_new_n8764__ = new_new_n8402__ & new_new_n8763__;
  assign new_new_n8765__ = ~new_new_n8402__ & ~new_new_n8763__;
  assign new_new_n8766__ = ~new_new_n8764__ & ~new_new_n8765__;
  assign new_new_n8767__ = ~pi069 & new_new_n8766__;
  assign new_new_n8768__ = pi069 & ~new_new_n8766__;
  assign new_new_n8769__ = ~new_new_n8347__ & ~new_new_n8348__;
  assign new_new_n8770__ = new_new_n8391__ & po026;
  assign new_new_n8771__ = ~pi067 & ~po026;
  assign new_new_n8772__ = ~new_new_n8770__ & ~new_new_n8771__;
  assign new_new_n8773__ = ~new_new_n8769__ & ~new_new_n8772__;
  assign new_new_n8774__ = new_new_n8769__ & new_new_n8772__;
  assign new_new_n8775__ = ~new_new_n8773__ & ~new_new_n8774__;
  assign new_new_n8776__ = ~pi068 & ~new_new_n8775__;
  assign new_new_n8777__ = pi068 & new_new_n8775__;
  assign new_new_n8778__ = ~new_new_n8361__ & ~new_new_n8389__;
  assign new_new_n8779__ = po026 & new_new_n8778__;
  assign new_new_n8780__ = new_new_n8388__ & ~new_new_n8779__;
  assign new_new_n8781__ = ~new_new_n8388__ & new_new_n8779__;
  assign new_new_n8782__ = ~new_new_n8780__ & ~new_new_n8781__;
  assign new_new_n8783__ = ~pi067 & ~new_new_n8782__;
  assign new_new_n8784__ = pi067 & new_new_n8782__;
  assign new_new_n8785__ = pi026 & po026;
  assign new_new_n8786__ = pi025 & ~pi065;
  assign new_new_n8787__ = new_new_n8785__ & ~new_new_n8786__;
  assign new_new_n8788__ = ~pi026 & ~po026;
  assign new_new_n8789__ = ~pi065 & ~new_new_n8788__;
  assign new_new_n8790__ = ~pi025 & ~new_new_n8789__;
  assign new_new_n8791__ = ~new_new_n8787__ & ~new_new_n8790__;
  assign new_new_n8792__ = pi064 & ~new_new_n8791__;
  assign new_new_n8793__ = pi064 & po026;
  assign new_new_n8794__ = ~pi026 & pi065;
  assign new_new_n8795__ = ~new_new_n8793__ & new_new_n8794__;
  assign new_new_n8796__ = ~new_new_n8792__ & ~new_new_n8795__;
  assign new_new_n8797__ = pi066 & ~new_new_n8796__;
  assign new_new_n8798__ = new_new_n426__ & ~po027;
  assign new_new_n8799__ = new_new_n8377__ & po026;
  assign new_new_n8800__ = ~new_new_n8798__ & ~new_new_n8799__;
  assign new_new_n8801__ = ~pi026 & ~new_new_n8800__;
  assign new_new_n8802__ = ~new_new_n332__ & po026;
  assign new_new_n8803__ = ~new_new_n8357__ & ~new_new_n8802__;
  assign new_new_n8804__ = pi065 & po026;
  assign new_new_n8805__ = po027 & ~new_new_n8804__;
  assign new_new_n8806__ = pi065 & ~new_new_n8357__;
  assign new_new_n8807__ = pi026 & ~new_new_n8806__;
  assign new_new_n8808__ = ~new_new_n8805__ & new_new_n8807__;
  assign new_new_n8809__ = ~new_new_n8801__ & ~new_new_n8803__;
  assign new_new_n8810__ = ~new_new_n8808__ & new_new_n8809__;
  assign new_new_n8811__ = ~pi027 & ~new_new_n8810__;
  assign new_new_n8812__ = ~new_new_n8357__ & ~new_new_n8804__;
  assign new_new_n8813__ = pi026 & ~new_new_n8368__;
  assign new_new_n8814__ = pi064 & ~new_new_n8813__;
  assign new_new_n8815__ = ~new_new_n8812__ & ~new_new_n8814__;
  assign new_new_n8816__ = ~pi065 & po026;
  assign new_new_n8817__ = ~po027 & ~new_new_n8816__;
  assign new_new_n8818__ = pi064 & ~new_new_n8785__;
  assign new_new_n8819__ = ~new_new_n8799__ & new_new_n8818__;
  assign new_new_n8820__ = ~new_new_n8817__ & new_new_n8819__;
  assign new_new_n8821__ = ~new_new_n8815__ & ~new_new_n8820__;
  assign new_new_n8822__ = pi027 & ~new_new_n8821__;
  assign new_new_n8823__ = ~new_new_n8811__ & ~new_new_n8822__;
  assign new_new_n8824__ = ~pi066 & new_new_n8796__;
  assign new_new_n8825__ = ~new_new_n8823__ & ~new_new_n8824__;
  assign new_new_n8826__ = ~new_new_n8797__ & ~new_new_n8825__;
  assign new_new_n8827__ = ~new_new_n8784__ & new_new_n8826__;
  assign new_new_n8828__ = ~new_new_n8783__ & ~new_new_n8827__;
  assign new_new_n8829__ = ~new_new_n8777__ & ~new_new_n8828__;
  assign new_new_n8830__ = ~new_new_n8776__ & ~new_new_n8829__;
  assign new_new_n8831__ = ~new_new_n8768__ & ~new_new_n8830__;
  assign new_new_n8832__ = ~new_new_n8767__ & ~new_new_n8831__;
  assign new_new_n8833__ = ~new_new_n8761__ & new_new_n8832__;
  assign new_new_n8834__ = ~new_new_n8760__ & ~new_new_n8833__;
  assign new_new_n8835__ = ~new_new_n8752__ & ~new_new_n8834__;
  assign new_new_n8836__ = ~new_new_n8751__ & ~new_new_n8835__;
  assign new_new_n8837__ = ~new_new_n8745__ & new_new_n8836__;
  assign new_new_n8838__ = ~new_new_n8744__ & ~new_new_n8837__;
  assign new_new_n8839__ = ~new_new_n8736__ & ~new_new_n8838__;
  assign new_new_n8840__ = ~new_new_n8735__ & ~new_new_n8839__;
  assign new_new_n8841__ = ~new_new_n8727__ & ~new_new_n8840__;
  assign new_new_n8842__ = ~new_new_n8726__ & ~new_new_n8841__;
  assign new_new_n8843__ = ~new_new_n8718__ & ~new_new_n8842__;
  assign new_new_n8844__ = ~new_new_n8717__ & ~new_new_n8843__;
  assign new_new_n8845__ = ~new_new_n8709__ & new_new_n8844__;
  assign new_new_n8846__ = ~new_new_n8708__ & ~new_new_n8845__;
  assign new_new_n8847__ = ~new_new_n8700__ & new_new_n8846__;
  assign new_new_n8848__ = ~new_new_n8699__ & ~new_new_n8847__;
  assign new_new_n8849__ = ~new_new_n8691__ & ~new_new_n8848__;
  assign new_new_n8850__ = ~new_new_n8690__ & ~new_new_n8849__;
  assign new_new_n8851__ = ~new_new_n8682__ & ~new_new_n8850__;
  assign new_new_n8852__ = ~new_new_n8681__ & ~new_new_n8851__;
  assign new_new_n8853__ = ~new_new_n8673__ & ~new_new_n8852__;
  assign new_new_n8854__ = ~new_new_n8672__ & ~new_new_n8853__;
  assign new_new_n8855__ = ~new_new_n8664__ & ~new_new_n8854__;
  assign new_new_n8856__ = ~new_new_n8663__ & ~new_new_n8855__;
  assign new_new_n8857__ = ~new_new_n8655__ & ~new_new_n8856__;
  assign new_new_n8858__ = ~new_new_n8654__ & ~new_new_n8857__;
  assign new_new_n8859__ = ~new_new_n8646__ & ~new_new_n8858__;
  assign new_new_n8860__ = ~new_new_n8645__ & ~new_new_n8859__;
  assign new_new_n8861__ = ~new_new_n8637__ & ~new_new_n8860__;
  assign new_new_n8862__ = ~new_new_n8636__ & ~new_new_n8861__;
  assign new_new_n8863__ = ~pi085 & new_new_n8627__;
  assign new_new_n8864__ = new_new_n8862__ & ~new_new_n8863__;
  assign new_new_n8865__ = ~new_new_n8628__ & ~new_new_n8864__;
  assign new_new_n8866__ = ~new_new_n8620__ & ~new_new_n8865__;
  assign new_new_n8867__ = ~new_new_n8619__ & ~new_new_n8866__;
  assign new_new_n8868__ = ~new_new_n8611__ & ~new_new_n8867__;
  assign new_new_n8869__ = ~new_new_n8610__ & ~new_new_n8868__;
  assign new_new_n8870__ = ~new_new_n8602__ & new_new_n8869__;
  assign new_new_n8871__ = ~new_new_n8601__ & ~new_new_n8870__;
  assign new_new_n8872__ = ~new_new_n8593__ & new_new_n8871__;
  assign new_new_n8873__ = ~new_new_n8592__ & ~new_new_n8872__;
  assign new_new_n8874__ = ~new_new_n8584__ & ~new_new_n8873__;
  assign new_new_n8875__ = ~new_new_n8583__ & ~new_new_n8874__;
  assign new_new_n8876__ = ~new_new_n8575__ & new_new_n8875__;
  assign new_new_n8877__ = ~new_new_n8574__ & ~new_new_n8876__;
  assign new_new_n8878__ = ~new_new_n8566__ & ~new_new_n8877__;
  assign new_new_n8879__ = ~new_new_n8565__ & ~new_new_n8878__;
  assign new_new_n8880__ = ~new_new_n8557__ & ~new_new_n8879__;
  assign new_new_n8881__ = ~new_new_n8556__ & ~new_new_n8880__;
  assign new_new_n8882__ = ~new_new_n8548__ & ~new_new_n8881__;
  assign new_new_n8883__ = ~new_new_n8547__ & ~new_new_n8882__;
  assign new_new_n8884__ = ~new_new_n8539__ & ~new_new_n8883__;
  assign new_new_n8885__ = ~new_new_n8538__ & ~new_new_n8884__;
  assign new_new_n8886__ = ~pi096 & ~new_new_n8885__;
  assign new_new_n8887__ = pi096 & new_new_n8885__;
  assign new_new_n8888__ = ~pi095 & ~new_new_n8465__;
  assign new_new_n8889__ = pi095 & new_new_n8465__;
  assign new_new_n8890__ = ~new_new_n8888__ & ~new_new_n8889__;
  assign new_new_n8891__ = po026 & new_new_n8890__;
  assign new_new_n8892__ = new_new_n8116__ & new_new_n8891__;
  assign new_new_n8893__ = ~new_new_n8116__ & ~new_new_n8891__;
  assign new_new_n8894__ = ~new_new_n8892__ & ~new_new_n8893__;
  assign new_new_n8895__ = ~new_new_n8887__ & ~new_new_n8894__;
  assign new_new_n8896__ = ~new_new_n8886__ & ~new_new_n8895__;
  assign new_new_n8897__ = ~new_new_n8530__ & ~new_new_n8896__;
  assign new_new_n8898__ = ~new_new_n8529__ & ~new_new_n8897__;
  assign new_new_n8899__ = ~new_new_n8521__ & ~new_new_n8898__;
  assign new_new_n8900__ = ~new_new_n8520__ & ~new_new_n8899__;
  assign new_new_n8901__ = ~new_new_n8512__ & ~new_new_n8900__;
  assign new_new_n8902__ = ~new_new_n8511__ & ~new_new_n8901__;
  assign new_new_n8903__ = ~new_new_n8503__ & ~new_new_n8902__;
  assign new_new_n8904__ = ~new_new_n8502__ & ~new_new_n8903__;
  assign new_new_n8905__ = ~new_new_n8489__ & new_new_n8904__;
  assign new_new_n8906__ = ~new_new_n8483__ & ~new_new_n8905__;
  assign new_new_n8907__ = pi102 & ~new_new_n8906__;
  assign new_new_n8908__ = new_new_n8070__ & ~new_new_n8907__;
  assign new_new_n8909__ = ~new_new_n8064__ & ~new_new_n8908__;
  assign new_new_n8910__ = ~new_new_n376__ & ~new_new_n8909__;
  assign new_new_n8911__ = new_new_n8063__ & ~po026;
  assign new_new_n8912__ = ~new_new_n376__ & ~new_new_n8911__;
  assign new_new_n8913__ = pi102 & new_new_n8912__;
  assign new_new_n8914__ = new_new_n8070__ & ~new_new_n8913__;
  assign new_new_n8915__ = ~pi101 & new_new_n8904__;
  assign new_new_n8916__ = pi101 & ~new_new_n8904__;
  assign new_new_n8917__ = ~new_new_n8915__ & ~new_new_n8916__;
  assign new_new_n8918__ = new_new_n8914__ & ~new_new_n8917__;
  assign new_new_n8919__ = ~new_new_n8488__ & ~new_new_n8918__;
  assign new_new_n8920__ = ~pi102 & ~new_new_n8912__;
  assign new_new_n8921__ = new_new_n8070__ & new_new_n8488__;
  assign new_new_n8922__ = new_new_n8920__ & new_new_n8921__;
  assign new_new_n8923__ = ~new_new_n8917__ & new_new_n8922__;
  assign new_new_n8924__ = ~new_new_n8919__ & ~new_new_n8923__;
  assign new_new_n8925__ = ~pi102 & ~new_new_n8924__;
  assign new_new_n8926__ = ~new_new_n8502__ & ~new_new_n8503__;
  assign new_new_n8927__ = ~new_new_n8906__ & ~new_new_n8920__;
  assign po025 = new_new_n8914__ & ~new_new_n8927__;
  assign new_new_n8929__ = ~new_new_n8902__ & po025;
  assign new_new_n8930__ = ~pi100 & ~po025;
  assign new_new_n8931__ = ~new_new_n8929__ & ~new_new_n8930__;
  assign new_new_n8932__ = new_new_n8926__ & new_new_n8931__;
  assign new_new_n8933__ = ~new_new_n8926__ & ~new_new_n8931__;
  assign new_new_n8934__ = ~new_new_n8932__ & ~new_new_n8933__;
  assign new_new_n8935__ = ~pi101 & ~new_new_n8934__;
  assign new_new_n8936__ = pi101 & new_new_n8934__;
  assign new_new_n8937__ = ~new_new_n8511__ & ~new_new_n8512__;
  assign new_new_n8938__ = ~new_new_n8900__ & po025;
  assign new_new_n8939__ = ~pi099 & ~po025;
  assign new_new_n8940__ = ~new_new_n8938__ & ~new_new_n8939__;
  assign new_new_n8941__ = new_new_n8937__ & ~new_new_n8940__;
  assign new_new_n8942__ = ~new_new_n8937__ & new_new_n8940__;
  assign new_new_n8943__ = ~new_new_n8941__ & ~new_new_n8942__;
  assign new_new_n8944__ = pi100 & ~new_new_n8943__;
  assign new_new_n8945__ = ~pi100 & new_new_n8943__;
  assign new_new_n8946__ = ~pi098 & ~new_new_n8898__;
  assign new_new_n8947__ = pi098 & new_new_n8898__;
  assign new_new_n8948__ = ~new_new_n8946__ & ~new_new_n8947__;
  assign new_new_n8949__ = po025 & new_new_n8948__;
  assign new_new_n8950__ = ~new_new_n8519__ & ~new_new_n8949__;
  assign new_new_n8951__ = new_new_n8519__ & new_new_n8949__;
  assign new_new_n8952__ = ~new_new_n8950__ & ~new_new_n8951__;
  assign new_new_n8953__ = ~pi099 & ~new_new_n8952__;
  assign new_new_n8954__ = pi099 & new_new_n8952__;
  assign new_new_n8955__ = ~new_new_n8529__ & ~new_new_n8530__;
  assign new_new_n8956__ = ~new_new_n8896__ & po025;
  assign new_new_n8957__ = ~pi097 & ~po025;
  assign new_new_n8958__ = ~new_new_n8956__ & ~new_new_n8957__;
  assign new_new_n8959__ = new_new_n8955__ & ~new_new_n8958__;
  assign new_new_n8960__ = ~new_new_n8955__ & new_new_n8958__;
  assign new_new_n8961__ = ~new_new_n8959__ & ~new_new_n8960__;
  assign new_new_n8962__ = pi098 & ~new_new_n8961__;
  assign new_new_n8963__ = ~pi098 & new_new_n8961__;
  assign new_new_n8964__ = ~new_new_n8886__ & ~new_new_n8887__;
  assign new_new_n8965__ = po025 & new_new_n8964__;
  assign new_new_n8966__ = new_new_n8894__ & ~new_new_n8965__;
  assign new_new_n8967__ = ~new_new_n8894__ & new_new_n8965__;
  assign new_new_n8968__ = ~new_new_n8966__ & ~new_new_n8967__;
  assign new_new_n8969__ = pi097 & ~new_new_n8968__;
  assign new_new_n8970__ = ~pi097 & new_new_n8968__;
  assign new_new_n8971__ = ~pi095 & ~new_new_n8883__;
  assign new_new_n8972__ = pi095 & new_new_n8883__;
  assign new_new_n8973__ = ~new_new_n8971__ & ~new_new_n8972__;
  assign new_new_n8974__ = po025 & new_new_n8973__;
  assign new_new_n8975__ = new_new_n8537__ & new_new_n8974__;
  assign new_new_n8976__ = ~new_new_n8537__ & ~new_new_n8974__;
  assign new_new_n8977__ = ~new_new_n8975__ & ~new_new_n8976__;
  assign new_new_n8978__ = ~pi096 & ~new_new_n8977__;
  assign new_new_n8979__ = pi096 & new_new_n8977__;
  assign new_new_n8980__ = ~pi094 & ~new_new_n8881__;
  assign new_new_n8981__ = pi094 & new_new_n8881__;
  assign new_new_n8982__ = ~new_new_n8980__ & ~new_new_n8981__;
  assign new_new_n8983__ = po025 & new_new_n8982__;
  assign new_new_n8984__ = new_new_n8546__ & new_new_n8983__;
  assign new_new_n8985__ = ~new_new_n8546__ & ~new_new_n8983__;
  assign new_new_n8986__ = ~new_new_n8984__ & ~new_new_n8985__;
  assign new_new_n8987__ = pi095 & new_new_n8986__;
  assign new_new_n8988__ = ~pi095 & ~new_new_n8986__;
  assign new_new_n8989__ = ~new_new_n8556__ & ~new_new_n8557__;
  assign new_new_n8990__ = ~new_new_n8879__ & po025;
  assign new_new_n8991__ = ~pi093 & ~po025;
  assign new_new_n8992__ = ~new_new_n8990__ & ~new_new_n8991__;
  assign new_new_n8993__ = new_new_n8989__ & ~new_new_n8992__;
  assign new_new_n8994__ = ~new_new_n8989__ & new_new_n8992__;
  assign new_new_n8995__ = ~new_new_n8993__ & ~new_new_n8994__;
  assign new_new_n8996__ = pi094 & ~new_new_n8995__;
  assign new_new_n8997__ = ~pi094 & new_new_n8995__;
  assign new_new_n8998__ = ~new_new_n8565__ & ~new_new_n8566__;
  assign new_new_n8999__ = ~new_new_n8877__ & po025;
  assign new_new_n9000__ = ~pi092 & ~po025;
  assign new_new_n9001__ = ~new_new_n8999__ & ~new_new_n9000__;
  assign new_new_n9002__ = ~new_new_n8998__ & ~new_new_n9001__;
  assign new_new_n9003__ = new_new_n8998__ & new_new_n9001__;
  assign new_new_n9004__ = ~new_new_n9002__ & ~new_new_n9003__;
  assign new_new_n9005__ = ~pi093 & ~new_new_n9004__;
  assign new_new_n9006__ = pi093 & new_new_n9004__;
  assign new_new_n9007__ = new_new_n8875__ & po025;
  assign new_new_n9008__ = ~pi091 & ~po025;
  assign new_new_n9009__ = ~new_new_n9007__ & ~new_new_n9008__;
  assign new_new_n9010__ = ~new_new_n8574__ & ~new_new_n8575__;
  assign new_new_n9011__ = ~new_new_n9009__ & ~new_new_n9010__;
  assign new_new_n9012__ = new_new_n9009__ & new_new_n9010__;
  assign new_new_n9013__ = ~new_new_n9011__ & ~new_new_n9012__;
  assign new_new_n9014__ = ~pi092 & ~new_new_n9013__;
  assign new_new_n9015__ = pi092 & new_new_n9013__;
  assign new_new_n9016__ = pi090 & ~new_new_n8873__;
  assign new_new_n9017__ = ~pi090 & new_new_n8873__;
  assign new_new_n9018__ = ~new_new_n9016__ & ~new_new_n9017__;
  assign new_new_n9019__ = po025 & new_new_n9018__;
  assign new_new_n9020__ = new_new_n8582__ & new_new_n9019__;
  assign new_new_n9021__ = ~new_new_n8582__ & ~new_new_n9019__;
  assign new_new_n9022__ = ~new_new_n9020__ & ~new_new_n9021__;
  assign new_new_n9023__ = ~pi091 & new_new_n9022__;
  assign new_new_n9024__ = pi091 & ~new_new_n9022__;
  assign new_new_n9025__ = ~new_new_n8592__ & ~new_new_n8593__;
  assign new_new_n9026__ = ~new_new_n8871__ & po025;
  assign new_new_n9027__ = ~pi089 & ~po025;
  assign new_new_n9028__ = ~new_new_n9026__ & ~new_new_n9027__;
  assign new_new_n9029__ = new_new_n9025__ & ~new_new_n9028__;
  assign new_new_n9030__ = ~new_new_n9025__ & new_new_n9028__;
  assign new_new_n9031__ = ~new_new_n9029__ & ~new_new_n9030__;
  assign new_new_n9032__ = ~pi090 & new_new_n9031__;
  assign new_new_n9033__ = pi090 & ~new_new_n9031__;
  assign new_new_n9034__ = ~new_new_n8869__ & po025;
  assign new_new_n9035__ = pi088 & ~po025;
  assign new_new_n9036__ = ~new_new_n9034__ & ~new_new_n9035__;
  assign new_new_n9037__ = ~new_new_n8601__ & ~new_new_n8602__;
  assign new_new_n9038__ = ~new_new_n9036__ & new_new_n9037__;
  assign new_new_n9039__ = new_new_n9036__ & ~new_new_n9037__;
  assign new_new_n9040__ = ~new_new_n9038__ & ~new_new_n9039__;
  assign new_new_n9041__ = ~pi089 & ~new_new_n9040__;
  assign new_new_n9042__ = pi089 & new_new_n9040__;
  assign new_new_n9043__ = ~new_new_n8867__ & po025;
  assign new_new_n9044__ = pi087 & ~po025;
  assign new_new_n9045__ = ~new_new_n9043__ & ~new_new_n9044__;
  assign new_new_n9046__ = ~new_new_n8610__ & ~new_new_n8611__;
  assign new_new_n9047__ = ~new_new_n9045__ & new_new_n9046__;
  assign new_new_n9048__ = new_new_n9045__ & ~new_new_n9046__;
  assign new_new_n9049__ = ~new_new_n9047__ & ~new_new_n9048__;
  assign new_new_n9050__ = ~pi088 & ~new_new_n9049__;
  assign new_new_n9051__ = pi088 & new_new_n9049__;
  assign new_new_n9052__ = ~new_new_n8619__ & ~new_new_n8620__;
  assign new_new_n9053__ = ~new_new_n8865__ & po025;
  assign new_new_n9054__ = pi086 & ~po025;
  assign new_new_n9055__ = ~new_new_n9053__ & ~new_new_n9054__;
  assign new_new_n9056__ = new_new_n9052__ & ~new_new_n9055__;
  assign new_new_n9057__ = ~new_new_n9052__ & new_new_n9055__;
  assign new_new_n9058__ = ~new_new_n9056__ & ~new_new_n9057__;
  assign new_new_n9059__ = pi087 & new_new_n9058__;
  assign new_new_n9060__ = ~pi087 & ~new_new_n9058__;
  assign new_new_n9061__ = ~new_new_n8628__ & ~new_new_n8863__;
  assign new_new_n9062__ = ~new_new_n8862__ & po025;
  assign new_new_n9063__ = ~pi085 & ~po025;
  assign new_new_n9064__ = ~new_new_n9062__ & ~new_new_n9063__;
  assign new_new_n9065__ = new_new_n9061__ & ~new_new_n9064__;
  assign new_new_n9066__ = ~new_new_n9061__ & new_new_n9064__;
  assign new_new_n9067__ = ~new_new_n9065__ & ~new_new_n9066__;
  assign new_new_n9068__ = pi086 & ~new_new_n9067__;
  assign new_new_n9069__ = ~pi086 & new_new_n9067__;
  assign new_new_n9070__ = ~new_new_n8636__ & ~new_new_n8637__;
  assign new_new_n9071__ = ~new_new_n8860__ & po025;
  assign new_new_n9072__ = ~pi084 & ~po025;
  assign new_new_n9073__ = ~new_new_n9071__ & ~new_new_n9072__;
  assign new_new_n9074__ = ~new_new_n9070__ & ~new_new_n9073__;
  assign new_new_n9075__ = new_new_n9070__ & new_new_n9073__;
  assign new_new_n9076__ = ~new_new_n9074__ & ~new_new_n9075__;
  assign new_new_n9077__ = pi085 & new_new_n9076__;
  assign new_new_n9078__ = ~pi085 & ~new_new_n9076__;
  assign new_new_n9079__ = ~new_new_n8645__ & ~new_new_n8646__;
  assign new_new_n9080__ = ~new_new_n8858__ & po025;
  assign new_new_n9081__ = ~pi083 & ~po025;
  assign new_new_n9082__ = ~new_new_n9080__ & ~new_new_n9081__;
  assign new_new_n9083__ = ~new_new_n9079__ & ~new_new_n9082__;
  assign new_new_n9084__ = new_new_n9079__ & new_new_n9082__;
  assign new_new_n9085__ = ~new_new_n9083__ & ~new_new_n9084__;
  assign new_new_n9086__ = pi084 & new_new_n9085__;
  assign new_new_n9087__ = ~pi084 & ~new_new_n9085__;
  assign new_new_n9088__ = ~pi082 & ~new_new_n8856__;
  assign new_new_n9089__ = pi082 & new_new_n8856__;
  assign new_new_n9090__ = ~new_new_n9088__ & ~new_new_n9089__;
  assign new_new_n9091__ = po025 & new_new_n9090__;
  assign new_new_n9092__ = ~new_new_n8653__ & ~new_new_n9091__;
  assign new_new_n9093__ = new_new_n8653__ & new_new_n9091__;
  assign new_new_n9094__ = ~new_new_n9092__ & ~new_new_n9093__;
  assign new_new_n9095__ = pi083 & new_new_n9094__;
  assign new_new_n9096__ = ~pi083 & ~new_new_n9094__;
  assign new_new_n9097__ = ~new_new_n8663__ & ~new_new_n8664__;
  assign new_new_n9098__ = ~new_new_n8854__ & po025;
  assign new_new_n9099__ = ~pi081 & ~po025;
  assign new_new_n9100__ = ~new_new_n9098__ & ~new_new_n9099__;
  assign new_new_n9101__ = new_new_n9097__ & ~new_new_n9100__;
  assign new_new_n9102__ = ~new_new_n9097__ & new_new_n9100__;
  assign new_new_n9103__ = ~new_new_n9101__ & ~new_new_n9102__;
  assign new_new_n9104__ = pi082 & ~new_new_n9103__;
  assign new_new_n9105__ = ~pi082 & new_new_n9103__;
  assign new_new_n9106__ = ~new_new_n8672__ & ~new_new_n8673__;
  assign new_new_n9107__ = ~new_new_n8852__ & po025;
  assign new_new_n9108__ = ~pi080 & ~po025;
  assign new_new_n9109__ = ~new_new_n9107__ & ~new_new_n9108__;
  assign new_new_n9110__ = new_new_n9106__ & ~new_new_n9109__;
  assign new_new_n9111__ = ~new_new_n9106__ & new_new_n9109__;
  assign new_new_n9112__ = ~new_new_n9110__ & ~new_new_n9111__;
  assign new_new_n9113__ = pi081 & ~new_new_n9112__;
  assign new_new_n9114__ = ~pi081 & new_new_n9112__;
  assign new_new_n9115__ = ~new_new_n8681__ & ~new_new_n8682__;
  assign new_new_n9116__ = ~new_new_n8850__ & po025;
  assign new_new_n9117__ = ~pi079 & ~po025;
  assign new_new_n9118__ = ~new_new_n9116__ & ~new_new_n9117__;
  assign new_new_n9119__ = new_new_n9115__ & ~new_new_n9118__;
  assign new_new_n9120__ = ~new_new_n9115__ & new_new_n9118__;
  assign new_new_n9121__ = ~new_new_n9119__ & ~new_new_n9120__;
  assign new_new_n9122__ = pi080 & ~new_new_n9121__;
  assign new_new_n9123__ = ~pi080 & new_new_n9121__;
  assign new_new_n9124__ = ~pi078 & ~new_new_n8848__;
  assign new_new_n9125__ = pi078 & new_new_n8848__;
  assign new_new_n9126__ = ~new_new_n9124__ & ~new_new_n9125__;
  assign new_new_n9127__ = po025 & new_new_n9126__;
  assign new_new_n9128__ = new_new_n8689__ & new_new_n9127__;
  assign new_new_n9129__ = ~new_new_n8689__ & ~new_new_n9127__;
  assign new_new_n9130__ = ~new_new_n9128__ & ~new_new_n9129__;
  assign new_new_n9131__ = ~pi079 & ~new_new_n9130__;
  assign new_new_n9132__ = pi079 & new_new_n9130__;
  assign new_new_n9133__ = ~new_new_n8699__ & ~new_new_n8700__;
  assign new_new_n9134__ = ~new_new_n8846__ & po025;
  assign new_new_n9135__ = pi077 & ~po025;
  assign new_new_n9136__ = ~new_new_n9134__ & ~new_new_n9135__;
  assign new_new_n9137__ = new_new_n9133__ & ~new_new_n9136__;
  assign new_new_n9138__ = ~new_new_n9133__ & new_new_n9136__;
  assign new_new_n9139__ = ~new_new_n9137__ & ~new_new_n9138__;
  assign new_new_n9140__ = ~pi078 & ~new_new_n9139__;
  assign new_new_n9141__ = pi078 & new_new_n9139__;
  assign new_new_n9142__ = ~new_new_n8708__ & ~new_new_n8709__;
  assign new_new_n9143__ = ~new_new_n8844__ & po025;
  assign new_new_n9144__ = ~pi076 & ~po025;
  assign new_new_n9145__ = ~new_new_n9143__ & ~new_new_n9144__;
  assign new_new_n9146__ = new_new_n9142__ & ~new_new_n9145__;
  assign new_new_n9147__ = ~new_new_n9142__ & new_new_n9145__;
  assign new_new_n9148__ = ~new_new_n9146__ & ~new_new_n9147__;
  assign new_new_n9149__ = pi077 & ~new_new_n9148__;
  assign new_new_n9150__ = ~pi077 & new_new_n9148__;
  assign new_new_n9151__ = ~new_new_n8717__ & ~new_new_n8718__;
  assign new_new_n9152__ = ~new_new_n8842__ & po025;
  assign new_new_n9153__ = ~pi075 & ~po025;
  assign new_new_n9154__ = ~new_new_n9152__ & ~new_new_n9153__;
  assign new_new_n9155__ = new_new_n9151__ & ~new_new_n9154__;
  assign new_new_n9156__ = ~new_new_n9151__ & new_new_n9154__;
  assign new_new_n9157__ = ~new_new_n9155__ & ~new_new_n9156__;
  assign new_new_n9158__ = pi076 & ~new_new_n9157__;
  assign new_new_n9159__ = ~pi076 & new_new_n9157__;
  assign new_new_n9160__ = ~new_new_n8726__ & ~new_new_n8727__;
  assign new_new_n9161__ = ~new_new_n8840__ & po025;
  assign new_new_n9162__ = ~pi074 & ~po025;
  assign new_new_n9163__ = ~new_new_n9161__ & ~new_new_n9162__;
  assign new_new_n9164__ = new_new_n9160__ & new_new_n9163__;
  assign new_new_n9165__ = ~new_new_n9160__ & ~new_new_n9163__;
  assign new_new_n9166__ = ~new_new_n9164__ & ~new_new_n9165__;
  assign new_new_n9167__ = ~pi075 & ~new_new_n9166__;
  assign new_new_n9168__ = pi075 & new_new_n9166__;
  assign new_new_n9169__ = ~new_new_n8735__ & ~new_new_n8736__;
  assign new_new_n9170__ = ~new_new_n8838__ & po025;
  assign new_new_n9171__ = ~pi073 & ~po025;
  assign new_new_n9172__ = ~new_new_n9170__ & ~new_new_n9171__;
  assign new_new_n9173__ = new_new_n9169__ & ~new_new_n9172__;
  assign new_new_n9174__ = ~new_new_n9169__ & new_new_n9172__;
  assign new_new_n9175__ = ~new_new_n9173__ & ~new_new_n9174__;
  assign new_new_n9176__ = ~pi074 & new_new_n9175__;
  assign new_new_n9177__ = pi074 & ~new_new_n9175__;
  assign new_new_n9178__ = ~new_new_n8836__ & po025;
  assign new_new_n9179__ = pi072 & ~po025;
  assign new_new_n9180__ = ~new_new_n9178__ & ~new_new_n9179__;
  assign new_new_n9181__ = ~new_new_n8744__ & ~new_new_n8745__;
  assign new_new_n9182__ = ~new_new_n9180__ & new_new_n9181__;
  assign new_new_n9183__ = new_new_n9180__ & ~new_new_n9181__;
  assign new_new_n9184__ = ~new_new_n9182__ & ~new_new_n9183__;
  assign new_new_n9185__ = ~pi073 & ~new_new_n9184__;
  assign new_new_n9186__ = pi073 & new_new_n9184__;
  assign new_new_n9187__ = ~new_new_n8751__ & ~new_new_n8752__;
  assign new_new_n9188__ = ~new_new_n8834__ & po025;
  assign new_new_n9189__ = pi071 & ~po025;
  assign new_new_n9190__ = ~new_new_n9188__ & ~new_new_n9189__;
  assign new_new_n9191__ = new_new_n9187__ & new_new_n9190__;
  assign new_new_n9192__ = ~new_new_n9187__ & ~new_new_n9190__;
  assign new_new_n9193__ = ~new_new_n9191__ & ~new_new_n9192__;
  assign new_new_n9194__ = pi072 & ~new_new_n9193__;
  assign new_new_n9195__ = ~pi072 & new_new_n9193__;
  assign new_new_n9196__ = new_new_n8832__ & po025;
  assign new_new_n9197__ = pi070 & ~po025;
  assign new_new_n9198__ = ~new_new_n9196__ & ~new_new_n9197__;
  assign new_new_n9199__ = ~new_new_n8760__ & ~new_new_n8761__;
  assign new_new_n9200__ = ~new_new_n9198__ & ~new_new_n9199__;
  assign new_new_n9201__ = new_new_n9198__ & new_new_n9199__;
  assign new_new_n9202__ = ~new_new_n9200__ & ~new_new_n9201__;
  assign new_new_n9203__ = pi071 & ~new_new_n9202__;
  assign new_new_n9204__ = ~pi071 & new_new_n9202__;
  assign new_new_n9205__ = ~new_new_n8776__ & ~new_new_n8777__;
  assign new_new_n9206__ = ~new_new_n8828__ & po025;
  assign new_new_n9207__ = ~pi068 & ~po025;
  assign new_new_n9208__ = ~new_new_n9206__ & ~new_new_n9207__;
  assign new_new_n9209__ = new_new_n9205__ & ~new_new_n9208__;
  assign new_new_n9210__ = ~new_new_n9205__ & new_new_n9208__;
  assign new_new_n9211__ = ~new_new_n9209__ & ~new_new_n9210__;
  assign new_new_n9212__ = pi069 & ~new_new_n9211__;
  assign new_new_n9213__ = ~pi069 & new_new_n9211__;
  assign new_new_n9214__ = ~new_new_n8797__ & po025;
  assign new_new_n9215__ = ~new_new_n8824__ & new_new_n9214__;
  assign new_new_n9216__ = new_new_n8823__ & ~new_new_n9215__;
  assign new_new_n9217__ = new_new_n8825__ & new_new_n9214__;
  assign new_new_n9218__ = ~new_new_n9216__ & ~new_new_n9217__;
  assign new_new_n9219__ = ~pi067 & ~new_new_n9218__;
  assign new_new_n9220__ = pi067 & new_new_n9218__;
  assign new_new_n9221__ = pi025 & po025;
  assign new_new_n9222__ = ~pi025 & ~po025;
  assign new_new_n9223__ = ~pi065 & ~new_new_n9221__;
  assign new_new_n9224__ = ~new_new_n9222__ & new_new_n9223__;
  assign new_new_n9225__ = ~pi024 & ~new_new_n9224__;
  assign new_new_n9226__ = pi065 & new_new_n9221__;
  assign new_new_n9227__ = ~new_new_n9225__ & ~new_new_n9226__;
  assign new_new_n9228__ = pi064 & ~new_new_n9227__;
  assign new_new_n9229__ = pi064 & po025;
  assign new_new_n9230__ = ~pi025 & pi065;
  assign new_new_n9231__ = ~new_new_n9229__ & new_new_n9230__;
  assign new_new_n9232__ = ~new_new_n9228__ & ~new_new_n9231__;
  assign new_new_n9233__ = pi066 & ~new_new_n9232__;
  assign new_new_n9234__ = new_new_n426__ & ~po026;
  assign new_new_n9235__ = new_new_n8816__ & po025;
  assign new_new_n9236__ = ~new_new_n9234__ & ~new_new_n9235__;
  assign new_new_n9237__ = ~pi025 & ~new_new_n9236__;
  assign new_new_n9238__ = ~new_new_n332__ & po025;
  assign new_new_n9239__ = ~new_new_n8793__ & ~new_new_n9238__;
  assign new_new_n9240__ = pi065 & po025;
  assign new_new_n9241__ = po026 & ~new_new_n9240__;
  assign new_new_n9242__ = pi065 & ~new_new_n8793__;
  assign new_new_n9243__ = pi025 & ~new_new_n9242__;
  assign new_new_n9244__ = ~new_new_n9241__ & new_new_n9243__;
  assign new_new_n9245__ = ~new_new_n9237__ & ~new_new_n9239__;
  assign new_new_n9246__ = ~new_new_n9244__ & new_new_n9245__;
  assign new_new_n9247__ = ~pi026 & ~new_new_n9246__;
  assign new_new_n9248__ = ~pi064 & ~new_new_n9240__;
  assign new_new_n9249__ = ~pi065 & po025;
  assign new_new_n9250__ = ~po026 & ~new_new_n9249__;
  assign new_new_n9251__ = ~new_new_n9221__ & ~new_new_n9235__;
  assign new_new_n9252__ = ~new_new_n9250__ & new_new_n9251__;
  assign new_new_n9253__ = pi064 & ~new_new_n9252__;
  assign new_new_n9254__ = ~new_new_n9248__ & ~new_new_n9253__;
  assign new_new_n9255__ = ~new_new_n8793__ & ~new_new_n9240__;
  assign new_new_n9256__ = pi025 & ~new_new_n8804__;
  assign new_new_n9257__ = ~new_new_n9255__ & new_new_n9256__;
  assign new_new_n9258__ = ~new_new_n9254__ & ~new_new_n9257__;
  assign new_new_n9259__ = pi026 & ~new_new_n9258__;
  assign new_new_n9260__ = ~new_new_n9247__ & ~new_new_n9259__;
  assign new_new_n9261__ = ~pi066 & new_new_n9232__;
  assign new_new_n9262__ = ~new_new_n9260__ & ~new_new_n9261__;
  assign new_new_n9263__ = ~new_new_n9233__ & ~new_new_n9262__;
  assign new_new_n9264__ = ~new_new_n9220__ & new_new_n9263__;
  assign new_new_n9265__ = ~new_new_n9219__ & ~new_new_n9264__;
  assign new_new_n9266__ = pi068 & new_new_n9265__;
  assign new_new_n9267__ = ~pi068 & ~new_new_n9265__;
  assign new_new_n9268__ = ~new_new_n8783__ & ~new_new_n8784__;
  assign new_new_n9269__ = new_new_n8826__ & po025;
  assign new_new_n9270__ = ~pi067 & ~po025;
  assign new_new_n9271__ = ~new_new_n9269__ & ~new_new_n9270__;
  assign new_new_n9272__ = ~new_new_n9268__ & ~new_new_n9271__;
  assign new_new_n9273__ = new_new_n9268__ & new_new_n9271__;
  assign new_new_n9274__ = ~new_new_n9272__ & ~new_new_n9273__;
  assign new_new_n9275__ = ~new_new_n9267__ & new_new_n9274__;
  assign new_new_n9276__ = ~new_new_n9266__ & ~new_new_n9275__;
  assign new_new_n9277__ = ~new_new_n9213__ & ~new_new_n9276__;
  assign new_new_n9278__ = ~new_new_n9212__ & ~new_new_n9277__;
  assign new_new_n9279__ = pi070 & ~new_new_n9278__;
  assign new_new_n9280__ = ~pi070 & new_new_n9278__;
  assign new_new_n9281__ = ~new_new_n8767__ & ~new_new_n8768__;
  assign new_new_n9282__ = ~new_new_n8830__ & po025;
  assign new_new_n9283__ = ~pi069 & ~po025;
  assign new_new_n9284__ = ~new_new_n9282__ & ~new_new_n9283__;
  assign new_new_n9285__ = new_new_n9281__ & ~new_new_n9284__;
  assign new_new_n9286__ = ~new_new_n9281__ & new_new_n9284__;
  assign new_new_n9287__ = ~new_new_n9285__ & ~new_new_n9286__;
  assign new_new_n9288__ = ~new_new_n9280__ & ~new_new_n9287__;
  assign new_new_n9289__ = ~new_new_n9279__ & ~new_new_n9288__;
  assign new_new_n9290__ = ~new_new_n9204__ & ~new_new_n9289__;
  assign new_new_n9291__ = ~new_new_n9203__ & ~new_new_n9290__;
  assign new_new_n9292__ = ~new_new_n9195__ & ~new_new_n9291__;
  assign new_new_n9293__ = ~new_new_n9194__ & ~new_new_n9292__;
  assign new_new_n9294__ = ~new_new_n9186__ & new_new_n9293__;
  assign new_new_n9295__ = ~new_new_n9185__ & ~new_new_n9294__;
  assign new_new_n9296__ = ~new_new_n9177__ & ~new_new_n9295__;
  assign new_new_n9297__ = ~new_new_n9176__ & ~new_new_n9296__;
  assign new_new_n9298__ = ~new_new_n9168__ & ~new_new_n9297__;
  assign new_new_n9299__ = ~new_new_n9167__ & ~new_new_n9298__;
  assign new_new_n9300__ = ~new_new_n9159__ & new_new_n9299__;
  assign new_new_n9301__ = ~new_new_n9158__ & ~new_new_n9300__;
  assign new_new_n9302__ = ~new_new_n9150__ & ~new_new_n9301__;
  assign new_new_n9303__ = ~new_new_n9149__ & ~new_new_n9302__;
  assign new_new_n9304__ = ~new_new_n9141__ & new_new_n9303__;
  assign new_new_n9305__ = ~new_new_n9140__ & ~new_new_n9304__;
  assign new_new_n9306__ = ~new_new_n9132__ & ~new_new_n9305__;
  assign new_new_n9307__ = ~new_new_n9131__ & ~new_new_n9306__;
  assign new_new_n9308__ = ~new_new_n9123__ & new_new_n9307__;
  assign new_new_n9309__ = ~new_new_n9122__ & ~new_new_n9308__;
  assign new_new_n9310__ = ~new_new_n9114__ & ~new_new_n9309__;
  assign new_new_n9311__ = ~new_new_n9113__ & ~new_new_n9310__;
  assign new_new_n9312__ = ~new_new_n9105__ & ~new_new_n9311__;
  assign new_new_n9313__ = ~new_new_n9104__ & ~new_new_n9312__;
  assign new_new_n9314__ = ~new_new_n9096__ & ~new_new_n9313__;
  assign new_new_n9315__ = ~new_new_n9095__ & ~new_new_n9314__;
  assign new_new_n9316__ = ~new_new_n9087__ & ~new_new_n9315__;
  assign new_new_n9317__ = ~new_new_n9086__ & ~new_new_n9316__;
  assign new_new_n9318__ = ~new_new_n9078__ & ~new_new_n9317__;
  assign new_new_n9319__ = ~new_new_n9077__ & ~new_new_n9318__;
  assign new_new_n9320__ = ~new_new_n9069__ & ~new_new_n9319__;
  assign new_new_n9321__ = ~new_new_n9068__ & ~new_new_n9320__;
  assign new_new_n9322__ = ~new_new_n9060__ & ~new_new_n9321__;
  assign new_new_n9323__ = ~new_new_n9059__ & ~new_new_n9322__;
  assign new_new_n9324__ = ~new_new_n9051__ & new_new_n9323__;
  assign new_new_n9325__ = ~new_new_n9050__ & ~new_new_n9324__;
  assign new_new_n9326__ = ~new_new_n9042__ & ~new_new_n9325__;
  assign new_new_n9327__ = ~new_new_n9041__ & ~new_new_n9326__;
  assign new_new_n9328__ = ~new_new_n9033__ & ~new_new_n9327__;
  assign new_new_n9329__ = ~new_new_n9032__ & ~new_new_n9328__;
  assign new_new_n9330__ = ~new_new_n9024__ & ~new_new_n9329__;
  assign new_new_n9331__ = ~new_new_n9023__ & ~new_new_n9330__;
  assign new_new_n9332__ = ~new_new_n9015__ & ~new_new_n9331__;
  assign new_new_n9333__ = ~new_new_n9014__ & ~new_new_n9332__;
  assign new_new_n9334__ = ~new_new_n9006__ & ~new_new_n9333__;
  assign new_new_n9335__ = ~new_new_n9005__ & ~new_new_n9334__;
  assign new_new_n9336__ = ~new_new_n8997__ & new_new_n9335__;
  assign new_new_n9337__ = ~new_new_n8996__ & ~new_new_n9336__;
  assign new_new_n9338__ = ~new_new_n8988__ & ~new_new_n9337__;
  assign new_new_n9339__ = ~new_new_n8987__ & ~new_new_n9338__;
  assign new_new_n9340__ = ~new_new_n8979__ & new_new_n9339__;
  assign new_new_n9341__ = ~new_new_n8978__ & ~new_new_n9340__;
  assign new_new_n9342__ = ~new_new_n8970__ & new_new_n9341__;
  assign new_new_n9343__ = ~new_new_n8969__ & ~new_new_n9342__;
  assign new_new_n9344__ = ~new_new_n8963__ & ~new_new_n9343__;
  assign new_new_n9345__ = ~new_new_n8962__ & ~new_new_n9344__;
  assign new_new_n9346__ = ~new_new_n8954__ & new_new_n9345__;
  assign new_new_n9347__ = ~new_new_n8953__ & ~new_new_n9346__;
  assign new_new_n9348__ = ~new_new_n8945__ & new_new_n9347__;
  assign new_new_n9349__ = ~new_new_n8944__ & ~new_new_n9348__;
  assign new_new_n9350__ = ~new_new_n8936__ & new_new_n9349__;
  assign new_new_n9351__ = ~new_new_n8935__ & ~new_new_n9350__;
  assign new_new_n9352__ = ~new_new_n8925__ & new_new_n9351__;
  assign new_new_n9353__ = pi102 & new_new_n8924__;
  assign new_new_n9354__ = pi103 & new_new_n8064__;
  assign new_new_n9355__ = ~new_new_n9353__ & ~new_new_n9354__;
  assign new_new_n9356__ = ~new_new_n9352__ & new_new_n9355__;
  assign new_new_n9357__ = ~pi103 & ~new_new_n8910__;
  assign new_new_n9358__ = ~new_new_n9356__ & ~new_new_n9357__;
  assign po024 = new_new_n8069__ & ~new_new_n9358__;
  assign new_new_n9360__ = ~new_new_n376__ & po024;
  assign new_new_n9361__ = ~new_new_n8910__ & ~new_new_n9360__;
  assign new_new_n9362__ = ~new_new_n8925__ & ~new_new_n9353__;
  assign new_new_n9363__ = ~new_new_n9351__ & po024;
  assign new_new_n9364__ = ~pi102 & ~po024;
  assign new_new_n9365__ = ~new_new_n9363__ & ~new_new_n9364__;
  assign new_new_n9366__ = new_new_n9362__ & ~new_new_n9365__;
  assign new_new_n9367__ = ~new_new_n9362__ & new_new_n9365__;
  assign new_new_n9368__ = ~new_new_n9366__ & ~new_new_n9367__;
  assign new_new_n9369__ = pi103 & ~new_new_n9368__;
  assign new_new_n9370__ = ~pi103 & new_new_n9368__;
  assign new_new_n9371__ = ~new_new_n9349__ & po024;
  assign new_new_n9372__ = pi101 & ~po024;
  assign new_new_n9373__ = ~new_new_n9371__ & ~new_new_n9372__;
  assign new_new_n9374__ = ~new_new_n8935__ & ~new_new_n8936__;
  assign new_new_n9375__ = ~new_new_n9373__ & new_new_n9374__;
  assign new_new_n9376__ = new_new_n9373__ & ~new_new_n9374__;
  assign new_new_n9377__ = ~new_new_n9375__ & ~new_new_n9376__;
  assign new_new_n9378__ = pi102 & new_new_n9377__;
  assign new_new_n9379__ = ~pi102 & ~new_new_n9377__;
  assign new_new_n9380__ = ~new_new_n8944__ & ~new_new_n8945__;
  assign new_new_n9381__ = ~new_new_n9347__ & po024;
  assign new_new_n9382__ = ~pi100 & ~po024;
  assign new_new_n9383__ = ~new_new_n9381__ & ~new_new_n9382__;
  assign new_new_n9384__ = new_new_n9380__ & ~new_new_n9383__;
  assign new_new_n9385__ = ~new_new_n9380__ & new_new_n9383__;
  assign new_new_n9386__ = ~new_new_n9384__ & ~new_new_n9385__;
  assign new_new_n9387__ = pi101 & ~new_new_n9386__;
  assign new_new_n9388__ = ~pi101 & new_new_n9386__;
  assign new_new_n9389__ = new_new_n9345__ & po024;
  assign new_new_n9390__ = ~pi099 & ~po024;
  assign new_new_n9391__ = ~new_new_n9389__ & ~new_new_n9390__;
  assign new_new_n9392__ = ~new_new_n8953__ & ~new_new_n8954__;
  assign new_new_n9393__ = ~new_new_n9391__ & ~new_new_n9392__;
  assign new_new_n9394__ = new_new_n9391__ & new_new_n9392__;
  assign new_new_n9395__ = ~new_new_n9393__ & ~new_new_n9394__;
  assign new_new_n9396__ = ~pi100 & ~new_new_n9395__;
  assign new_new_n9397__ = pi100 & new_new_n9395__;
  assign new_new_n9398__ = ~new_new_n8962__ & ~new_new_n8963__;
  assign new_new_n9399__ = ~new_new_n9343__ & po024;
  assign new_new_n9400__ = pi098 & ~po024;
  assign new_new_n9401__ = ~new_new_n9399__ & ~new_new_n9400__;
  assign new_new_n9402__ = new_new_n9398__ & new_new_n9401__;
  assign new_new_n9403__ = ~new_new_n9398__ & ~new_new_n9401__;
  assign new_new_n9404__ = ~new_new_n9402__ & ~new_new_n9403__;
  assign new_new_n9405__ = pi099 & ~new_new_n9404__;
  assign new_new_n9406__ = ~pi099 & new_new_n9404__;
  assign new_new_n9407__ = new_new_n9341__ & po024;
  assign new_new_n9408__ = pi097 & ~po024;
  assign new_new_n9409__ = ~new_new_n9407__ & ~new_new_n9408__;
  assign new_new_n9410__ = ~new_new_n8969__ & ~new_new_n8970__;
  assign new_new_n9411__ = ~new_new_n9409__ & ~new_new_n9410__;
  assign new_new_n9412__ = new_new_n9409__ & new_new_n9410__;
  assign new_new_n9413__ = ~new_new_n9411__ & ~new_new_n9412__;
  assign new_new_n9414__ = pi098 & ~new_new_n9413__;
  assign new_new_n9415__ = ~pi098 & new_new_n9413__;
  assign new_new_n9416__ = ~new_new_n8978__ & ~new_new_n8979__;
  assign new_new_n9417__ = new_new_n9339__ & po024;
  assign new_new_n9418__ = ~pi096 & ~po024;
  assign new_new_n9419__ = ~new_new_n9417__ & ~new_new_n9418__;
  assign new_new_n9420__ = ~new_new_n9416__ & ~new_new_n9419__;
  assign new_new_n9421__ = new_new_n9416__ & new_new_n9419__;
  assign new_new_n9422__ = ~new_new_n9420__ & ~new_new_n9421__;
  assign new_new_n9423__ = ~pi097 & ~new_new_n9422__;
  assign new_new_n9424__ = pi097 & new_new_n9422__;
  assign new_new_n9425__ = new_new_n9337__ & po024;
  assign new_new_n9426__ = ~pi095 & ~po024;
  assign new_new_n9427__ = ~new_new_n9425__ & ~new_new_n9426__;
  assign new_new_n9428__ = ~new_new_n8987__ & ~new_new_n8988__;
  assign new_new_n9429__ = ~new_new_n9427__ & ~new_new_n9428__;
  assign new_new_n9430__ = new_new_n9427__ & new_new_n9428__;
  assign new_new_n9431__ = ~new_new_n9429__ & ~new_new_n9430__;
  assign new_new_n9432__ = ~pi096 & ~new_new_n9431__;
  assign new_new_n9433__ = pi096 & new_new_n9431__;
  assign new_new_n9434__ = new_new_n9335__ & po024;
  assign new_new_n9435__ = pi094 & ~po024;
  assign new_new_n9436__ = ~new_new_n9434__ & ~new_new_n9435__;
  assign new_new_n9437__ = ~new_new_n8996__ & ~new_new_n8997__;
  assign new_new_n9438__ = ~new_new_n9436__ & ~new_new_n9437__;
  assign new_new_n9439__ = new_new_n9436__ & new_new_n9437__;
  assign new_new_n9440__ = ~new_new_n9438__ & ~new_new_n9439__;
  assign new_new_n9441__ = pi095 & ~new_new_n9440__;
  assign new_new_n9442__ = ~pi095 & new_new_n9440__;
  assign new_new_n9443__ = ~new_new_n9005__ & ~new_new_n9006__;
  assign new_new_n9444__ = ~new_new_n9333__ & po024;
  assign new_new_n9445__ = ~pi093 & ~po024;
  assign new_new_n9446__ = ~new_new_n9444__ & ~new_new_n9445__;
  assign new_new_n9447__ = ~new_new_n9443__ & ~new_new_n9446__;
  assign new_new_n9448__ = new_new_n9443__ & new_new_n9446__;
  assign new_new_n9449__ = ~new_new_n9447__ & ~new_new_n9448__;
  assign new_new_n9450__ = pi094 & new_new_n9449__;
  assign new_new_n9451__ = ~pi094 & ~new_new_n9449__;
  assign new_new_n9452__ = ~new_new_n9014__ & ~new_new_n9015__;
  assign new_new_n9453__ = ~new_new_n9331__ & po024;
  assign new_new_n9454__ = ~pi092 & ~po024;
  assign new_new_n9455__ = ~new_new_n9453__ & ~new_new_n9454__;
  assign new_new_n9456__ = new_new_n9452__ & ~new_new_n9455__;
  assign new_new_n9457__ = ~new_new_n9452__ & new_new_n9455__;
  assign new_new_n9458__ = ~new_new_n9456__ & ~new_new_n9457__;
  assign new_new_n9459__ = pi093 & ~new_new_n9458__;
  assign new_new_n9460__ = ~pi093 & new_new_n9458__;
  assign new_new_n9461__ = ~new_new_n9023__ & ~new_new_n9024__;
  assign new_new_n9462__ = ~new_new_n9329__ & po024;
  assign new_new_n9463__ = ~pi091 & ~po024;
  assign new_new_n9464__ = ~new_new_n9462__ & ~new_new_n9463__;
  assign new_new_n9465__ = new_new_n9461__ & ~new_new_n9464__;
  assign new_new_n9466__ = ~new_new_n9461__ & new_new_n9464__;
  assign new_new_n9467__ = ~new_new_n9465__ & ~new_new_n9466__;
  assign new_new_n9468__ = ~pi092 & new_new_n9467__;
  assign new_new_n9469__ = pi092 & ~new_new_n9467__;
  assign new_new_n9470__ = ~new_new_n9032__ & ~new_new_n9033__;
  assign new_new_n9471__ = ~new_new_n9327__ & po024;
  assign new_new_n9472__ = ~pi090 & ~po024;
  assign new_new_n9473__ = ~new_new_n9471__ & ~new_new_n9472__;
  assign new_new_n9474__ = new_new_n9470__ & ~new_new_n9473__;
  assign new_new_n9475__ = ~new_new_n9470__ & new_new_n9473__;
  assign new_new_n9476__ = ~new_new_n9474__ & ~new_new_n9475__;
  assign new_new_n9477__ = ~pi091 & new_new_n9476__;
  assign new_new_n9478__ = pi091 & ~new_new_n9476__;
  assign new_new_n9479__ = ~pi089 & ~new_new_n9325__;
  assign new_new_n9480__ = pi089 & new_new_n9325__;
  assign new_new_n9481__ = ~new_new_n9479__ & ~new_new_n9480__;
  assign new_new_n9482__ = po024 & new_new_n9481__;
  assign new_new_n9483__ = new_new_n9040__ & new_new_n9482__;
  assign new_new_n9484__ = ~new_new_n9040__ & ~new_new_n9482__;
  assign new_new_n9485__ = ~new_new_n9483__ & ~new_new_n9484__;
  assign new_new_n9486__ = ~pi090 & ~new_new_n9485__;
  assign new_new_n9487__ = pi090 & new_new_n9485__;
  assign new_new_n9488__ = ~new_new_n9323__ & po024;
  assign new_new_n9489__ = pi088 & ~po024;
  assign new_new_n9490__ = ~new_new_n9488__ & ~new_new_n9489__;
  assign new_new_n9491__ = ~new_new_n9050__ & ~new_new_n9051__;
  assign new_new_n9492__ = ~new_new_n9490__ & new_new_n9491__;
  assign new_new_n9493__ = new_new_n9490__ & ~new_new_n9491__;
  assign new_new_n9494__ = ~new_new_n9492__ & ~new_new_n9493__;
  assign new_new_n9495__ = ~pi089 & ~new_new_n9494__;
  assign new_new_n9496__ = pi089 & new_new_n9494__;
  assign new_new_n9497__ = ~new_new_n9321__ & po024;
  assign new_new_n9498__ = pi087 & ~po024;
  assign new_new_n9499__ = ~new_new_n9497__ & ~new_new_n9498__;
  assign new_new_n9500__ = ~new_new_n9059__ & ~new_new_n9060__;
  assign new_new_n9501__ = ~new_new_n9499__ & new_new_n9500__;
  assign new_new_n9502__ = new_new_n9499__ & ~new_new_n9500__;
  assign new_new_n9503__ = ~new_new_n9501__ & ~new_new_n9502__;
  assign new_new_n9504__ = ~pi088 & ~new_new_n9503__;
  assign new_new_n9505__ = pi088 & new_new_n9503__;
  assign new_new_n9506__ = ~new_new_n9068__ & ~new_new_n9069__;
  assign new_new_n9507__ = ~new_new_n9319__ & po024;
  assign new_new_n9508__ = pi086 & ~po024;
  assign new_new_n9509__ = ~new_new_n9507__ & ~new_new_n9508__;
  assign new_new_n9510__ = new_new_n9506__ & ~new_new_n9509__;
  assign new_new_n9511__ = ~new_new_n9506__ & new_new_n9509__;
  assign new_new_n9512__ = ~new_new_n9510__ & ~new_new_n9511__;
  assign new_new_n9513__ = ~pi087 & ~new_new_n9512__;
  assign new_new_n9514__ = pi087 & new_new_n9512__;
  assign new_new_n9515__ = ~new_new_n9317__ & po024;
  assign new_new_n9516__ = pi085 & ~po024;
  assign new_new_n9517__ = ~new_new_n9515__ & ~new_new_n9516__;
  assign new_new_n9518__ = ~new_new_n9077__ & ~new_new_n9078__;
  assign new_new_n9519__ = ~new_new_n9517__ & new_new_n9518__;
  assign new_new_n9520__ = new_new_n9517__ & ~new_new_n9518__;
  assign new_new_n9521__ = ~new_new_n9519__ & ~new_new_n9520__;
  assign new_new_n9522__ = ~pi086 & ~new_new_n9521__;
  assign new_new_n9523__ = pi086 & new_new_n9521__;
  assign new_new_n9524__ = ~new_new_n9315__ & po024;
  assign new_new_n9525__ = pi084 & ~po024;
  assign new_new_n9526__ = ~new_new_n9524__ & ~new_new_n9525__;
  assign new_new_n9527__ = ~new_new_n9086__ & ~new_new_n9087__;
  assign new_new_n9528__ = ~new_new_n9526__ & new_new_n9527__;
  assign new_new_n9529__ = new_new_n9526__ & ~new_new_n9527__;
  assign new_new_n9530__ = ~new_new_n9528__ & ~new_new_n9529__;
  assign new_new_n9531__ = ~pi085 & ~new_new_n9530__;
  assign new_new_n9532__ = pi085 & new_new_n9530__;
  assign new_new_n9533__ = ~new_new_n9095__ & ~new_new_n9096__;
  assign new_new_n9534__ = ~new_new_n9313__ & po024;
  assign new_new_n9535__ = pi083 & ~po024;
  assign new_new_n9536__ = ~new_new_n9534__ & ~new_new_n9535__;
  assign new_new_n9537__ = new_new_n9533__ & ~new_new_n9536__;
  assign new_new_n9538__ = ~new_new_n9533__ & new_new_n9536__;
  assign new_new_n9539__ = ~new_new_n9537__ & ~new_new_n9538__;
  assign new_new_n9540__ = ~pi084 & ~new_new_n9539__;
  assign new_new_n9541__ = pi084 & new_new_n9539__;
  assign new_new_n9542__ = pi082 & ~new_new_n9311__;
  assign new_new_n9543__ = ~pi082 & new_new_n9311__;
  assign new_new_n9544__ = ~new_new_n9542__ & ~new_new_n9543__;
  assign new_new_n9545__ = po024 & new_new_n9544__;
  assign new_new_n9546__ = ~new_new_n9103__ & ~new_new_n9545__;
  assign new_new_n9547__ = new_new_n9103__ & new_new_n9545__;
  assign new_new_n9548__ = ~new_new_n9546__ & ~new_new_n9547__;
  assign new_new_n9549__ = ~pi083 & new_new_n9548__;
  assign new_new_n9550__ = pi083 & ~new_new_n9548__;
  assign new_new_n9551__ = ~new_new_n9113__ & ~new_new_n9114__;
  assign new_new_n9552__ = ~new_new_n9309__ & po024;
  assign new_new_n9553__ = pi081 & ~po024;
  assign new_new_n9554__ = ~new_new_n9552__ & ~new_new_n9553__;
  assign new_new_n9555__ = new_new_n9551__ & ~new_new_n9554__;
  assign new_new_n9556__ = ~new_new_n9551__ & new_new_n9554__;
  assign new_new_n9557__ = ~new_new_n9555__ & ~new_new_n9556__;
  assign new_new_n9558__ = ~pi082 & ~new_new_n9557__;
  assign new_new_n9559__ = pi082 & new_new_n9557__;
  assign new_new_n9560__ = ~new_new_n9122__ & ~new_new_n9123__;
  assign new_new_n9561__ = ~new_new_n9307__ & po024;
  assign new_new_n9562__ = ~pi080 & ~po024;
  assign new_new_n9563__ = ~new_new_n9561__ & ~new_new_n9562__;
  assign new_new_n9564__ = new_new_n9560__ & ~new_new_n9563__;
  assign new_new_n9565__ = ~new_new_n9560__ & new_new_n9563__;
  assign new_new_n9566__ = ~new_new_n9564__ & ~new_new_n9565__;
  assign new_new_n9567__ = pi081 & ~new_new_n9566__;
  assign new_new_n9568__ = ~pi081 & new_new_n9566__;
  assign new_new_n9569__ = ~new_new_n9131__ & ~new_new_n9132__;
  assign new_new_n9570__ = ~new_new_n9305__ & po024;
  assign new_new_n9571__ = ~pi079 & ~po024;
  assign new_new_n9572__ = ~new_new_n9570__ & ~new_new_n9571__;
  assign new_new_n9573__ = new_new_n9569__ & ~new_new_n9572__;
  assign new_new_n9574__ = ~new_new_n9569__ & new_new_n9572__;
  assign new_new_n9575__ = ~new_new_n9573__ & ~new_new_n9574__;
  assign new_new_n9576__ = pi080 & ~new_new_n9575__;
  assign new_new_n9577__ = ~pi080 & new_new_n9575__;
  assign new_new_n9578__ = ~new_new_n9303__ & po024;
  assign new_new_n9579__ = pi078 & ~po024;
  assign new_new_n9580__ = ~new_new_n9578__ & ~new_new_n9579__;
  assign new_new_n9581__ = ~new_new_n9140__ & ~new_new_n9141__;
  assign new_new_n9582__ = ~new_new_n9580__ & new_new_n9581__;
  assign new_new_n9583__ = new_new_n9580__ & ~new_new_n9581__;
  assign new_new_n9584__ = ~new_new_n9582__ & ~new_new_n9583__;
  assign new_new_n9585__ = ~pi079 & ~new_new_n9584__;
  assign new_new_n9586__ = pi079 & new_new_n9584__;
  assign new_new_n9587__ = ~new_new_n9149__ & ~new_new_n9150__;
  assign new_new_n9588__ = ~new_new_n9301__ & po024;
  assign new_new_n9589__ = pi077 & ~po024;
  assign new_new_n9590__ = ~new_new_n9588__ & ~new_new_n9589__;
  assign new_new_n9591__ = new_new_n9587__ & ~new_new_n9590__;
  assign new_new_n9592__ = ~new_new_n9587__ & new_new_n9590__;
  assign new_new_n9593__ = ~new_new_n9591__ & ~new_new_n9592__;
  assign new_new_n9594__ = pi078 & new_new_n9593__;
  assign new_new_n9595__ = ~pi078 & ~new_new_n9593__;
  assign new_new_n9596__ = ~new_new_n9158__ & ~new_new_n9159__;
  assign new_new_n9597__ = ~new_new_n9299__ & po024;
  assign new_new_n9598__ = ~pi076 & ~po024;
  assign new_new_n9599__ = ~new_new_n9597__ & ~new_new_n9598__;
  assign new_new_n9600__ = new_new_n9596__ & ~new_new_n9599__;
  assign new_new_n9601__ = ~new_new_n9596__ & new_new_n9599__;
  assign new_new_n9602__ = ~new_new_n9600__ & ~new_new_n9601__;
  assign new_new_n9603__ = pi077 & ~new_new_n9602__;
  assign new_new_n9604__ = ~pi077 & new_new_n9602__;
  assign new_new_n9605__ = ~pi075 & ~new_new_n9297__;
  assign new_new_n9606__ = pi075 & new_new_n9297__;
  assign new_new_n9607__ = ~new_new_n9605__ & ~new_new_n9606__;
  assign new_new_n9608__ = po024 & new_new_n9607__;
  assign new_new_n9609__ = new_new_n9166__ & new_new_n9608__;
  assign new_new_n9610__ = ~new_new_n9166__ & ~new_new_n9608__;
  assign new_new_n9611__ = ~new_new_n9609__ & ~new_new_n9610__;
  assign new_new_n9612__ = ~pi076 & ~new_new_n9611__;
  assign new_new_n9613__ = pi076 & new_new_n9611__;
  assign new_new_n9614__ = ~new_new_n9176__ & ~new_new_n9177__;
  assign new_new_n9615__ = ~new_new_n9295__ & po024;
  assign new_new_n9616__ = ~pi074 & ~po024;
  assign new_new_n9617__ = ~new_new_n9615__ & ~new_new_n9616__;
  assign new_new_n9618__ = new_new_n9614__ & ~new_new_n9617__;
  assign new_new_n9619__ = ~new_new_n9614__ & new_new_n9617__;
  assign new_new_n9620__ = ~new_new_n9618__ & ~new_new_n9619__;
  assign new_new_n9621__ = pi075 & ~new_new_n9620__;
  assign new_new_n9622__ = ~new_new_n9293__ & po024;
  assign new_new_n9623__ = pi073 & ~po024;
  assign new_new_n9624__ = ~new_new_n9622__ & ~new_new_n9623__;
  assign new_new_n9625__ = ~new_new_n9185__ & ~new_new_n9186__;
  assign new_new_n9626__ = ~new_new_n9624__ & new_new_n9625__;
  assign new_new_n9627__ = new_new_n9624__ & ~new_new_n9625__;
  assign new_new_n9628__ = ~new_new_n9626__ & ~new_new_n9627__;
  assign new_new_n9629__ = ~pi074 & ~new_new_n9628__;
  assign new_new_n9630__ = pi074 & new_new_n9628__;
  assign new_new_n9631__ = ~new_new_n9194__ & ~new_new_n9195__;
  assign new_new_n9632__ = pi072 & ~po024;
  assign new_new_n9633__ = ~new_new_n9291__ & po024;
  assign new_new_n9634__ = ~new_new_n9632__ & ~new_new_n9633__;
  assign new_new_n9635__ = new_new_n9631__ & new_new_n9634__;
  assign new_new_n9636__ = ~new_new_n9631__ & ~new_new_n9634__;
  assign new_new_n9637__ = ~new_new_n9635__ & ~new_new_n9636__;
  assign new_new_n9638__ = ~pi073 & new_new_n9637__;
  assign new_new_n9639__ = pi073 & ~new_new_n9637__;
  assign new_new_n9640__ = ~new_new_n9203__ & ~new_new_n9204__;
  assign new_new_n9641__ = ~new_new_n9289__ & po024;
  assign new_new_n9642__ = pi071 & ~po024;
  assign new_new_n9643__ = ~new_new_n9641__ & ~new_new_n9642__;
  assign new_new_n9644__ = new_new_n9640__ & ~new_new_n9643__;
  assign new_new_n9645__ = ~new_new_n9640__ & new_new_n9643__;
  assign new_new_n9646__ = ~new_new_n9644__ & ~new_new_n9645__;
  assign new_new_n9647__ = ~pi072 & ~new_new_n9646__;
  assign new_new_n9648__ = pi072 & new_new_n9646__;
  assign new_new_n9649__ = ~new_new_n9279__ & ~new_new_n9280__;
  assign new_new_n9650__ = po024 & new_new_n9649__;
  assign new_new_n9651__ = ~new_new_n9287__ & ~new_new_n9650__;
  assign new_new_n9652__ = new_new_n9287__ & new_new_n9650__;
  assign new_new_n9653__ = ~new_new_n9651__ & ~new_new_n9652__;
  assign new_new_n9654__ = pi071 & ~new_new_n9653__;
  assign new_new_n9655__ = ~pi071 & new_new_n9653__;
  assign new_new_n9656__ = ~new_new_n9212__ & ~new_new_n9213__;
  assign new_new_n9657__ = ~new_new_n9276__ & po024;
  assign new_new_n9658__ = pi069 & ~po024;
  assign new_new_n9659__ = ~new_new_n9657__ & ~new_new_n9658__;
  assign new_new_n9660__ = new_new_n9656__ & new_new_n9659__;
  assign new_new_n9661__ = ~new_new_n9656__ & ~new_new_n9659__;
  assign new_new_n9662__ = ~new_new_n9660__ & ~new_new_n9661__;
  assign new_new_n9663__ = ~pi070 & new_new_n9662__;
  assign new_new_n9664__ = pi070 & ~new_new_n9662__;
  assign new_new_n9665__ = ~new_new_n9266__ & ~new_new_n9267__;
  assign new_new_n9666__ = po024 & new_new_n9665__;
  assign new_new_n9667__ = ~new_new_n9274__ & ~new_new_n9666__;
  assign new_new_n9668__ = new_new_n9274__ & new_new_n9666__;
  assign new_new_n9669__ = ~new_new_n9667__ & ~new_new_n9668__;
  assign new_new_n9670__ = pi069 & new_new_n9669__;
  assign new_new_n9671__ = ~new_new_n9219__ & ~new_new_n9220__;
  assign new_new_n9672__ = ~new_new_n9263__ & po024;
  assign new_new_n9673__ = pi067 & ~po024;
  assign new_new_n9674__ = ~new_new_n9672__ & ~new_new_n9673__;
  assign new_new_n9675__ = new_new_n9671__ & ~new_new_n9674__;
  assign new_new_n9676__ = ~new_new_n9671__ & new_new_n9674__;
  assign new_new_n9677__ = ~new_new_n9675__ & ~new_new_n9676__;
  assign new_new_n9678__ = ~pi068 & ~new_new_n9677__;
  assign new_new_n9679__ = pi068 & new_new_n9677__;
  assign new_new_n9680__ = ~new_new_n9233__ & po024;
  assign new_new_n9681__ = ~new_new_n9261__ & new_new_n9680__;
  assign new_new_n9682__ = new_new_n9260__ & ~new_new_n9681__;
  assign new_new_n9683__ = new_new_n9262__ & new_new_n9680__;
  assign new_new_n9684__ = ~new_new_n9682__ & ~new_new_n9683__;
  assign new_new_n9685__ = ~pi067 & ~new_new_n9684__;
  assign new_new_n9686__ = pi067 & new_new_n9684__;
  assign new_new_n9687__ = pi024 & po024;
  assign new_new_n9688__ = pi023 & ~pi065;
  assign new_new_n9689__ = new_new_n9687__ & ~new_new_n9688__;
  assign new_new_n9690__ = ~pi024 & ~po024;
  assign new_new_n9691__ = ~pi065 & ~new_new_n9690__;
  assign new_new_n9692__ = ~pi023 & ~new_new_n9691__;
  assign new_new_n9693__ = ~new_new_n9689__ & ~new_new_n9692__;
  assign new_new_n9694__ = pi064 & ~new_new_n9693__;
  assign new_new_n9695__ = pi064 & po024;
  assign new_new_n9696__ = ~pi024 & pi065;
  assign new_new_n9697__ = ~new_new_n9695__ & new_new_n9696__;
  assign new_new_n9698__ = ~new_new_n9694__ & ~new_new_n9697__;
  assign new_new_n9699__ = pi066 & ~new_new_n9698__;
  assign new_new_n9700__ = ~pi066 & new_new_n9698__;
  assign new_new_n9701__ = new_new_n426__ & ~po025;
  assign new_new_n9702__ = new_new_n9249__ & po024;
  assign new_new_n9703__ = ~new_new_n9701__ & ~new_new_n9702__;
  assign new_new_n9704__ = ~pi024 & ~new_new_n9703__;
  assign new_new_n9705__ = ~new_new_n332__ & po024;
  assign new_new_n9706__ = ~new_new_n9229__ & ~new_new_n9705__;
  assign new_new_n9707__ = pi065 & po024;
  assign new_new_n9708__ = po025 & ~new_new_n9707__;
  assign new_new_n9709__ = pi065 & ~new_new_n9229__;
  assign new_new_n9710__ = pi024 & ~new_new_n9709__;
  assign new_new_n9711__ = ~new_new_n9708__ & new_new_n9710__;
  assign new_new_n9712__ = ~new_new_n9704__ & ~new_new_n9706__;
  assign new_new_n9713__ = ~new_new_n9711__ & new_new_n9712__;
  assign new_new_n9714__ = ~pi025 & ~new_new_n9713__;
  assign new_new_n9715__ = ~new_new_n9229__ & ~new_new_n9707__;
  assign new_new_n9716__ = pi024 & ~new_new_n9240__;
  assign new_new_n9717__ = pi064 & ~new_new_n9716__;
  assign new_new_n9718__ = ~new_new_n9715__ & ~new_new_n9717__;
  assign new_new_n9719__ = ~pi065 & po024;
  assign new_new_n9720__ = ~po025 & ~new_new_n9719__;
  assign new_new_n9721__ = pi064 & ~new_new_n9687__;
  assign new_new_n9722__ = ~new_new_n9702__ & new_new_n9721__;
  assign new_new_n9723__ = ~new_new_n9720__ & new_new_n9722__;
  assign new_new_n9724__ = ~new_new_n9718__ & ~new_new_n9723__;
  assign new_new_n9725__ = pi025 & ~new_new_n9724__;
  assign new_new_n9726__ = ~new_new_n9714__ & ~new_new_n9725__;
  assign new_new_n9727__ = ~new_new_n9700__ & ~new_new_n9726__;
  assign new_new_n9728__ = ~new_new_n9699__ & ~new_new_n9727__;
  assign new_new_n9729__ = ~new_new_n9686__ & new_new_n9728__;
  assign new_new_n9730__ = ~new_new_n9685__ & ~new_new_n9729__;
  assign new_new_n9731__ = ~new_new_n9679__ & ~new_new_n9730__;
  assign new_new_n9732__ = ~new_new_n9678__ & ~new_new_n9731__;
  assign new_new_n9733__ = ~new_new_n9670__ & ~new_new_n9732__;
  assign new_new_n9734__ = ~pi069 & ~new_new_n9669__;
  assign new_new_n9735__ = ~new_new_n9733__ & ~new_new_n9734__;
  assign new_new_n9736__ = ~new_new_n9664__ & ~new_new_n9735__;
  assign new_new_n9737__ = ~new_new_n9663__ & ~new_new_n9736__;
  assign new_new_n9738__ = ~new_new_n9655__ & new_new_n9737__;
  assign new_new_n9739__ = ~new_new_n9654__ & ~new_new_n9738__;
  assign new_new_n9740__ = ~new_new_n9648__ & new_new_n9739__;
  assign new_new_n9741__ = ~new_new_n9647__ & ~new_new_n9740__;
  assign new_new_n9742__ = ~new_new_n9639__ & ~new_new_n9741__;
  assign new_new_n9743__ = ~new_new_n9638__ & ~new_new_n9742__;
  assign new_new_n9744__ = ~new_new_n9630__ & ~new_new_n9743__;
  assign new_new_n9745__ = ~new_new_n9629__ & ~new_new_n9744__;
  assign new_new_n9746__ = ~pi075 & new_new_n9620__;
  assign new_new_n9747__ = new_new_n9745__ & ~new_new_n9746__;
  assign new_new_n9748__ = ~new_new_n9621__ & ~new_new_n9747__;
  assign new_new_n9749__ = ~new_new_n9613__ & new_new_n9748__;
  assign new_new_n9750__ = ~new_new_n9612__ & ~new_new_n9749__;
  assign new_new_n9751__ = ~new_new_n9604__ & new_new_n9750__;
  assign new_new_n9752__ = ~new_new_n9603__ & ~new_new_n9751__;
  assign new_new_n9753__ = ~new_new_n9595__ & ~new_new_n9752__;
  assign new_new_n9754__ = ~new_new_n9594__ & ~new_new_n9753__;
  assign new_new_n9755__ = ~new_new_n9586__ & new_new_n9754__;
  assign new_new_n9756__ = ~new_new_n9585__ & ~new_new_n9755__;
  assign new_new_n9757__ = ~new_new_n9577__ & new_new_n9756__;
  assign new_new_n9758__ = ~new_new_n9576__ & ~new_new_n9757__;
  assign new_new_n9759__ = ~new_new_n9568__ & ~new_new_n9758__;
  assign new_new_n9760__ = ~new_new_n9567__ & ~new_new_n9759__;
  assign new_new_n9761__ = ~new_new_n9559__ & new_new_n9760__;
  assign new_new_n9762__ = ~new_new_n9558__ & ~new_new_n9761__;
  assign new_new_n9763__ = ~new_new_n9550__ & ~new_new_n9762__;
  assign new_new_n9764__ = ~new_new_n9549__ & ~new_new_n9763__;
  assign new_new_n9765__ = ~new_new_n9541__ & ~new_new_n9764__;
  assign new_new_n9766__ = ~new_new_n9540__ & ~new_new_n9765__;
  assign new_new_n9767__ = ~new_new_n9532__ & ~new_new_n9766__;
  assign new_new_n9768__ = ~new_new_n9531__ & ~new_new_n9767__;
  assign new_new_n9769__ = ~new_new_n9523__ & ~new_new_n9768__;
  assign new_new_n9770__ = ~new_new_n9522__ & ~new_new_n9769__;
  assign new_new_n9771__ = ~new_new_n9514__ & ~new_new_n9770__;
  assign new_new_n9772__ = ~new_new_n9513__ & ~new_new_n9771__;
  assign new_new_n9773__ = ~new_new_n9505__ & ~new_new_n9772__;
  assign new_new_n9774__ = ~new_new_n9504__ & ~new_new_n9773__;
  assign new_new_n9775__ = ~new_new_n9496__ & ~new_new_n9774__;
  assign new_new_n9776__ = ~new_new_n9495__ & ~new_new_n9775__;
  assign new_new_n9777__ = ~new_new_n9487__ & ~new_new_n9776__;
  assign new_new_n9778__ = ~new_new_n9486__ & ~new_new_n9777__;
  assign new_new_n9779__ = ~new_new_n9478__ & ~new_new_n9778__;
  assign new_new_n9780__ = ~new_new_n9477__ & ~new_new_n9779__;
  assign new_new_n9781__ = ~new_new_n9469__ & ~new_new_n9780__;
  assign new_new_n9782__ = ~new_new_n9468__ & ~new_new_n9781__;
  assign new_new_n9783__ = ~new_new_n9460__ & new_new_n9782__;
  assign new_new_n9784__ = ~new_new_n9459__ & ~new_new_n9783__;
  assign new_new_n9785__ = ~new_new_n9451__ & ~new_new_n9784__;
  assign new_new_n9786__ = ~new_new_n9450__ & ~new_new_n9785__;
  assign new_new_n9787__ = ~new_new_n9442__ & ~new_new_n9786__;
  assign new_new_n9788__ = ~new_new_n9441__ & ~new_new_n9787__;
  assign new_new_n9789__ = ~new_new_n9433__ & new_new_n9788__;
  assign new_new_n9790__ = ~new_new_n9432__ & ~new_new_n9789__;
  assign new_new_n9791__ = ~new_new_n9424__ & ~new_new_n9790__;
  assign new_new_n9792__ = ~new_new_n9423__ & ~new_new_n9791__;
  assign new_new_n9793__ = ~new_new_n9415__ & new_new_n9792__;
  assign new_new_n9794__ = ~new_new_n9414__ & ~new_new_n9793__;
  assign new_new_n9795__ = ~new_new_n9406__ & ~new_new_n9794__;
  assign new_new_n9796__ = ~new_new_n9405__ & ~new_new_n9795__;
  assign new_new_n9797__ = ~new_new_n9397__ & new_new_n9796__;
  assign new_new_n9798__ = ~new_new_n9396__ & ~new_new_n9797__;
  assign new_new_n9799__ = ~new_new_n9388__ & new_new_n9798__;
  assign new_new_n9800__ = ~new_new_n9387__ & ~new_new_n9799__;
  assign new_new_n9801__ = ~new_new_n9379__ & ~new_new_n9800__;
  assign new_new_n9802__ = ~new_new_n9378__ & ~new_new_n9801__;
  assign new_new_n9803__ = ~new_new_n9370__ & ~new_new_n9802__;
  assign new_new_n9804__ = ~new_new_n9369__ & ~new_new_n9803__;
  assign new_new_n9805__ = pi104 & ~new_new_n9804__;
  assign new_new_n9806__ = ~new_new_n376__ & new_new_n8068__;
  assign new_new_n9807__ = ~new_new_n9805__ & new_new_n9806__;
  assign new_new_n9808__ = new_new_n9361__ & ~new_new_n9807__;
  assign new_new_n9809__ = ~new_new_n9369__ & ~new_new_n9370__;
  assign new_new_n9810__ = ~pi104 & new_new_n9361__;
  assign new_new_n9811__ = ~new_new_n9804__ & ~new_new_n9810__;
  assign new_new_n9812__ = pi104 & ~new_new_n9361__;
  assign new_new_n9813__ = new_new_n8068__ & ~new_new_n9812__;
  assign po023 = ~new_new_n9811__ & new_new_n9813__;
  assign new_new_n9815__ = ~new_new_n9802__ & po023;
  assign new_new_n9816__ = pi103 & ~po023;
  assign new_new_n9817__ = ~new_new_n9815__ & ~new_new_n9816__;
  assign new_new_n9818__ = new_new_n9809__ & ~new_new_n9817__;
  assign new_new_n9819__ = ~new_new_n9809__ & new_new_n9817__;
  assign new_new_n9820__ = ~new_new_n9818__ & ~new_new_n9819__;
  assign new_new_n9821__ = pi104 & new_new_n9820__;
  assign new_new_n9822__ = ~pi104 & ~new_new_n9820__;
  assign new_new_n9823__ = ~new_new_n9821__ & ~new_new_n9822__;
  assign new_new_n9824__ = ~new_new_n9800__ & po023;
  assign new_new_n9825__ = pi102 & ~po023;
  assign new_new_n9826__ = ~new_new_n9824__ & ~new_new_n9825__;
  assign new_new_n9827__ = ~new_new_n9378__ & ~new_new_n9379__;
  assign new_new_n9828__ = ~new_new_n9826__ & new_new_n9827__;
  assign new_new_n9829__ = new_new_n9826__ & ~new_new_n9827__;
  assign new_new_n9830__ = ~new_new_n9828__ & ~new_new_n9829__;
  assign new_new_n9831__ = pi103 & new_new_n9830__;
  assign new_new_n9832__ = ~pi103 & ~new_new_n9830__;
  assign new_new_n9833__ = ~new_new_n9387__ & ~new_new_n9388__;
  assign new_new_n9834__ = ~new_new_n9798__ & po023;
  assign new_new_n9835__ = ~pi101 & ~po023;
  assign new_new_n9836__ = ~new_new_n9834__ & ~new_new_n9835__;
  assign new_new_n9837__ = new_new_n9833__ & ~new_new_n9836__;
  assign new_new_n9838__ = ~new_new_n9833__ & new_new_n9836__;
  assign new_new_n9839__ = ~new_new_n9837__ & ~new_new_n9838__;
  assign new_new_n9840__ = pi102 & ~new_new_n9839__;
  assign new_new_n9841__ = ~pi102 & new_new_n9839__;
  assign new_new_n9842__ = new_new_n9796__ & po023;
  assign new_new_n9843__ = ~pi100 & ~po023;
  assign new_new_n9844__ = ~new_new_n9842__ & ~new_new_n9843__;
  assign new_new_n9845__ = ~new_new_n9396__ & ~new_new_n9397__;
  assign new_new_n9846__ = ~new_new_n9844__ & ~new_new_n9845__;
  assign new_new_n9847__ = new_new_n9844__ & new_new_n9845__;
  assign new_new_n9848__ = ~new_new_n9846__ & ~new_new_n9847__;
  assign new_new_n9849__ = pi101 & new_new_n9848__;
  assign new_new_n9850__ = ~pi101 & ~new_new_n9848__;
  assign new_new_n9851__ = pi099 & ~new_new_n9794__;
  assign new_new_n9852__ = ~pi099 & new_new_n9794__;
  assign new_new_n9853__ = ~new_new_n9851__ & ~new_new_n9852__;
  assign new_new_n9854__ = po023 & new_new_n9853__;
  assign new_new_n9855__ = new_new_n9404__ & new_new_n9854__;
  assign new_new_n9856__ = ~new_new_n9404__ & ~new_new_n9854__;
  assign new_new_n9857__ = ~new_new_n9855__ & ~new_new_n9856__;
  assign new_new_n9858__ = pi100 & ~new_new_n9857__;
  assign new_new_n9859__ = ~pi100 & new_new_n9857__;
  assign new_new_n9860__ = ~new_new_n9414__ & ~new_new_n9415__;
  assign new_new_n9861__ = ~new_new_n9792__ & po023;
  assign new_new_n9862__ = ~pi098 & ~po023;
  assign new_new_n9863__ = ~new_new_n9861__ & ~new_new_n9862__;
  assign new_new_n9864__ = new_new_n9860__ & ~new_new_n9863__;
  assign new_new_n9865__ = ~new_new_n9860__ & new_new_n9863__;
  assign new_new_n9866__ = ~new_new_n9864__ & ~new_new_n9865__;
  assign new_new_n9867__ = ~pi099 & new_new_n9866__;
  assign new_new_n9868__ = pi099 & ~new_new_n9866__;
  assign new_new_n9869__ = ~pi097 & ~new_new_n9790__;
  assign new_new_n9870__ = pi097 & new_new_n9790__;
  assign new_new_n9871__ = ~new_new_n9869__ & ~new_new_n9870__;
  assign new_new_n9872__ = po023 & new_new_n9871__;
  assign new_new_n9873__ = new_new_n9422__ & new_new_n9872__;
  assign new_new_n9874__ = ~new_new_n9422__ & ~new_new_n9872__;
  assign new_new_n9875__ = ~new_new_n9873__ & ~new_new_n9874__;
  assign new_new_n9876__ = ~pi098 & ~new_new_n9875__;
  assign new_new_n9877__ = pi098 & new_new_n9875__;
  assign new_new_n9878__ = new_new_n9788__ & po023;
  assign new_new_n9879__ = ~pi096 & ~po023;
  assign new_new_n9880__ = ~new_new_n9878__ & ~new_new_n9879__;
  assign new_new_n9881__ = ~new_new_n9432__ & ~new_new_n9433__;
  assign new_new_n9882__ = ~new_new_n9880__ & ~new_new_n9881__;
  assign new_new_n9883__ = new_new_n9880__ & new_new_n9881__;
  assign new_new_n9884__ = ~new_new_n9882__ & ~new_new_n9883__;
  assign new_new_n9885__ = ~pi097 & ~new_new_n9884__;
  assign new_new_n9886__ = pi097 & new_new_n9884__;
  assign new_new_n9887__ = ~new_new_n9441__ & ~new_new_n9442__;
  assign new_new_n9888__ = ~new_new_n9786__ & po023;
  assign new_new_n9889__ = pi095 & ~po023;
  assign new_new_n9890__ = ~new_new_n9888__ & ~new_new_n9889__;
  assign new_new_n9891__ = new_new_n9887__ & ~new_new_n9890__;
  assign new_new_n9892__ = ~new_new_n9887__ & new_new_n9890__;
  assign new_new_n9893__ = ~new_new_n9891__ & ~new_new_n9892__;
  assign new_new_n9894__ = ~pi096 & ~new_new_n9893__;
  assign new_new_n9895__ = pi096 & new_new_n9893__;
  assign new_new_n9896__ = ~new_new_n9784__ & po023;
  assign new_new_n9897__ = pi094 & ~po023;
  assign new_new_n9898__ = ~new_new_n9896__ & ~new_new_n9897__;
  assign new_new_n9899__ = ~new_new_n9450__ & ~new_new_n9451__;
  assign new_new_n9900__ = ~new_new_n9898__ & new_new_n9899__;
  assign new_new_n9901__ = new_new_n9898__ & ~new_new_n9899__;
  assign new_new_n9902__ = ~new_new_n9900__ & ~new_new_n9901__;
  assign new_new_n9903__ = pi095 & new_new_n9902__;
  assign new_new_n9904__ = ~pi095 & ~new_new_n9902__;
  assign new_new_n9905__ = ~new_new_n9459__ & ~new_new_n9460__;
  assign new_new_n9906__ = ~new_new_n9782__ & po023;
  assign new_new_n9907__ = ~pi093 & ~po023;
  assign new_new_n9908__ = ~new_new_n9906__ & ~new_new_n9907__;
  assign new_new_n9909__ = new_new_n9905__ & ~new_new_n9908__;
  assign new_new_n9910__ = ~new_new_n9905__ & new_new_n9908__;
  assign new_new_n9911__ = ~new_new_n9909__ & ~new_new_n9910__;
  assign new_new_n9912__ = pi094 & ~new_new_n9911__;
  assign new_new_n9913__ = ~pi094 & new_new_n9911__;
  assign new_new_n9914__ = ~new_new_n9468__ & ~new_new_n9469__;
  assign new_new_n9915__ = ~new_new_n9780__ & po023;
  assign new_new_n9916__ = ~pi092 & ~po023;
  assign new_new_n9917__ = ~new_new_n9915__ & ~new_new_n9916__;
  assign new_new_n9918__ = new_new_n9914__ & ~new_new_n9917__;
  assign new_new_n9919__ = ~new_new_n9914__ & new_new_n9917__;
  assign new_new_n9920__ = ~new_new_n9918__ & ~new_new_n9919__;
  assign new_new_n9921__ = pi093 & ~new_new_n9920__;
  assign new_new_n9922__ = ~pi093 & new_new_n9920__;
  assign new_new_n9923__ = ~new_new_n9477__ & ~new_new_n9478__;
  assign new_new_n9924__ = ~new_new_n9778__ & po023;
  assign new_new_n9925__ = ~pi091 & ~po023;
  assign new_new_n9926__ = ~new_new_n9924__ & ~new_new_n9925__;
  assign new_new_n9927__ = new_new_n9923__ & ~new_new_n9926__;
  assign new_new_n9928__ = ~new_new_n9923__ & new_new_n9926__;
  assign new_new_n9929__ = ~new_new_n9927__ & ~new_new_n9928__;
  assign new_new_n9930__ = pi092 & ~new_new_n9929__;
  assign new_new_n9931__ = ~pi092 & new_new_n9929__;
  assign new_new_n9932__ = ~pi090 & ~new_new_n9776__;
  assign new_new_n9933__ = pi090 & new_new_n9776__;
  assign new_new_n9934__ = ~new_new_n9932__ & ~new_new_n9933__;
  assign new_new_n9935__ = po023 & new_new_n9934__;
  assign new_new_n9936__ = ~new_new_n9485__ & ~new_new_n9935__;
  assign new_new_n9937__ = new_new_n9485__ & new_new_n9935__;
  assign new_new_n9938__ = ~new_new_n9936__ & ~new_new_n9937__;
  assign new_new_n9939__ = ~pi091 & ~new_new_n9938__;
  assign new_new_n9940__ = pi091 & new_new_n9938__;
  assign new_new_n9941__ = ~new_new_n9495__ & ~new_new_n9496__;
  assign new_new_n9942__ = ~new_new_n9774__ & po023;
  assign new_new_n9943__ = ~pi089 & ~po023;
  assign new_new_n9944__ = ~new_new_n9942__ & ~new_new_n9943__;
  assign new_new_n9945__ = new_new_n9941__ & ~new_new_n9944__;
  assign new_new_n9946__ = ~new_new_n9941__ & new_new_n9944__;
  assign new_new_n9947__ = ~new_new_n9945__ & ~new_new_n9946__;
  assign new_new_n9948__ = pi090 & ~new_new_n9947__;
  assign new_new_n9949__ = ~pi090 & new_new_n9947__;
  assign new_new_n9950__ = ~new_new_n9504__ & ~new_new_n9505__;
  assign new_new_n9951__ = ~new_new_n9772__ & po023;
  assign new_new_n9952__ = ~pi088 & ~po023;
  assign new_new_n9953__ = ~new_new_n9951__ & ~new_new_n9952__;
  assign new_new_n9954__ = ~new_new_n9950__ & ~new_new_n9953__;
  assign new_new_n9955__ = new_new_n9950__ & new_new_n9953__;
  assign new_new_n9956__ = ~new_new_n9954__ & ~new_new_n9955__;
  assign new_new_n9957__ = ~pi089 & ~new_new_n9956__;
  assign new_new_n9958__ = pi089 & new_new_n9956__;
  assign new_new_n9959__ = ~pi087 & ~new_new_n9770__;
  assign new_new_n9960__ = pi087 & new_new_n9770__;
  assign new_new_n9961__ = ~new_new_n9959__ & ~new_new_n9960__;
  assign new_new_n9962__ = po023 & new_new_n9961__;
  assign new_new_n9963__ = new_new_n9512__ & new_new_n9962__;
  assign new_new_n9964__ = ~new_new_n9512__ & ~new_new_n9962__;
  assign new_new_n9965__ = ~new_new_n9963__ & ~new_new_n9964__;
  assign new_new_n9966__ = ~pi088 & ~new_new_n9965__;
  assign new_new_n9967__ = pi088 & new_new_n9965__;
  assign new_new_n9968__ = ~new_new_n9522__ & ~new_new_n9523__;
  assign new_new_n9969__ = ~new_new_n9768__ & po023;
  assign new_new_n9970__ = ~pi086 & ~po023;
  assign new_new_n9971__ = ~new_new_n9969__ & ~new_new_n9970__;
  assign new_new_n9972__ = ~new_new_n9968__ & ~new_new_n9971__;
  assign new_new_n9973__ = new_new_n9968__ & new_new_n9971__;
  assign new_new_n9974__ = ~new_new_n9972__ & ~new_new_n9973__;
  assign new_new_n9975__ = ~pi087 & ~new_new_n9974__;
  assign new_new_n9976__ = pi087 & new_new_n9974__;
  assign new_new_n9977__ = ~pi085 & ~new_new_n9766__;
  assign new_new_n9978__ = pi085 & new_new_n9766__;
  assign new_new_n9979__ = ~new_new_n9977__ & ~new_new_n9978__;
  assign new_new_n9980__ = po023 & new_new_n9979__;
  assign new_new_n9981__ = new_new_n9530__ & new_new_n9980__;
  assign new_new_n9982__ = ~new_new_n9530__ & ~new_new_n9980__;
  assign new_new_n9983__ = ~new_new_n9981__ & ~new_new_n9982__;
  assign new_new_n9984__ = ~pi086 & ~new_new_n9983__;
  assign new_new_n9985__ = pi086 & new_new_n9983__;
  assign new_new_n9986__ = ~pi084 & ~new_new_n9764__;
  assign new_new_n9987__ = pi084 & new_new_n9764__;
  assign new_new_n9988__ = ~new_new_n9986__ & ~new_new_n9987__;
  assign new_new_n9989__ = po023 & new_new_n9988__;
  assign new_new_n9990__ = new_new_n9539__ & new_new_n9989__;
  assign new_new_n9991__ = ~new_new_n9539__ & ~new_new_n9989__;
  assign new_new_n9992__ = ~new_new_n9990__ & ~new_new_n9991__;
  assign new_new_n9993__ = ~pi085 & ~new_new_n9992__;
  assign new_new_n9994__ = pi085 & new_new_n9992__;
  assign new_new_n9995__ = ~new_new_n9549__ & ~new_new_n9550__;
  assign new_new_n9996__ = ~new_new_n9762__ & po023;
  assign new_new_n9997__ = ~pi083 & ~po023;
  assign new_new_n9998__ = ~new_new_n9996__ & ~new_new_n9997__;
  assign new_new_n9999__ = new_new_n9995__ & ~new_new_n9998__;
  assign new_new_n10000__ = ~new_new_n9995__ & new_new_n9998__;
  assign new_new_n10001__ = ~new_new_n9999__ & ~new_new_n10000__;
  assign new_new_n10002__ = ~pi084 & new_new_n10001__;
  assign new_new_n10003__ = pi084 & ~new_new_n10001__;
  assign new_new_n10004__ = ~new_new_n9760__ & po023;
  assign new_new_n10005__ = pi082 & ~po023;
  assign new_new_n10006__ = ~new_new_n10004__ & ~new_new_n10005__;
  assign new_new_n10007__ = ~new_new_n9558__ & ~new_new_n9559__;
  assign new_new_n10008__ = ~new_new_n10006__ & new_new_n10007__;
  assign new_new_n10009__ = new_new_n10006__ & ~new_new_n10007__;
  assign new_new_n10010__ = ~new_new_n10008__ & ~new_new_n10009__;
  assign new_new_n10011__ = ~pi083 & ~new_new_n10010__;
  assign new_new_n10012__ = pi083 & new_new_n10010__;
  assign new_new_n10013__ = ~new_new_n9567__ & ~new_new_n9568__;
  assign new_new_n10014__ = ~new_new_n9758__ & po023;
  assign new_new_n10015__ = pi081 & ~po023;
  assign new_new_n10016__ = ~new_new_n10014__ & ~new_new_n10015__;
  assign new_new_n10017__ = new_new_n10013__ & ~new_new_n10016__;
  assign new_new_n10018__ = ~new_new_n10013__ & new_new_n10016__;
  assign new_new_n10019__ = ~new_new_n10017__ & ~new_new_n10018__;
  assign new_new_n10020__ = ~pi082 & ~new_new_n10019__;
  assign new_new_n10021__ = pi082 & new_new_n10019__;
  assign new_new_n10022__ = ~new_new_n9576__ & ~new_new_n9577__;
  assign new_new_n10023__ = ~new_new_n9756__ & po023;
  assign new_new_n10024__ = ~pi080 & ~po023;
  assign new_new_n10025__ = ~new_new_n10023__ & ~new_new_n10024__;
  assign new_new_n10026__ = new_new_n10022__ & ~new_new_n10025__;
  assign new_new_n10027__ = ~new_new_n10022__ & new_new_n10025__;
  assign new_new_n10028__ = ~new_new_n10026__ & ~new_new_n10027__;
  assign new_new_n10029__ = ~pi081 & new_new_n10028__;
  assign new_new_n10030__ = pi081 & ~new_new_n10028__;
  assign new_new_n10031__ = ~new_new_n9585__ & ~new_new_n9586__;
  assign new_new_n10032__ = ~new_new_n9754__ & po023;
  assign new_new_n10033__ = pi079 & ~po023;
  assign new_new_n10034__ = ~new_new_n10032__ & ~new_new_n10033__;
  assign new_new_n10035__ = new_new_n10031__ & ~new_new_n10034__;
  assign new_new_n10036__ = ~new_new_n10031__ & new_new_n10034__;
  assign new_new_n10037__ = ~new_new_n10035__ & ~new_new_n10036__;
  assign new_new_n10038__ = ~pi080 & ~new_new_n10037__;
  assign new_new_n10039__ = pi080 & new_new_n10037__;
  assign new_new_n10040__ = ~new_new_n9752__ & po023;
  assign new_new_n10041__ = pi078 & ~po023;
  assign new_new_n10042__ = ~new_new_n10040__ & ~new_new_n10041__;
  assign new_new_n10043__ = ~new_new_n9594__ & ~new_new_n9595__;
  assign new_new_n10044__ = ~new_new_n10042__ & new_new_n10043__;
  assign new_new_n10045__ = new_new_n10042__ & ~new_new_n10043__;
  assign new_new_n10046__ = ~new_new_n10044__ & ~new_new_n10045__;
  assign new_new_n10047__ = ~pi079 & ~new_new_n10046__;
  assign new_new_n10048__ = pi079 & new_new_n10046__;
  assign new_new_n10049__ = ~new_new_n9603__ & ~new_new_n9604__;
  assign new_new_n10050__ = ~new_new_n9750__ & po023;
  assign new_new_n10051__ = ~pi077 & ~po023;
  assign new_new_n10052__ = ~new_new_n10050__ & ~new_new_n10051__;
  assign new_new_n10053__ = new_new_n10049__ & ~new_new_n10052__;
  assign new_new_n10054__ = ~new_new_n10049__ & new_new_n10052__;
  assign new_new_n10055__ = ~new_new_n10053__ & ~new_new_n10054__;
  assign new_new_n10056__ = pi078 & ~new_new_n10055__;
  assign new_new_n10057__ = ~pi078 & new_new_n10055__;
  assign new_new_n10058__ = ~new_new_n9748__ & po023;
  assign new_new_n10059__ = pi076 & ~po023;
  assign new_new_n10060__ = ~new_new_n10058__ & ~new_new_n10059__;
  assign new_new_n10061__ = ~new_new_n9612__ & ~new_new_n9613__;
  assign new_new_n10062__ = ~new_new_n10060__ & new_new_n10061__;
  assign new_new_n10063__ = new_new_n10060__ & ~new_new_n10061__;
  assign new_new_n10064__ = ~new_new_n10062__ & ~new_new_n10063__;
  assign new_new_n10065__ = pi077 & new_new_n10064__;
  assign new_new_n10066__ = ~pi077 & ~new_new_n10064__;
  assign new_new_n10067__ = ~new_new_n9621__ & ~new_new_n9746__;
  assign new_new_n10068__ = ~new_new_n9745__ & po023;
  assign new_new_n10069__ = ~pi075 & ~po023;
  assign new_new_n10070__ = ~new_new_n10068__ & ~new_new_n10069__;
  assign new_new_n10071__ = new_new_n10067__ & ~new_new_n10070__;
  assign new_new_n10072__ = ~new_new_n10067__ & new_new_n10070__;
  assign new_new_n10073__ = ~new_new_n10071__ & ~new_new_n10072__;
  assign new_new_n10074__ = pi076 & ~new_new_n10073__;
  assign new_new_n10075__ = ~pi076 & new_new_n10073__;
  assign new_new_n10076__ = ~pi074 & ~new_new_n9743__;
  assign new_new_n10077__ = pi074 & new_new_n9743__;
  assign new_new_n10078__ = ~new_new_n10076__ & ~new_new_n10077__;
  assign new_new_n10079__ = po023 & new_new_n10078__;
  assign new_new_n10080__ = new_new_n9628__ & new_new_n10079__;
  assign new_new_n10081__ = ~new_new_n9628__ & ~new_new_n10079__;
  assign new_new_n10082__ = ~new_new_n10080__ & ~new_new_n10081__;
  assign new_new_n10083__ = ~pi075 & ~new_new_n10082__;
  assign new_new_n10084__ = pi075 & new_new_n10082__;
  assign new_new_n10085__ = ~new_new_n9638__ & ~new_new_n9639__;
  assign new_new_n10086__ = ~new_new_n9741__ & po023;
  assign new_new_n10087__ = ~pi073 & ~po023;
  assign new_new_n10088__ = ~new_new_n10086__ & ~new_new_n10087__;
  assign new_new_n10089__ = new_new_n10085__ & ~new_new_n10088__;
  assign new_new_n10090__ = ~new_new_n10085__ & new_new_n10088__;
  assign new_new_n10091__ = ~new_new_n10089__ & ~new_new_n10090__;
  assign new_new_n10092__ = ~pi074 & new_new_n10091__;
  assign new_new_n10093__ = pi074 & ~new_new_n10091__;
  assign new_new_n10094__ = ~new_new_n9739__ & po023;
  assign new_new_n10095__ = pi072 & ~po023;
  assign new_new_n10096__ = ~new_new_n10094__ & ~new_new_n10095__;
  assign new_new_n10097__ = ~new_new_n9647__ & ~new_new_n9648__;
  assign new_new_n10098__ = ~new_new_n10096__ & new_new_n10097__;
  assign new_new_n10099__ = new_new_n10096__ & ~new_new_n10097__;
  assign new_new_n10100__ = ~new_new_n10098__ & ~new_new_n10099__;
  assign new_new_n10101__ = ~pi073 & ~new_new_n10100__;
  assign new_new_n10102__ = pi073 & new_new_n10100__;
  assign new_new_n10103__ = ~new_new_n9654__ & ~new_new_n9655__;
  assign new_new_n10104__ = ~new_new_n9737__ & po023;
  assign new_new_n10105__ = ~pi071 & ~po023;
  assign new_new_n10106__ = ~new_new_n10104__ & ~new_new_n10105__;
  assign new_new_n10107__ = new_new_n10103__ & new_new_n10106__;
  assign new_new_n10108__ = ~new_new_n10103__ & ~new_new_n10106__;
  assign new_new_n10109__ = ~new_new_n10107__ & ~new_new_n10108__;
  assign new_new_n10110__ = pi072 & new_new_n10109__;
  assign new_new_n10111__ = ~pi072 & ~new_new_n10109__;
  assign new_new_n10112__ = new_new_n9735__ & po023;
  assign new_new_n10113__ = pi070 & ~po023;
  assign new_new_n10114__ = ~new_new_n10112__ & ~new_new_n10113__;
  assign new_new_n10115__ = ~new_new_n9663__ & ~new_new_n9664__;
  assign new_new_n10116__ = ~new_new_n10114__ & ~new_new_n10115__;
  assign new_new_n10117__ = new_new_n10114__ & new_new_n10115__;
  assign new_new_n10118__ = ~new_new_n10116__ & ~new_new_n10117__;
  assign new_new_n10119__ = pi071 & ~new_new_n10118__;
  assign new_new_n10120__ = ~pi071 & new_new_n10118__;
  assign new_new_n10121__ = ~new_new_n9670__ & ~new_new_n9734__;
  assign new_new_n10122__ = ~new_new_n9732__ & po023;
  assign new_new_n10123__ = ~pi069 & ~po023;
  assign new_new_n10124__ = ~new_new_n10122__ & ~new_new_n10123__;
  assign new_new_n10125__ = new_new_n10121__ & ~new_new_n10124__;
  assign new_new_n10126__ = ~new_new_n10121__ & new_new_n10124__;
  assign new_new_n10127__ = ~new_new_n10125__ & ~new_new_n10126__;
  assign new_new_n10128__ = pi070 & ~new_new_n10127__;
  assign new_new_n10129__ = ~pi070 & new_new_n10127__;
  assign new_new_n10130__ = ~new_new_n9678__ & ~new_new_n9679__;
  assign new_new_n10131__ = ~new_new_n9730__ & po023;
  assign new_new_n10132__ = ~pi068 & ~po023;
  assign new_new_n10133__ = ~new_new_n10131__ & ~new_new_n10132__;
  assign new_new_n10134__ = new_new_n10130__ & ~new_new_n10133__;
  assign new_new_n10135__ = ~new_new_n10130__ & new_new_n10133__;
  assign new_new_n10136__ = ~new_new_n10134__ & ~new_new_n10135__;
  assign new_new_n10137__ = pi069 & ~new_new_n10136__;
  assign new_new_n10138__ = ~pi069 & new_new_n10136__;
  assign new_new_n10139__ = ~new_new_n9699__ & ~new_new_n9700__;
  assign new_new_n10140__ = po023 & new_new_n10139__;
  assign new_new_n10141__ = new_new_n9726__ & ~new_new_n10140__;
  assign new_new_n10142__ = ~new_new_n9726__ & new_new_n10140__;
  assign new_new_n10143__ = ~new_new_n10141__ & ~new_new_n10142__;
  assign new_new_n10144__ = ~pi067 & ~new_new_n10143__;
  assign new_new_n10145__ = pi067 & new_new_n10143__;
  assign new_new_n10146__ = ~pi022 & pi064;
  assign new_new_n10147__ = pi064 & po023;
  assign new_new_n10148__ = ~pi023 & ~new_new_n10147__;
  assign new_new_n10149__ = pi023 & po023;
  assign new_new_n10150__ = pi064 & new_new_n10149__;
  assign new_new_n10151__ = ~new_new_n10148__ & ~new_new_n10150__;
  assign new_new_n10152__ = pi065 & ~new_new_n10151__;
  assign new_new_n10153__ = ~new_new_n10146__ & ~new_new_n10152__;
  assign new_new_n10154__ = ~pi065 & new_new_n10151__;
  assign new_new_n10155__ = ~new_new_n10153__ & ~new_new_n10154__;
  assign new_new_n10156__ = ~pi066 & ~new_new_n10155__;
  assign new_new_n10157__ = pi066 & new_new_n10155__;
  assign new_new_n10158__ = new_new_n426__ & ~po024;
  assign new_new_n10159__ = new_new_n9719__ & po023;
  assign new_new_n10160__ = ~new_new_n10158__ & ~new_new_n10159__;
  assign new_new_n10161__ = ~pi023 & ~new_new_n10160__;
  assign new_new_n10162__ = ~new_new_n332__ & po023;
  assign new_new_n10163__ = ~new_new_n9695__ & ~new_new_n10162__;
  assign new_new_n10164__ = pi065 & po023;
  assign new_new_n10165__ = po024 & ~new_new_n10164__;
  assign new_new_n10166__ = pi065 & ~new_new_n9695__;
  assign new_new_n10167__ = pi023 & ~new_new_n10166__;
  assign new_new_n10168__ = ~new_new_n10165__ & new_new_n10167__;
  assign new_new_n10169__ = ~new_new_n10161__ & ~new_new_n10163__;
  assign new_new_n10170__ = ~new_new_n10168__ & new_new_n10169__;
  assign new_new_n10171__ = ~pi024 & ~new_new_n10170__;
  assign new_new_n10172__ = ~new_new_n9695__ & ~new_new_n10164__;
  assign new_new_n10173__ = pi023 & ~new_new_n9707__;
  assign new_new_n10174__ = pi064 & ~new_new_n10173__;
  assign new_new_n10175__ = ~new_new_n10172__ & ~new_new_n10174__;
  assign new_new_n10176__ = pi064 & ~new_new_n10149__;
  assign new_new_n10177__ = ~pi065 & po023;
  assign new_new_n10178__ = ~po024 & ~new_new_n10177__;
  assign new_new_n10179__ = ~new_new_n10159__ & new_new_n10176__;
  assign new_new_n10180__ = ~new_new_n10178__ & new_new_n10179__;
  assign new_new_n10181__ = ~new_new_n10175__ & ~new_new_n10180__;
  assign new_new_n10182__ = pi024 & ~new_new_n10181__;
  assign new_new_n10183__ = ~new_new_n10171__ & ~new_new_n10182__;
  assign new_new_n10184__ = ~new_new_n10157__ & new_new_n10183__;
  assign new_new_n10185__ = ~new_new_n10156__ & ~new_new_n10184__;
  assign new_new_n10186__ = ~new_new_n10145__ & ~new_new_n10185__;
  assign new_new_n10187__ = ~new_new_n10144__ & ~new_new_n10186__;
  assign new_new_n10188__ = pi068 & new_new_n10187__;
  assign new_new_n10189__ = ~pi068 & ~new_new_n10187__;
  assign new_new_n10190__ = ~new_new_n9685__ & ~new_new_n9686__;
  assign new_new_n10191__ = ~new_new_n9728__ & po023;
  assign new_new_n10192__ = pi067 & ~po023;
  assign new_new_n10193__ = ~new_new_n10191__ & ~new_new_n10192__;
  assign new_new_n10194__ = new_new_n10190__ & ~new_new_n10193__;
  assign new_new_n10195__ = ~new_new_n10190__ & new_new_n10193__;
  assign new_new_n10196__ = ~new_new_n10194__ & ~new_new_n10195__;
  assign new_new_n10197__ = ~new_new_n10189__ & new_new_n10196__;
  assign new_new_n10198__ = ~new_new_n10188__ & ~new_new_n10197__;
  assign new_new_n10199__ = ~new_new_n10138__ & ~new_new_n10198__;
  assign new_new_n10200__ = ~new_new_n10137__ & ~new_new_n10199__;
  assign new_new_n10201__ = ~new_new_n10129__ & ~new_new_n10200__;
  assign new_new_n10202__ = ~new_new_n10128__ & ~new_new_n10201__;
  assign new_new_n10203__ = ~new_new_n10120__ & ~new_new_n10202__;
  assign new_new_n10204__ = ~new_new_n10119__ & ~new_new_n10203__;
  assign new_new_n10205__ = ~new_new_n10111__ & ~new_new_n10204__;
  assign new_new_n10206__ = ~new_new_n10110__ & ~new_new_n10205__;
  assign new_new_n10207__ = ~new_new_n10102__ & new_new_n10206__;
  assign new_new_n10208__ = ~new_new_n10101__ & ~new_new_n10207__;
  assign new_new_n10209__ = ~new_new_n10093__ & ~new_new_n10208__;
  assign new_new_n10210__ = ~new_new_n10092__ & ~new_new_n10209__;
  assign new_new_n10211__ = ~new_new_n10084__ & ~new_new_n10210__;
  assign new_new_n10212__ = ~new_new_n10083__ & ~new_new_n10211__;
  assign new_new_n10213__ = ~new_new_n10075__ & new_new_n10212__;
  assign new_new_n10214__ = ~new_new_n10074__ & ~new_new_n10213__;
  assign new_new_n10215__ = ~new_new_n10066__ & ~new_new_n10214__;
  assign new_new_n10216__ = ~new_new_n10065__ & ~new_new_n10215__;
  assign new_new_n10217__ = ~new_new_n10057__ & ~new_new_n10216__;
  assign new_new_n10218__ = ~new_new_n10056__ & ~new_new_n10217__;
  assign new_new_n10219__ = ~new_new_n10048__ & new_new_n10218__;
  assign new_new_n10220__ = ~new_new_n10047__ & ~new_new_n10219__;
  assign new_new_n10221__ = ~new_new_n10039__ & ~new_new_n10220__;
  assign new_new_n10222__ = ~new_new_n10038__ & ~new_new_n10221__;
  assign new_new_n10223__ = ~new_new_n10030__ & ~new_new_n10222__;
  assign new_new_n10224__ = ~new_new_n10029__ & ~new_new_n10223__;
  assign new_new_n10225__ = ~new_new_n10021__ & ~new_new_n10224__;
  assign new_new_n10226__ = ~new_new_n10020__ & ~new_new_n10225__;
  assign new_new_n10227__ = ~new_new_n10012__ & ~new_new_n10226__;
  assign new_new_n10228__ = ~new_new_n10011__ & ~new_new_n10227__;
  assign new_new_n10229__ = ~new_new_n10003__ & ~new_new_n10228__;
  assign new_new_n10230__ = ~new_new_n10002__ & ~new_new_n10229__;
  assign new_new_n10231__ = ~new_new_n9994__ & ~new_new_n10230__;
  assign new_new_n10232__ = ~new_new_n9993__ & ~new_new_n10231__;
  assign new_new_n10233__ = ~new_new_n9985__ & ~new_new_n10232__;
  assign new_new_n10234__ = ~new_new_n9984__ & ~new_new_n10233__;
  assign new_new_n10235__ = ~new_new_n9976__ & ~new_new_n10234__;
  assign new_new_n10236__ = ~new_new_n9975__ & ~new_new_n10235__;
  assign new_new_n10237__ = ~new_new_n9967__ & ~new_new_n10236__;
  assign new_new_n10238__ = ~new_new_n9966__ & ~new_new_n10237__;
  assign new_new_n10239__ = ~new_new_n9958__ & ~new_new_n10238__;
  assign new_new_n10240__ = ~new_new_n9957__ & ~new_new_n10239__;
  assign new_new_n10241__ = ~new_new_n9949__ & new_new_n10240__;
  assign new_new_n10242__ = ~new_new_n9948__ & ~new_new_n10241__;
  assign new_new_n10243__ = ~new_new_n9940__ & new_new_n10242__;
  assign new_new_n10244__ = ~new_new_n9939__ & ~new_new_n10243__;
  assign new_new_n10245__ = ~new_new_n9931__ & new_new_n10244__;
  assign new_new_n10246__ = ~new_new_n9930__ & ~new_new_n10245__;
  assign new_new_n10247__ = ~new_new_n9922__ & ~new_new_n10246__;
  assign new_new_n10248__ = ~new_new_n9921__ & ~new_new_n10247__;
  assign new_new_n10249__ = ~new_new_n9913__ & ~new_new_n10248__;
  assign new_new_n10250__ = ~new_new_n9912__ & ~new_new_n10249__;
  assign new_new_n10251__ = ~new_new_n9904__ & ~new_new_n10250__;
  assign new_new_n10252__ = ~new_new_n9903__ & ~new_new_n10251__;
  assign new_new_n10253__ = ~new_new_n9895__ & new_new_n10252__;
  assign new_new_n10254__ = ~new_new_n9894__ & ~new_new_n10253__;
  assign new_new_n10255__ = ~new_new_n9886__ & ~new_new_n10254__;
  assign new_new_n10256__ = ~new_new_n9885__ & ~new_new_n10255__;
  assign new_new_n10257__ = ~new_new_n9877__ & ~new_new_n10256__;
  assign new_new_n10258__ = ~new_new_n9876__ & ~new_new_n10257__;
  assign new_new_n10259__ = ~new_new_n9868__ & ~new_new_n10258__;
  assign new_new_n10260__ = ~new_new_n9867__ & ~new_new_n10259__;
  assign new_new_n10261__ = ~new_new_n9859__ & new_new_n10260__;
  assign new_new_n10262__ = ~new_new_n9858__ & ~new_new_n10261__;
  assign new_new_n10263__ = ~new_new_n9850__ & ~new_new_n10262__;
  assign new_new_n10264__ = ~new_new_n9849__ & ~new_new_n10263__;
  assign new_new_n10265__ = ~new_new_n9841__ & ~new_new_n10264__;
  assign new_new_n10266__ = ~new_new_n9840__ & ~new_new_n10265__;
  assign new_new_n10267__ = ~new_new_n9832__ & ~new_new_n10266__;
  assign new_new_n10268__ = ~new_new_n9831__ & ~new_new_n10267__;
  assign new_new_n10269__ = ~new_new_n9821__ & new_new_n10268__;
  assign new_new_n10270__ = ~new_new_n9822__ & ~new_new_n10269__;
  assign new_new_n10271__ = ~pi105 & ~new_new_n10270__;
  assign new_new_n10272__ = ~new_new_n9808__ & ~new_new_n10271__;
  assign new_new_n10273__ = pi105 & new_new_n10270__;
  assign new_new_n10274__ = ~pi106 & new_new_n279__;
  assign new_new_n10275__ = ~new_new_n10273__ & new_new_n10274__;
  assign po022 = ~new_new_n10272__ & new_new_n10275__;
  assign new_new_n10277__ = pi104 & ~po022;
  assign new_new_n10278__ = ~new_new_n10268__ & po022;
  assign new_new_n10279__ = ~new_new_n10277__ & ~new_new_n10278__;
  assign new_new_n10280__ = new_new_n9823__ & ~new_new_n10279__;
  assign new_new_n10281__ = ~new_new_n9823__ & new_new_n10279__;
  assign new_new_n10282__ = ~new_new_n10280__ & ~new_new_n10281__;
  assign new_new_n10283__ = pi105 & new_new_n10282__;
  assign new_new_n10284__ = ~pi105 & ~new_new_n10282__;
  assign new_new_n10285__ = ~new_new_n10266__ & po022;
  assign new_new_n10286__ = pi103 & ~po022;
  assign new_new_n10287__ = ~new_new_n10285__ & ~new_new_n10286__;
  assign new_new_n10288__ = ~new_new_n9831__ & ~new_new_n9832__;
  assign new_new_n10289__ = ~new_new_n10287__ & new_new_n10288__;
  assign new_new_n10290__ = new_new_n10287__ & ~new_new_n10288__;
  assign new_new_n10291__ = ~new_new_n10289__ & ~new_new_n10290__;
  assign new_new_n10292__ = ~pi104 & ~new_new_n10291__;
  assign new_new_n10293__ = pi104 & new_new_n10291__;
  assign new_new_n10294__ = pi102 & ~new_new_n10264__;
  assign new_new_n10295__ = ~pi102 & new_new_n10264__;
  assign new_new_n10296__ = ~new_new_n10294__ & ~new_new_n10295__;
  assign new_new_n10297__ = po022 & new_new_n10296__;
  assign new_new_n10298__ = new_new_n9839__ & new_new_n10297__;
  assign new_new_n10299__ = ~new_new_n9839__ & ~new_new_n10297__;
  assign new_new_n10300__ = ~new_new_n10298__ & ~new_new_n10299__;
  assign new_new_n10301__ = pi103 & ~new_new_n10300__;
  assign new_new_n10302__ = ~pi103 & new_new_n10300__;
  assign new_new_n10303__ = ~new_new_n9849__ & ~new_new_n9850__;
  assign new_new_n10304__ = new_new_n10262__ & po022;
  assign new_new_n10305__ = ~pi101 & ~po022;
  assign new_new_n10306__ = ~new_new_n10304__ & ~new_new_n10305__;
  assign new_new_n10307__ = ~new_new_n10303__ & ~new_new_n10306__;
  assign new_new_n10308__ = new_new_n10303__ & new_new_n10306__;
  assign new_new_n10309__ = ~new_new_n10307__ & ~new_new_n10308__;
  assign new_new_n10310__ = pi102 & new_new_n10309__;
  assign new_new_n10311__ = ~pi102 & ~new_new_n10309__;
  assign new_new_n10312__ = new_new_n10260__ & po022;
  assign new_new_n10313__ = pi100 & ~po022;
  assign new_new_n10314__ = ~new_new_n10312__ & ~new_new_n10313__;
  assign new_new_n10315__ = ~new_new_n9858__ & ~new_new_n9859__;
  assign new_new_n10316__ = ~new_new_n10314__ & ~new_new_n10315__;
  assign new_new_n10317__ = new_new_n10314__ & new_new_n10315__;
  assign new_new_n10318__ = ~new_new_n10316__ & ~new_new_n10317__;
  assign new_new_n10319__ = pi101 & ~new_new_n10318__;
  assign new_new_n10320__ = ~pi101 & new_new_n10318__;
  assign new_new_n10321__ = ~new_new_n9867__ & ~new_new_n9868__;
  assign new_new_n10322__ = ~new_new_n10258__ & po022;
  assign new_new_n10323__ = ~pi099 & ~po022;
  assign new_new_n10324__ = ~new_new_n10322__ & ~new_new_n10323__;
  assign new_new_n10325__ = new_new_n10321__ & ~new_new_n10324__;
  assign new_new_n10326__ = ~new_new_n10321__ & new_new_n10324__;
  assign new_new_n10327__ = ~new_new_n10325__ & ~new_new_n10326__;
  assign new_new_n10328__ = pi100 & ~new_new_n10327__;
  assign new_new_n10329__ = ~pi100 & new_new_n10327__;
  assign new_new_n10330__ = ~new_new_n9876__ & ~new_new_n9877__;
  assign new_new_n10331__ = ~new_new_n10256__ & po022;
  assign new_new_n10332__ = ~pi098 & ~po022;
  assign new_new_n10333__ = ~new_new_n10331__ & ~new_new_n10332__;
  assign new_new_n10334__ = new_new_n10330__ & ~new_new_n10333__;
  assign new_new_n10335__ = ~new_new_n10330__ & new_new_n10333__;
  assign new_new_n10336__ = ~new_new_n10334__ & ~new_new_n10335__;
  assign new_new_n10337__ = pi099 & ~new_new_n10336__;
  assign new_new_n10338__ = ~pi099 & new_new_n10336__;
  assign new_new_n10339__ = ~new_new_n9885__ & ~new_new_n9886__;
  assign new_new_n10340__ = ~new_new_n10254__ & po022;
  assign new_new_n10341__ = ~pi097 & ~po022;
  assign new_new_n10342__ = ~new_new_n10340__ & ~new_new_n10341__;
  assign new_new_n10343__ = new_new_n10339__ & ~new_new_n10342__;
  assign new_new_n10344__ = ~new_new_n10339__ & new_new_n10342__;
  assign new_new_n10345__ = ~new_new_n10343__ & ~new_new_n10344__;
  assign new_new_n10346__ = pi098 & ~new_new_n10345__;
  assign new_new_n10347__ = ~pi098 & new_new_n10345__;
  assign new_new_n10348__ = ~new_new_n9894__ & ~new_new_n9895__;
  assign new_new_n10349__ = pi096 & ~po022;
  assign new_new_n10350__ = ~new_new_n10252__ & po022;
  assign new_new_n10351__ = ~new_new_n10349__ & ~new_new_n10350__;
  assign new_new_n10352__ = new_new_n10348__ & ~new_new_n10351__;
  assign new_new_n10353__ = ~new_new_n10348__ & new_new_n10351__;
  assign new_new_n10354__ = ~new_new_n10352__ & ~new_new_n10353__;
  assign new_new_n10355__ = pi097 & new_new_n10354__;
  assign new_new_n10356__ = ~pi097 & ~new_new_n10354__;
  assign new_new_n10357__ = ~new_new_n10250__ & po022;
  assign new_new_n10358__ = pi095 & ~po022;
  assign new_new_n10359__ = ~new_new_n10357__ & ~new_new_n10358__;
  assign new_new_n10360__ = ~new_new_n9903__ & ~new_new_n9904__;
  assign new_new_n10361__ = ~new_new_n10359__ & new_new_n10360__;
  assign new_new_n10362__ = new_new_n10359__ & ~new_new_n10360__;
  assign new_new_n10363__ = ~new_new_n10361__ & ~new_new_n10362__;
  assign new_new_n10364__ = pi096 & new_new_n10363__;
  assign new_new_n10365__ = ~pi096 & ~new_new_n10363__;
  assign new_new_n10366__ = ~new_new_n9912__ & ~new_new_n9913__;
  assign new_new_n10367__ = ~new_new_n10248__ & po022;
  assign new_new_n10368__ = pi094 & ~po022;
  assign new_new_n10369__ = ~new_new_n10367__ & ~new_new_n10368__;
  assign new_new_n10370__ = new_new_n10366__ & new_new_n10369__;
  assign new_new_n10371__ = ~new_new_n10366__ & ~new_new_n10369__;
  assign new_new_n10372__ = ~new_new_n10370__ & ~new_new_n10371__;
  assign new_new_n10373__ = pi095 & ~new_new_n10372__;
  assign new_new_n10374__ = ~pi095 & new_new_n10372__;
  assign new_new_n10375__ = pi093 & ~new_new_n10246__;
  assign new_new_n10376__ = ~pi093 & new_new_n10246__;
  assign new_new_n10377__ = ~new_new_n10375__ & ~new_new_n10376__;
  assign new_new_n10378__ = po022 & new_new_n10377__;
  assign new_new_n10379__ = ~new_new_n9920__ & ~new_new_n10378__;
  assign new_new_n10380__ = new_new_n9920__ & new_new_n10378__;
  assign new_new_n10381__ = ~new_new_n10379__ & ~new_new_n10380__;
  assign new_new_n10382__ = pi094 & ~new_new_n10381__;
  assign new_new_n10383__ = ~pi094 & new_new_n10381__;
  assign new_new_n10384__ = ~new_new_n9930__ & ~new_new_n9931__;
  assign new_new_n10385__ = ~new_new_n10244__ & po022;
  assign new_new_n10386__ = ~pi092 & ~po022;
  assign new_new_n10387__ = ~new_new_n10385__ & ~new_new_n10386__;
  assign new_new_n10388__ = new_new_n10384__ & new_new_n10387__;
  assign new_new_n10389__ = ~new_new_n10384__ & ~new_new_n10387__;
  assign new_new_n10390__ = ~new_new_n10388__ & ~new_new_n10389__;
  assign new_new_n10391__ = ~pi093 & ~new_new_n10390__;
  assign new_new_n10392__ = pi093 & new_new_n10390__;
  assign new_new_n10393__ = new_new_n10242__ & po022;
  assign new_new_n10394__ = ~pi091 & ~po022;
  assign new_new_n10395__ = ~new_new_n10393__ & ~new_new_n10394__;
  assign new_new_n10396__ = ~new_new_n9939__ & ~new_new_n9940__;
  assign new_new_n10397__ = ~new_new_n10395__ & ~new_new_n10396__;
  assign new_new_n10398__ = new_new_n10395__ & new_new_n10396__;
  assign new_new_n10399__ = ~new_new_n10397__ & ~new_new_n10398__;
  assign new_new_n10400__ = ~pi092 & ~new_new_n10399__;
  assign new_new_n10401__ = pi092 & new_new_n10399__;
  assign new_new_n10402__ = ~new_new_n9948__ & ~new_new_n9949__;
  assign new_new_n10403__ = ~new_new_n10240__ & po022;
  assign new_new_n10404__ = ~pi090 & ~po022;
  assign new_new_n10405__ = ~new_new_n10403__ & ~new_new_n10404__;
  assign new_new_n10406__ = new_new_n10402__ & ~new_new_n10405__;
  assign new_new_n10407__ = ~new_new_n10402__ & new_new_n10405__;
  assign new_new_n10408__ = ~new_new_n10406__ & ~new_new_n10407__;
  assign new_new_n10409__ = pi091 & ~new_new_n10408__;
  assign new_new_n10410__ = ~pi091 & new_new_n10408__;
  assign new_new_n10411__ = ~pi089 & ~new_new_n10238__;
  assign new_new_n10412__ = pi089 & new_new_n10238__;
  assign new_new_n10413__ = ~new_new_n10411__ & ~new_new_n10412__;
  assign new_new_n10414__ = po022 & new_new_n10413__;
  assign new_new_n10415__ = ~new_new_n9956__ & new_new_n10414__;
  assign new_new_n10416__ = new_new_n9956__ & ~new_new_n10414__;
  assign new_new_n10417__ = ~new_new_n10415__ & ~new_new_n10416__;
  assign new_new_n10418__ = pi090 & ~new_new_n10417__;
  assign new_new_n10419__ = ~pi090 & new_new_n10417__;
  assign new_new_n10420__ = ~pi088 & ~new_new_n10236__;
  assign new_new_n10421__ = pi088 & new_new_n10236__;
  assign new_new_n10422__ = ~new_new_n10420__ & ~new_new_n10421__;
  assign new_new_n10423__ = po022 & new_new_n10422__;
  assign new_new_n10424__ = new_new_n9965__ & new_new_n10423__;
  assign new_new_n10425__ = ~new_new_n9965__ & ~new_new_n10423__;
  assign new_new_n10426__ = ~new_new_n10424__ & ~new_new_n10425__;
  assign new_new_n10427__ = pi089 & new_new_n10426__;
  assign new_new_n10428__ = ~pi089 & ~new_new_n10426__;
  assign new_new_n10429__ = ~pi087 & ~new_new_n10234__;
  assign new_new_n10430__ = pi087 & new_new_n10234__;
  assign new_new_n10431__ = ~new_new_n10429__ & ~new_new_n10430__;
  assign new_new_n10432__ = po022 & new_new_n10431__;
  assign new_new_n10433__ = ~new_new_n9974__ & new_new_n10432__;
  assign new_new_n10434__ = new_new_n9974__ & ~new_new_n10432__;
  assign new_new_n10435__ = ~new_new_n10433__ & ~new_new_n10434__;
  assign new_new_n10436__ = pi088 & ~new_new_n10435__;
  assign new_new_n10437__ = ~pi088 & new_new_n10435__;
  assign new_new_n10438__ = ~new_new_n9984__ & ~new_new_n9985__;
  assign new_new_n10439__ = ~new_new_n10232__ & po022;
  assign new_new_n10440__ = ~pi086 & ~po022;
  assign new_new_n10441__ = ~new_new_n10439__ & ~new_new_n10440__;
  assign new_new_n10442__ = new_new_n10438__ & ~new_new_n10441__;
  assign new_new_n10443__ = ~new_new_n10438__ & new_new_n10441__;
  assign new_new_n10444__ = ~new_new_n10442__ & ~new_new_n10443__;
  assign new_new_n10445__ = pi087 & ~new_new_n10444__;
  assign new_new_n10446__ = ~pi087 & new_new_n10444__;
  assign new_new_n10447__ = ~pi085 & ~new_new_n10230__;
  assign new_new_n10448__ = pi085 & new_new_n10230__;
  assign new_new_n10449__ = ~new_new_n10447__ & ~new_new_n10448__;
  assign new_new_n10450__ = po022 & new_new_n10449__;
  assign new_new_n10451__ = new_new_n9992__ & new_new_n10450__;
  assign new_new_n10452__ = ~new_new_n9992__ & ~new_new_n10450__;
  assign new_new_n10453__ = ~new_new_n10451__ & ~new_new_n10452__;
  assign new_new_n10454__ = ~pi086 & ~new_new_n10453__;
  assign new_new_n10455__ = pi086 & new_new_n10453__;
  assign new_new_n10456__ = ~new_new_n10002__ & ~new_new_n10003__;
  assign new_new_n10457__ = ~new_new_n10228__ & po022;
  assign new_new_n10458__ = ~pi084 & ~po022;
  assign new_new_n10459__ = ~new_new_n10457__ & ~new_new_n10458__;
  assign new_new_n10460__ = new_new_n10456__ & ~new_new_n10459__;
  assign new_new_n10461__ = ~new_new_n10456__ & new_new_n10459__;
  assign new_new_n10462__ = ~new_new_n10460__ & ~new_new_n10461__;
  assign new_new_n10463__ = ~pi085 & new_new_n10462__;
  assign new_new_n10464__ = pi085 & ~new_new_n10462__;
  assign new_new_n10465__ = ~pi083 & ~new_new_n10226__;
  assign new_new_n10466__ = pi083 & new_new_n10226__;
  assign new_new_n10467__ = ~new_new_n10465__ & ~new_new_n10466__;
  assign new_new_n10468__ = po022 & new_new_n10467__;
  assign new_new_n10469__ = new_new_n10010__ & new_new_n10468__;
  assign new_new_n10470__ = ~new_new_n10010__ & ~new_new_n10468__;
  assign new_new_n10471__ = ~new_new_n10469__ & ~new_new_n10470__;
  assign new_new_n10472__ = ~pi084 & ~new_new_n10471__;
  assign new_new_n10473__ = pi084 & new_new_n10471__;
  assign new_new_n10474__ = ~pi082 & ~new_new_n10224__;
  assign new_new_n10475__ = pi082 & new_new_n10224__;
  assign new_new_n10476__ = ~new_new_n10474__ & ~new_new_n10475__;
  assign new_new_n10477__ = po022 & new_new_n10476__;
  assign new_new_n10478__ = new_new_n10019__ & new_new_n10477__;
  assign new_new_n10479__ = ~new_new_n10019__ & ~new_new_n10477__;
  assign new_new_n10480__ = ~new_new_n10478__ & ~new_new_n10479__;
  assign new_new_n10481__ = ~pi083 & ~new_new_n10480__;
  assign new_new_n10482__ = pi083 & new_new_n10480__;
  assign new_new_n10483__ = ~new_new_n10029__ & ~new_new_n10030__;
  assign new_new_n10484__ = ~new_new_n10222__ & po022;
  assign new_new_n10485__ = ~pi081 & ~po022;
  assign new_new_n10486__ = ~new_new_n10484__ & ~new_new_n10485__;
  assign new_new_n10487__ = new_new_n10483__ & ~new_new_n10486__;
  assign new_new_n10488__ = ~new_new_n10483__ & new_new_n10486__;
  assign new_new_n10489__ = ~new_new_n10487__ & ~new_new_n10488__;
  assign new_new_n10490__ = ~pi082 & new_new_n10489__;
  assign new_new_n10491__ = pi082 & ~new_new_n10489__;
  assign new_new_n10492__ = ~pi080 & ~new_new_n10220__;
  assign new_new_n10493__ = pi080 & new_new_n10220__;
  assign new_new_n10494__ = ~new_new_n10492__ & ~new_new_n10493__;
  assign new_new_n10495__ = po022 & new_new_n10494__;
  assign new_new_n10496__ = new_new_n10037__ & new_new_n10495__;
  assign new_new_n10497__ = ~new_new_n10037__ & ~new_new_n10495__;
  assign new_new_n10498__ = ~new_new_n10496__ & ~new_new_n10497__;
  assign new_new_n10499__ = ~pi081 & ~new_new_n10498__;
  assign new_new_n10500__ = pi081 & new_new_n10498__;
  assign new_new_n10501__ = ~new_new_n10218__ & po022;
  assign new_new_n10502__ = pi079 & ~po022;
  assign new_new_n10503__ = ~new_new_n10501__ & ~new_new_n10502__;
  assign new_new_n10504__ = ~new_new_n10047__ & ~new_new_n10048__;
  assign new_new_n10505__ = ~new_new_n10503__ & new_new_n10504__;
  assign new_new_n10506__ = new_new_n10503__ & ~new_new_n10504__;
  assign new_new_n10507__ = ~new_new_n10505__ & ~new_new_n10506__;
  assign new_new_n10508__ = ~pi080 & ~new_new_n10507__;
  assign new_new_n10509__ = pi080 & new_new_n10507__;
  assign new_new_n10510__ = pi078 & ~new_new_n10216__;
  assign new_new_n10511__ = ~pi078 & new_new_n10216__;
  assign new_new_n10512__ = ~new_new_n10510__ & ~new_new_n10511__;
  assign new_new_n10513__ = po022 & new_new_n10512__;
  assign new_new_n10514__ = new_new_n10055__ & new_new_n10513__;
  assign new_new_n10515__ = ~new_new_n10055__ & ~new_new_n10513__;
  assign new_new_n10516__ = ~new_new_n10514__ & ~new_new_n10515__;
  assign new_new_n10517__ = ~pi079 & new_new_n10516__;
  assign new_new_n10518__ = pi079 & ~new_new_n10516__;
  assign new_new_n10519__ = ~new_new_n10065__ & ~new_new_n10066__;
  assign new_new_n10520__ = pi077 & ~po022;
  assign new_new_n10521__ = ~new_new_n10214__ & po022;
  assign new_new_n10522__ = ~new_new_n10520__ & ~new_new_n10521__;
  assign new_new_n10523__ = new_new_n10519__ & ~new_new_n10522__;
  assign new_new_n10524__ = ~new_new_n10519__ & new_new_n10522__;
  assign new_new_n10525__ = ~new_new_n10523__ & ~new_new_n10524__;
  assign new_new_n10526__ = ~pi078 & ~new_new_n10525__;
  assign new_new_n10527__ = pi078 & new_new_n10525__;
  assign new_new_n10528__ = ~new_new_n10074__ & ~new_new_n10075__;
  assign new_new_n10529__ = ~new_new_n10212__ & po022;
  assign new_new_n10530__ = ~pi076 & ~po022;
  assign new_new_n10531__ = ~new_new_n10529__ & ~new_new_n10530__;
  assign new_new_n10532__ = new_new_n10528__ & ~new_new_n10531__;
  assign new_new_n10533__ = ~new_new_n10528__ & new_new_n10531__;
  assign new_new_n10534__ = ~new_new_n10532__ & ~new_new_n10533__;
  assign new_new_n10535__ = ~pi077 & new_new_n10534__;
  assign new_new_n10536__ = pi077 & ~new_new_n10534__;
  assign new_new_n10537__ = ~pi075 & ~new_new_n10210__;
  assign new_new_n10538__ = pi075 & new_new_n10210__;
  assign new_new_n10539__ = ~new_new_n10537__ & ~new_new_n10538__;
  assign new_new_n10540__ = po022 & new_new_n10539__;
  assign new_new_n10541__ = new_new_n10082__ & new_new_n10540__;
  assign new_new_n10542__ = ~new_new_n10082__ & ~new_new_n10540__;
  assign new_new_n10543__ = ~new_new_n10541__ & ~new_new_n10542__;
  assign new_new_n10544__ = ~pi076 & ~new_new_n10543__;
  assign new_new_n10545__ = pi076 & new_new_n10543__;
  assign new_new_n10546__ = ~new_new_n10092__ & ~new_new_n10093__;
  assign new_new_n10547__ = ~new_new_n10208__ & po022;
  assign new_new_n10548__ = ~pi074 & ~po022;
  assign new_new_n10549__ = ~new_new_n10547__ & ~new_new_n10548__;
  assign new_new_n10550__ = new_new_n10546__ & ~new_new_n10549__;
  assign new_new_n10551__ = ~new_new_n10546__ & new_new_n10549__;
  assign new_new_n10552__ = ~new_new_n10550__ & ~new_new_n10551__;
  assign new_new_n10553__ = ~pi075 & new_new_n10552__;
  assign new_new_n10554__ = pi075 & ~new_new_n10552__;
  assign new_new_n10555__ = ~new_new_n10206__ & po022;
  assign new_new_n10556__ = pi073 & ~po022;
  assign new_new_n10557__ = ~new_new_n10555__ & ~new_new_n10556__;
  assign new_new_n10558__ = ~new_new_n10101__ & ~new_new_n10102__;
  assign new_new_n10559__ = ~new_new_n10557__ & new_new_n10558__;
  assign new_new_n10560__ = new_new_n10557__ & ~new_new_n10558__;
  assign new_new_n10561__ = ~new_new_n10559__ & ~new_new_n10560__;
  assign new_new_n10562__ = ~pi074 & ~new_new_n10561__;
  assign new_new_n10563__ = pi074 & new_new_n10561__;
  assign new_new_n10564__ = ~new_new_n10204__ & po022;
  assign new_new_n10565__ = pi072 & ~po022;
  assign new_new_n10566__ = ~new_new_n10564__ & ~new_new_n10565__;
  assign new_new_n10567__ = ~new_new_n10110__ & ~new_new_n10111__;
  assign new_new_n10568__ = ~new_new_n10566__ & new_new_n10567__;
  assign new_new_n10569__ = new_new_n10566__ & ~new_new_n10567__;
  assign new_new_n10570__ = ~new_new_n10568__ & ~new_new_n10569__;
  assign new_new_n10571__ = ~pi073 & ~new_new_n10570__;
  assign new_new_n10572__ = pi073 & new_new_n10570__;
  assign new_new_n10573__ = ~new_new_n10119__ & ~new_new_n10120__;
  assign new_new_n10574__ = ~new_new_n10202__ & po022;
  assign new_new_n10575__ = pi071 & ~po022;
  assign new_new_n10576__ = ~new_new_n10574__ & ~new_new_n10575__;
  assign new_new_n10577__ = new_new_n10573__ & ~new_new_n10576__;
  assign new_new_n10578__ = ~new_new_n10573__ & new_new_n10576__;
  assign new_new_n10579__ = ~new_new_n10577__ & ~new_new_n10578__;
  assign new_new_n10580__ = pi072 & new_new_n10579__;
  assign new_new_n10581__ = ~pi072 & ~new_new_n10579__;
  assign new_new_n10582__ = pi070 & ~new_new_n10200__;
  assign new_new_n10583__ = ~pi070 & new_new_n10200__;
  assign new_new_n10584__ = ~new_new_n10582__ & ~new_new_n10583__;
  assign new_new_n10585__ = po022 & new_new_n10584__;
  assign new_new_n10586__ = ~new_new_n10127__ & ~new_new_n10585__;
  assign new_new_n10587__ = new_new_n10127__ & new_new_n10585__;
  assign new_new_n10588__ = ~new_new_n10586__ & ~new_new_n10587__;
  assign new_new_n10589__ = pi071 & ~new_new_n10588__;
  assign new_new_n10590__ = ~pi071 & new_new_n10588__;
  assign new_new_n10591__ = ~new_new_n10137__ & ~new_new_n10138__;
  assign new_new_n10592__ = pi069 & ~po022;
  assign new_new_n10593__ = ~new_new_n10198__ & po022;
  assign new_new_n10594__ = ~new_new_n10592__ & ~new_new_n10593__;
  assign new_new_n10595__ = new_new_n10591__ & ~new_new_n10594__;
  assign new_new_n10596__ = ~new_new_n10591__ & new_new_n10594__;
  assign new_new_n10597__ = ~new_new_n10595__ & ~new_new_n10596__;
  assign new_new_n10598__ = pi070 & new_new_n10597__;
  assign new_new_n10599__ = ~pi070 & ~new_new_n10597__;
  assign new_new_n10600__ = ~new_new_n10188__ & ~new_new_n10189__;
  assign new_new_n10601__ = po022 & new_new_n10600__;
  assign new_new_n10602__ = ~new_new_n10196__ & ~new_new_n10601__;
  assign new_new_n10603__ = new_new_n10196__ & new_new_n10601__;
  assign new_new_n10604__ = ~new_new_n10602__ & ~new_new_n10603__;
  assign new_new_n10605__ = pi069 & new_new_n10604__;
  assign new_new_n10606__ = ~pi069 & ~new_new_n10604__;
  assign new_new_n10607__ = ~new_new_n10144__ & ~new_new_n10145__;
  assign new_new_n10608__ = ~new_new_n10185__ & po022;
  assign new_new_n10609__ = ~pi067 & ~po022;
  assign new_new_n10610__ = ~new_new_n10608__ & ~new_new_n10609__;
  assign new_new_n10611__ = new_new_n10607__ & ~new_new_n10610__;
  assign new_new_n10612__ = ~new_new_n10607__ & new_new_n10610__;
  assign new_new_n10613__ = ~new_new_n10611__ & ~new_new_n10612__;
  assign new_new_n10614__ = pi068 & ~new_new_n10613__;
  assign new_new_n10615__ = ~pi068 & new_new_n10613__;
  assign new_new_n10616__ = ~pi021 & pi065;
  assign new_new_n10617__ = pi065 & new_new_n10151__;
  assign new_new_n10618__ = ~pi065 & ~new_new_n10151__;
  assign new_new_n10619__ = ~new_new_n10617__ & ~new_new_n10618__;
  assign new_new_n10620__ = new_new_n10146__ & ~new_new_n10616__;
  assign new_new_n10621__ = ~new_new_n10619__ & new_new_n10620__;
  assign new_new_n10622__ = pi022 & new_new_n403__;
  assign new_new_n10623__ = ~new_new_n10151__ & new_new_n10622__;
  assign new_new_n10624__ = ~new_new_n10621__ & ~new_new_n10623__;
  assign new_new_n10625__ = po022 & ~new_new_n10624__;
  assign new_new_n10626__ = pi022 & ~po022;
  assign new_new_n10627__ = ~new_new_n332__ & ~new_new_n10626__;
  assign new_new_n10628__ = ~new_new_n426__ & ~new_new_n10627__;
  assign new_new_n10629__ = pi065 & po022;
  assign new_new_n10630__ = ~pi065 & ~po022;
  assign new_new_n10631__ = ~pi022 & ~new_new_n10630__;
  assign new_new_n10632__ = pi021 & ~new_new_n10629__;
  assign new_new_n10633__ = ~new_new_n10631__ & new_new_n10632__;
  assign new_new_n10634__ = ~new_new_n10628__ & ~new_new_n10633__;
  assign new_new_n10635__ = new_new_n10151__ & ~new_new_n10634__;
  assign new_new_n10636__ = ~pi023 & ~po023;
  assign new_new_n10637__ = new_new_n10176__ & ~new_new_n10636__;
  assign new_new_n10638__ = pi023 & ~pi064;
  assign new_new_n10639__ = po022 & ~new_new_n10638__;
  assign new_new_n10640__ = ~po022 & new_new_n10638__;
  assign new_new_n10641__ = ~pi022 & pi065;
  assign new_new_n10642__ = ~new_new_n10637__ & new_new_n10641__;
  assign new_new_n10643__ = ~new_new_n10639__ & new_new_n10642__;
  assign new_new_n10644__ = ~new_new_n10640__ & new_new_n10643__;
  assign new_new_n10645__ = pi021 & ~pi065;
  assign new_new_n10646__ = pi022 & po022;
  assign new_new_n10647__ = ~new_new_n10619__ & ~new_new_n10645__;
  assign new_new_n10648__ = new_new_n10646__ & new_new_n10647__;
  assign new_new_n10649__ = ~pi065 & po022;
  assign new_new_n10650__ = pi065 & ~po022;
  assign new_new_n10651__ = pi022 & ~new_new_n10650__;
  assign new_new_n10652__ = ~pi021 & ~new_new_n10151__;
  assign new_new_n10653__ = ~new_new_n10649__ & new_new_n10652__;
  assign new_new_n10654__ = ~new_new_n10651__ & new_new_n10653__;
  assign new_new_n10655__ = ~new_new_n10648__ & ~new_new_n10654__;
  assign new_new_n10656__ = pi064 & ~new_new_n10655__;
  assign new_new_n10657__ = ~pi066 & ~new_new_n10644__;
  assign new_new_n10658__ = ~new_new_n10656__ & new_new_n10657__;
  assign new_new_n10659__ = ~new_new_n10625__ & ~new_new_n10635__;
  assign new_new_n10660__ = ~new_new_n10658__ & new_new_n10659__;
  assign new_new_n10661__ = pi067 & new_new_n10660__;
  assign new_new_n10662__ = ~pi067 & ~new_new_n10660__;
  assign new_new_n10663__ = ~new_new_n10156__ & ~new_new_n10157__;
  assign new_new_n10664__ = po022 & new_new_n10663__;
  assign new_new_n10665__ = new_new_n10183__ & ~new_new_n10664__;
  assign new_new_n10666__ = ~new_new_n10183__ & new_new_n10664__;
  assign new_new_n10667__ = ~new_new_n10665__ & ~new_new_n10666__;
  assign new_new_n10668__ = ~new_new_n10662__ & new_new_n10667__;
  assign new_new_n10669__ = ~new_new_n10661__ & ~new_new_n10668__;
  assign new_new_n10670__ = ~new_new_n10615__ & ~new_new_n10669__;
  assign new_new_n10671__ = ~new_new_n10614__ & ~new_new_n10670__;
  assign new_new_n10672__ = ~new_new_n10606__ & ~new_new_n10671__;
  assign new_new_n10673__ = ~new_new_n10605__ & ~new_new_n10672__;
  assign new_new_n10674__ = ~new_new_n10599__ & ~new_new_n10673__;
  assign new_new_n10675__ = ~new_new_n10598__ & ~new_new_n10674__;
  assign new_new_n10676__ = ~new_new_n10590__ & ~new_new_n10675__;
  assign new_new_n10677__ = ~new_new_n10589__ & ~new_new_n10676__;
  assign new_new_n10678__ = ~new_new_n10581__ & ~new_new_n10677__;
  assign new_new_n10679__ = ~new_new_n10580__ & ~new_new_n10678__;
  assign new_new_n10680__ = ~new_new_n10572__ & new_new_n10679__;
  assign new_new_n10681__ = ~new_new_n10571__ & ~new_new_n10680__;
  assign new_new_n10682__ = ~new_new_n10563__ & ~new_new_n10681__;
  assign new_new_n10683__ = ~new_new_n10562__ & ~new_new_n10682__;
  assign new_new_n10684__ = ~new_new_n10554__ & ~new_new_n10683__;
  assign new_new_n10685__ = ~new_new_n10553__ & ~new_new_n10684__;
  assign new_new_n10686__ = ~new_new_n10545__ & ~new_new_n10685__;
  assign new_new_n10687__ = ~new_new_n10544__ & ~new_new_n10686__;
  assign new_new_n10688__ = ~new_new_n10536__ & ~new_new_n10687__;
  assign new_new_n10689__ = ~new_new_n10535__ & ~new_new_n10688__;
  assign new_new_n10690__ = ~new_new_n10527__ & ~new_new_n10689__;
  assign new_new_n10691__ = ~new_new_n10526__ & ~new_new_n10690__;
  assign new_new_n10692__ = ~new_new_n10518__ & ~new_new_n10691__;
  assign new_new_n10693__ = ~new_new_n10517__ & ~new_new_n10692__;
  assign new_new_n10694__ = ~new_new_n10509__ & ~new_new_n10693__;
  assign new_new_n10695__ = ~new_new_n10508__ & ~new_new_n10694__;
  assign new_new_n10696__ = ~new_new_n10500__ & ~new_new_n10695__;
  assign new_new_n10697__ = ~new_new_n10499__ & ~new_new_n10696__;
  assign new_new_n10698__ = ~new_new_n10491__ & ~new_new_n10697__;
  assign new_new_n10699__ = ~new_new_n10490__ & ~new_new_n10698__;
  assign new_new_n10700__ = ~new_new_n10482__ & ~new_new_n10699__;
  assign new_new_n10701__ = ~new_new_n10481__ & ~new_new_n10700__;
  assign new_new_n10702__ = ~new_new_n10473__ & ~new_new_n10701__;
  assign new_new_n10703__ = ~new_new_n10472__ & ~new_new_n10702__;
  assign new_new_n10704__ = ~new_new_n10464__ & ~new_new_n10703__;
  assign new_new_n10705__ = ~new_new_n10463__ & ~new_new_n10704__;
  assign new_new_n10706__ = ~new_new_n10455__ & ~new_new_n10705__;
  assign new_new_n10707__ = ~new_new_n10454__ & ~new_new_n10706__;
  assign new_new_n10708__ = ~new_new_n10446__ & new_new_n10707__;
  assign new_new_n10709__ = ~new_new_n10445__ & ~new_new_n10708__;
  assign new_new_n10710__ = ~new_new_n10437__ & ~new_new_n10709__;
  assign new_new_n10711__ = ~new_new_n10436__ & ~new_new_n10710__;
  assign new_new_n10712__ = ~new_new_n10428__ & ~new_new_n10711__;
  assign new_new_n10713__ = ~new_new_n10427__ & ~new_new_n10712__;
  assign new_new_n10714__ = ~new_new_n10419__ & ~new_new_n10713__;
  assign new_new_n10715__ = ~new_new_n10418__ & ~new_new_n10714__;
  assign new_new_n10716__ = ~new_new_n10410__ & ~new_new_n10715__;
  assign new_new_n10717__ = ~new_new_n10409__ & ~new_new_n10716__;
  assign new_new_n10718__ = ~new_new_n10401__ & new_new_n10717__;
  assign new_new_n10719__ = ~new_new_n10400__ & ~new_new_n10718__;
  assign new_new_n10720__ = ~new_new_n10392__ & ~new_new_n10719__;
  assign new_new_n10721__ = ~new_new_n10391__ & ~new_new_n10720__;
  assign new_new_n10722__ = ~new_new_n10383__ & new_new_n10721__;
  assign new_new_n10723__ = ~new_new_n10382__ & ~new_new_n10722__;
  assign new_new_n10724__ = ~new_new_n10374__ & ~new_new_n10723__;
  assign new_new_n10725__ = ~new_new_n10373__ & ~new_new_n10724__;
  assign new_new_n10726__ = ~new_new_n10365__ & ~new_new_n10725__;
  assign new_new_n10727__ = ~new_new_n10364__ & ~new_new_n10726__;
  assign new_new_n10728__ = ~new_new_n10356__ & ~new_new_n10727__;
  assign new_new_n10729__ = ~new_new_n10355__ & ~new_new_n10728__;
  assign new_new_n10730__ = ~new_new_n10347__ & ~new_new_n10729__;
  assign new_new_n10731__ = ~new_new_n10346__ & ~new_new_n10730__;
  assign new_new_n10732__ = ~new_new_n10338__ & ~new_new_n10731__;
  assign new_new_n10733__ = ~new_new_n10337__ & ~new_new_n10732__;
  assign new_new_n10734__ = ~new_new_n10329__ & ~new_new_n10733__;
  assign new_new_n10735__ = ~new_new_n10328__ & ~new_new_n10734__;
  assign new_new_n10736__ = ~new_new_n10320__ & ~new_new_n10735__;
  assign new_new_n10737__ = ~new_new_n10319__ & ~new_new_n10736__;
  assign new_new_n10738__ = ~new_new_n10311__ & ~new_new_n10737__;
  assign new_new_n10739__ = ~new_new_n10310__ & ~new_new_n10738__;
  assign new_new_n10740__ = ~new_new_n10302__ & ~new_new_n10739__;
  assign new_new_n10741__ = ~new_new_n10301__ & ~new_new_n10740__;
  assign new_new_n10742__ = ~new_new_n10293__ & new_new_n10741__;
  assign new_new_n10743__ = ~new_new_n10292__ & ~new_new_n10742__;
  assign new_new_n10744__ = ~new_new_n10284__ & new_new_n10743__;
  assign new_new_n10745__ = ~new_new_n10283__ & ~new_new_n10744__;
  assign new_new_n10746__ = pi106 & ~new_new_n10745__;
  assign new_new_n10747__ = ~new_new_n10271__ & ~new_new_n10273__;
  assign new_new_n10748__ = ~pi106 & ~new_new_n10747__;
  assign new_new_n10749__ = new_new_n10745__ & new_new_n10748__;
  assign new_new_n10750__ = new_new_n279__ & ~new_new_n10746__;
  assign new_new_n10751__ = ~new_new_n10749__ & new_new_n10750__;
  assign new_new_n10752__ = new_new_n9808__ & ~new_new_n10751__;
  assign new_new_n10753__ = ~pi109 & new_new_n8066__;
  assign new_new_n10754__ = pi106 & ~new_new_n9808__;
  assign new_new_n10755__ = new_new_n10745__ & ~new_new_n10754__;
  assign new_new_n10756__ = ~pi106 & new_new_n9808__;
  assign new_new_n10757__ = ~new_new_n10747__ & new_new_n10756__;
  assign new_new_n10758__ = ~new_new_n10755__ & ~new_new_n10757__;
  assign po021 = new_new_n279__ & ~new_new_n10758__;
  assign new_new_n10760__ = ~new_new_n10741__ & po021;
  assign new_new_n10761__ = pi104 & ~po021;
  assign new_new_n10762__ = ~new_new_n10760__ & ~new_new_n10761__;
  assign new_new_n10763__ = ~new_new_n10292__ & ~new_new_n10293__;
  assign new_new_n10764__ = ~new_new_n10762__ & new_new_n10763__;
  assign new_new_n10765__ = new_new_n10762__ & ~new_new_n10763__;
  assign new_new_n10766__ = ~new_new_n10764__ & ~new_new_n10765__;
  assign new_new_n10767__ = pi105 & new_new_n10766__;
  assign new_new_n10768__ = ~pi105 & ~new_new_n10766__;
  assign new_new_n10769__ = ~new_new_n10767__ & ~new_new_n10768__;
  assign new_new_n10770__ = ~new_new_n10739__ & po021;
  assign new_new_n10771__ = pi103 & ~po021;
  assign new_new_n10772__ = ~new_new_n10770__ & ~new_new_n10771__;
  assign new_new_n10773__ = ~new_new_n10301__ & ~new_new_n10302__;
  assign new_new_n10774__ = ~new_new_n10772__ & new_new_n10773__;
  assign new_new_n10775__ = new_new_n10772__ & ~new_new_n10773__;
  assign new_new_n10776__ = ~new_new_n10774__ & ~new_new_n10775__;
  assign new_new_n10777__ = ~pi104 & ~new_new_n10776__;
  assign new_new_n10778__ = pi104 & new_new_n10776__;
  assign new_new_n10779__ = ~new_new_n10310__ & ~new_new_n10311__;
  assign new_new_n10780__ = new_new_n10737__ & po021;
  assign new_new_n10781__ = ~pi102 & ~po021;
  assign new_new_n10782__ = ~new_new_n10780__ & ~new_new_n10781__;
  assign new_new_n10783__ = ~new_new_n10779__ & ~new_new_n10782__;
  assign new_new_n10784__ = new_new_n10779__ & new_new_n10782__;
  assign new_new_n10785__ = ~new_new_n10783__ & ~new_new_n10784__;
  assign new_new_n10786__ = ~pi103 & ~new_new_n10785__;
  assign new_new_n10787__ = pi103 & new_new_n10785__;
  assign new_new_n10788__ = ~new_new_n10733__ & po021;
  assign new_new_n10789__ = pi100 & ~po021;
  assign new_new_n10790__ = ~new_new_n10788__ & ~new_new_n10789__;
  assign new_new_n10791__ = ~new_new_n10328__ & ~new_new_n10329__;
  assign new_new_n10792__ = new_new_n10790__ & new_new_n10791__;
  assign new_new_n10793__ = ~new_new_n10790__ & ~new_new_n10791__;
  assign new_new_n10794__ = ~new_new_n10792__ & ~new_new_n10793__;
  assign new_new_n10795__ = pi101 & ~new_new_n10794__;
  assign new_new_n10796__ = ~pi101 & new_new_n10794__;
  assign new_new_n10797__ = ~new_new_n10337__ & ~new_new_n10338__;
  assign new_new_n10798__ = pi099 & ~po021;
  assign new_new_n10799__ = ~new_new_n10731__ & po021;
  assign new_new_n10800__ = ~new_new_n10798__ & ~new_new_n10799__;
  assign new_new_n10801__ = new_new_n10797__ & new_new_n10800__;
  assign new_new_n10802__ = ~new_new_n10797__ & ~new_new_n10800__;
  assign new_new_n10803__ = ~new_new_n10801__ & ~new_new_n10802__;
  assign new_new_n10804__ = pi100 & ~new_new_n10803__;
  assign new_new_n10805__ = ~pi100 & new_new_n10803__;
  assign new_new_n10806__ = ~new_new_n10346__ & ~new_new_n10347__;
  assign new_new_n10807__ = ~new_new_n10729__ & po021;
  assign new_new_n10808__ = pi098 & ~po021;
  assign new_new_n10809__ = ~new_new_n10807__ & ~new_new_n10808__;
  assign new_new_n10810__ = new_new_n10806__ & new_new_n10809__;
  assign new_new_n10811__ = ~new_new_n10806__ & ~new_new_n10809__;
  assign new_new_n10812__ = ~new_new_n10810__ & ~new_new_n10811__;
  assign new_new_n10813__ = ~pi099 & new_new_n10812__;
  assign new_new_n10814__ = pi099 & ~new_new_n10812__;
  assign new_new_n10815__ = new_new_n10727__ & po021;
  assign new_new_n10816__ = ~pi097 & ~po021;
  assign new_new_n10817__ = ~new_new_n10815__ & ~new_new_n10816__;
  assign new_new_n10818__ = ~new_new_n10355__ & ~new_new_n10356__;
  assign new_new_n10819__ = ~new_new_n10817__ & ~new_new_n10818__;
  assign new_new_n10820__ = new_new_n10817__ & new_new_n10818__;
  assign new_new_n10821__ = ~new_new_n10819__ & ~new_new_n10820__;
  assign new_new_n10822__ = ~pi098 & ~new_new_n10821__;
  assign new_new_n10823__ = pi098 & new_new_n10821__;
  assign new_new_n10824__ = new_new_n10725__ & po021;
  assign new_new_n10825__ = ~pi096 & ~po021;
  assign new_new_n10826__ = ~new_new_n10824__ & ~new_new_n10825__;
  assign new_new_n10827__ = ~new_new_n10364__ & ~new_new_n10365__;
  assign new_new_n10828__ = ~new_new_n10826__ & ~new_new_n10827__;
  assign new_new_n10829__ = new_new_n10826__ & new_new_n10827__;
  assign new_new_n10830__ = ~new_new_n10828__ & ~new_new_n10829__;
  assign new_new_n10831__ = ~pi097 & ~new_new_n10830__;
  assign new_new_n10832__ = pi097 & new_new_n10830__;
  assign new_new_n10833__ = pi095 & ~new_new_n10723__;
  assign new_new_n10834__ = ~pi095 & new_new_n10723__;
  assign new_new_n10835__ = ~new_new_n10833__ & ~new_new_n10834__;
  assign new_new_n10836__ = po021 & new_new_n10835__;
  assign new_new_n10837__ = new_new_n10372__ & new_new_n10836__;
  assign new_new_n10838__ = ~new_new_n10372__ & ~new_new_n10836__;
  assign new_new_n10839__ = ~new_new_n10837__ & ~new_new_n10838__;
  assign new_new_n10840__ = pi096 & ~new_new_n10839__;
  assign new_new_n10841__ = ~pi096 & new_new_n10839__;
  assign new_new_n10842__ = ~new_new_n10382__ & ~new_new_n10383__;
  assign new_new_n10843__ = ~new_new_n10721__ & po021;
  assign new_new_n10844__ = ~pi094 & ~po021;
  assign new_new_n10845__ = ~new_new_n10843__ & ~new_new_n10844__;
  assign new_new_n10846__ = new_new_n10842__ & new_new_n10845__;
  assign new_new_n10847__ = ~new_new_n10842__ & ~new_new_n10845__;
  assign new_new_n10848__ = ~new_new_n10846__ & ~new_new_n10847__;
  assign new_new_n10849__ = ~pi095 & ~new_new_n10848__;
  assign new_new_n10850__ = pi095 & new_new_n10848__;
  assign new_new_n10851__ = ~new_new_n10391__ & ~new_new_n10392__;
  assign new_new_n10852__ = ~new_new_n10719__ & po021;
  assign new_new_n10853__ = ~pi093 & ~po021;
  assign new_new_n10854__ = ~new_new_n10852__ & ~new_new_n10853__;
  assign new_new_n10855__ = ~new_new_n10851__ & ~new_new_n10854__;
  assign new_new_n10856__ = new_new_n10851__ & new_new_n10854__;
  assign new_new_n10857__ = ~new_new_n10855__ & ~new_new_n10856__;
  assign new_new_n10858__ = ~pi094 & ~new_new_n10857__;
  assign new_new_n10859__ = pi094 & new_new_n10857__;
  assign new_new_n10860__ = new_new_n10717__ & po021;
  assign new_new_n10861__ = ~pi092 & ~po021;
  assign new_new_n10862__ = ~new_new_n10860__ & ~new_new_n10861__;
  assign new_new_n10863__ = ~new_new_n10400__ & ~new_new_n10401__;
  assign new_new_n10864__ = ~new_new_n10862__ & ~new_new_n10863__;
  assign new_new_n10865__ = new_new_n10862__ & new_new_n10863__;
  assign new_new_n10866__ = ~new_new_n10864__ & ~new_new_n10865__;
  assign new_new_n10867__ = ~pi093 & ~new_new_n10866__;
  assign new_new_n10868__ = pi093 & new_new_n10866__;
  assign new_new_n10869__ = pi091 & ~new_new_n10715__;
  assign new_new_n10870__ = ~pi091 & new_new_n10715__;
  assign new_new_n10871__ = ~new_new_n10869__ & ~new_new_n10870__;
  assign new_new_n10872__ = po021 & new_new_n10871__;
  assign new_new_n10873__ = new_new_n10408__ & new_new_n10872__;
  assign new_new_n10874__ = ~new_new_n10408__ & ~new_new_n10872__;
  assign new_new_n10875__ = ~new_new_n10873__ & ~new_new_n10874__;
  assign new_new_n10876__ = pi092 & ~new_new_n10875__;
  assign new_new_n10877__ = ~pi092 & new_new_n10875__;
  assign new_new_n10878__ = ~new_new_n10418__ & ~new_new_n10419__;
  assign new_new_n10879__ = ~new_new_n10713__ & po021;
  assign new_new_n10880__ = pi090 & ~po021;
  assign new_new_n10881__ = ~new_new_n10879__ & ~new_new_n10880__;
  assign new_new_n10882__ = new_new_n10878__ & ~new_new_n10881__;
  assign new_new_n10883__ = ~new_new_n10878__ & new_new_n10881__;
  assign new_new_n10884__ = ~new_new_n10882__ & ~new_new_n10883__;
  assign new_new_n10885__ = ~pi091 & ~new_new_n10884__;
  assign new_new_n10886__ = pi091 & new_new_n10884__;
  assign new_new_n10887__ = ~new_new_n10711__ & po021;
  assign new_new_n10888__ = pi089 & ~po021;
  assign new_new_n10889__ = ~new_new_n10887__ & ~new_new_n10888__;
  assign new_new_n10890__ = ~new_new_n10427__ & ~new_new_n10428__;
  assign new_new_n10891__ = ~new_new_n10889__ & new_new_n10890__;
  assign new_new_n10892__ = new_new_n10889__ & ~new_new_n10890__;
  assign new_new_n10893__ = ~new_new_n10891__ & ~new_new_n10892__;
  assign new_new_n10894__ = ~pi090 & ~new_new_n10893__;
  assign new_new_n10895__ = pi090 & new_new_n10893__;
  assign new_new_n10896__ = ~new_new_n10436__ & ~new_new_n10437__;
  assign new_new_n10897__ = ~new_new_n10709__ & po021;
  assign new_new_n10898__ = pi088 & ~po021;
  assign new_new_n10899__ = ~new_new_n10897__ & ~new_new_n10898__;
  assign new_new_n10900__ = new_new_n10896__ & ~new_new_n10899__;
  assign new_new_n10901__ = ~new_new_n10896__ & new_new_n10899__;
  assign new_new_n10902__ = ~new_new_n10900__ & ~new_new_n10901__;
  assign new_new_n10903__ = ~pi089 & ~new_new_n10902__;
  assign new_new_n10904__ = pi089 & new_new_n10902__;
  assign new_new_n10905__ = ~new_new_n10445__ & ~new_new_n10446__;
  assign new_new_n10906__ = ~new_new_n10707__ & po021;
  assign new_new_n10907__ = ~pi087 & ~po021;
  assign new_new_n10908__ = ~new_new_n10906__ & ~new_new_n10907__;
  assign new_new_n10909__ = new_new_n10905__ & ~new_new_n10908__;
  assign new_new_n10910__ = ~new_new_n10905__ & new_new_n10908__;
  assign new_new_n10911__ = ~new_new_n10909__ & ~new_new_n10910__;
  assign new_new_n10912__ = ~pi088 & new_new_n10911__;
  assign new_new_n10913__ = pi088 & ~new_new_n10911__;
  assign new_new_n10914__ = ~pi086 & ~new_new_n10705__;
  assign new_new_n10915__ = pi086 & new_new_n10705__;
  assign new_new_n10916__ = ~new_new_n10914__ & ~new_new_n10915__;
  assign new_new_n10917__ = po021 & new_new_n10916__;
  assign new_new_n10918__ = ~new_new_n10453__ & ~new_new_n10917__;
  assign new_new_n10919__ = new_new_n10453__ & new_new_n10917__;
  assign new_new_n10920__ = ~new_new_n10918__ & ~new_new_n10919__;
  assign new_new_n10921__ = ~pi087 & ~new_new_n10920__;
  assign new_new_n10922__ = pi087 & new_new_n10920__;
  assign new_new_n10923__ = ~new_new_n10463__ & ~new_new_n10464__;
  assign new_new_n10924__ = ~new_new_n10703__ & po021;
  assign new_new_n10925__ = ~pi085 & ~po021;
  assign new_new_n10926__ = ~new_new_n10924__ & ~new_new_n10925__;
  assign new_new_n10927__ = new_new_n10923__ & ~new_new_n10926__;
  assign new_new_n10928__ = ~new_new_n10923__ & new_new_n10926__;
  assign new_new_n10929__ = ~new_new_n10927__ & ~new_new_n10928__;
  assign new_new_n10930__ = ~pi086 & new_new_n10929__;
  assign new_new_n10931__ = pi086 & ~new_new_n10929__;
  assign new_new_n10932__ = ~pi084 & ~new_new_n10701__;
  assign new_new_n10933__ = pi084 & new_new_n10701__;
  assign new_new_n10934__ = ~new_new_n10932__ & ~new_new_n10933__;
  assign new_new_n10935__ = po021 & new_new_n10934__;
  assign new_new_n10936__ = new_new_n10471__ & new_new_n10935__;
  assign new_new_n10937__ = ~new_new_n10471__ & ~new_new_n10935__;
  assign new_new_n10938__ = ~new_new_n10936__ & ~new_new_n10937__;
  assign new_new_n10939__ = ~pi085 & ~new_new_n10938__;
  assign new_new_n10940__ = pi085 & new_new_n10938__;
  assign new_new_n10941__ = ~pi083 & ~new_new_n10699__;
  assign new_new_n10942__ = pi083 & new_new_n10699__;
  assign new_new_n10943__ = ~new_new_n10941__ & ~new_new_n10942__;
  assign new_new_n10944__ = po021 & new_new_n10943__;
  assign new_new_n10945__ = new_new_n10480__ & new_new_n10944__;
  assign new_new_n10946__ = ~new_new_n10480__ & ~new_new_n10944__;
  assign new_new_n10947__ = ~new_new_n10945__ & ~new_new_n10946__;
  assign new_new_n10948__ = ~pi084 & ~new_new_n10947__;
  assign new_new_n10949__ = pi084 & new_new_n10947__;
  assign new_new_n10950__ = ~new_new_n10490__ & ~new_new_n10491__;
  assign new_new_n10951__ = ~new_new_n10697__ & po021;
  assign new_new_n10952__ = ~pi082 & ~po021;
  assign new_new_n10953__ = ~new_new_n10951__ & ~new_new_n10952__;
  assign new_new_n10954__ = new_new_n10950__ & ~new_new_n10953__;
  assign new_new_n10955__ = ~new_new_n10950__ & new_new_n10953__;
  assign new_new_n10956__ = ~new_new_n10954__ & ~new_new_n10955__;
  assign new_new_n10957__ = pi083 & ~new_new_n10956__;
  assign new_new_n10958__ = ~pi083 & new_new_n10956__;
  assign new_new_n10959__ = ~pi081 & ~new_new_n10695__;
  assign new_new_n10960__ = pi081 & new_new_n10695__;
  assign new_new_n10961__ = ~new_new_n10959__ & ~new_new_n10960__;
  assign new_new_n10962__ = po021 & new_new_n10961__;
  assign new_new_n10963__ = new_new_n10498__ & new_new_n10962__;
  assign new_new_n10964__ = ~new_new_n10498__ & ~new_new_n10962__;
  assign new_new_n10965__ = ~new_new_n10963__ & ~new_new_n10964__;
  assign new_new_n10966__ = ~pi082 & ~new_new_n10965__;
  assign new_new_n10967__ = pi082 & new_new_n10965__;
  assign new_new_n10968__ = ~pi080 & ~new_new_n10693__;
  assign new_new_n10969__ = pi080 & new_new_n10693__;
  assign new_new_n10970__ = ~new_new_n10968__ & ~new_new_n10969__;
  assign new_new_n10971__ = po021 & new_new_n10970__;
  assign new_new_n10972__ = new_new_n10507__ & new_new_n10971__;
  assign new_new_n10973__ = ~new_new_n10507__ & ~new_new_n10971__;
  assign new_new_n10974__ = ~new_new_n10972__ & ~new_new_n10973__;
  assign new_new_n10975__ = ~pi081 & ~new_new_n10974__;
  assign new_new_n10976__ = pi081 & new_new_n10974__;
  assign new_new_n10977__ = ~new_new_n10517__ & ~new_new_n10518__;
  assign new_new_n10978__ = ~new_new_n10691__ & po021;
  assign new_new_n10979__ = ~pi079 & ~po021;
  assign new_new_n10980__ = ~new_new_n10978__ & ~new_new_n10979__;
  assign new_new_n10981__ = new_new_n10977__ & ~new_new_n10980__;
  assign new_new_n10982__ = ~new_new_n10977__ & new_new_n10980__;
  assign new_new_n10983__ = ~new_new_n10981__ & ~new_new_n10982__;
  assign new_new_n10984__ = pi080 & ~new_new_n10983__;
  assign new_new_n10985__ = ~pi080 & new_new_n10983__;
  assign new_new_n10986__ = ~pi078 & ~new_new_n10689__;
  assign new_new_n10987__ = pi078 & new_new_n10689__;
  assign new_new_n10988__ = ~new_new_n10986__ & ~new_new_n10987__;
  assign new_new_n10989__ = po021 & new_new_n10988__;
  assign new_new_n10990__ = new_new_n10525__ & new_new_n10989__;
  assign new_new_n10991__ = ~new_new_n10525__ & ~new_new_n10989__;
  assign new_new_n10992__ = ~new_new_n10990__ & ~new_new_n10991__;
  assign new_new_n10993__ = pi079 & new_new_n10992__;
  assign new_new_n10994__ = ~pi079 & ~new_new_n10992__;
  assign new_new_n10995__ = ~new_new_n10535__ & ~new_new_n10536__;
  assign new_new_n10996__ = ~new_new_n10687__ & po021;
  assign new_new_n10997__ = ~pi077 & ~po021;
  assign new_new_n10998__ = ~new_new_n10996__ & ~new_new_n10997__;
  assign new_new_n10999__ = new_new_n10995__ & ~new_new_n10998__;
  assign new_new_n11000__ = ~new_new_n10995__ & new_new_n10998__;
  assign new_new_n11001__ = ~new_new_n10999__ & ~new_new_n11000__;
  assign new_new_n11002__ = pi078 & ~new_new_n11001__;
  assign new_new_n11003__ = ~pi078 & new_new_n11001__;
  assign new_new_n11004__ = ~new_new_n10544__ & ~new_new_n10545__;
  assign new_new_n11005__ = ~new_new_n10685__ & po021;
  assign new_new_n11006__ = ~pi076 & ~po021;
  assign new_new_n11007__ = ~new_new_n11005__ & ~new_new_n11006__;
  assign new_new_n11008__ = new_new_n11004__ & ~new_new_n11007__;
  assign new_new_n11009__ = ~new_new_n11004__ & new_new_n11007__;
  assign new_new_n11010__ = ~new_new_n11008__ & ~new_new_n11009__;
  assign new_new_n11011__ = ~pi077 & new_new_n11010__;
  assign new_new_n11012__ = pi077 & ~new_new_n11010__;
  assign new_new_n11013__ = ~new_new_n10553__ & ~new_new_n10554__;
  assign new_new_n11014__ = ~new_new_n10683__ & po021;
  assign new_new_n11015__ = ~pi075 & ~po021;
  assign new_new_n11016__ = ~new_new_n11014__ & ~new_new_n11015__;
  assign new_new_n11017__ = new_new_n11013__ & ~new_new_n11016__;
  assign new_new_n11018__ = ~new_new_n11013__ & new_new_n11016__;
  assign new_new_n11019__ = ~new_new_n11017__ & ~new_new_n11018__;
  assign new_new_n11020__ = ~pi076 & new_new_n11019__;
  assign new_new_n11021__ = pi076 & ~new_new_n11019__;
  assign new_new_n11022__ = ~pi074 & ~new_new_n10681__;
  assign new_new_n11023__ = pi074 & new_new_n10681__;
  assign new_new_n11024__ = ~new_new_n11022__ & ~new_new_n11023__;
  assign new_new_n11025__ = po021 & new_new_n11024__;
  assign new_new_n11026__ = new_new_n10561__ & new_new_n11025__;
  assign new_new_n11027__ = ~new_new_n10561__ & ~new_new_n11025__;
  assign new_new_n11028__ = ~new_new_n11026__ & ~new_new_n11027__;
  assign new_new_n11029__ = ~pi075 & ~new_new_n11028__;
  assign new_new_n11030__ = pi075 & new_new_n11028__;
  assign new_new_n11031__ = ~new_new_n10571__ & ~new_new_n10572__;
  assign new_new_n11032__ = new_new_n10679__ & po021;
  assign new_new_n11033__ = ~pi073 & ~po021;
  assign new_new_n11034__ = ~new_new_n11032__ & ~new_new_n11033__;
  assign new_new_n11035__ = ~new_new_n11031__ & ~new_new_n11034__;
  assign new_new_n11036__ = new_new_n11031__ & new_new_n11034__;
  assign new_new_n11037__ = ~new_new_n11035__ & ~new_new_n11036__;
  assign new_new_n11038__ = ~pi074 & ~new_new_n11037__;
  assign new_new_n11039__ = pi074 & new_new_n11037__;
  assign new_new_n11040__ = new_new_n10677__ & po021;
  assign new_new_n11041__ = ~pi072 & ~po021;
  assign new_new_n11042__ = ~new_new_n11040__ & ~new_new_n11041__;
  assign new_new_n11043__ = ~new_new_n10580__ & ~new_new_n10581__;
  assign new_new_n11044__ = ~new_new_n11042__ & ~new_new_n11043__;
  assign new_new_n11045__ = new_new_n11042__ & new_new_n11043__;
  assign new_new_n11046__ = ~new_new_n11044__ & ~new_new_n11045__;
  assign new_new_n11047__ = ~pi073 & ~new_new_n11046__;
  assign new_new_n11048__ = pi073 & new_new_n11046__;
  assign new_new_n11049__ = ~new_new_n10589__ & ~new_new_n10590__;
  assign new_new_n11050__ = ~new_new_n10675__ & po021;
  assign new_new_n11051__ = pi071 & ~po021;
  assign new_new_n11052__ = ~new_new_n11050__ & ~new_new_n11051__;
  assign new_new_n11053__ = new_new_n11049__ & ~new_new_n11052__;
  assign new_new_n11054__ = ~new_new_n11049__ & new_new_n11052__;
  assign new_new_n11055__ = ~new_new_n11053__ & ~new_new_n11054__;
  assign new_new_n11056__ = ~pi072 & ~new_new_n11055__;
  assign new_new_n11057__ = pi072 & new_new_n11055__;
  assign new_new_n11058__ = ~new_new_n10673__ & po021;
  assign new_new_n11059__ = pi070 & ~po021;
  assign new_new_n11060__ = ~new_new_n11058__ & ~new_new_n11059__;
  assign new_new_n11061__ = ~new_new_n10598__ & ~new_new_n10599__;
  assign new_new_n11062__ = ~new_new_n11060__ & new_new_n11061__;
  assign new_new_n11063__ = new_new_n11060__ & ~new_new_n11061__;
  assign new_new_n11064__ = ~new_new_n11062__ & ~new_new_n11063__;
  assign new_new_n11065__ = ~pi071 & ~new_new_n11064__;
  assign new_new_n11066__ = pi071 & new_new_n11064__;
  assign new_new_n11067__ = ~new_new_n10605__ & ~new_new_n10606__;
  assign new_new_n11068__ = new_new_n10671__ & po021;
  assign new_new_n11069__ = ~pi069 & ~po021;
  assign new_new_n11070__ = ~new_new_n11068__ & ~new_new_n11069__;
  assign new_new_n11071__ = ~new_new_n11067__ & ~new_new_n11070__;
  assign new_new_n11072__ = new_new_n11067__ & new_new_n11070__;
  assign new_new_n11073__ = ~new_new_n11071__ & ~new_new_n11072__;
  assign new_new_n11074__ = ~new_new_n10614__ & ~new_new_n10615__;
  assign new_new_n11075__ = ~new_new_n10669__ & po021;
  assign new_new_n11076__ = pi068 & ~po021;
  assign new_new_n11077__ = ~new_new_n11075__ & ~new_new_n11076__;
  assign new_new_n11078__ = new_new_n11074__ & new_new_n11077__;
  assign new_new_n11079__ = ~new_new_n11074__ & ~new_new_n11077__;
  assign new_new_n11080__ = ~new_new_n11078__ & ~new_new_n11079__;
  assign new_new_n11081__ = pi069 & ~new_new_n11080__;
  assign new_new_n11082__ = ~pi069 & new_new_n11080__;
  assign new_new_n11083__ = ~new_new_n10661__ & ~new_new_n10662__;
  assign new_new_n11084__ = po021 & new_new_n11083__;
  assign new_new_n11085__ = ~pi065 & ~new_new_n10149__;
  assign new_new_n11086__ = ~new_new_n10636__ & new_new_n11085__;
  assign new_new_n11087__ = ~pi022 & ~new_new_n11086__;
  assign new_new_n11088__ = pi065 & new_new_n10149__;
  assign new_new_n11089__ = ~new_new_n11087__ & ~new_new_n11088__;
  assign new_new_n11090__ = pi064 & ~new_new_n11089__;
  assign new_new_n11091__ = pi065 & new_new_n10148__;
  assign new_new_n11092__ = ~new_new_n11090__ & ~new_new_n11091__;
  assign new_new_n11093__ = ~pi066 & ~new_new_n11092__;
  assign new_new_n11094__ = pi066 & new_new_n11092__;
  assign new_new_n11095__ = ~new_new_n11093__ & ~new_new_n11094__;
  assign new_new_n11096__ = po022 & ~new_new_n11095__;
  assign new_new_n11097__ = new_new_n10183__ & ~new_new_n11096__;
  assign new_new_n11098__ = ~new_new_n10183__ & new_new_n11096__;
  assign new_new_n11099__ = ~new_new_n11097__ & ~new_new_n11098__;
  assign new_new_n11100__ = new_new_n11084__ & new_new_n11099__;
  assign new_new_n11101__ = ~new_new_n11084__ & ~new_new_n11099__;
  assign new_new_n11102__ = ~new_new_n11100__ & ~new_new_n11101__;
  assign new_new_n11103__ = ~pi068 & ~new_new_n11102__;
  assign new_new_n11104__ = pi068 & new_new_n11102__;
  assign new_new_n11105__ = ~pi065 & ~po023;
  assign new_new_n11106__ = new_new_n10147__ & new_new_n10629__;
  assign new_new_n11107__ = ~new_new_n11105__ & ~new_new_n11106__;
  assign new_new_n11108__ = pi022 & ~new_new_n11107__;
  assign new_new_n11109__ = ~new_new_n332__ & po022;
  assign new_new_n11110__ = ~new_new_n10147__ & ~new_new_n11109__;
  assign new_new_n11111__ = po023 & ~po022;
  assign new_new_n11112__ = ~new_new_n426__ & ~po023;
  assign new_new_n11113__ = ~pi022 & ~new_new_n10164__;
  assign new_new_n11114__ = ~new_new_n11112__ & new_new_n11113__;
  assign new_new_n11115__ = ~new_new_n11111__ & new_new_n11114__;
  assign new_new_n11116__ = ~new_new_n11110__ & ~new_new_n11115__;
  assign new_new_n11117__ = ~new_new_n11108__ & new_new_n11116__;
  assign new_new_n11118__ = ~pi023 & ~new_new_n11117__;
  assign new_new_n11119__ = ~new_new_n10164__ & ~new_new_n11105__;
  assign new_new_n11120__ = new_new_n10631__ & ~new_new_n11119__;
  assign new_new_n11121__ = ~new_new_n11111__ & ~new_new_n11120__;
  assign new_new_n11122__ = pi064 & ~new_new_n11121__;
  assign new_new_n11123__ = ~new_new_n10147__ & ~new_new_n10629__;
  assign new_new_n11124__ = pi022 & ~new_new_n10164__;
  assign new_new_n11125__ = pi064 & ~new_new_n11124__;
  assign new_new_n11126__ = ~new_new_n11123__ & ~new_new_n11125__;
  assign new_new_n11127__ = ~new_new_n11122__ & ~new_new_n11126__;
  assign new_new_n11128__ = pi023 & ~new_new_n11127__;
  assign new_new_n11129__ = ~new_new_n11118__ & ~new_new_n11128__;
  assign new_new_n11130__ = pi021 & ~new_new_n10646__;
  assign new_new_n11131__ = pi065 & ~new_new_n11130__;
  assign new_new_n11132__ = ~pi022 & po022;
  assign new_new_n11133__ = ~pi021 & ~new_new_n10626__;
  assign new_new_n11134__ = ~new_new_n11132__ & new_new_n11133__;
  assign new_new_n11135__ = ~new_new_n11131__ & ~new_new_n11134__;
  assign new_new_n11136__ = pi064 & ~new_new_n11135__;
  assign new_new_n11137__ = pi064 & po022;
  assign new_new_n11138__ = new_new_n10641__ & ~new_new_n11137__;
  assign new_new_n11139__ = ~new_new_n11136__ & ~new_new_n11138__;
  assign new_new_n11140__ = ~pi066 & new_new_n11139__;
  assign new_new_n11141__ = pi066 & ~new_new_n11139__;
  assign new_new_n11142__ = ~new_new_n11140__ & ~new_new_n11141__;
  assign new_new_n11143__ = po021 & new_new_n11142__;
  assign new_new_n11144__ = new_new_n11129__ & ~new_new_n11143__;
  assign new_new_n11145__ = ~new_new_n11129__ & new_new_n11143__;
  assign new_new_n11146__ = ~new_new_n11144__ & ~new_new_n11145__;
  assign new_new_n11147__ = ~pi067 & ~new_new_n11146__;
  assign new_new_n11148__ = pi067 & new_new_n11146__;
  assign new_new_n11149__ = ~pi021 & ~po021;
  assign new_new_n11150__ = ~pi065 & ~new_new_n11149__;
  assign new_new_n11151__ = ~pi020 & ~new_new_n11150__;
  assign new_new_n11152__ = pi020 & ~pi065;
  assign new_new_n11153__ = pi021 & ~new_new_n11152__;
  assign new_new_n11154__ = po021 & new_new_n11153__;
  assign new_new_n11155__ = ~new_new_n11151__ & ~new_new_n11154__;
  assign new_new_n11156__ = pi064 & ~new_new_n11155__;
  assign new_new_n11157__ = pi064 & po021;
  assign new_new_n11158__ = ~pi021 & ~new_new_n11157__;
  assign new_new_n11159__ = pi065 & new_new_n11158__;
  assign new_new_n11160__ = ~new_new_n11156__ & ~new_new_n11159__;
  assign new_new_n11161__ = ~pi066 & new_new_n11160__;
  assign new_new_n11162__ = pi066 & ~new_new_n11160__;
  assign new_new_n11163__ = new_new_n403__ & po021;
  assign new_new_n11164__ = po022 & new_new_n10758__;
  assign new_new_n11165__ = ~pi065 & ~po021;
  assign new_new_n11166__ = ~new_new_n10629__ & ~new_new_n10630__;
  assign new_new_n11167__ = ~pi021 & ~new_new_n11166__;
  assign new_new_n11168__ = ~new_new_n11165__ & new_new_n11167__;
  assign new_new_n11169__ = ~new_new_n11164__ & ~new_new_n11168__;
  assign new_new_n11170__ = pi064 & ~new_new_n11169__;
  assign new_new_n11171__ = pi065 & po021;
  assign new_new_n11172__ = ~new_new_n11137__ & ~new_new_n11171__;
  assign new_new_n11173__ = new_new_n10632__ & ~new_new_n11172__;
  assign new_new_n11174__ = ~new_new_n11163__ & ~new_new_n11173__;
  assign new_new_n11175__ = ~new_new_n11170__ & new_new_n11174__;
  assign new_new_n11176__ = ~pi022 & ~new_new_n11175__;
  assign new_new_n11177__ = pi022 & new_new_n11175__;
  assign new_new_n11178__ = ~new_new_n11176__ & ~new_new_n11177__;
  assign new_new_n11179__ = ~new_new_n11162__ & ~new_new_n11178__;
  assign new_new_n11180__ = ~new_new_n11161__ & ~new_new_n11179__;
  assign new_new_n11181__ = ~new_new_n11148__ & ~new_new_n11180__;
  assign new_new_n11182__ = ~new_new_n11147__ & ~new_new_n11181__;
  assign new_new_n11183__ = ~new_new_n11104__ & ~new_new_n11182__;
  assign new_new_n11184__ = ~new_new_n11103__ & ~new_new_n11183__;
  assign new_new_n11185__ = ~new_new_n11082__ & new_new_n11184__;
  assign new_new_n11186__ = ~new_new_n11081__ & ~new_new_n11185__;
  assign new_new_n11187__ = ~pi070 & new_new_n11186__;
  assign new_new_n11188__ = new_new_n11073__ & ~new_new_n11187__;
  assign new_new_n11189__ = pi070 & ~new_new_n11186__;
  assign new_new_n11190__ = ~new_new_n11188__ & ~new_new_n11189__;
  assign new_new_n11191__ = ~new_new_n11066__ & new_new_n11190__;
  assign new_new_n11192__ = ~new_new_n11065__ & ~new_new_n11191__;
  assign new_new_n11193__ = ~new_new_n11057__ & ~new_new_n11192__;
  assign new_new_n11194__ = ~new_new_n11056__ & ~new_new_n11193__;
  assign new_new_n11195__ = ~new_new_n11048__ & ~new_new_n11194__;
  assign new_new_n11196__ = ~new_new_n11047__ & ~new_new_n11195__;
  assign new_new_n11197__ = ~new_new_n11039__ & ~new_new_n11196__;
  assign new_new_n11198__ = ~new_new_n11038__ & ~new_new_n11197__;
  assign new_new_n11199__ = ~new_new_n11030__ & ~new_new_n11198__;
  assign new_new_n11200__ = ~new_new_n11029__ & ~new_new_n11199__;
  assign new_new_n11201__ = ~new_new_n11021__ & ~new_new_n11200__;
  assign new_new_n11202__ = ~new_new_n11020__ & ~new_new_n11201__;
  assign new_new_n11203__ = ~new_new_n11012__ & ~new_new_n11202__;
  assign new_new_n11204__ = ~new_new_n11011__ & ~new_new_n11203__;
  assign new_new_n11205__ = ~new_new_n11003__ & new_new_n11204__;
  assign new_new_n11206__ = ~new_new_n11002__ & ~new_new_n11205__;
  assign new_new_n11207__ = ~new_new_n10994__ & ~new_new_n11206__;
  assign new_new_n11208__ = ~new_new_n10993__ & ~new_new_n11207__;
  assign new_new_n11209__ = ~new_new_n10985__ & ~new_new_n11208__;
  assign new_new_n11210__ = ~new_new_n10984__ & ~new_new_n11209__;
  assign new_new_n11211__ = ~new_new_n10976__ & new_new_n11210__;
  assign new_new_n11212__ = ~new_new_n10975__ & ~new_new_n11211__;
  assign new_new_n11213__ = ~new_new_n10967__ & ~new_new_n11212__;
  assign new_new_n11214__ = ~new_new_n10966__ & ~new_new_n11213__;
  assign new_new_n11215__ = ~new_new_n10958__ & new_new_n11214__;
  assign new_new_n11216__ = ~new_new_n10957__ & ~new_new_n11215__;
  assign new_new_n11217__ = ~new_new_n10949__ & new_new_n11216__;
  assign new_new_n11218__ = ~new_new_n10948__ & ~new_new_n11217__;
  assign new_new_n11219__ = ~new_new_n10940__ & ~new_new_n11218__;
  assign new_new_n11220__ = ~new_new_n10939__ & ~new_new_n11219__;
  assign new_new_n11221__ = ~new_new_n10931__ & ~new_new_n11220__;
  assign new_new_n11222__ = ~new_new_n10930__ & ~new_new_n11221__;
  assign new_new_n11223__ = ~new_new_n10922__ & ~new_new_n11222__;
  assign new_new_n11224__ = ~new_new_n10921__ & ~new_new_n11223__;
  assign new_new_n11225__ = ~new_new_n10913__ & ~new_new_n11224__;
  assign new_new_n11226__ = ~new_new_n10912__ & ~new_new_n11225__;
  assign new_new_n11227__ = ~new_new_n10904__ & ~new_new_n11226__;
  assign new_new_n11228__ = ~new_new_n10903__ & ~new_new_n11227__;
  assign new_new_n11229__ = ~new_new_n10895__ & ~new_new_n11228__;
  assign new_new_n11230__ = ~new_new_n10894__ & ~new_new_n11229__;
  assign new_new_n11231__ = ~new_new_n10886__ & ~new_new_n11230__;
  assign new_new_n11232__ = ~new_new_n10885__ & ~new_new_n11231__;
  assign new_new_n11233__ = ~new_new_n10877__ & new_new_n11232__;
  assign new_new_n11234__ = ~new_new_n10876__ & ~new_new_n11233__;
  assign new_new_n11235__ = ~new_new_n10868__ & new_new_n11234__;
  assign new_new_n11236__ = ~new_new_n10867__ & ~new_new_n11235__;
  assign new_new_n11237__ = ~new_new_n10859__ & ~new_new_n11236__;
  assign new_new_n11238__ = ~new_new_n10858__ & ~new_new_n11237__;
  assign new_new_n11239__ = ~new_new_n10850__ & ~new_new_n11238__;
  assign new_new_n11240__ = ~new_new_n10849__ & ~new_new_n11239__;
  assign new_new_n11241__ = ~new_new_n10841__ & new_new_n11240__;
  assign new_new_n11242__ = ~new_new_n10840__ & ~new_new_n11241__;
  assign new_new_n11243__ = ~new_new_n10832__ & new_new_n11242__;
  assign new_new_n11244__ = ~new_new_n10831__ & ~new_new_n11243__;
  assign new_new_n11245__ = ~new_new_n10823__ & ~new_new_n11244__;
  assign new_new_n11246__ = ~new_new_n10822__ & ~new_new_n11245__;
  assign new_new_n11247__ = ~new_new_n10814__ & ~new_new_n11246__;
  assign new_new_n11248__ = ~new_new_n10813__ & ~new_new_n11247__;
  assign new_new_n11249__ = ~new_new_n10805__ & new_new_n11248__;
  assign new_new_n11250__ = ~new_new_n10804__ & ~new_new_n11249__;
  assign new_new_n11251__ = ~new_new_n10796__ & ~new_new_n11250__;
  assign new_new_n11252__ = ~new_new_n10795__ & ~new_new_n11251__;
  assign new_new_n11253__ = ~pi102 & new_new_n11252__;
  assign new_new_n11254__ = pi102 & ~new_new_n11252__;
  assign new_new_n11255__ = ~new_new_n10735__ & po021;
  assign new_new_n11256__ = pi101 & ~po021;
  assign new_new_n11257__ = ~new_new_n11255__ & ~new_new_n11256__;
  assign new_new_n11258__ = ~new_new_n10319__ & ~new_new_n10320__;
  assign new_new_n11259__ = ~new_new_n11257__ & new_new_n11258__;
  assign new_new_n11260__ = new_new_n11257__ & ~new_new_n11258__;
  assign new_new_n11261__ = ~new_new_n11259__ & ~new_new_n11260__;
  assign new_new_n11262__ = ~new_new_n11254__ & ~new_new_n11261__;
  assign new_new_n11263__ = ~new_new_n11253__ & ~new_new_n11262__;
  assign new_new_n11264__ = ~new_new_n10787__ & ~new_new_n11263__;
  assign new_new_n11265__ = ~new_new_n10786__ & ~new_new_n11264__;
  assign new_new_n11266__ = ~new_new_n10778__ & ~new_new_n11265__;
  assign new_new_n11267__ = ~new_new_n10777__ & ~new_new_n11266__;
  assign new_new_n11268__ = ~pi107 & new_new_n10752__;
  assign new_new_n11269__ = ~pi105 & ~new_new_n10743__;
  assign new_new_n11270__ = pi105 & new_new_n10743__;
  assign new_new_n11271__ = ~new_new_n11269__ & ~new_new_n11270__;
  assign new_new_n11272__ = po021 & new_new_n11271__;
  assign new_new_n11273__ = new_new_n10282__ & new_new_n11272__;
  assign new_new_n11274__ = ~new_new_n10282__ & ~new_new_n11272__;
  assign new_new_n11275__ = ~new_new_n11273__ & ~new_new_n11274__;
  assign new_new_n11276__ = ~pi106 & ~new_new_n11275__;
  assign new_new_n11277__ = pi106 & new_new_n11275__;
  assign new_new_n11278__ = ~new_new_n10767__ & ~new_new_n11267__;
  assign new_new_n11279__ = ~new_new_n10768__ & ~new_new_n11278__;
  assign new_new_n11280__ = ~new_new_n11277__ & ~new_new_n11279__;
  assign new_new_n11281__ = ~new_new_n11276__ & ~new_new_n11280__;
  assign new_new_n11282__ = ~new_new_n11268__ & new_new_n11281__;
  assign new_new_n11283__ = pi107 & ~new_new_n9808__;
  assign new_new_n11284__ = ~pi108 & new_new_n10753__;
  assign new_new_n11285__ = ~new_new_n11283__ & new_new_n11284__;
  assign po020 = ~new_new_n11282__ & new_new_n11285__;
  assign new_new_n11287__ = ~new_new_n11267__ & po020;
  assign new_new_n11288__ = ~pi105 & ~po020;
  assign new_new_n11289__ = ~new_new_n11287__ & ~new_new_n11288__;
  assign new_new_n11290__ = new_new_n10769__ & ~new_new_n11289__;
  assign new_new_n11291__ = ~new_new_n10769__ & new_new_n11289__;
  assign new_new_n11292__ = ~new_new_n11290__ & ~new_new_n11291__;
  assign new_new_n11293__ = pi106 & ~new_new_n11292__;
  assign new_new_n11294__ = ~pi106 & new_new_n11292__;
  assign new_new_n11295__ = ~pi104 & ~new_new_n11265__;
  assign new_new_n11296__ = pi104 & new_new_n11265__;
  assign new_new_n11297__ = ~new_new_n11295__ & ~new_new_n11296__;
  assign new_new_n11298__ = po020 & new_new_n11297__;
  assign new_new_n11299__ = new_new_n10776__ & new_new_n11298__;
  assign new_new_n11300__ = ~new_new_n10776__ & ~new_new_n11298__;
  assign new_new_n11301__ = ~new_new_n11299__ & ~new_new_n11300__;
  assign new_new_n11302__ = pi105 & new_new_n11301__;
  assign new_new_n11303__ = ~pi105 & ~new_new_n11301__;
  assign new_new_n11304__ = ~new_new_n10786__ & ~new_new_n10787__;
  assign new_new_n11305__ = ~new_new_n11263__ & po020;
  assign new_new_n11306__ = ~pi103 & ~po020;
  assign new_new_n11307__ = ~new_new_n11305__ & ~new_new_n11306__;
  assign new_new_n11308__ = new_new_n11304__ & ~new_new_n11307__;
  assign new_new_n11309__ = ~new_new_n11304__ & new_new_n11307__;
  assign new_new_n11310__ = ~new_new_n11308__ & ~new_new_n11309__;
  assign new_new_n11311__ = pi104 & ~new_new_n11310__;
  assign new_new_n11312__ = ~pi104 & new_new_n11310__;
  assign new_new_n11313__ = ~new_new_n11253__ & ~new_new_n11254__;
  assign new_new_n11314__ = po020 & new_new_n11313__;
  assign new_new_n11315__ = new_new_n11261__ & new_new_n11314__;
  assign new_new_n11316__ = ~new_new_n11261__ & ~new_new_n11314__;
  assign new_new_n11317__ = ~new_new_n11315__ & ~new_new_n11316__;
  assign new_new_n11318__ = ~pi103 & ~new_new_n11317__;
  assign new_new_n11319__ = pi103 & new_new_n11317__;
  assign new_new_n11320__ = pi101 & ~new_new_n11250__;
  assign new_new_n11321__ = ~pi101 & new_new_n11250__;
  assign new_new_n11322__ = ~new_new_n11320__ & ~new_new_n11321__;
  assign new_new_n11323__ = po020 & new_new_n11322__;
  assign new_new_n11324__ = new_new_n10794__ & new_new_n11323__;
  assign new_new_n11325__ = ~new_new_n10794__ & ~new_new_n11323__;
  assign new_new_n11326__ = ~new_new_n11324__ & ~new_new_n11325__;
  assign new_new_n11327__ = pi102 & ~new_new_n11326__;
  assign new_new_n11328__ = ~pi102 & new_new_n11326__;
  assign new_new_n11329__ = ~new_new_n10804__ & ~new_new_n10805__;
  assign new_new_n11330__ = ~new_new_n11248__ & po020;
  assign new_new_n11331__ = ~pi100 & ~po020;
  assign new_new_n11332__ = ~new_new_n11330__ & ~new_new_n11331__;
  assign new_new_n11333__ = new_new_n11329__ & ~new_new_n11332__;
  assign new_new_n11334__ = ~new_new_n11329__ & new_new_n11332__;
  assign new_new_n11335__ = ~new_new_n11333__ & ~new_new_n11334__;
  assign new_new_n11336__ = pi101 & ~new_new_n11335__;
  assign new_new_n11337__ = ~pi101 & new_new_n11335__;
  assign new_new_n11338__ = ~new_new_n10813__ & ~new_new_n10814__;
  assign new_new_n11339__ = ~new_new_n11246__ & po020;
  assign new_new_n11340__ = ~pi099 & ~po020;
  assign new_new_n11341__ = ~new_new_n11339__ & ~new_new_n11340__;
  assign new_new_n11342__ = new_new_n11338__ & ~new_new_n11341__;
  assign new_new_n11343__ = ~new_new_n11338__ & new_new_n11341__;
  assign new_new_n11344__ = ~new_new_n11342__ & ~new_new_n11343__;
  assign new_new_n11345__ = pi100 & ~new_new_n11344__;
  assign new_new_n11346__ = ~pi100 & new_new_n11344__;
  assign new_new_n11347__ = ~pi098 & ~new_new_n11244__;
  assign new_new_n11348__ = pi098 & new_new_n11244__;
  assign new_new_n11349__ = ~new_new_n11347__ & ~new_new_n11348__;
  assign new_new_n11350__ = po020 & new_new_n11349__;
  assign new_new_n11351__ = new_new_n10821__ & ~new_new_n11350__;
  assign new_new_n11352__ = ~new_new_n10821__ & new_new_n11350__;
  assign new_new_n11353__ = ~new_new_n11351__ & ~new_new_n11352__;
  assign new_new_n11354__ = pi099 & ~new_new_n11353__;
  assign new_new_n11355__ = ~pi099 & new_new_n11353__;
  assign new_new_n11356__ = ~new_new_n11242__ & po020;
  assign new_new_n11357__ = pi097 & ~po020;
  assign new_new_n11358__ = ~new_new_n11356__ & ~new_new_n11357__;
  assign new_new_n11359__ = ~new_new_n10831__ & ~new_new_n10832__;
  assign new_new_n11360__ = ~new_new_n11358__ & new_new_n11359__;
  assign new_new_n11361__ = new_new_n11358__ & ~new_new_n11359__;
  assign new_new_n11362__ = ~new_new_n11360__ & ~new_new_n11361__;
  assign new_new_n11363__ = ~pi098 & ~new_new_n11362__;
  assign new_new_n11364__ = pi098 & new_new_n11362__;
  assign new_new_n11365__ = ~new_new_n10840__ & ~new_new_n10841__;
  assign new_new_n11366__ = ~new_new_n11240__ & po020;
  assign new_new_n11367__ = ~pi096 & ~po020;
  assign new_new_n11368__ = ~new_new_n11366__ & ~new_new_n11367__;
  assign new_new_n11369__ = new_new_n11365__ & ~new_new_n11368__;
  assign new_new_n11370__ = ~new_new_n11365__ & new_new_n11368__;
  assign new_new_n11371__ = ~new_new_n11369__ & ~new_new_n11370__;
  assign new_new_n11372__ = ~pi097 & new_new_n11371__;
  assign new_new_n11373__ = pi097 & ~new_new_n11371__;
  assign new_new_n11374__ = ~pi095 & ~new_new_n11238__;
  assign new_new_n11375__ = pi095 & new_new_n11238__;
  assign new_new_n11376__ = ~new_new_n11374__ & ~new_new_n11375__;
  assign new_new_n11377__ = po020 & new_new_n11376__;
  assign new_new_n11378__ = new_new_n10848__ & new_new_n11377__;
  assign new_new_n11379__ = ~new_new_n10848__ & ~new_new_n11377__;
  assign new_new_n11380__ = ~new_new_n11378__ & ~new_new_n11379__;
  assign new_new_n11381__ = ~pi096 & ~new_new_n11380__;
  assign new_new_n11382__ = pi096 & new_new_n11380__;
  assign new_new_n11383__ = ~new_new_n10858__ & ~new_new_n10859__;
  assign new_new_n11384__ = ~new_new_n11236__ & po020;
  assign new_new_n11385__ = ~pi094 & ~po020;
  assign new_new_n11386__ = ~new_new_n11384__ & ~new_new_n11385__;
  assign new_new_n11387__ = ~new_new_n11383__ & ~new_new_n11386__;
  assign new_new_n11388__ = new_new_n11383__ & new_new_n11386__;
  assign new_new_n11389__ = ~new_new_n11387__ & ~new_new_n11388__;
  assign new_new_n11390__ = ~pi095 & ~new_new_n11389__;
  assign new_new_n11391__ = pi095 & new_new_n11389__;
  assign new_new_n11392__ = new_new_n11234__ & po020;
  assign new_new_n11393__ = ~pi093 & ~po020;
  assign new_new_n11394__ = ~new_new_n11392__ & ~new_new_n11393__;
  assign new_new_n11395__ = ~new_new_n10867__ & ~new_new_n10868__;
  assign new_new_n11396__ = ~new_new_n11394__ & ~new_new_n11395__;
  assign new_new_n11397__ = new_new_n11394__ & new_new_n11395__;
  assign new_new_n11398__ = ~new_new_n11396__ & ~new_new_n11397__;
  assign new_new_n11399__ = pi094 & new_new_n11398__;
  assign new_new_n11400__ = ~pi094 & ~new_new_n11398__;
  assign new_new_n11401__ = ~new_new_n10876__ & ~new_new_n10877__;
  assign new_new_n11402__ = ~new_new_n11232__ & po020;
  assign new_new_n11403__ = ~pi092 & ~po020;
  assign new_new_n11404__ = ~new_new_n11402__ & ~new_new_n11403__;
  assign new_new_n11405__ = new_new_n11401__ & ~new_new_n11404__;
  assign new_new_n11406__ = ~new_new_n11401__ & new_new_n11404__;
  assign new_new_n11407__ = ~new_new_n11405__ & ~new_new_n11406__;
  assign new_new_n11408__ = pi093 & ~new_new_n11407__;
  assign new_new_n11409__ = ~pi093 & new_new_n11407__;
  assign new_new_n11410__ = ~new_new_n10885__ & ~new_new_n10886__;
  assign new_new_n11411__ = ~new_new_n11230__ & po020;
  assign new_new_n11412__ = ~pi091 & ~po020;
  assign new_new_n11413__ = ~new_new_n11411__ & ~new_new_n11412__;
  assign new_new_n11414__ = new_new_n11410__ & ~new_new_n11413__;
  assign new_new_n11415__ = ~new_new_n11410__ & new_new_n11413__;
  assign new_new_n11416__ = ~new_new_n11414__ & ~new_new_n11415__;
  assign new_new_n11417__ = ~pi092 & new_new_n11416__;
  assign new_new_n11418__ = pi092 & ~new_new_n11416__;
  assign new_new_n11419__ = ~pi090 & ~new_new_n11228__;
  assign new_new_n11420__ = pi090 & new_new_n11228__;
  assign new_new_n11421__ = ~new_new_n11419__ & ~new_new_n11420__;
  assign new_new_n11422__ = po020 & new_new_n11421__;
  assign new_new_n11423__ = new_new_n10893__ & new_new_n11422__;
  assign new_new_n11424__ = ~new_new_n10893__ & ~new_new_n11422__;
  assign new_new_n11425__ = ~new_new_n11423__ & ~new_new_n11424__;
  assign new_new_n11426__ = ~pi091 & ~new_new_n11425__;
  assign new_new_n11427__ = pi091 & new_new_n11425__;
  assign new_new_n11428__ = ~pi089 & ~new_new_n11226__;
  assign new_new_n11429__ = pi089 & new_new_n11226__;
  assign new_new_n11430__ = ~new_new_n11428__ & ~new_new_n11429__;
  assign new_new_n11431__ = po020 & new_new_n11430__;
  assign new_new_n11432__ = new_new_n10902__ & new_new_n11431__;
  assign new_new_n11433__ = ~new_new_n10902__ & ~new_new_n11431__;
  assign new_new_n11434__ = ~new_new_n11432__ & ~new_new_n11433__;
  assign new_new_n11435__ = ~pi090 & ~new_new_n11434__;
  assign new_new_n11436__ = pi090 & new_new_n11434__;
  assign new_new_n11437__ = ~new_new_n10912__ & ~new_new_n10913__;
  assign new_new_n11438__ = ~new_new_n11224__ & po020;
  assign new_new_n11439__ = ~pi088 & ~po020;
  assign new_new_n11440__ = ~new_new_n11438__ & ~new_new_n11439__;
  assign new_new_n11441__ = new_new_n11437__ & ~new_new_n11440__;
  assign new_new_n11442__ = ~new_new_n11437__ & new_new_n11440__;
  assign new_new_n11443__ = ~new_new_n11441__ & ~new_new_n11442__;
  assign new_new_n11444__ = pi089 & ~new_new_n11443__;
  assign new_new_n11445__ = ~pi089 & new_new_n11443__;
  assign new_new_n11446__ = ~new_new_n10921__ & ~new_new_n10922__;
  assign new_new_n11447__ = ~new_new_n11222__ & po020;
  assign new_new_n11448__ = ~pi087 & ~po020;
  assign new_new_n11449__ = ~new_new_n11447__ & ~new_new_n11448__;
  assign new_new_n11450__ = new_new_n11446__ & ~new_new_n11449__;
  assign new_new_n11451__ = ~new_new_n11446__ & new_new_n11449__;
  assign new_new_n11452__ = ~new_new_n11450__ & ~new_new_n11451__;
  assign new_new_n11453__ = pi088 & ~new_new_n11452__;
  assign new_new_n11454__ = ~pi088 & new_new_n11452__;
  assign new_new_n11455__ = ~new_new_n10930__ & ~new_new_n10931__;
  assign new_new_n11456__ = ~new_new_n11220__ & po020;
  assign new_new_n11457__ = ~pi086 & ~po020;
  assign new_new_n11458__ = ~new_new_n11456__ & ~new_new_n11457__;
  assign new_new_n11459__ = new_new_n11455__ & ~new_new_n11458__;
  assign new_new_n11460__ = ~new_new_n11455__ & new_new_n11458__;
  assign new_new_n11461__ = ~new_new_n11459__ & ~new_new_n11460__;
  assign new_new_n11462__ = pi087 & ~new_new_n11461__;
  assign new_new_n11463__ = ~pi087 & new_new_n11461__;
  assign new_new_n11464__ = ~new_new_n10939__ & ~new_new_n10940__;
  assign new_new_n11465__ = ~new_new_n11218__ & po020;
  assign new_new_n11466__ = ~pi085 & ~po020;
  assign new_new_n11467__ = ~new_new_n11465__ & ~new_new_n11466__;
  assign new_new_n11468__ = new_new_n11464__ & ~new_new_n11467__;
  assign new_new_n11469__ = ~new_new_n11464__ & new_new_n11467__;
  assign new_new_n11470__ = ~new_new_n11468__ & ~new_new_n11469__;
  assign new_new_n11471__ = ~pi086 & new_new_n11470__;
  assign new_new_n11472__ = pi086 & ~new_new_n11470__;
  assign new_new_n11473__ = ~new_new_n11216__ & po020;
  assign new_new_n11474__ = pi084 & ~po020;
  assign new_new_n11475__ = ~new_new_n11473__ & ~new_new_n11474__;
  assign new_new_n11476__ = ~new_new_n10948__ & ~new_new_n10949__;
  assign new_new_n11477__ = ~new_new_n11475__ & new_new_n11476__;
  assign new_new_n11478__ = new_new_n11475__ & ~new_new_n11476__;
  assign new_new_n11479__ = ~new_new_n11477__ & ~new_new_n11478__;
  assign new_new_n11480__ = ~pi085 & ~new_new_n11479__;
  assign new_new_n11481__ = pi085 & new_new_n11479__;
  assign new_new_n11482__ = ~new_new_n10957__ & ~new_new_n10958__;
  assign new_new_n11483__ = ~new_new_n11214__ & po020;
  assign new_new_n11484__ = ~pi083 & ~po020;
  assign new_new_n11485__ = ~new_new_n11483__ & ~new_new_n11484__;
  assign new_new_n11486__ = new_new_n11482__ & ~new_new_n11485__;
  assign new_new_n11487__ = ~new_new_n11482__ & new_new_n11485__;
  assign new_new_n11488__ = ~new_new_n11486__ & ~new_new_n11487__;
  assign new_new_n11489__ = ~pi084 & new_new_n11488__;
  assign new_new_n11490__ = pi084 & ~new_new_n11488__;
  assign new_new_n11491__ = ~pi082 & ~new_new_n11212__;
  assign new_new_n11492__ = pi082 & new_new_n11212__;
  assign new_new_n11493__ = ~new_new_n11491__ & ~new_new_n11492__;
  assign new_new_n11494__ = po020 & new_new_n11493__;
  assign new_new_n11495__ = new_new_n10965__ & new_new_n11494__;
  assign new_new_n11496__ = ~new_new_n10965__ & ~new_new_n11494__;
  assign new_new_n11497__ = ~new_new_n11495__ & ~new_new_n11496__;
  assign new_new_n11498__ = ~pi083 & ~new_new_n11497__;
  assign new_new_n11499__ = pi083 & new_new_n11497__;
  assign new_new_n11500__ = ~new_new_n11210__ & po020;
  assign new_new_n11501__ = pi081 & ~po020;
  assign new_new_n11502__ = ~new_new_n11500__ & ~new_new_n11501__;
  assign new_new_n11503__ = ~new_new_n10975__ & ~new_new_n10976__;
  assign new_new_n11504__ = ~new_new_n11502__ & new_new_n11503__;
  assign new_new_n11505__ = new_new_n11502__ & ~new_new_n11503__;
  assign new_new_n11506__ = ~new_new_n11504__ & ~new_new_n11505__;
  assign new_new_n11507__ = ~pi082 & ~new_new_n11506__;
  assign new_new_n11508__ = pi082 & new_new_n11506__;
  assign new_new_n11509__ = pi080 & ~new_new_n11208__;
  assign new_new_n11510__ = ~pi080 & new_new_n11208__;
  assign new_new_n11511__ = ~new_new_n11509__ & ~new_new_n11510__;
  assign new_new_n11512__ = po020 & new_new_n11511__;
  assign new_new_n11513__ = new_new_n10983__ & new_new_n11512__;
  assign new_new_n11514__ = ~new_new_n10983__ & ~new_new_n11512__;
  assign new_new_n11515__ = ~new_new_n11513__ & ~new_new_n11514__;
  assign new_new_n11516__ = pi081 & ~new_new_n11515__;
  assign new_new_n11517__ = ~pi081 & new_new_n11515__;
  assign new_new_n11518__ = ~new_new_n11206__ & po020;
  assign new_new_n11519__ = pi079 & ~po020;
  assign new_new_n11520__ = ~new_new_n11518__ & ~new_new_n11519__;
  assign new_new_n11521__ = ~new_new_n10993__ & ~new_new_n10994__;
  assign new_new_n11522__ = ~new_new_n11520__ & new_new_n11521__;
  assign new_new_n11523__ = new_new_n11520__ & ~new_new_n11521__;
  assign new_new_n11524__ = ~new_new_n11522__ & ~new_new_n11523__;
  assign new_new_n11525__ = ~pi080 & ~new_new_n11524__;
  assign new_new_n11526__ = pi080 & new_new_n11524__;
  assign new_new_n11527__ = ~new_new_n11002__ & ~new_new_n11003__;
  assign new_new_n11528__ = ~new_new_n11204__ & po020;
  assign new_new_n11529__ = ~pi078 & ~po020;
  assign new_new_n11530__ = ~new_new_n11528__ & ~new_new_n11529__;
  assign new_new_n11531__ = new_new_n11527__ & new_new_n11530__;
  assign new_new_n11532__ = ~new_new_n11527__ & ~new_new_n11530__;
  assign new_new_n11533__ = ~new_new_n11531__ & ~new_new_n11532__;
  assign new_new_n11534__ = pi079 & new_new_n11533__;
  assign new_new_n11535__ = ~pi079 & ~new_new_n11533__;
  assign new_new_n11536__ = new_new_n11202__ & po020;
  assign new_new_n11537__ = pi077 & ~po020;
  assign new_new_n11538__ = ~new_new_n11536__ & ~new_new_n11537__;
  assign new_new_n11539__ = ~new_new_n11011__ & ~new_new_n11012__;
  assign new_new_n11540__ = ~new_new_n11538__ & ~new_new_n11539__;
  assign new_new_n11541__ = new_new_n11538__ & new_new_n11539__;
  assign new_new_n11542__ = ~new_new_n11540__ & ~new_new_n11541__;
  assign new_new_n11543__ = ~pi078 & new_new_n11542__;
  assign new_new_n11544__ = new_new_n11200__ & po020;
  assign new_new_n11545__ = pi076 & ~po020;
  assign new_new_n11546__ = ~new_new_n11544__ & ~new_new_n11545__;
  assign new_new_n11547__ = ~new_new_n11020__ & ~new_new_n11021__;
  assign new_new_n11548__ = ~new_new_n11546__ & ~new_new_n11547__;
  assign new_new_n11549__ = new_new_n11546__ & new_new_n11547__;
  assign new_new_n11550__ = ~new_new_n11548__ & ~new_new_n11549__;
  assign new_new_n11551__ = pi077 & ~new_new_n11550__;
  assign new_new_n11552__ = ~pi077 & new_new_n11550__;
  assign new_new_n11553__ = ~new_new_n11029__ & ~new_new_n11030__;
  assign new_new_n11554__ = ~new_new_n11198__ & po020;
  assign new_new_n11555__ = ~pi075 & ~po020;
  assign new_new_n11556__ = ~new_new_n11554__ & ~new_new_n11555__;
  assign new_new_n11557__ = ~new_new_n11553__ & ~new_new_n11556__;
  assign new_new_n11558__ = new_new_n11553__ & new_new_n11556__;
  assign new_new_n11559__ = ~new_new_n11557__ & ~new_new_n11558__;
  assign new_new_n11560__ = ~pi076 & ~new_new_n11559__;
  assign new_new_n11561__ = pi076 & new_new_n11559__;
  assign new_new_n11562__ = ~new_new_n11038__ & ~new_new_n11039__;
  assign new_new_n11563__ = ~new_new_n11196__ & po020;
  assign new_new_n11564__ = ~pi074 & ~po020;
  assign new_new_n11565__ = ~new_new_n11563__ & ~new_new_n11564__;
  assign new_new_n11566__ = new_new_n11562__ & ~new_new_n11565__;
  assign new_new_n11567__ = ~new_new_n11562__ & new_new_n11565__;
  assign new_new_n11568__ = ~new_new_n11566__ & ~new_new_n11567__;
  assign new_new_n11569__ = ~pi075 & new_new_n11568__;
  assign new_new_n11570__ = pi075 & ~new_new_n11568__;
  assign new_new_n11571__ = ~pi073 & ~new_new_n11194__;
  assign new_new_n11572__ = pi073 & new_new_n11194__;
  assign new_new_n11573__ = ~new_new_n11571__ & ~new_new_n11572__;
  assign new_new_n11574__ = po020 & new_new_n11573__;
  assign new_new_n11575__ = ~new_new_n11046__ & new_new_n11574__;
  assign new_new_n11576__ = new_new_n11046__ & ~new_new_n11574__;
  assign new_new_n11577__ = ~new_new_n11575__ & ~new_new_n11576__;
  assign new_new_n11578__ = ~pi074 & new_new_n11577__;
  assign new_new_n11579__ = pi074 & ~new_new_n11577__;
  assign new_new_n11580__ = ~pi072 & ~new_new_n11192__;
  assign new_new_n11581__ = pi072 & new_new_n11192__;
  assign new_new_n11582__ = ~new_new_n11580__ & ~new_new_n11581__;
  assign new_new_n11583__ = po020 & new_new_n11582__;
  assign new_new_n11584__ = new_new_n11055__ & new_new_n11583__;
  assign new_new_n11585__ = ~new_new_n11055__ & ~new_new_n11583__;
  assign new_new_n11586__ = ~new_new_n11584__ & ~new_new_n11585__;
  assign new_new_n11587__ = ~pi073 & ~new_new_n11586__;
  assign new_new_n11588__ = pi073 & new_new_n11586__;
  assign new_new_n11589__ = ~new_new_n11190__ & po020;
  assign new_new_n11590__ = pi071 & ~po020;
  assign new_new_n11591__ = ~new_new_n11589__ & ~new_new_n11590__;
  assign new_new_n11592__ = ~new_new_n11065__ & ~new_new_n11066__;
  assign new_new_n11593__ = ~new_new_n11591__ & new_new_n11592__;
  assign new_new_n11594__ = new_new_n11591__ & ~new_new_n11592__;
  assign new_new_n11595__ = ~new_new_n11593__ & ~new_new_n11594__;
  assign new_new_n11596__ = ~pi072 & ~new_new_n11595__;
  assign new_new_n11597__ = pi072 & new_new_n11595__;
  assign new_new_n11598__ = ~new_new_n11187__ & ~new_new_n11189__;
  assign new_new_n11599__ = po020 & new_new_n11598__;
  assign new_new_n11600__ = ~new_new_n11073__ & ~new_new_n11599__;
  assign new_new_n11601__ = new_new_n11073__ & new_new_n11599__;
  assign new_new_n11602__ = ~new_new_n11600__ & ~new_new_n11601__;
  assign new_new_n11603__ = ~pi071 & ~new_new_n11602__;
  assign new_new_n11604__ = pi071 & new_new_n11602__;
  assign new_new_n11605__ = ~new_new_n11081__ & ~new_new_n11082__;
  assign new_new_n11606__ = ~new_new_n11184__ & po020;
  assign new_new_n11607__ = ~pi069 & ~po020;
  assign new_new_n11608__ = ~new_new_n11606__ & ~new_new_n11607__;
  assign new_new_n11609__ = new_new_n11605__ & ~new_new_n11608__;
  assign new_new_n11610__ = ~new_new_n11605__ & new_new_n11608__;
  assign new_new_n11611__ = ~new_new_n11609__ & ~new_new_n11610__;
  assign new_new_n11612__ = pi070 & ~new_new_n11611__;
  assign new_new_n11613__ = ~pi070 & new_new_n11611__;
  assign new_new_n11614__ = ~new_new_n11161__ & ~new_new_n11162__;
  assign new_new_n11615__ = po020 & new_new_n11614__;
  assign new_new_n11616__ = ~new_new_n11178__ & ~new_new_n11615__;
  assign new_new_n11617__ = new_new_n11178__ & new_new_n11615__;
  assign new_new_n11618__ = ~new_new_n11616__ & ~new_new_n11617__;
  assign new_new_n11619__ = ~pi067 & ~new_new_n11618__;
  assign new_new_n11620__ = pi067 & new_new_n11618__;
  assign new_new_n11621__ = pi020 & po020;
  assign new_new_n11622__ = pi021 & pi064;
  assign new_new_n11623__ = new_new_n275__ & new_new_n11622__;
  assign new_new_n11624__ = new_new_n10753__ & new_new_n11623__;
  assign new_new_n11625__ = ~new_new_n10758__ & new_new_n11624__;
  assign new_new_n11626__ = ~new_new_n11158__ & ~new_new_n11625__;
  assign new_new_n11627__ = pi065 & new_new_n11626__;
  assign new_new_n11628__ = ~pi065 & ~new_new_n11626__;
  assign new_new_n11629__ = ~pi019 & new_new_n11628__;
  assign new_new_n11630__ = ~new_new_n11627__ & ~new_new_n11629__;
  assign new_new_n11631__ = new_new_n11621__ & ~new_new_n11630__;
  assign new_new_n11632__ = ~pi020 & pi065;
  assign new_new_n11633__ = po020 & ~new_new_n11632__;
  assign new_new_n11634__ = ~pi019 & ~new_new_n11152__;
  assign new_new_n11635__ = ~new_new_n11626__ & new_new_n11634__;
  assign new_new_n11636__ = ~new_new_n11633__ & new_new_n11635__;
  assign new_new_n11637__ = ~new_new_n11631__ & ~new_new_n11636__;
  assign new_new_n11638__ = pi064 & ~new_new_n11637__;
  assign new_new_n11639__ = po020 & ~new_new_n11626__;
  assign new_new_n11640__ = pi064 & po020;
  assign new_new_n11641__ = new_new_n11632__ & ~new_new_n11640__;
  assign new_new_n11642__ = ~po020 & new_new_n11626__;
  assign new_new_n11643__ = ~new_new_n11639__ & ~new_new_n11642__;
  assign new_new_n11644__ = new_new_n11641__ & new_new_n11643__;
  assign new_new_n11645__ = ~pi066 & ~new_new_n11644__;
  assign new_new_n11646__ = ~new_new_n11638__ & new_new_n11645__;
  assign new_new_n11647__ = pi065 & po020;
  assign new_new_n11648__ = pi019 & ~new_new_n11647__;
  assign new_new_n11649__ = ~pi065 & ~po020;
  assign new_new_n11650__ = ~pi020 & ~new_new_n11649__;
  assign new_new_n11651__ = new_new_n11648__ & ~new_new_n11650__;
  assign new_new_n11652__ = pi020 & ~po020;
  assign new_new_n11653__ = ~new_new_n426__ & new_new_n11652__;
  assign new_new_n11654__ = ~new_new_n332__ & ~new_new_n11653__;
  assign new_new_n11655__ = ~new_new_n11651__ & new_new_n11654__;
  assign new_new_n11656__ = new_new_n11626__ & ~new_new_n11655__;
  assign new_new_n11657__ = new_new_n403__ & ~new_new_n11626__;
  assign new_new_n11658__ = pi020 & ~new_new_n11657__;
  assign new_new_n11659__ = pi019 & new_new_n11627__;
  assign new_new_n11660__ = ~new_new_n11628__ & ~new_new_n11659__;
  assign new_new_n11661__ = pi064 & ~new_new_n11660__;
  assign new_new_n11662__ = ~pi020 & ~new_new_n11661__;
  assign new_new_n11663__ = ~new_new_n11658__ & ~new_new_n11662__;
  assign new_new_n11664__ = po020 & new_new_n11663__;
  assign new_new_n11665__ = ~new_new_n11646__ & ~new_new_n11664__;
  assign new_new_n11666__ = ~new_new_n11656__ & new_new_n11665__;
  assign new_new_n11667__ = ~new_new_n11620__ & ~new_new_n11666__;
  assign new_new_n11668__ = ~new_new_n11619__ & ~new_new_n11667__;
  assign new_new_n11669__ = pi068 & new_new_n11668__;
  assign new_new_n11670__ = ~new_new_n11147__ & ~new_new_n11148__;
  assign new_new_n11671__ = ~new_new_n11180__ & po020;
  assign new_new_n11672__ = ~pi067 & ~po020;
  assign new_new_n11673__ = ~new_new_n11671__ & ~new_new_n11672__;
  assign new_new_n11674__ = new_new_n11670__ & ~new_new_n11673__;
  assign new_new_n11675__ = ~new_new_n11670__ & new_new_n11673__;
  assign new_new_n11676__ = ~new_new_n11674__ & ~new_new_n11675__;
  assign new_new_n11677__ = ~new_new_n11669__ & new_new_n11676__;
  assign new_new_n11678__ = ~pi068 & ~new_new_n11668__;
  assign new_new_n11679__ = ~new_new_n11677__ & ~new_new_n11678__;
  assign new_new_n11680__ = pi069 & new_new_n11679__;
  assign new_new_n11681__ = ~pi069 & ~new_new_n11679__;
  assign new_new_n11682__ = ~new_new_n11103__ & ~new_new_n11104__;
  assign new_new_n11683__ = ~new_new_n11182__ & po020;
  assign new_new_n11684__ = ~pi068 & ~po020;
  assign new_new_n11685__ = ~new_new_n11683__ & ~new_new_n11684__;
  assign new_new_n11686__ = new_new_n11682__ & ~new_new_n11685__;
  assign new_new_n11687__ = ~new_new_n11682__ & new_new_n11685__;
  assign new_new_n11688__ = ~new_new_n11686__ & ~new_new_n11687__;
  assign new_new_n11689__ = ~new_new_n11681__ & ~new_new_n11688__;
  assign new_new_n11690__ = ~new_new_n11680__ & ~new_new_n11689__;
  assign new_new_n11691__ = ~new_new_n11613__ & ~new_new_n11690__;
  assign new_new_n11692__ = ~new_new_n11612__ & ~new_new_n11691__;
  assign new_new_n11693__ = ~new_new_n11604__ & new_new_n11692__;
  assign new_new_n11694__ = ~new_new_n11603__ & ~new_new_n11693__;
  assign new_new_n11695__ = ~new_new_n11597__ & ~new_new_n11694__;
  assign new_new_n11696__ = ~new_new_n11596__ & ~new_new_n11695__;
  assign new_new_n11697__ = ~new_new_n11588__ & ~new_new_n11696__;
  assign new_new_n11698__ = ~new_new_n11587__ & ~new_new_n11697__;
  assign new_new_n11699__ = ~new_new_n11579__ & ~new_new_n11698__;
  assign new_new_n11700__ = ~new_new_n11578__ & ~new_new_n11699__;
  assign new_new_n11701__ = ~new_new_n11570__ & ~new_new_n11700__;
  assign new_new_n11702__ = ~new_new_n11569__ & ~new_new_n11701__;
  assign new_new_n11703__ = ~new_new_n11561__ & ~new_new_n11702__;
  assign new_new_n11704__ = ~new_new_n11560__ & ~new_new_n11703__;
  assign new_new_n11705__ = ~new_new_n11552__ & new_new_n11704__;
  assign new_new_n11706__ = ~new_new_n11551__ & ~new_new_n11705__;
  assign new_new_n11707__ = ~new_new_n11543__ & ~new_new_n11706__;
  assign new_new_n11708__ = pi078 & ~new_new_n11542__;
  assign new_new_n11709__ = ~new_new_n11707__ & ~new_new_n11708__;
  assign new_new_n11710__ = ~new_new_n11535__ & ~new_new_n11709__;
  assign new_new_n11711__ = ~new_new_n11534__ & ~new_new_n11710__;
  assign new_new_n11712__ = ~new_new_n11526__ & new_new_n11711__;
  assign new_new_n11713__ = ~new_new_n11525__ & ~new_new_n11712__;
  assign new_new_n11714__ = ~new_new_n11517__ & new_new_n11713__;
  assign new_new_n11715__ = ~new_new_n11516__ & ~new_new_n11714__;
  assign new_new_n11716__ = ~new_new_n11508__ & new_new_n11715__;
  assign new_new_n11717__ = ~new_new_n11507__ & ~new_new_n11716__;
  assign new_new_n11718__ = ~new_new_n11499__ & ~new_new_n11717__;
  assign new_new_n11719__ = ~new_new_n11498__ & ~new_new_n11718__;
  assign new_new_n11720__ = ~new_new_n11490__ & ~new_new_n11719__;
  assign new_new_n11721__ = ~new_new_n11489__ & ~new_new_n11720__;
  assign new_new_n11722__ = ~new_new_n11481__ & ~new_new_n11721__;
  assign new_new_n11723__ = ~new_new_n11480__ & ~new_new_n11722__;
  assign new_new_n11724__ = ~new_new_n11472__ & ~new_new_n11723__;
  assign new_new_n11725__ = ~new_new_n11471__ & ~new_new_n11724__;
  assign new_new_n11726__ = ~new_new_n11463__ & new_new_n11725__;
  assign new_new_n11727__ = ~new_new_n11462__ & ~new_new_n11726__;
  assign new_new_n11728__ = ~new_new_n11454__ & ~new_new_n11727__;
  assign new_new_n11729__ = ~new_new_n11453__ & ~new_new_n11728__;
  assign new_new_n11730__ = ~new_new_n11445__ & ~new_new_n11729__;
  assign new_new_n11731__ = ~new_new_n11444__ & ~new_new_n11730__;
  assign new_new_n11732__ = ~new_new_n11436__ & new_new_n11731__;
  assign new_new_n11733__ = ~new_new_n11435__ & ~new_new_n11732__;
  assign new_new_n11734__ = ~new_new_n11427__ & ~new_new_n11733__;
  assign new_new_n11735__ = ~new_new_n11426__ & ~new_new_n11734__;
  assign new_new_n11736__ = ~new_new_n11418__ & ~new_new_n11735__;
  assign new_new_n11737__ = ~new_new_n11417__ & ~new_new_n11736__;
  assign new_new_n11738__ = ~new_new_n11409__ & new_new_n11737__;
  assign new_new_n11739__ = ~new_new_n11408__ & ~new_new_n11738__;
  assign new_new_n11740__ = ~new_new_n11400__ & ~new_new_n11739__;
  assign new_new_n11741__ = ~new_new_n11399__ & ~new_new_n11740__;
  assign new_new_n11742__ = ~new_new_n11391__ & new_new_n11741__;
  assign new_new_n11743__ = ~new_new_n11390__ & ~new_new_n11742__;
  assign new_new_n11744__ = ~new_new_n11382__ & ~new_new_n11743__;
  assign new_new_n11745__ = ~new_new_n11381__ & ~new_new_n11744__;
  assign new_new_n11746__ = ~new_new_n11373__ & ~new_new_n11745__;
  assign new_new_n11747__ = ~new_new_n11372__ & ~new_new_n11746__;
  assign new_new_n11748__ = ~new_new_n11364__ & ~new_new_n11747__;
  assign new_new_n11749__ = ~new_new_n11363__ & ~new_new_n11748__;
  assign new_new_n11750__ = ~new_new_n11355__ & new_new_n11749__;
  assign new_new_n11751__ = ~new_new_n11354__ & ~new_new_n11750__;
  assign new_new_n11752__ = ~new_new_n11346__ & ~new_new_n11751__;
  assign new_new_n11753__ = ~new_new_n11345__ & ~new_new_n11752__;
  assign new_new_n11754__ = ~new_new_n11337__ & ~new_new_n11753__;
  assign new_new_n11755__ = ~new_new_n11336__ & ~new_new_n11754__;
  assign new_new_n11756__ = ~new_new_n11328__ & ~new_new_n11755__;
  assign new_new_n11757__ = ~new_new_n11327__ & ~new_new_n11756__;
  assign new_new_n11758__ = ~new_new_n11319__ & new_new_n11757__;
  assign new_new_n11759__ = ~new_new_n11318__ & ~new_new_n11758__;
  assign new_new_n11760__ = ~new_new_n11312__ & new_new_n11759__;
  assign new_new_n11761__ = ~new_new_n11311__ & ~new_new_n11760__;
  assign new_new_n11762__ = ~new_new_n11303__ & ~new_new_n11761__;
  assign new_new_n11763__ = ~new_new_n11302__ & ~new_new_n11762__;
  assign new_new_n11764__ = ~new_new_n11294__ & ~new_new_n11763__;
  assign new_new_n11765__ = ~new_new_n11293__ & ~new_new_n11764__;
  assign new_new_n11766__ = ~pi107 & new_new_n11765__;
  assign new_new_n11767__ = pi107 & ~new_new_n11765__;
  assign new_new_n11768__ = ~pi106 & ~new_new_n11279__;
  assign new_new_n11769__ = pi106 & new_new_n11279__;
  assign new_new_n11770__ = ~new_new_n11768__ & ~new_new_n11769__;
  assign new_new_n11771__ = po020 & new_new_n11770__;
  assign new_new_n11772__ = new_new_n11275__ & new_new_n11771__;
  assign new_new_n11773__ = ~new_new_n11275__ & ~new_new_n11771__;
  assign new_new_n11774__ = ~new_new_n11772__ & ~new_new_n11773__;
  assign new_new_n11775__ = ~new_new_n11767__ & ~new_new_n11774__;
  assign new_new_n11776__ = ~new_new_n11766__ & ~new_new_n11775__;
  assign new_new_n11777__ = pi108 & new_new_n11776__;
  assign new_new_n11778__ = pi107 & ~new_new_n11281__;
  assign new_new_n11779__ = ~pi107 & new_new_n11281__;
  assign new_new_n11780__ = ~pi108 & ~new_new_n11778__;
  assign new_new_n11781__ = ~new_new_n11779__ & new_new_n11780__;
  assign new_new_n11782__ = ~new_new_n11776__ & new_new_n11781__;
  assign new_new_n11783__ = new_new_n10753__ & ~new_new_n11777__;
  assign new_new_n11784__ = ~new_new_n11782__ & new_new_n11783__;
  assign new_new_n11785__ = new_new_n10752__ & ~new_new_n11784__;
  assign new_new_n11786__ = pi108 & ~new_new_n9808__;
  assign new_new_n11787__ = ~new_new_n11776__ & ~new_new_n11786__;
  assign new_new_n11788__ = new_new_n10752__ & new_new_n11781__;
  assign new_new_n11789__ = ~new_new_n11787__ & ~new_new_n11788__;
  assign po019 = new_new_n10753__ & ~new_new_n11789__;
  assign new_new_n11791__ = ~new_new_n11766__ & ~new_new_n11767__;
  assign new_new_n11792__ = po019 & new_new_n11791__;
  assign new_new_n11793__ = ~new_new_n11774__ & ~new_new_n11792__;
  assign new_new_n11794__ = new_new_n11774__ & new_new_n11792__;
  assign new_new_n11795__ = ~new_new_n11793__ & ~new_new_n11794__;
  assign new_new_n11796__ = ~pi108 & ~new_new_n11795__;
  assign new_new_n11797__ = pi108 & new_new_n11795__;
  assign new_new_n11798__ = pi106 & ~new_new_n11763__;
  assign new_new_n11799__ = ~pi106 & new_new_n11763__;
  assign new_new_n11800__ = ~new_new_n11798__ & ~new_new_n11799__;
  assign new_new_n11801__ = po019 & new_new_n11800__;
  assign new_new_n11802__ = new_new_n11292__ & new_new_n11801__;
  assign new_new_n11803__ = ~new_new_n11292__ & ~new_new_n11801__;
  assign new_new_n11804__ = ~new_new_n11802__ & ~new_new_n11803__;
  assign new_new_n11805__ = pi107 & ~new_new_n11804__;
  assign new_new_n11806__ = ~pi107 & new_new_n11804__;
  assign new_new_n11807__ = ~new_new_n11761__ & po019;
  assign new_new_n11808__ = pi105 & ~po019;
  assign new_new_n11809__ = ~new_new_n11807__ & ~new_new_n11808__;
  assign new_new_n11810__ = ~new_new_n11302__ & ~new_new_n11303__;
  assign new_new_n11811__ = ~new_new_n11809__ & new_new_n11810__;
  assign new_new_n11812__ = new_new_n11809__ & ~new_new_n11810__;
  assign new_new_n11813__ = ~new_new_n11811__ & ~new_new_n11812__;
  assign new_new_n11814__ = ~pi106 & ~new_new_n11813__;
  assign new_new_n11815__ = pi106 & new_new_n11813__;
  assign new_new_n11816__ = ~new_new_n11311__ & ~new_new_n11312__;
  assign new_new_n11817__ = ~new_new_n11759__ & po019;
  assign new_new_n11818__ = ~pi104 & ~po019;
  assign new_new_n11819__ = ~new_new_n11817__ & ~new_new_n11818__;
  assign new_new_n11820__ = new_new_n11816__ & ~new_new_n11819__;
  assign new_new_n11821__ = ~new_new_n11816__ & new_new_n11819__;
  assign new_new_n11822__ = ~new_new_n11820__ & ~new_new_n11821__;
  assign new_new_n11823__ = pi105 & ~new_new_n11822__;
  assign new_new_n11824__ = ~pi105 & new_new_n11822__;
  assign new_new_n11825__ = ~new_new_n11757__ & po019;
  assign new_new_n11826__ = pi103 & ~po019;
  assign new_new_n11827__ = ~new_new_n11825__ & ~new_new_n11826__;
  assign new_new_n11828__ = ~new_new_n11318__ & ~new_new_n11319__;
  assign new_new_n11829__ = ~new_new_n11827__ & new_new_n11828__;
  assign new_new_n11830__ = new_new_n11827__ & ~new_new_n11828__;
  assign new_new_n11831__ = ~new_new_n11829__ & ~new_new_n11830__;
  assign new_new_n11832__ = pi104 & new_new_n11831__;
  assign new_new_n11833__ = ~pi104 & ~new_new_n11831__;
  assign new_new_n11834__ = pi102 & ~new_new_n11755__;
  assign new_new_n11835__ = ~pi102 & new_new_n11755__;
  assign new_new_n11836__ = ~new_new_n11834__ & ~new_new_n11835__;
  assign new_new_n11837__ = po019 & new_new_n11836__;
  assign new_new_n11838__ = ~new_new_n11326__ & new_new_n11837__;
  assign new_new_n11839__ = new_new_n11326__ & ~new_new_n11837__;
  assign new_new_n11840__ = ~new_new_n11838__ & ~new_new_n11839__;
  assign new_new_n11841__ = pi103 & new_new_n11840__;
  assign new_new_n11842__ = ~pi103 & ~new_new_n11840__;
  assign new_new_n11843__ = pi101 & ~new_new_n11753__;
  assign new_new_n11844__ = ~pi101 & new_new_n11753__;
  assign new_new_n11845__ = ~new_new_n11843__ & ~new_new_n11844__;
  assign new_new_n11846__ = po019 & new_new_n11845__;
  assign new_new_n11847__ = ~new_new_n11335__ & ~new_new_n11846__;
  assign new_new_n11848__ = new_new_n11335__ & new_new_n11846__;
  assign new_new_n11849__ = ~new_new_n11847__ & ~new_new_n11848__;
  assign new_new_n11850__ = pi102 & ~new_new_n11849__;
  assign new_new_n11851__ = ~pi102 & new_new_n11849__;
  assign new_new_n11852__ = ~new_new_n11345__ & ~new_new_n11346__;
  assign new_new_n11853__ = ~new_new_n11751__ & po019;
  assign new_new_n11854__ = pi100 & ~po019;
  assign new_new_n11855__ = ~new_new_n11853__ & ~new_new_n11854__;
  assign new_new_n11856__ = new_new_n11852__ & new_new_n11855__;
  assign new_new_n11857__ = ~new_new_n11852__ & ~new_new_n11855__;
  assign new_new_n11858__ = ~new_new_n11856__ & ~new_new_n11857__;
  assign new_new_n11859__ = pi101 & ~new_new_n11858__;
  assign new_new_n11860__ = ~pi101 & new_new_n11858__;
  assign new_new_n11861__ = new_new_n11749__ & po019;
  assign new_new_n11862__ = pi099 & ~po019;
  assign new_new_n11863__ = ~new_new_n11861__ & ~new_new_n11862__;
  assign new_new_n11864__ = ~new_new_n11354__ & ~new_new_n11355__;
  assign new_new_n11865__ = ~new_new_n11863__ & ~new_new_n11864__;
  assign new_new_n11866__ = new_new_n11863__ & new_new_n11864__;
  assign new_new_n11867__ = ~new_new_n11865__ & ~new_new_n11866__;
  assign new_new_n11868__ = pi100 & ~new_new_n11867__;
  assign new_new_n11869__ = ~pi100 & new_new_n11867__;
  assign new_new_n11870__ = ~new_new_n11363__ & ~new_new_n11364__;
  assign new_new_n11871__ = ~new_new_n11747__ & po019;
  assign new_new_n11872__ = ~pi098 & ~po019;
  assign new_new_n11873__ = ~new_new_n11871__ & ~new_new_n11872__;
  assign new_new_n11874__ = new_new_n11870__ & ~new_new_n11873__;
  assign new_new_n11875__ = ~new_new_n11870__ & new_new_n11873__;
  assign new_new_n11876__ = ~new_new_n11874__ & ~new_new_n11875__;
  assign new_new_n11877__ = pi099 & ~new_new_n11876__;
  assign new_new_n11878__ = ~pi099 & new_new_n11876__;
  assign new_new_n11879__ = ~new_new_n11372__ & ~new_new_n11373__;
  assign new_new_n11880__ = ~new_new_n11745__ & po019;
  assign new_new_n11881__ = ~pi097 & ~po019;
  assign new_new_n11882__ = ~new_new_n11880__ & ~new_new_n11881__;
  assign new_new_n11883__ = new_new_n11879__ & ~new_new_n11882__;
  assign new_new_n11884__ = ~new_new_n11879__ & new_new_n11882__;
  assign new_new_n11885__ = ~new_new_n11883__ & ~new_new_n11884__;
  assign new_new_n11886__ = pi098 & ~new_new_n11885__;
  assign new_new_n11887__ = ~pi098 & new_new_n11885__;
  assign new_new_n11888__ = ~pi096 & ~new_new_n11743__;
  assign new_new_n11889__ = pi096 & new_new_n11743__;
  assign new_new_n11890__ = ~new_new_n11888__ & ~new_new_n11889__;
  assign new_new_n11891__ = po019 & new_new_n11890__;
  assign new_new_n11892__ = new_new_n11380__ & new_new_n11891__;
  assign new_new_n11893__ = ~new_new_n11380__ & ~new_new_n11891__;
  assign new_new_n11894__ = ~new_new_n11892__ & ~new_new_n11893__;
  assign new_new_n11895__ = ~pi097 & ~new_new_n11894__;
  assign new_new_n11896__ = pi097 & new_new_n11894__;
  assign new_new_n11897__ = ~new_new_n11741__ & po019;
  assign new_new_n11898__ = pi095 & ~po019;
  assign new_new_n11899__ = ~new_new_n11897__ & ~new_new_n11898__;
  assign new_new_n11900__ = ~new_new_n11390__ & ~new_new_n11391__;
  assign new_new_n11901__ = ~new_new_n11899__ & new_new_n11900__;
  assign new_new_n11902__ = new_new_n11899__ & ~new_new_n11900__;
  assign new_new_n11903__ = ~new_new_n11901__ & ~new_new_n11902__;
  assign new_new_n11904__ = ~pi096 & ~new_new_n11903__;
  assign new_new_n11905__ = pi096 & new_new_n11903__;
  assign new_new_n11906__ = ~new_new_n11739__ & po019;
  assign new_new_n11907__ = pi094 & ~po019;
  assign new_new_n11908__ = ~new_new_n11906__ & ~new_new_n11907__;
  assign new_new_n11909__ = ~new_new_n11399__ & ~new_new_n11400__;
  assign new_new_n11910__ = ~new_new_n11908__ & new_new_n11909__;
  assign new_new_n11911__ = new_new_n11908__ & ~new_new_n11909__;
  assign new_new_n11912__ = ~new_new_n11910__ & ~new_new_n11911__;
  assign new_new_n11913__ = pi095 & new_new_n11912__;
  assign new_new_n11914__ = ~pi095 & ~new_new_n11912__;
  assign new_new_n11915__ = ~new_new_n11408__ & ~new_new_n11409__;
  assign new_new_n11916__ = ~new_new_n11737__ & po019;
  assign new_new_n11917__ = ~pi093 & ~po019;
  assign new_new_n11918__ = ~new_new_n11916__ & ~new_new_n11917__;
  assign new_new_n11919__ = new_new_n11915__ & ~new_new_n11918__;
  assign new_new_n11920__ = ~new_new_n11915__ & new_new_n11918__;
  assign new_new_n11921__ = ~new_new_n11919__ & ~new_new_n11920__;
  assign new_new_n11922__ = pi094 & ~new_new_n11921__;
  assign new_new_n11923__ = ~pi094 & new_new_n11921__;
  assign new_new_n11924__ = ~new_new_n11417__ & ~new_new_n11418__;
  assign new_new_n11925__ = ~new_new_n11735__ & po019;
  assign new_new_n11926__ = ~pi092 & ~po019;
  assign new_new_n11927__ = ~new_new_n11925__ & ~new_new_n11926__;
  assign new_new_n11928__ = new_new_n11924__ & ~new_new_n11927__;
  assign new_new_n11929__ = ~new_new_n11924__ & new_new_n11927__;
  assign new_new_n11930__ = ~new_new_n11928__ & ~new_new_n11929__;
  assign new_new_n11931__ = pi093 & ~new_new_n11930__;
  assign new_new_n11932__ = ~pi093 & new_new_n11930__;
  assign new_new_n11933__ = ~pi091 & ~new_new_n11733__;
  assign new_new_n11934__ = pi091 & new_new_n11733__;
  assign new_new_n11935__ = ~new_new_n11933__ & ~new_new_n11934__;
  assign new_new_n11936__ = po019 & new_new_n11935__;
  assign new_new_n11937__ = ~new_new_n11425__ & ~new_new_n11936__;
  assign new_new_n11938__ = new_new_n11425__ & new_new_n11936__;
  assign new_new_n11939__ = ~new_new_n11937__ & ~new_new_n11938__;
  assign new_new_n11940__ = pi092 & new_new_n11939__;
  assign new_new_n11941__ = ~pi092 & ~new_new_n11939__;
  assign new_new_n11942__ = ~new_new_n11731__ & po019;
  assign new_new_n11943__ = pi090 & ~po019;
  assign new_new_n11944__ = ~new_new_n11942__ & ~new_new_n11943__;
  assign new_new_n11945__ = ~new_new_n11435__ & ~new_new_n11436__;
  assign new_new_n11946__ = ~new_new_n11944__ & new_new_n11945__;
  assign new_new_n11947__ = new_new_n11944__ & ~new_new_n11945__;
  assign new_new_n11948__ = ~new_new_n11946__ & ~new_new_n11947__;
  assign new_new_n11949__ = pi091 & new_new_n11948__;
  assign new_new_n11950__ = ~pi091 & ~new_new_n11948__;
  assign new_new_n11951__ = pi089 & ~new_new_n11729__;
  assign new_new_n11952__ = ~pi089 & new_new_n11729__;
  assign new_new_n11953__ = ~new_new_n11951__ & ~new_new_n11952__;
  assign new_new_n11954__ = po019 & new_new_n11953__;
  assign new_new_n11955__ = ~new_new_n11443__ & ~new_new_n11954__;
  assign new_new_n11956__ = new_new_n11443__ & new_new_n11954__;
  assign new_new_n11957__ = ~new_new_n11955__ & ~new_new_n11956__;
  assign new_new_n11958__ = pi090 & ~new_new_n11957__;
  assign new_new_n11959__ = ~pi090 & new_new_n11957__;
  assign new_new_n11960__ = ~new_new_n11453__ & ~new_new_n11454__;
  assign new_new_n11961__ = ~new_new_n11727__ & po019;
  assign new_new_n11962__ = pi088 & ~po019;
  assign new_new_n11963__ = ~new_new_n11961__ & ~new_new_n11962__;
  assign new_new_n11964__ = new_new_n11960__ & ~new_new_n11963__;
  assign new_new_n11965__ = ~new_new_n11960__ & new_new_n11963__;
  assign new_new_n11966__ = ~new_new_n11964__ & ~new_new_n11965__;
  assign new_new_n11967__ = pi089 & new_new_n11966__;
  assign new_new_n11968__ = ~pi089 & ~new_new_n11966__;
  assign new_new_n11969__ = ~new_new_n11462__ & ~new_new_n11463__;
  assign new_new_n11970__ = ~new_new_n11725__ & po019;
  assign new_new_n11971__ = ~pi087 & ~po019;
  assign new_new_n11972__ = ~new_new_n11970__ & ~new_new_n11971__;
  assign new_new_n11973__ = new_new_n11969__ & ~new_new_n11972__;
  assign new_new_n11974__ = ~new_new_n11969__ & new_new_n11972__;
  assign new_new_n11975__ = ~new_new_n11973__ & ~new_new_n11974__;
  assign new_new_n11976__ = pi088 & ~new_new_n11975__;
  assign new_new_n11977__ = ~pi088 & new_new_n11975__;
  assign new_new_n11978__ = ~new_new_n11471__ & ~new_new_n11472__;
  assign new_new_n11979__ = ~new_new_n11723__ & po019;
  assign new_new_n11980__ = ~pi086 & ~po019;
  assign new_new_n11981__ = ~new_new_n11979__ & ~new_new_n11980__;
  assign new_new_n11982__ = new_new_n11978__ & ~new_new_n11981__;
  assign new_new_n11983__ = ~new_new_n11978__ & new_new_n11981__;
  assign new_new_n11984__ = ~new_new_n11982__ & ~new_new_n11983__;
  assign new_new_n11985__ = ~pi087 & new_new_n11984__;
  assign new_new_n11986__ = pi087 & ~new_new_n11984__;
  assign new_new_n11987__ = ~pi085 & ~new_new_n11721__;
  assign new_new_n11988__ = pi085 & new_new_n11721__;
  assign new_new_n11989__ = ~new_new_n11987__ & ~new_new_n11988__;
  assign new_new_n11990__ = po019 & new_new_n11989__;
  assign new_new_n11991__ = new_new_n11479__ & new_new_n11990__;
  assign new_new_n11992__ = ~new_new_n11479__ & ~new_new_n11990__;
  assign new_new_n11993__ = ~new_new_n11991__ & ~new_new_n11992__;
  assign new_new_n11994__ = ~pi086 & ~new_new_n11993__;
  assign new_new_n11995__ = pi086 & new_new_n11993__;
  assign new_new_n11996__ = ~new_new_n11489__ & ~new_new_n11490__;
  assign new_new_n11997__ = ~new_new_n11719__ & po019;
  assign new_new_n11998__ = ~pi084 & ~po019;
  assign new_new_n11999__ = ~new_new_n11997__ & ~new_new_n11998__;
  assign new_new_n12000__ = new_new_n11996__ & ~new_new_n11999__;
  assign new_new_n12001__ = ~new_new_n11996__ & new_new_n11999__;
  assign new_new_n12002__ = ~new_new_n12000__ & ~new_new_n12001__;
  assign new_new_n12003__ = pi085 & ~new_new_n12002__;
  assign new_new_n12004__ = ~pi085 & new_new_n12002__;
  assign new_new_n12005__ = ~new_new_n11498__ & ~new_new_n11499__;
  assign new_new_n12006__ = ~new_new_n11717__ & po019;
  assign new_new_n12007__ = ~pi083 & ~po019;
  assign new_new_n12008__ = ~new_new_n12006__ & ~new_new_n12007__;
  assign new_new_n12009__ = new_new_n12005__ & ~new_new_n12008__;
  assign new_new_n12010__ = ~new_new_n12005__ & new_new_n12008__;
  assign new_new_n12011__ = ~new_new_n12009__ & ~new_new_n12010__;
  assign new_new_n12012__ = pi084 & ~new_new_n12011__;
  assign new_new_n12013__ = ~pi084 & new_new_n12011__;
  assign new_new_n12014__ = ~new_new_n11507__ & ~new_new_n11508__;
  assign new_new_n12015__ = ~new_new_n11715__ & po019;
  assign new_new_n12016__ = pi082 & ~po019;
  assign new_new_n12017__ = ~new_new_n12015__ & ~new_new_n12016__;
  assign new_new_n12018__ = new_new_n12014__ & ~new_new_n12017__;
  assign new_new_n12019__ = ~new_new_n12014__ & new_new_n12017__;
  assign new_new_n12020__ = ~new_new_n12018__ & ~new_new_n12019__;
  assign new_new_n12021__ = ~pi083 & ~new_new_n12020__;
  assign new_new_n12022__ = pi083 & new_new_n12020__;
  assign new_new_n12023__ = ~new_new_n11516__ & ~new_new_n11517__;
  assign new_new_n12024__ = ~new_new_n11713__ & po019;
  assign new_new_n12025__ = ~pi081 & ~po019;
  assign new_new_n12026__ = ~new_new_n12024__ & ~new_new_n12025__;
  assign new_new_n12027__ = new_new_n12023__ & ~new_new_n12026__;
  assign new_new_n12028__ = ~new_new_n12023__ & new_new_n12026__;
  assign new_new_n12029__ = ~new_new_n12027__ & ~new_new_n12028__;
  assign new_new_n12030__ = ~pi082 & new_new_n12029__;
  assign new_new_n12031__ = pi082 & ~new_new_n12029__;
  assign new_new_n12032__ = ~new_new_n11525__ & ~new_new_n11526__;
  assign new_new_n12033__ = new_new_n11711__ & po019;
  assign new_new_n12034__ = ~pi080 & ~po019;
  assign new_new_n12035__ = ~new_new_n12033__ & ~new_new_n12034__;
  assign new_new_n12036__ = ~new_new_n12032__ & ~new_new_n12035__;
  assign new_new_n12037__ = new_new_n12032__ & new_new_n12035__;
  assign new_new_n12038__ = ~new_new_n12036__ & ~new_new_n12037__;
  assign new_new_n12039__ = ~pi081 & ~new_new_n12038__;
  assign new_new_n12040__ = pi081 & new_new_n12038__;
  assign new_new_n12041__ = new_new_n11709__ & po019;
  assign new_new_n12042__ = ~pi079 & ~po019;
  assign new_new_n12043__ = ~new_new_n12041__ & ~new_new_n12042__;
  assign new_new_n12044__ = ~new_new_n11534__ & ~new_new_n11535__;
  assign new_new_n12045__ = ~new_new_n12043__ & ~new_new_n12044__;
  assign new_new_n12046__ = new_new_n12043__ & new_new_n12044__;
  assign new_new_n12047__ = ~new_new_n12045__ & ~new_new_n12046__;
  assign new_new_n12048__ = ~pi080 & ~new_new_n12047__;
  assign new_new_n12049__ = pi080 & new_new_n12047__;
  assign new_new_n12050__ = ~new_new_n11543__ & ~new_new_n11708__;
  assign new_new_n12051__ = ~new_new_n11706__ & po019;
  assign new_new_n12052__ = pi078 & ~po019;
  assign new_new_n12053__ = ~new_new_n12051__ & ~new_new_n12052__;
  assign new_new_n12054__ = new_new_n12050__ & new_new_n12053__;
  assign new_new_n12055__ = ~new_new_n12050__ & ~new_new_n12053__;
  assign new_new_n12056__ = ~new_new_n12054__ & ~new_new_n12055__;
  assign new_new_n12057__ = pi079 & ~new_new_n12056__;
  assign new_new_n12058__ = ~pi079 & new_new_n12056__;
  assign new_new_n12059__ = new_new_n11704__ & po019;
  assign new_new_n12060__ = pi077 & ~po019;
  assign new_new_n12061__ = ~new_new_n12059__ & ~new_new_n12060__;
  assign new_new_n12062__ = ~new_new_n11551__ & ~new_new_n11552__;
  assign new_new_n12063__ = ~new_new_n12061__ & ~new_new_n12062__;
  assign new_new_n12064__ = new_new_n12061__ & new_new_n12062__;
  assign new_new_n12065__ = ~new_new_n12063__ & ~new_new_n12064__;
  assign new_new_n12066__ = pi078 & ~new_new_n12065__;
  assign new_new_n12067__ = ~pi078 & new_new_n12065__;
  assign new_new_n12068__ = ~new_new_n11560__ & ~new_new_n11561__;
  assign new_new_n12069__ = ~new_new_n11702__ & po019;
  assign new_new_n12070__ = ~pi076 & ~po019;
  assign new_new_n12071__ = ~new_new_n12069__ & ~new_new_n12070__;
  assign new_new_n12072__ = new_new_n12068__ & ~new_new_n12071__;
  assign new_new_n12073__ = ~new_new_n12068__ & new_new_n12071__;
  assign new_new_n12074__ = ~new_new_n12072__ & ~new_new_n12073__;
  assign new_new_n12075__ = pi077 & ~new_new_n12074__;
  assign new_new_n12076__ = ~pi077 & new_new_n12074__;
  assign new_new_n12077__ = ~new_new_n11569__ & ~new_new_n11570__;
  assign new_new_n12078__ = ~new_new_n11700__ & po019;
  assign new_new_n12079__ = ~pi075 & ~po019;
  assign new_new_n12080__ = ~new_new_n12078__ & ~new_new_n12079__;
  assign new_new_n12081__ = new_new_n12077__ & ~new_new_n12080__;
  assign new_new_n12082__ = ~new_new_n12077__ & new_new_n12080__;
  assign new_new_n12083__ = ~new_new_n12081__ & ~new_new_n12082__;
  assign new_new_n12084__ = pi076 & ~new_new_n12083__;
  assign new_new_n12085__ = ~pi076 & new_new_n12083__;
  assign new_new_n12086__ = ~new_new_n11578__ & ~new_new_n11579__;
  assign new_new_n12087__ = ~new_new_n11698__ & po019;
  assign new_new_n12088__ = ~pi074 & ~po019;
  assign new_new_n12089__ = ~new_new_n12087__ & ~new_new_n12088__;
  assign new_new_n12090__ = new_new_n12086__ & ~new_new_n12089__;
  assign new_new_n12091__ = ~new_new_n12086__ & new_new_n12089__;
  assign new_new_n12092__ = ~new_new_n12090__ & ~new_new_n12091__;
  assign new_new_n12093__ = pi075 & ~new_new_n12092__;
  assign new_new_n12094__ = ~pi075 & new_new_n12092__;
  assign new_new_n12095__ = ~pi073 & ~new_new_n11696__;
  assign new_new_n12096__ = pi073 & new_new_n11696__;
  assign new_new_n12097__ = ~new_new_n12095__ & ~new_new_n12096__;
  assign new_new_n12098__ = po019 & new_new_n12097__;
  assign new_new_n12099__ = new_new_n11586__ & new_new_n12098__;
  assign new_new_n12100__ = ~new_new_n11586__ & ~new_new_n12098__;
  assign new_new_n12101__ = ~new_new_n12099__ & ~new_new_n12100__;
  assign new_new_n12102__ = ~pi074 & ~new_new_n12101__;
  assign new_new_n12103__ = pi074 & new_new_n12101__;
  assign new_new_n12104__ = ~new_new_n11596__ & ~new_new_n11597__;
  assign new_new_n12105__ = ~new_new_n11694__ & po019;
  assign new_new_n12106__ = ~pi072 & ~po019;
  assign new_new_n12107__ = ~new_new_n12105__ & ~new_new_n12106__;
  assign new_new_n12108__ = ~new_new_n12104__ & ~new_new_n12107__;
  assign new_new_n12109__ = new_new_n12104__ & new_new_n12107__;
  assign new_new_n12110__ = ~new_new_n12108__ & ~new_new_n12109__;
  assign new_new_n12111__ = ~pi073 & ~new_new_n12110__;
  assign new_new_n12112__ = pi073 & new_new_n12110__;
  assign new_new_n12113__ = new_new_n11692__ & po019;
  assign new_new_n12114__ = ~pi071 & ~po019;
  assign new_new_n12115__ = ~new_new_n12113__ & ~new_new_n12114__;
  assign new_new_n12116__ = ~new_new_n11603__ & ~new_new_n11604__;
  assign new_new_n12117__ = ~new_new_n12115__ & ~new_new_n12116__;
  assign new_new_n12118__ = new_new_n12115__ & new_new_n12116__;
  assign new_new_n12119__ = ~new_new_n12117__ & ~new_new_n12118__;
  assign new_new_n12120__ = ~pi072 & ~new_new_n12119__;
  assign new_new_n12121__ = pi072 & new_new_n12119__;
  assign new_new_n12122__ = ~new_new_n11612__ & ~new_new_n11613__;
  assign new_new_n12123__ = ~new_new_n11690__ & po019;
  assign new_new_n12124__ = pi070 & ~po019;
  assign new_new_n12125__ = ~new_new_n12123__ & ~new_new_n12124__;
  assign new_new_n12126__ = new_new_n12122__ & new_new_n12125__;
  assign new_new_n12127__ = ~new_new_n12122__ & ~new_new_n12125__;
  assign new_new_n12128__ = ~new_new_n12126__ & ~new_new_n12127__;
  assign new_new_n12129__ = pi071 & ~new_new_n12128__;
  assign new_new_n12130__ = ~pi071 & new_new_n12128__;
  assign new_new_n12131__ = ~new_new_n11680__ & ~new_new_n11681__;
  assign new_new_n12132__ = po019 & new_new_n12131__;
  assign new_new_n12133__ = new_new_n11688__ & new_new_n12132__;
  assign new_new_n12134__ = ~new_new_n11688__ & ~new_new_n12132__;
  assign new_new_n12135__ = ~new_new_n12133__ & ~new_new_n12134__;
  assign new_new_n12136__ = pi070 & ~new_new_n12135__;
  assign new_new_n12137__ = ~pi070 & new_new_n12135__;
  assign new_new_n12138__ = ~new_new_n11669__ & ~new_new_n11678__;
  assign new_new_n12139__ = po019 & new_new_n12138__;
  assign new_new_n12140__ = ~new_new_n11676__ & ~new_new_n12139__;
  assign new_new_n12141__ = new_new_n11676__ & new_new_n12139__;
  assign new_new_n12142__ = ~new_new_n12140__ & ~new_new_n12141__;
  assign new_new_n12143__ = pi069 & ~new_new_n12142__;
  assign new_new_n12144__ = ~pi069 & new_new_n12142__;
  assign new_new_n12145__ = new_new_n426__ & ~po021;
  assign new_new_n12146__ = ~pi065 & po020;
  assign new_new_n12147__ = po021 & new_new_n12146__;
  assign new_new_n12148__ = ~new_new_n12145__ & ~new_new_n12147__;
  assign new_new_n12149__ = ~pi020 & ~new_new_n12148__;
  assign new_new_n12150__ = new_new_n11157__ & new_new_n11647__;
  assign new_new_n12151__ = ~new_new_n11165__ & ~new_new_n12150__;
  assign new_new_n12152__ = pi020 & ~new_new_n12151__;
  assign new_new_n12153__ = ~new_new_n332__ & po020;
  assign new_new_n12154__ = ~new_new_n11157__ & ~new_new_n12153__;
  assign new_new_n12155__ = ~new_new_n12149__ & ~new_new_n12154__;
  assign new_new_n12156__ = ~new_new_n12152__ & new_new_n12155__;
  assign new_new_n12157__ = ~pi021 & ~new_new_n12156__;
  assign new_new_n12158__ = ~new_new_n11157__ & ~new_new_n11647__;
  assign new_new_n12159__ = pi020 & ~new_new_n11171__;
  assign new_new_n12160__ = pi064 & ~new_new_n12159__;
  assign new_new_n12161__ = ~new_new_n12158__ & ~new_new_n12160__;
  assign new_new_n12162__ = ~po021 & ~new_new_n12146__;
  assign new_new_n12163__ = pi064 & ~new_new_n11621__;
  assign new_new_n12164__ = ~new_new_n12147__ & new_new_n12163__;
  assign new_new_n12165__ = ~new_new_n12162__ & new_new_n12164__;
  assign new_new_n12166__ = ~new_new_n12161__ & ~new_new_n12165__;
  assign new_new_n12167__ = pi021 & ~new_new_n12166__;
  assign new_new_n12168__ = ~new_new_n12157__ & ~new_new_n12167__;
  assign new_new_n12169__ = pi019 & ~new_new_n11621__;
  assign new_new_n12170__ = pi065 & ~new_new_n12169__;
  assign new_new_n12171__ = ~pi020 & po020;
  assign new_new_n12172__ = ~pi019 & ~new_new_n11652__;
  assign new_new_n12173__ = ~new_new_n12171__ & new_new_n12172__;
  assign new_new_n12174__ = ~new_new_n12170__ & ~new_new_n12173__;
  assign new_new_n12175__ = pi064 & ~new_new_n12174__;
  assign new_new_n12176__ = ~new_new_n11641__ & ~new_new_n12175__;
  assign new_new_n12177__ = pi066 & ~new_new_n12176__;
  assign new_new_n12178__ = ~pi066 & new_new_n12176__;
  assign new_new_n12179__ = ~new_new_n12177__ & ~new_new_n12178__;
  assign new_new_n12180__ = po019 & new_new_n12179__;
  assign new_new_n12181__ = ~new_new_n12168__ & new_new_n12180__;
  assign new_new_n12182__ = new_new_n12168__ & ~new_new_n12180__;
  assign new_new_n12183__ = ~new_new_n12181__ & ~new_new_n12182__;
  assign new_new_n12184__ = ~pi067 & ~new_new_n12183__;
  assign new_new_n12185__ = pi067 & new_new_n12183__;
  assign new_new_n12186__ = pi019 & po019;
  assign new_new_n12187__ = pi018 & ~pi065;
  assign new_new_n12188__ = new_new_n12186__ & ~new_new_n12187__;
  assign new_new_n12189__ = ~pi019 & ~po019;
  assign new_new_n12190__ = ~pi065 & ~new_new_n12189__;
  assign new_new_n12191__ = ~pi018 & ~new_new_n12190__;
  assign new_new_n12192__ = ~new_new_n12188__ & ~new_new_n12191__;
  assign new_new_n12193__ = pi064 & ~new_new_n12192__;
  assign new_new_n12194__ = pi064 & po019;
  assign new_new_n12195__ = ~pi019 & pi065;
  assign new_new_n12196__ = ~new_new_n12194__ & new_new_n12195__;
  assign new_new_n12197__ = ~new_new_n12193__ & ~new_new_n12196__;
  assign new_new_n12198__ = pi066 & ~new_new_n12197__;
  assign new_new_n12199__ = pi065 & po019;
  assign new_new_n12200__ = new_new_n11640__ & new_new_n12199__;
  assign new_new_n12201__ = ~new_new_n11649__ & ~new_new_n12200__;
  assign new_new_n12202__ = pi019 & ~new_new_n12201__;
  assign new_new_n12203__ = po019 & new_new_n12146__;
  assign new_new_n12204__ = new_new_n426__ & ~po020;
  assign new_new_n12205__ = ~new_new_n12203__ & ~new_new_n12204__;
  assign new_new_n12206__ = ~pi019 & ~new_new_n12205__;
  assign new_new_n12207__ = ~new_new_n332__ & po019;
  assign new_new_n12208__ = ~new_new_n11640__ & ~new_new_n12207__;
  assign new_new_n12209__ = ~new_new_n12206__ & ~new_new_n12208__;
  assign new_new_n12210__ = ~new_new_n12202__ & new_new_n12209__;
  assign new_new_n12211__ = ~pi020 & ~new_new_n12210__;
  assign new_new_n12212__ = ~new_new_n11640__ & ~new_new_n12199__;
  assign new_new_n12213__ = pi064 & ~new_new_n11648__;
  assign new_new_n12214__ = ~new_new_n12212__ & ~new_new_n12213__;
  assign new_new_n12215__ = ~pi065 & po019;
  assign new_new_n12216__ = ~po020 & ~new_new_n12215__;
  assign new_new_n12217__ = pi064 & ~new_new_n12186__;
  assign new_new_n12218__ = ~new_new_n12203__ & new_new_n12217__;
  assign new_new_n12219__ = ~new_new_n12216__ & new_new_n12218__;
  assign new_new_n12220__ = ~new_new_n12214__ & ~new_new_n12219__;
  assign new_new_n12221__ = pi020 & ~new_new_n12220__;
  assign new_new_n12222__ = ~new_new_n12211__ & ~new_new_n12221__;
  assign new_new_n12223__ = ~pi066 & new_new_n12197__;
  assign new_new_n12224__ = ~new_new_n12222__ & ~new_new_n12223__;
  assign new_new_n12225__ = ~new_new_n12198__ & ~new_new_n12224__;
  assign new_new_n12226__ = ~new_new_n12185__ & new_new_n12225__;
  assign new_new_n12227__ = ~new_new_n12184__ & ~new_new_n12226__;
  assign new_new_n12228__ = ~pi068 & ~new_new_n12227__;
  assign new_new_n12229__ = pi068 & new_new_n12227__;
  assign new_new_n12230__ = ~pi067 & ~new_new_n11666__;
  assign new_new_n12231__ = pi067 & new_new_n11666__;
  assign new_new_n12232__ = ~new_new_n12230__ & ~new_new_n12231__;
  assign new_new_n12233__ = po019 & new_new_n12232__;
  assign new_new_n12234__ = new_new_n11618__ & new_new_n12233__;
  assign new_new_n12235__ = ~new_new_n11618__ & ~new_new_n12233__;
  assign new_new_n12236__ = ~new_new_n12234__ & ~new_new_n12235__;
  assign new_new_n12237__ = ~new_new_n12229__ & ~new_new_n12236__;
  assign new_new_n12238__ = ~new_new_n12228__ & ~new_new_n12237__;
  assign new_new_n12239__ = ~new_new_n12144__ & new_new_n12238__;
  assign new_new_n12240__ = ~new_new_n12143__ & ~new_new_n12239__;
  assign new_new_n12241__ = ~new_new_n12137__ & ~new_new_n12240__;
  assign new_new_n12242__ = ~new_new_n12136__ & ~new_new_n12241__;
  assign new_new_n12243__ = ~new_new_n12130__ & ~new_new_n12242__;
  assign new_new_n12244__ = ~new_new_n12129__ & ~new_new_n12243__;
  assign new_new_n12245__ = ~new_new_n12121__ & new_new_n12244__;
  assign new_new_n12246__ = ~new_new_n12120__ & ~new_new_n12245__;
  assign new_new_n12247__ = ~new_new_n12112__ & ~new_new_n12246__;
  assign new_new_n12248__ = ~new_new_n12111__ & ~new_new_n12247__;
  assign new_new_n12249__ = ~new_new_n12103__ & ~new_new_n12248__;
  assign new_new_n12250__ = ~new_new_n12102__ & ~new_new_n12249__;
  assign new_new_n12251__ = ~new_new_n12094__ & new_new_n12250__;
  assign new_new_n12252__ = ~new_new_n12093__ & ~new_new_n12251__;
  assign new_new_n12253__ = ~new_new_n12085__ & ~new_new_n12252__;
  assign new_new_n12254__ = ~new_new_n12084__ & ~new_new_n12253__;
  assign new_new_n12255__ = ~new_new_n12076__ & ~new_new_n12254__;
  assign new_new_n12256__ = ~new_new_n12075__ & ~new_new_n12255__;
  assign new_new_n12257__ = ~new_new_n12067__ & ~new_new_n12256__;
  assign new_new_n12258__ = ~new_new_n12066__ & ~new_new_n12257__;
  assign new_new_n12259__ = ~new_new_n12058__ & ~new_new_n12258__;
  assign new_new_n12260__ = ~new_new_n12057__ & ~new_new_n12259__;
  assign new_new_n12261__ = ~new_new_n12049__ & new_new_n12260__;
  assign new_new_n12262__ = ~new_new_n12048__ & ~new_new_n12261__;
  assign new_new_n12263__ = ~new_new_n12040__ & ~new_new_n12262__;
  assign new_new_n12264__ = ~new_new_n12039__ & ~new_new_n12263__;
  assign new_new_n12265__ = ~new_new_n12031__ & ~new_new_n12264__;
  assign new_new_n12266__ = ~new_new_n12030__ & ~new_new_n12265__;
  assign new_new_n12267__ = ~new_new_n12022__ & ~new_new_n12266__;
  assign new_new_n12268__ = ~new_new_n12021__ & ~new_new_n12267__;
  assign new_new_n12269__ = ~new_new_n12013__ & new_new_n12268__;
  assign new_new_n12270__ = ~new_new_n12012__ & ~new_new_n12269__;
  assign new_new_n12271__ = ~new_new_n12004__ & ~new_new_n12270__;
  assign new_new_n12272__ = ~new_new_n12003__ & ~new_new_n12271__;
  assign new_new_n12273__ = ~new_new_n11995__ & new_new_n12272__;
  assign new_new_n12274__ = ~new_new_n11994__ & ~new_new_n12273__;
  assign new_new_n12275__ = ~new_new_n11986__ & ~new_new_n12274__;
  assign new_new_n12276__ = ~new_new_n11985__ & ~new_new_n12275__;
  assign new_new_n12277__ = ~new_new_n11977__ & new_new_n12276__;
  assign new_new_n12278__ = ~new_new_n11976__ & ~new_new_n12277__;
  assign new_new_n12279__ = ~new_new_n11968__ & ~new_new_n12278__;
  assign new_new_n12280__ = ~new_new_n11967__ & ~new_new_n12279__;
  assign new_new_n12281__ = ~new_new_n11959__ & ~new_new_n12280__;
  assign new_new_n12282__ = ~new_new_n11958__ & ~new_new_n12281__;
  assign new_new_n12283__ = ~new_new_n11950__ & ~new_new_n12282__;
  assign new_new_n12284__ = ~new_new_n11949__ & ~new_new_n12283__;
  assign new_new_n12285__ = ~new_new_n11941__ & ~new_new_n12284__;
  assign new_new_n12286__ = ~new_new_n11940__ & ~new_new_n12285__;
  assign new_new_n12287__ = ~new_new_n11932__ & ~new_new_n12286__;
  assign new_new_n12288__ = ~new_new_n11931__ & ~new_new_n12287__;
  assign new_new_n12289__ = ~new_new_n11923__ & ~new_new_n12288__;
  assign new_new_n12290__ = ~new_new_n11922__ & ~new_new_n12289__;
  assign new_new_n12291__ = ~new_new_n11914__ & ~new_new_n12290__;
  assign new_new_n12292__ = ~new_new_n11913__ & ~new_new_n12291__;
  assign new_new_n12293__ = ~new_new_n11905__ & new_new_n12292__;
  assign new_new_n12294__ = ~new_new_n11904__ & ~new_new_n12293__;
  assign new_new_n12295__ = ~new_new_n11896__ & ~new_new_n12294__;
  assign new_new_n12296__ = ~new_new_n11895__ & ~new_new_n12295__;
  assign new_new_n12297__ = ~new_new_n11887__ & new_new_n12296__;
  assign new_new_n12298__ = ~new_new_n11886__ & ~new_new_n12297__;
  assign new_new_n12299__ = ~new_new_n11878__ & ~new_new_n12298__;
  assign new_new_n12300__ = ~new_new_n11877__ & ~new_new_n12299__;
  assign new_new_n12301__ = ~new_new_n11869__ & ~new_new_n12300__;
  assign new_new_n12302__ = ~new_new_n11868__ & ~new_new_n12301__;
  assign new_new_n12303__ = ~new_new_n11860__ & ~new_new_n12302__;
  assign new_new_n12304__ = ~new_new_n11859__ & ~new_new_n12303__;
  assign new_new_n12305__ = ~new_new_n11851__ & ~new_new_n12304__;
  assign new_new_n12306__ = ~new_new_n11850__ & ~new_new_n12305__;
  assign new_new_n12307__ = ~new_new_n11842__ & ~new_new_n12306__;
  assign new_new_n12308__ = ~new_new_n11841__ & ~new_new_n12307__;
  assign new_new_n12309__ = ~new_new_n11833__ & ~new_new_n12308__;
  assign new_new_n12310__ = ~new_new_n11832__ & ~new_new_n12309__;
  assign new_new_n12311__ = ~new_new_n11824__ & ~new_new_n12310__;
  assign new_new_n12312__ = ~new_new_n11823__ & ~new_new_n12311__;
  assign new_new_n12313__ = ~new_new_n11815__ & new_new_n12312__;
  assign new_new_n12314__ = ~new_new_n11814__ & ~new_new_n12313__;
  assign new_new_n12315__ = ~new_new_n11806__ & new_new_n12314__;
  assign new_new_n12316__ = ~new_new_n11805__ & ~new_new_n12315__;
  assign new_new_n12317__ = ~new_new_n11797__ & new_new_n12316__;
  assign new_new_n12318__ = ~new_new_n11796__ & ~new_new_n12317__;
  assign new_new_n12319__ = pi109 & new_new_n12318__;
  assign new_new_n12320__ = ~pi109 & ~new_new_n12318__;
  assign new_new_n12321__ = new_new_n8066__ & ~new_new_n12319__;
  assign new_new_n12322__ = ~new_new_n12320__ & new_new_n12321__;
  assign new_new_n12323__ = new_new_n11785__ & ~new_new_n12322__;
  assign new_new_n12324__ = ~pi109 & new_new_n11785__;
  assign new_new_n12325__ = new_new_n12318__ & ~new_new_n12324__;
  assign new_new_n12326__ = pi109 & ~new_new_n9808__;
  assign new_new_n12327__ = new_new_n8066__ & ~new_new_n12326__;
  assign po018 = ~new_new_n12325__ & new_new_n12327__;
  assign new_new_n12329__ = new_new_n12316__ & po018;
  assign new_new_n12330__ = ~pi108 & ~po018;
  assign new_new_n12331__ = ~new_new_n12329__ & ~new_new_n12330__;
  assign new_new_n12332__ = ~new_new_n11796__ & ~new_new_n11797__;
  assign new_new_n12333__ = ~new_new_n12331__ & ~new_new_n12332__;
  assign new_new_n12334__ = new_new_n12331__ & new_new_n12332__;
  assign new_new_n12335__ = ~new_new_n12333__ & ~new_new_n12334__;
  assign new_new_n12336__ = ~pi109 & ~new_new_n12335__;
  assign new_new_n12337__ = pi109 & new_new_n12335__;
  assign new_new_n12338__ = ~new_new_n11805__ & ~new_new_n11806__;
  assign new_new_n12339__ = ~new_new_n12314__ & po018;
  assign new_new_n12340__ = ~pi107 & ~po018;
  assign new_new_n12341__ = ~new_new_n12339__ & ~new_new_n12340__;
  assign new_new_n12342__ = new_new_n12338__ & ~new_new_n12341__;
  assign new_new_n12343__ = ~new_new_n12338__ & new_new_n12341__;
  assign new_new_n12344__ = ~new_new_n12342__ & ~new_new_n12343__;
  assign new_new_n12345__ = pi108 & ~new_new_n12344__;
  assign new_new_n12346__ = ~pi108 & new_new_n12344__;
  assign new_new_n12347__ = ~new_new_n12312__ & po018;
  assign new_new_n12348__ = pi106 & ~po018;
  assign new_new_n12349__ = ~new_new_n12347__ & ~new_new_n12348__;
  assign new_new_n12350__ = ~new_new_n11814__ & ~new_new_n11815__;
  assign new_new_n12351__ = ~new_new_n12349__ & new_new_n12350__;
  assign new_new_n12352__ = new_new_n12349__ & ~new_new_n12350__;
  assign new_new_n12353__ = ~new_new_n12351__ & ~new_new_n12352__;
  assign new_new_n12354__ = pi107 & new_new_n12353__;
  assign new_new_n12355__ = ~pi107 & ~new_new_n12353__;
  assign new_new_n12356__ = pi105 & ~new_new_n12310__;
  assign new_new_n12357__ = ~pi105 & new_new_n12310__;
  assign new_new_n12358__ = ~new_new_n12356__ & ~new_new_n12357__;
  assign new_new_n12359__ = po018 & new_new_n12358__;
  assign new_new_n12360__ = new_new_n11822__ & new_new_n12359__;
  assign new_new_n12361__ = ~new_new_n11822__ & ~new_new_n12359__;
  assign new_new_n12362__ = ~new_new_n12360__ & ~new_new_n12361__;
  assign new_new_n12363__ = pi106 & ~new_new_n12362__;
  assign new_new_n12364__ = ~pi106 & new_new_n12362__;
  assign new_new_n12365__ = ~new_new_n12308__ & po018;
  assign new_new_n12366__ = pi104 & ~po018;
  assign new_new_n12367__ = ~new_new_n12365__ & ~new_new_n12366__;
  assign new_new_n12368__ = ~new_new_n11832__ & ~new_new_n11833__;
  assign new_new_n12369__ = ~new_new_n12367__ & new_new_n12368__;
  assign new_new_n12370__ = new_new_n12367__ & ~new_new_n12368__;
  assign new_new_n12371__ = ~new_new_n12369__ & ~new_new_n12370__;
  assign new_new_n12372__ = ~pi105 & ~new_new_n12371__;
  assign new_new_n12373__ = pi105 & new_new_n12371__;
  assign new_new_n12374__ = ~new_new_n11841__ & ~new_new_n11842__;
  assign new_new_n12375__ = new_new_n12306__ & po018;
  assign new_new_n12376__ = ~pi103 & ~po018;
  assign new_new_n12377__ = ~new_new_n12375__ & ~new_new_n12376__;
  assign new_new_n12378__ = ~new_new_n12374__ & ~new_new_n12377__;
  assign new_new_n12379__ = new_new_n12374__ & new_new_n12377__;
  assign new_new_n12380__ = ~new_new_n12378__ & ~new_new_n12379__;
  assign new_new_n12381__ = ~pi104 & ~new_new_n12380__;
  assign new_new_n12382__ = pi104 & new_new_n12380__;
  assign new_new_n12383__ = ~new_new_n12304__ & po018;
  assign new_new_n12384__ = pi102 & ~po018;
  assign new_new_n12385__ = ~new_new_n12383__ & ~new_new_n12384__;
  assign new_new_n12386__ = ~new_new_n11850__ & ~new_new_n11851__;
  assign new_new_n12387__ = ~new_new_n12385__ & new_new_n12386__;
  assign new_new_n12388__ = new_new_n12385__ & ~new_new_n12386__;
  assign new_new_n12389__ = ~new_new_n12387__ & ~new_new_n12388__;
  assign new_new_n12390__ = ~pi103 & ~new_new_n12389__;
  assign new_new_n12391__ = pi103 & new_new_n12389__;
  assign new_new_n12392__ = ~pi101 & ~new_new_n12302__;
  assign new_new_n12393__ = pi101 & new_new_n12302__;
  assign new_new_n12394__ = ~new_new_n12392__ & ~new_new_n12393__;
  assign new_new_n12395__ = po018 & ~new_new_n12394__;
  assign new_new_n12396__ = new_new_n11858__ & new_new_n12395__;
  assign new_new_n12397__ = ~new_new_n11858__ & ~new_new_n12395__;
  assign new_new_n12398__ = ~new_new_n12396__ & ~new_new_n12397__;
  assign new_new_n12399__ = pi102 & ~new_new_n12398__;
  assign new_new_n12400__ = ~pi102 & new_new_n12398__;
  assign new_new_n12401__ = ~new_new_n12300__ & po018;
  assign new_new_n12402__ = pi100 & ~po018;
  assign new_new_n12403__ = ~new_new_n12401__ & ~new_new_n12402__;
  assign new_new_n12404__ = ~new_new_n11868__ & ~new_new_n11869__;
  assign new_new_n12405__ = ~new_new_n12403__ & new_new_n12404__;
  assign new_new_n12406__ = new_new_n12403__ & ~new_new_n12404__;
  assign new_new_n12407__ = ~new_new_n12405__ & ~new_new_n12406__;
  assign new_new_n12408__ = pi101 & new_new_n12407__;
  assign new_new_n12409__ = ~pi101 & ~new_new_n12407__;
  assign new_new_n12410__ = pi099 & ~new_new_n12298__;
  assign new_new_n12411__ = ~pi099 & new_new_n12298__;
  assign new_new_n12412__ = ~new_new_n12410__ & ~new_new_n12411__;
  assign new_new_n12413__ = po018 & new_new_n12412__;
  assign new_new_n12414__ = new_new_n11876__ & new_new_n12413__;
  assign new_new_n12415__ = ~new_new_n11876__ & ~new_new_n12413__;
  assign new_new_n12416__ = ~new_new_n12414__ & ~new_new_n12415__;
  assign new_new_n12417__ = pi100 & ~new_new_n12416__;
  assign new_new_n12418__ = ~pi100 & new_new_n12416__;
  assign new_new_n12419__ = ~new_new_n11886__ & ~new_new_n11887__;
  assign new_new_n12420__ = ~new_new_n12296__ & po018;
  assign new_new_n12421__ = ~pi098 & ~po018;
  assign new_new_n12422__ = ~new_new_n12420__ & ~new_new_n12421__;
  assign new_new_n12423__ = new_new_n12419__ & ~new_new_n12422__;
  assign new_new_n12424__ = ~new_new_n12419__ & new_new_n12422__;
  assign new_new_n12425__ = ~new_new_n12423__ & ~new_new_n12424__;
  assign new_new_n12426__ = pi099 & ~new_new_n12425__;
  assign new_new_n12427__ = ~pi099 & new_new_n12425__;
  assign new_new_n12428__ = ~new_new_n11895__ & ~new_new_n11896__;
  assign new_new_n12429__ = ~new_new_n12294__ & po018;
  assign new_new_n12430__ = ~pi097 & ~po018;
  assign new_new_n12431__ = ~new_new_n12429__ & ~new_new_n12430__;
  assign new_new_n12432__ = new_new_n12428__ & ~new_new_n12431__;
  assign new_new_n12433__ = ~new_new_n12428__ & new_new_n12431__;
  assign new_new_n12434__ = ~new_new_n12432__ & ~new_new_n12433__;
  assign new_new_n12435__ = pi098 & ~new_new_n12434__;
  assign new_new_n12436__ = ~pi098 & new_new_n12434__;
  assign new_new_n12437__ = ~new_new_n11904__ & ~new_new_n11905__;
  assign new_new_n12438__ = pi096 & ~po018;
  assign new_new_n12439__ = ~new_new_n12292__ & po018;
  assign new_new_n12440__ = ~new_new_n12438__ & ~new_new_n12439__;
  assign new_new_n12441__ = new_new_n12437__ & ~new_new_n12440__;
  assign new_new_n12442__ = ~new_new_n12437__ & new_new_n12440__;
  assign new_new_n12443__ = ~new_new_n12441__ & ~new_new_n12442__;
  assign new_new_n12444__ = ~pi097 & ~new_new_n12443__;
  assign new_new_n12445__ = pi097 & new_new_n12443__;
  assign new_new_n12446__ = ~new_new_n12290__ & po018;
  assign new_new_n12447__ = pi095 & ~po018;
  assign new_new_n12448__ = ~new_new_n12446__ & ~new_new_n12447__;
  assign new_new_n12449__ = ~new_new_n11913__ & ~new_new_n11914__;
  assign new_new_n12450__ = ~new_new_n12448__ & new_new_n12449__;
  assign new_new_n12451__ = new_new_n12448__ & ~new_new_n12449__;
  assign new_new_n12452__ = ~new_new_n12450__ & ~new_new_n12451__;
  assign new_new_n12453__ = ~pi096 & ~new_new_n12452__;
  assign new_new_n12454__ = pi096 & new_new_n12452__;
  assign new_new_n12455__ = pi094 & ~new_new_n12288__;
  assign new_new_n12456__ = ~pi094 & new_new_n12288__;
  assign new_new_n12457__ = ~new_new_n12455__ & ~new_new_n12456__;
  assign new_new_n12458__ = po018 & new_new_n12457__;
  assign new_new_n12459__ = new_new_n11921__ & new_new_n12458__;
  assign new_new_n12460__ = ~new_new_n11921__ & ~new_new_n12458__;
  assign new_new_n12461__ = ~new_new_n12459__ & ~new_new_n12460__;
  assign new_new_n12462__ = pi095 & ~new_new_n12461__;
  assign new_new_n12463__ = ~pi095 & new_new_n12461__;
  assign new_new_n12464__ = ~new_new_n12286__ & po018;
  assign new_new_n12465__ = pi093 & ~po018;
  assign new_new_n12466__ = ~new_new_n12464__ & ~new_new_n12465__;
  assign new_new_n12467__ = ~new_new_n11931__ & ~new_new_n11932__;
  assign new_new_n12468__ = ~new_new_n12466__ & new_new_n12467__;
  assign new_new_n12469__ = new_new_n12466__ & ~new_new_n12467__;
  assign new_new_n12470__ = ~new_new_n12468__ & ~new_new_n12469__;
  assign new_new_n12471__ = ~pi094 & ~new_new_n12470__;
  assign new_new_n12472__ = pi094 & new_new_n12470__;
  assign new_new_n12473__ = ~new_new_n11940__ & ~new_new_n11941__;
  assign new_new_n12474__ = new_new_n12284__ & po018;
  assign new_new_n12475__ = ~pi092 & ~po018;
  assign new_new_n12476__ = ~new_new_n12474__ & ~new_new_n12475__;
  assign new_new_n12477__ = ~new_new_n12473__ & ~new_new_n12476__;
  assign new_new_n12478__ = new_new_n12473__ & new_new_n12476__;
  assign new_new_n12479__ = ~new_new_n12477__ & ~new_new_n12478__;
  assign new_new_n12480__ = ~pi093 & ~new_new_n12479__;
  assign new_new_n12481__ = pi093 & new_new_n12479__;
  assign new_new_n12482__ = new_new_n12282__ & po018;
  assign new_new_n12483__ = ~pi091 & ~po018;
  assign new_new_n12484__ = ~new_new_n12482__ & ~new_new_n12483__;
  assign new_new_n12485__ = ~new_new_n11949__ & ~new_new_n11950__;
  assign new_new_n12486__ = ~new_new_n12484__ & ~new_new_n12485__;
  assign new_new_n12487__ = new_new_n12484__ & new_new_n12485__;
  assign new_new_n12488__ = ~new_new_n12486__ & ~new_new_n12487__;
  assign new_new_n12489__ = ~pi092 & ~new_new_n12488__;
  assign new_new_n12490__ = pi092 & new_new_n12488__;
  assign new_new_n12491__ = ~new_new_n11958__ & ~new_new_n11959__;
  assign new_new_n12492__ = pi090 & ~po018;
  assign new_new_n12493__ = ~new_new_n12280__ & po018;
  assign new_new_n12494__ = ~new_new_n12492__ & ~new_new_n12493__;
  assign new_new_n12495__ = new_new_n12491__ & ~new_new_n12494__;
  assign new_new_n12496__ = ~new_new_n12491__ & new_new_n12494__;
  assign new_new_n12497__ = ~new_new_n12495__ & ~new_new_n12496__;
  assign new_new_n12498__ = pi091 & new_new_n12497__;
  assign new_new_n12499__ = ~pi091 & ~new_new_n12497__;
  assign new_new_n12500__ = ~new_new_n11967__ & ~new_new_n11968__;
  assign new_new_n12501__ = pi089 & ~po018;
  assign new_new_n12502__ = ~new_new_n12278__ & po018;
  assign new_new_n12503__ = ~new_new_n12501__ & ~new_new_n12502__;
  assign new_new_n12504__ = new_new_n12500__ & ~new_new_n12503__;
  assign new_new_n12505__ = ~new_new_n12500__ & new_new_n12503__;
  assign new_new_n12506__ = ~new_new_n12504__ & ~new_new_n12505__;
  assign new_new_n12507__ = pi090 & new_new_n12506__;
  assign new_new_n12508__ = ~pi090 & ~new_new_n12506__;
  assign new_new_n12509__ = ~new_new_n11976__ & ~new_new_n11977__;
  assign new_new_n12510__ = ~new_new_n12276__ & po018;
  assign new_new_n12511__ = ~pi088 & ~po018;
  assign new_new_n12512__ = ~new_new_n12510__ & ~new_new_n12511__;
  assign new_new_n12513__ = new_new_n12509__ & ~new_new_n12512__;
  assign new_new_n12514__ = ~new_new_n12509__ & new_new_n12512__;
  assign new_new_n12515__ = ~new_new_n12513__ & ~new_new_n12514__;
  assign new_new_n12516__ = pi089 & ~new_new_n12515__;
  assign new_new_n12517__ = ~pi089 & new_new_n12515__;
  assign new_new_n12518__ = ~new_new_n11985__ & ~new_new_n11986__;
  assign new_new_n12519__ = ~new_new_n12274__ & po018;
  assign new_new_n12520__ = ~pi087 & ~po018;
  assign new_new_n12521__ = ~new_new_n12519__ & ~new_new_n12520__;
  assign new_new_n12522__ = new_new_n12518__ & ~new_new_n12521__;
  assign new_new_n12523__ = ~new_new_n12518__ & new_new_n12521__;
  assign new_new_n12524__ = ~new_new_n12522__ & ~new_new_n12523__;
  assign new_new_n12525__ = pi088 & ~new_new_n12524__;
  assign new_new_n12526__ = ~pi088 & new_new_n12524__;
  assign new_new_n12527__ = ~new_new_n11994__ & ~new_new_n11995__;
  assign new_new_n12528__ = ~new_new_n12272__ & po018;
  assign new_new_n12529__ = pi086 & ~po018;
  assign new_new_n12530__ = ~new_new_n12528__ & ~new_new_n12529__;
  assign new_new_n12531__ = new_new_n12527__ & ~new_new_n12530__;
  assign new_new_n12532__ = ~new_new_n12527__ & new_new_n12530__;
  assign new_new_n12533__ = ~new_new_n12531__ & ~new_new_n12532__;
  assign new_new_n12534__ = pi087 & new_new_n12533__;
  assign new_new_n12535__ = ~pi087 & ~new_new_n12533__;
  assign new_new_n12536__ = pi085 & ~new_new_n12270__;
  assign new_new_n12537__ = ~pi085 & new_new_n12270__;
  assign new_new_n12538__ = ~new_new_n12536__ & ~new_new_n12537__;
  assign new_new_n12539__ = po018 & new_new_n12538__;
  assign new_new_n12540__ = new_new_n12002__ & new_new_n12539__;
  assign new_new_n12541__ = ~new_new_n12002__ & ~new_new_n12539__;
  assign new_new_n12542__ = ~new_new_n12540__ & ~new_new_n12541__;
  assign new_new_n12543__ = pi086 & ~new_new_n12542__;
  assign new_new_n12544__ = ~pi086 & new_new_n12542__;
  assign new_new_n12545__ = ~new_new_n12012__ & ~new_new_n12013__;
  assign new_new_n12546__ = ~new_new_n12268__ & po018;
  assign new_new_n12547__ = ~pi084 & ~po018;
  assign new_new_n12548__ = ~new_new_n12546__ & ~new_new_n12547__;
  assign new_new_n12549__ = new_new_n12545__ & ~new_new_n12548__;
  assign new_new_n12550__ = ~new_new_n12545__ & new_new_n12548__;
  assign new_new_n12551__ = ~new_new_n12549__ & ~new_new_n12550__;
  assign new_new_n12552__ = pi085 & ~new_new_n12551__;
  assign new_new_n12553__ = ~pi085 & new_new_n12551__;
  assign new_new_n12554__ = ~new_new_n12021__ & ~new_new_n12022__;
  assign new_new_n12555__ = ~new_new_n12266__ & po018;
  assign new_new_n12556__ = ~pi083 & ~po018;
  assign new_new_n12557__ = ~new_new_n12555__ & ~new_new_n12556__;
  assign new_new_n12558__ = ~new_new_n12554__ & ~new_new_n12557__;
  assign new_new_n12559__ = new_new_n12554__ & new_new_n12557__;
  assign new_new_n12560__ = ~new_new_n12558__ & ~new_new_n12559__;
  assign new_new_n12561__ = pi084 & new_new_n12560__;
  assign new_new_n12562__ = ~pi084 & ~new_new_n12560__;
  assign new_new_n12563__ = new_new_n12264__ & po018;
  assign new_new_n12564__ = pi082 & ~po018;
  assign new_new_n12565__ = ~new_new_n12563__ & ~new_new_n12564__;
  assign new_new_n12566__ = ~new_new_n12030__ & ~new_new_n12031__;
  assign new_new_n12567__ = ~new_new_n12565__ & ~new_new_n12566__;
  assign new_new_n12568__ = new_new_n12565__ & new_new_n12566__;
  assign new_new_n12569__ = ~new_new_n12567__ & ~new_new_n12568__;
  assign new_new_n12570__ = pi083 & ~new_new_n12569__;
  assign new_new_n12571__ = ~pi083 & new_new_n12569__;
  assign new_new_n12572__ = ~new_new_n12039__ & ~new_new_n12040__;
  assign new_new_n12573__ = ~new_new_n12262__ & po018;
  assign new_new_n12574__ = ~pi081 & ~po018;
  assign new_new_n12575__ = ~new_new_n12573__ & ~new_new_n12574__;
  assign new_new_n12576__ = new_new_n12572__ & ~new_new_n12575__;
  assign new_new_n12577__ = ~new_new_n12572__ & new_new_n12575__;
  assign new_new_n12578__ = ~new_new_n12576__ & ~new_new_n12577__;
  assign new_new_n12579__ = pi082 & ~new_new_n12578__;
  assign new_new_n12580__ = ~pi082 & new_new_n12578__;
  assign new_new_n12581__ = ~new_new_n12260__ & po018;
  assign new_new_n12582__ = pi080 & ~po018;
  assign new_new_n12583__ = ~new_new_n12581__ & ~new_new_n12582__;
  assign new_new_n12584__ = ~new_new_n12048__ & ~new_new_n12049__;
  assign new_new_n12585__ = ~new_new_n12583__ & new_new_n12584__;
  assign new_new_n12586__ = new_new_n12583__ & ~new_new_n12584__;
  assign new_new_n12587__ = ~new_new_n12585__ & ~new_new_n12586__;
  assign new_new_n12588__ = ~pi081 & ~new_new_n12587__;
  assign new_new_n12589__ = pi081 & new_new_n12587__;
  assign new_new_n12590__ = ~pi079 & ~new_new_n12258__;
  assign new_new_n12591__ = pi079 & new_new_n12258__;
  assign new_new_n12592__ = ~new_new_n12590__ & ~new_new_n12591__;
  assign new_new_n12593__ = po018 & ~new_new_n12592__;
  assign new_new_n12594__ = new_new_n12056__ & new_new_n12593__;
  assign new_new_n12595__ = ~new_new_n12056__ & ~new_new_n12593__;
  assign new_new_n12596__ = ~new_new_n12594__ & ~new_new_n12595__;
  assign new_new_n12597__ = ~pi080 & new_new_n12596__;
  assign new_new_n12598__ = pi080 & ~new_new_n12596__;
  assign new_new_n12599__ = ~new_new_n12066__ & ~new_new_n12067__;
  assign new_new_n12600__ = ~new_new_n12256__ & po018;
  assign new_new_n12601__ = pi078 & ~po018;
  assign new_new_n12602__ = ~new_new_n12600__ & ~new_new_n12601__;
  assign new_new_n12603__ = new_new_n12599__ & ~new_new_n12602__;
  assign new_new_n12604__ = ~new_new_n12599__ & new_new_n12602__;
  assign new_new_n12605__ = ~new_new_n12603__ & ~new_new_n12604__;
  assign new_new_n12606__ = ~pi079 & ~new_new_n12605__;
  assign new_new_n12607__ = pi079 & new_new_n12605__;
  assign new_new_n12608__ = pi077 & ~new_new_n12254__;
  assign new_new_n12609__ = ~pi077 & new_new_n12254__;
  assign new_new_n12610__ = ~new_new_n12608__ & ~new_new_n12609__;
  assign new_new_n12611__ = po018 & new_new_n12610__;
  assign new_new_n12612__ = new_new_n12074__ & new_new_n12611__;
  assign new_new_n12613__ = ~new_new_n12074__ & ~new_new_n12611__;
  assign new_new_n12614__ = ~new_new_n12612__ & ~new_new_n12613__;
  assign new_new_n12615__ = pi078 & ~new_new_n12614__;
  assign new_new_n12616__ = ~pi078 & new_new_n12614__;
  assign new_new_n12617__ = pi076 & ~new_new_n12252__;
  assign new_new_n12618__ = ~pi076 & new_new_n12252__;
  assign new_new_n12619__ = ~new_new_n12617__ & ~new_new_n12618__;
  assign new_new_n12620__ = po018 & new_new_n12619__;
  assign new_new_n12621__ = new_new_n12083__ & new_new_n12620__;
  assign new_new_n12622__ = ~new_new_n12083__ & ~new_new_n12620__;
  assign new_new_n12623__ = ~new_new_n12621__ & ~new_new_n12622__;
  assign new_new_n12624__ = ~pi077 & new_new_n12623__;
  assign new_new_n12625__ = pi077 & ~new_new_n12623__;
  assign new_new_n12626__ = ~new_new_n12093__ & ~new_new_n12094__;
  assign new_new_n12627__ = ~new_new_n12250__ & po018;
  assign new_new_n12628__ = ~pi075 & ~po018;
  assign new_new_n12629__ = ~new_new_n12627__ & ~new_new_n12628__;
  assign new_new_n12630__ = new_new_n12626__ & ~new_new_n12629__;
  assign new_new_n12631__ = ~new_new_n12626__ & new_new_n12629__;
  assign new_new_n12632__ = ~new_new_n12630__ & ~new_new_n12631__;
  assign new_new_n12633__ = ~pi076 & new_new_n12632__;
  assign new_new_n12634__ = pi076 & ~new_new_n12632__;
  assign new_new_n12635__ = ~new_new_n12102__ & ~new_new_n12103__;
  assign new_new_n12636__ = ~new_new_n12248__ & po018;
  assign new_new_n12637__ = ~pi074 & ~po018;
  assign new_new_n12638__ = ~new_new_n12636__ & ~new_new_n12637__;
  assign new_new_n12639__ = new_new_n12635__ & ~new_new_n12638__;
  assign new_new_n12640__ = ~new_new_n12635__ & new_new_n12638__;
  assign new_new_n12641__ = ~new_new_n12639__ & ~new_new_n12640__;
  assign new_new_n12642__ = ~pi075 & new_new_n12641__;
  assign new_new_n12643__ = pi075 & ~new_new_n12641__;
  assign new_new_n12644__ = ~new_new_n12111__ & ~new_new_n12112__;
  assign new_new_n12645__ = ~new_new_n12246__ & po018;
  assign new_new_n12646__ = ~pi073 & ~po018;
  assign new_new_n12647__ = ~new_new_n12645__ & ~new_new_n12646__;
  assign new_new_n12648__ = ~new_new_n12644__ & ~new_new_n12647__;
  assign new_new_n12649__ = new_new_n12644__ & new_new_n12647__;
  assign new_new_n12650__ = ~new_new_n12648__ & ~new_new_n12649__;
  assign new_new_n12651__ = ~pi074 & ~new_new_n12650__;
  assign new_new_n12652__ = pi074 & new_new_n12650__;
  assign new_new_n12653__ = new_new_n12244__ & po018;
  assign new_new_n12654__ = ~pi072 & ~po018;
  assign new_new_n12655__ = ~new_new_n12653__ & ~new_new_n12654__;
  assign new_new_n12656__ = ~new_new_n12120__ & ~new_new_n12121__;
  assign new_new_n12657__ = ~new_new_n12655__ & ~new_new_n12656__;
  assign new_new_n12658__ = new_new_n12655__ & new_new_n12656__;
  assign new_new_n12659__ = ~new_new_n12657__ & ~new_new_n12658__;
  assign new_new_n12660__ = pi073 & new_new_n12659__;
  assign new_new_n12661__ = ~pi073 & ~new_new_n12659__;
  assign new_new_n12662__ = pi071 & ~new_new_n12242__;
  assign new_new_n12663__ = ~pi071 & new_new_n12242__;
  assign new_new_n12664__ = ~new_new_n12662__ & ~new_new_n12663__;
  assign new_new_n12665__ = po018 & new_new_n12664__;
  assign new_new_n12666__ = new_new_n12128__ & new_new_n12665__;
  assign new_new_n12667__ = ~new_new_n12128__ & ~new_new_n12665__;
  assign new_new_n12668__ = ~new_new_n12666__ & ~new_new_n12667__;
  assign new_new_n12669__ = pi072 & ~new_new_n12668__;
  assign new_new_n12670__ = ~pi072 & new_new_n12668__;
  assign new_new_n12671__ = ~new_new_n12136__ & ~new_new_n12137__;
  assign new_new_n12672__ = pi070 & ~po018;
  assign new_new_n12673__ = ~new_new_n12240__ & po018;
  assign new_new_n12674__ = ~new_new_n12672__ & ~new_new_n12673__;
  assign new_new_n12675__ = new_new_n12671__ & new_new_n12674__;
  assign new_new_n12676__ = ~new_new_n12671__ & ~new_new_n12674__;
  assign new_new_n12677__ = ~new_new_n12675__ & ~new_new_n12676__;
  assign new_new_n12678__ = ~pi071 & new_new_n12677__;
  assign new_new_n12679__ = pi071 & ~new_new_n12677__;
  assign new_new_n12680__ = new_new_n12238__ & po018;
  assign new_new_n12681__ = pi069 & ~po018;
  assign new_new_n12682__ = ~new_new_n12680__ & ~new_new_n12681__;
  assign new_new_n12683__ = ~new_new_n12143__ & ~new_new_n12144__;
  assign new_new_n12684__ = ~new_new_n12682__ & ~new_new_n12683__;
  assign new_new_n12685__ = new_new_n12682__ & new_new_n12683__;
  assign new_new_n12686__ = ~new_new_n12684__ & ~new_new_n12685__;
  assign new_new_n12687__ = ~pi070 & new_new_n12686__;
  assign new_new_n12688__ = pi070 & ~new_new_n12686__;
  assign new_new_n12689__ = ~new_new_n12228__ & ~new_new_n12229__;
  assign new_new_n12690__ = po018 & new_new_n12689__;
  assign new_new_n12691__ = new_new_n12236__ & new_new_n12690__;
  assign new_new_n12692__ = ~new_new_n12236__ & ~new_new_n12690__;
  assign new_new_n12693__ = ~new_new_n12691__ & ~new_new_n12692__;
  assign new_new_n12694__ = ~pi069 & ~new_new_n12693__;
  assign new_new_n12695__ = pi069 & new_new_n12693__;
  assign new_new_n12696__ = ~new_new_n12184__ & ~new_new_n12185__;
  assign new_new_n12697__ = ~new_new_n12225__ & po018;
  assign new_new_n12698__ = pi067 & ~po018;
  assign new_new_n12699__ = ~new_new_n12697__ & ~new_new_n12698__;
  assign new_new_n12700__ = new_new_n12696__ & ~new_new_n12699__;
  assign new_new_n12701__ = ~new_new_n12696__ & new_new_n12699__;
  assign new_new_n12702__ = ~new_new_n12700__ & ~new_new_n12701__;
  assign new_new_n12703__ = ~pi068 & ~new_new_n12702__;
  assign new_new_n12704__ = pi068 & new_new_n12702__;
  assign new_new_n12705__ = ~new_new_n12198__ & po018;
  assign new_new_n12706__ = ~new_new_n12223__ & new_new_n12705__;
  assign new_new_n12707__ = new_new_n12222__ & ~new_new_n12706__;
  assign new_new_n12708__ = new_new_n12224__ & new_new_n12705__;
  assign new_new_n12709__ = ~new_new_n12707__ & ~new_new_n12708__;
  assign new_new_n12710__ = ~pi067 & ~new_new_n12709__;
  assign new_new_n12711__ = pi067 & new_new_n12709__;
  assign new_new_n12712__ = ~pi017 & pi064;
  assign new_new_n12713__ = ~pi065 & ~new_new_n12712__;
  assign new_new_n12714__ = pi064 & po018;
  assign new_new_n12715__ = ~pi018 & ~new_new_n12714__;
  assign new_new_n12716__ = ~new_new_n12713__ & new_new_n12715__;
  assign new_new_n12717__ = ~pi017 & pi065;
  assign new_new_n12718__ = pi017 & ~pi065;
  assign new_new_n12719__ = pi018 & ~new_new_n12718__;
  assign new_new_n12720__ = po018 & new_new_n12719__;
  assign new_new_n12721__ = ~new_new_n12717__ & ~new_new_n12720__;
  assign new_new_n12722__ = pi064 & ~new_new_n12721__;
  assign new_new_n12723__ = ~new_new_n12716__ & ~new_new_n12722__;
  assign new_new_n12724__ = ~pi065 & ~po019;
  assign new_new_n12725__ = pi065 & po018;
  assign new_new_n12726__ = new_new_n12194__ & new_new_n12725__;
  assign new_new_n12727__ = ~new_new_n12724__ & ~new_new_n12726__;
  assign new_new_n12728__ = pi018 & ~new_new_n12727__;
  assign new_new_n12729__ = ~new_new_n332__ & po018;
  assign new_new_n12730__ = ~new_new_n12194__ & ~new_new_n12729__;
  assign new_new_n12731__ = po019 & ~po018;
  assign new_new_n12732__ = ~new_new_n426__ & ~po019;
  assign new_new_n12733__ = ~pi018 & ~new_new_n12199__;
  assign new_new_n12734__ = ~new_new_n12732__ & new_new_n12733__;
  assign new_new_n12735__ = ~new_new_n12731__ & new_new_n12734__;
  assign new_new_n12736__ = ~new_new_n12730__ & ~new_new_n12735__;
  assign new_new_n12737__ = ~new_new_n12728__ & new_new_n12736__;
  assign new_new_n12738__ = ~pi019 & ~new_new_n12737__;
  assign new_new_n12739__ = po018 & new_new_n12724__;
  assign new_new_n12740__ = ~new_new_n12199__ & ~new_new_n12739__;
  assign new_new_n12741__ = ~pi018 & ~new_new_n12740__;
  assign new_new_n12742__ = ~new_new_n12731__ & ~new_new_n12741__;
  assign new_new_n12743__ = pi064 & ~new_new_n12742__;
  assign new_new_n12744__ = ~new_new_n12194__ & ~new_new_n12725__;
  assign new_new_n12745__ = pi018 & ~new_new_n12199__;
  assign new_new_n12746__ = pi064 & ~new_new_n12745__;
  assign new_new_n12747__ = ~new_new_n12744__ & ~new_new_n12746__;
  assign new_new_n12748__ = ~new_new_n12743__ & ~new_new_n12747__;
  assign new_new_n12749__ = pi019 & ~new_new_n12748__;
  assign new_new_n12750__ = ~new_new_n12738__ & ~new_new_n12749__;
  assign new_new_n12751__ = new_new_n12723__ & new_new_n12750__;
  assign new_new_n12752__ = pi066 & ~new_new_n12751__;
  assign new_new_n12753__ = ~new_new_n12723__ & ~new_new_n12750__;
  assign new_new_n12754__ = ~new_new_n12752__ & ~new_new_n12753__;
  assign new_new_n12755__ = ~new_new_n12711__ & new_new_n12754__;
  assign new_new_n12756__ = ~new_new_n12710__ & ~new_new_n12755__;
  assign new_new_n12757__ = ~new_new_n12704__ & ~new_new_n12756__;
  assign new_new_n12758__ = ~new_new_n12703__ & ~new_new_n12757__;
  assign new_new_n12759__ = ~new_new_n12695__ & ~new_new_n12758__;
  assign new_new_n12760__ = ~new_new_n12694__ & ~new_new_n12759__;
  assign new_new_n12761__ = ~new_new_n12688__ & ~new_new_n12760__;
  assign new_new_n12762__ = ~new_new_n12687__ & ~new_new_n12761__;
  assign new_new_n12763__ = ~new_new_n12679__ & ~new_new_n12762__;
  assign new_new_n12764__ = ~new_new_n12678__ & ~new_new_n12763__;
  assign new_new_n12765__ = ~new_new_n12670__ & new_new_n12764__;
  assign new_new_n12766__ = ~new_new_n12669__ & ~new_new_n12765__;
  assign new_new_n12767__ = ~new_new_n12661__ & ~new_new_n12766__;
  assign new_new_n12768__ = ~new_new_n12660__ & ~new_new_n12767__;
  assign new_new_n12769__ = ~new_new_n12652__ & new_new_n12768__;
  assign new_new_n12770__ = ~new_new_n12651__ & ~new_new_n12769__;
  assign new_new_n12771__ = ~new_new_n12643__ & ~new_new_n12770__;
  assign new_new_n12772__ = ~new_new_n12642__ & ~new_new_n12771__;
  assign new_new_n12773__ = ~new_new_n12634__ & ~new_new_n12772__;
  assign new_new_n12774__ = ~new_new_n12633__ & ~new_new_n12773__;
  assign new_new_n12775__ = ~new_new_n12625__ & ~new_new_n12774__;
  assign new_new_n12776__ = ~new_new_n12624__ & ~new_new_n12775__;
  assign new_new_n12777__ = ~new_new_n12616__ & new_new_n12776__;
  assign new_new_n12778__ = ~new_new_n12615__ & ~new_new_n12777__;
  assign new_new_n12779__ = ~new_new_n12607__ & new_new_n12778__;
  assign new_new_n12780__ = ~new_new_n12606__ & ~new_new_n12779__;
  assign new_new_n12781__ = ~new_new_n12598__ & ~new_new_n12780__;
  assign new_new_n12782__ = ~new_new_n12597__ & ~new_new_n12781__;
  assign new_new_n12783__ = ~new_new_n12589__ & ~new_new_n12782__;
  assign new_new_n12784__ = ~new_new_n12588__ & ~new_new_n12783__;
  assign new_new_n12785__ = ~new_new_n12580__ & new_new_n12784__;
  assign new_new_n12786__ = ~new_new_n12579__ & ~new_new_n12785__;
  assign new_new_n12787__ = ~new_new_n12571__ & ~new_new_n12786__;
  assign new_new_n12788__ = ~new_new_n12570__ & ~new_new_n12787__;
  assign new_new_n12789__ = ~new_new_n12562__ & ~new_new_n12788__;
  assign new_new_n12790__ = ~new_new_n12561__ & ~new_new_n12789__;
  assign new_new_n12791__ = ~new_new_n12553__ & ~new_new_n12790__;
  assign new_new_n12792__ = ~new_new_n12552__ & ~new_new_n12791__;
  assign new_new_n12793__ = ~new_new_n12544__ & ~new_new_n12792__;
  assign new_new_n12794__ = ~new_new_n12543__ & ~new_new_n12793__;
  assign new_new_n12795__ = ~new_new_n12535__ & ~new_new_n12794__;
  assign new_new_n12796__ = ~new_new_n12534__ & ~new_new_n12795__;
  assign new_new_n12797__ = ~new_new_n12526__ & ~new_new_n12796__;
  assign new_new_n12798__ = ~new_new_n12525__ & ~new_new_n12797__;
  assign new_new_n12799__ = ~new_new_n12517__ & ~new_new_n12798__;
  assign new_new_n12800__ = ~new_new_n12516__ & ~new_new_n12799__;
  assign new_new_n12801__ = ~new_new_n12508__ & ~new_new_n12800__;
  assign new_new_n12802__ = ~new_new_n12507__ & ~new_new_n12801__;
  assign new_new_n12803__ = ~new_new_n12499__ & ~new_new_n12802__;
  assign new_new_n12804__ = ~new_new_n12498__ & ~new_new_n12803__;
  assign new_new_n12805__ = ~new_new_n12490__ & new_new_n12804__;
  assign new_new_n12806__ = ~new_new_n12489__ & ~new_new_n12805__;
  assign new_new_n12807__ = ~new_new_n12481__ & ~new_new_n12806__;
  assign new_new_n12808__ = ~new_new_n12480__ & ~new_new_n12807__;
  assign new_new_n12809__ = ~new_new_n12472__ & ~new_new_n12808__;
  assign new_new_n12810__ = ~new_new_n12471__ & ~new_new_n12809__;
  assign new_new_n12811__ = ~new_new_n12463__ & new_new_n12810__;
  assign new_new_n12812__ = ~new_new_n12462__ & ~new_new_n12811__;
  assign new_new_n12813__ = ~new_new_n12454__ & new_new_n12812__;
  assign new_new_n12814__ = ~new_new_n12453__ & ~new_new_n12813__;
  assign new_new_n12815__ = ~new_new_n12445__ & ~new_new_n12814__;
  assign new_new_n12816__ = ~new_new_n12444__ & ~new_new_n12815__;
  assign new_new_n12817__ = ~new_new_n12436__ & new_new_n12816__;
  assign new_new_n12818__ = ~new_new_n12435__ & ~new_new_n12817__;
  assign new_new_n12819__ = ~new_new_n12427__ & ~new_new_n12818__;
  assign new_new_n12820__ = ~new_new_n12426__ & ~new_new_n12819__;
  assign new_new_n12821__ = ~new_new_n12418__ & ~new_new_n12820__;
  assign new_new_n12822__ = ~new_new_n12417__ & ~new_new_n12821__;
  assign new_new_n12823__ = ~new_new_n12409__ & ~new_new_n12822__;
  assign new_new_n12824__ = ~new_new_n12408__ & ~new_new_n12823__;
  assign new_new_n12825__ = ~new_new_n12400__ & ~new_new_n12824__;
  assign new_new_n12826__ = ~new_new_n12399__ & ~new_new_n12825__;
  assign new_new_n12827__ = ~new_new_n12391__ & new_new_n12826__;
  assign new_new_n12828__ = ~new_new_n12390__ & ~new_new_n12827__;
  assign new_new_n12829__ = ~new_new_n12382__ & ~new_new_n12828__;
  assign new_new_n12830__ = ~new_new_n12381__ & ~new_new_n12829__;
  assign new_new_n12831__ = ~new_new_n12373__ & ~new_new_n12830__;
  assign new_new_n12832__ = ~new_new_n12372__ & ~new_new_n12831__;
  assign new_new_n12833__ = ~new_new_n12364__ & new_new_n12832__;
  assign new_new_n12834__ = ~new_new_n12363__ & ~new_new_n12833__;
  assign new_new_n12835__ = ~new_new_n12355__ & ~new_new_n12834__;
  assign new_new_n12836__ = ~new_new_n12354__ & ~new_new_n12835__;
  assign new_new_n12837__ = ~new_new_n12346__ & ~new_new_n12836__;
  assign new_new_n12838__ = ~new_new_n12345__ & ~new_new_n12837__;
  assign new_new_n12839__ = ~new_new_n12337__ & new_new_n12838__;
  assign new_new_n12840__ = ~new_new_n12336__ & ~new_new_n12839__;
  assign new_new_n12841__ = pi110 & new_new_n12840__;
  assign new_new_n12842__ = ~pi110 & ~new_new_n12840__;
  assign new_new_n12843__ = new_new_n8065__ & ~new_new_n12841__;
  assign new_new_n12844__ = ~new_new_n12842__ & new_new_n12843__;
  assign new_new_n12845__ = new_new_n12323__ & ~new_new_n12844__;
  assign new_new_n12846__ = ~pi116 & new_new_n269__;
  assign new_new_n12847__ = ~pi115 & new_new_n12846__;
  assign new_new_n12848__ = ~pi114 & new_new_n12847__;
  assign new_new_n12849__ = ~pi113 & new_new_n12848__;
  assign new_new_n12850__ = ~new_new_n12323__ & ~new_new_n12842__;
  assign po017 = new_new_n12843__ & ~new_new_n12850__;
  assign new_new_n12852__ = pi108 & ~new_new_n12836__;
  assign new_new_n12853__ = ~pi108 & new_new_n12836__;
  assign new_new_n12854__ = ~new_new_n12852__ & ~new_new_n12853__;
  assign new_new_n12855__ = po017 & new_new_n12854__;
  assign new_new_n12856__ = new_new_n12344__ & new_new_n12855__;
  assign new_new_n12857__ = ~new_new_n12344__ & ~new_new_n12855__;
  assign new_new_n12858__ = ~new_new_n12856__ & ~new_new_n12857__;
  assign new_new_n12859__ = pi111 & ~new_new_n12323__;
  assign new_new_n12860__ = new_new_n274__ & ~new_new_n12859__;
  assign new_new_n12861__ = ~pi111 & new_new_n12845__;
  assign new_new_n12862__ = new_new_n12838__ & po017;
  assign new_new_n12863__ = ~pi109 & ~po017;
  assign new_new_n12864__ = ~new_new_n12862__ & ~new_new_n12863__;
  assign new_new_n12865__ = ~new_new_n12336__ & ~new_new_n12337__;
  assign new_new_n12866__ = ~new_new_n12864__ & ~new_new_n12865__;
  assign new_new_n12867__ = new_new_n12864__ & new_new_n12865__;
  assign new_new_n12868__ = ~new_new_n12866__ & ~new_new_n12867__;
  assign new_new_n12869__ = ~pi110 & ~new_new_n12868__;
  assign new_new_n12870__ = pi110 & new_new_n12868__;
  assign new_new_n12871__ = pi109 & ~new_new_n12858__;
  assign new_new_n12872__ = ~pi109 & new_new_n12858__;
  assign new_new_n12873__ = ~new_new_n12354__ & ~new_new_n12355__;
  assign new_new_n12874__ = pi107 & ~po017;
  assign new_new_n12875__ = ~new_new_n12834__ & po017;
  assign new_new_n12876__ = ~new_new_n12874__ & ~new_new_n12875__;
  assign new_new_n12877__ = new_new_n12873__ & ~new_new_n12876__;
  assign new_new_n12878__ = ~new_new_n12873__ & new_new_n12876__;
  assign new_new_n12879__ = ~new_new_n12877__ & ~new_new_n12878__;
  assign new_new_n12880__ = pi108 & new_new_n12879__;
  assign new_new_n12881__ = ~pi108 & ~new_new_n12879__;
  assign new_new_n12882__ = ~new_new_n12363__ & ~new_new_n12364__;
  assign new_new_n12883__ = ~new_new_n12832__ & po017;
  assign new_new_n12884__ = ~pi106 & ~po017;
  assign new_new_n12885__ = ~new_new_n12883__ & ~new_new_n12884__;
  assign new_new_n12886__ = new_new_n12882__ & ~new_new_n12885__;
  assign new_new_n12887__ = ~new_new_n12882__ & new_new_n12885__;
  assign new_new_n12888__ = ~new_new_n12886__ & ~new_new_n12887__;
  assign new_new_n12889__ = pi107 & ~new_new_n12888__;
  assign new_new_n12890__ = ~pi107 & new_new_n12888__;
  assign new_new_n12891__ = ~new_new_n12372__ & ~new_new_n12373__;
  assign new_new_n12892__ = ~new_new_n12830__ & po017;
  assign new_new_n12893__ = ~pi105 & ~po017;
  assign new_new_n12894__ = ~new_new_n12892__ & ~new_new_n12893__;
  assign new_new_n12895__ = ~new_new_n12891__ & ~new_new_n12894__;
  assign new_new_n12896__ = new_new_n12891__ & new_new_n12894__;
  assign new_new_n12897__ = ~new_new_n12895__ & ~new_new_n12896__;
  assign new_new_n12898__ = pi106 & new_new_n12897__;
  assign new_new_n12899__ = ~pi106 & ~new_new_n12897__;
  assign new_new_n12900__ = ~new_new_n12381__ & ~new_new_n12382__;
  assign new_new_n12901__ = ~new_new_n12828__ & po017;
  assign new_new_n12902__ = ~pi104 & ~po017;
  assign new_new_n12903__ = ~new_new_n12901__ & ~new_new_n12902__;
  assign new_new_n12904__ = new_new_n12900__ & ~new_new_n12903__;
  assign new_new_n12905__ = ~new_new_n12900__ & new_new_n12903__;
  assign new_new_n12906__ = ~new_new_n12904__ & ~new_new_n12905__;
  assign new_new_n12907__ = pi105 & ~new_new_n12906__;
  assign new_new_n12908__ = ~pi105 & new_new_n12906__;
  assign new_new_n12909__ = ~new_new_n12399__ & ~new_new_n12400__;
  assign new_new_n12910__ = pi102 & ~po017;
  assign new_new_n12911__ = ~new_new_n12824__ & po017;
  assign new_new_n12912__ = ~new_new_n12910__ & ~new_new_n12911__;
  assign new_new_n12913__ = new_new_n12909__ & ~new_new_n12912__;
  assign new_new_n12914__ = ~new_new_n12909__ & new_new_n12912__;
  assign new_new_n12915__ = ~new_new_n12913__ & ~new_new_n12914__;
  assign new_new_n12916__ = ~pi103 & ~new_new_n12915__;
  assign new_new_n12917__ = pi103 & new_new_n12915__;
  assign new_new_n12918__ = ~new_new_n12822__ & po017;
  assign new_new_n12919__ = pi101 & ~po017;
  assign new_new_n12920__ = ~new_new_n12918__ & ~new_new_n12919__;
  assign new_new_n12921__ = ~new_new_n12408__ & ~new_new_n12409__;
  assign new_new_n12922__ = ~new_new_n12920__ & new_new_n12921__;
  assign new_new_n12923__ = new_new_n12920__ & ~new_new_n12921__;
  assign new_new_n12924__ = ~new_new_n12922__ & ~new_new_n12923__;
  assign new_new_n12925__ = ~pi102 & ~new_new_n12924__;
  assign new_new_n12926__ = pi102 & new_new_n12924__;
  assign new_new_n12927__ = ~new_new_n12417__ & ~new_new_n12418__;
  assign new_new_n12928__ = ~new_new_n12820__ & po017;
  assign new_new_n12929__ = pi100 & ~po017;
  assign new_new_n12930__ = ~new_new_n12928__ & ~new_new_n12929__;
  assign new_new_n12931__ = new_new_n12927__ & new_new_n12930__;
  assign new_new_n12932__ = ~new_new_n12927__ & ~new_new_n12930__;
  assign new_new_n12933__ = ~new_new_n12931__ & ~new_new_n12932__;
  assign new_new_n12934__ = ~pi101 & new_new_n12933__;
  assign new_new_n12935__ = pi101 & ~new_new_n12933__;
  assign new_new_n12936__ = pi099 & ~new_new_n12818__;
  assign new_new_n12937__ = ~pi099 & new_new_n12818__;
  assign new_new_n12938__ = ~new_new_n12936__ & ~new_new_n12937__;
  assign new_new_n12939__ = po017 & new_new_n12938__;
  assign new_new_n12940__ = new_new_n12425__ & new_new_n12939__;
  assign new_new_n12941__ = ~new_new_n12425__ & ~new_new_n12939__;
  assign new_new_n12942__ = ~new_new_n12940__ & ~new_new_n12941__;
  assign new_new_n12943__ = ~pi100 & new_new_n12942__;
  assign new_new_n12944__ = pi100 & ~new_new_n12942__;
  assign new_new_n12945__ = ~new_new_n12435__ & ~new_new_n12436__;
  assign new_new_n12946__ = ~new_new_n12816__ & po017;
  assign new_new_n12947__ = ~pi098 & ~po017;
  assign new_new_n12948__ = ~new_new_n12946__ & ~new_new_n12947__;
  assign new_new_n12949__ = new_new_n12945__ & ~new_new_n12948__;
  assign new_new_n12950__ = ~new_new_n12945__ & new_new_n12948__;
  assign new_new_n12951__ = ~new_new_n12949__ & ~new_new_n12950__;
  assign new_new_n12952__ = ~pi099 & new_new_n12951__;
  assign new_new_n12953__ = pi099 & ~new_new_n12951__;
  assign new_new_n12954__ = ~pi097 & ~new_new_n12814__;
  assign new_new_n12955__ = pi097 & new_new_n12814__;
  assign new_new_n12956__ = ~new_new_n12954__ & ~new_new_n12955__;
  assign new_new_n12957__ = po017 & new_new_n12956__;
  assign new_new_n12958__ = new_new_n12443__ & new_new_n12957__;
  assign new_new_n12959__ = ~new_new_n12443__ & ~new_new_n12957__;
  assign new_new_n12960__ = ~new_new_n12958__ & ~new_new_n12959__;
  assign new_new_n12961__ = ~pi098 & ~new_new_n12960__;
  assign new_new_n12962__ = pi098 & new_new_n12960__;
  assign new_new_n12963__ = ~new_new_n12453__ & ~new_new_n12454__;
  assign new_new_n12964__ = pi096 & ~po017;
  assign new_new_n12965__ = ~new_new_n12812__ & po017;
  assign new_new_n12966__ = ~new_new_n12964__ & ~new_new_n12965__;
  assign new_new_n12967__ = new_new_n12963__ & ~new_new_n12966__;
  assign new_new_n12968__ = ~new_new_n12963__ & new_new_n12966__;
  assign new_new_n12969__ = ~new_new_n12967__ & ~new_new_n12968__;
  assign new_new_n12970__ = ~pi097 & ~new_new_n12969__;
  assign new_new_n12971__ = pi097 & new_new_n12969__;
  assign new_new_n12972__ = new_new_n12810__ & po017;
  assign new_new_n12973__ = pi095 & ~po017;
  assign new_new_n12974__ = ~new_new_n12972__ & ~new_new_n12973__;
  assign new_new_n12975__ = ~new_new_n12462__ & ~new_new_n12463__;
  assign new_new_n12976__ = ~new_new_n12974__ & ~new_new_n12975__;
  assign new_new_n12977__ = new_new_n12974__ & new_new_n12975__;
  assign new_new_n12978__ = ~new_new_n12976__ & ~new_new_n12977__;
  assign new_new_n12979__ = pi096 & ~new_new_n12978__;
  assign new_new_n12980__ = ~pi096 & new_new_n12978__;
  assign new_new_n12981__ = ~pi094 & ~new_new_n12808__;
  assign new_new_n12982__ = pi094 & new_new_n12808__;
  assign new_new_n12983__ = ~new_new_n12981__ & ~new_new_n12982__;
  assign new_new_n12984__ = po017 & new_new_n12983__;
  assign new_new_n12985__ = new_new_n12470__ & new_new_n12984__;
  assign new_new_n12986__ = ~new_new_n12470__ & ~new_new_n12984__;
  assign new_new_n12987__ = ~new_new_n12985__ & ~new_new_n12986__;
  assign new_new_n12988__ = ~pi095 & ~new_new_n12987__;
  assign new_new_n12989__ = pi095 & new_new_n12987__;
  assign new_new_n12990__ = ~new_new_n12480__ & ~new_new_n12481__;
  assign new_new_n12991__ = ~new_new_n12806__ & po017;
  assign new_new_n12992__ = ~pi093 & ~po017;
  assign new_new_n12993__ = ~new_new_n12991__ & ~new_new_n12992__;
  assign new_new_n12994__ = new_new_n12990__ & ~new_new_n12993__;
  assign new_new_n12995__ = ~new_new_n12990__ & new_new_n12993__;
  assign new_new_n12996__ = ~new_new_n12994__ & ~new_new_n12995__;
  assign new_new_n12997__ = ~pi094 & new_new_n12996__;
  assign new_new_n12998__ = pi094 & ~new_new_n12996__;
  assign new_new_n12999__ = ~new_new_n12489__ & ~new_new_n12490__;
  assign new_new_n13000__ = pi092 & ~po017;
  assign new_new_n13001__ = ~new_new_n12804__ & po017;
  assign new_new_n13002__ = ~new_new_n13000__ & ~new_new_n13001__;
  assign new_new_n13003__ = new_new_n12999__ & ~new_new_n13002__;
  assign new_new_n13004__ = ~new_new_n12999__ & new_new_n13002__;
  assign new_new_n13005__ = ~new_new_n13003__ & ~new_new_n13004__;
  assign new_new_n13006__ = ~pi093 & ~new_new_n13005__;
  assign new_new_n13007__ = pi093 & new_new_n13005__;
  assign new_new_n13008__ = ~new_new_n12802__ & po017;
  assign new_new_n13009__ = pi091 & ~po017;
  assign new_new_n13010__ = ~new_new_n13008__ & ~new_new_n13009__;
  assign new_new_n13011__ = ~new_new_n12498__ & ~new_new_n12499__;
  assign new_new_n13012__ = ~new_new_n13010__ & new_new_n13011__;
  assign new_new_n13013__ = new_new_n13010__ & ~new_new_n13011__;
  assign new_new_n13014__ = ~new_new_n13012__ & ~new_new_n13013__;
  assign new_new_n13015__ = ~pi092 & ~new_new_n13014__;
  assign new_new_n13016__ = pi092 & new_new_n13014__;
  assign new_new_n13017__ = ~new_new_n12507__ & ~new_new_n12508__;
  assign new_new_n13018__ = new_new_n12800__ & po017;
  assign new_new_n13019__ = ~pi090 & ~po017;
  assign new_new_n13020__ = ~new_new_n13018__ & ~new_new_n13019__;
  assign new_new_n13021__ = ~new_new_n13017__ & ~new_new_n13020__;
  assign new_new_n13022__ = new_new_n13017__ & new_new_n13020__;
  assign new_new_n13023__ = ~new_new_n13021__ & ~new_new_n13022__;
  assign new_new_n13024__ = ~pi091 & ~new_new_n13023__;
  assign new_new_n13025__ = pi091 & new_new_n13023__;
  assign new_new_n13026__ = pi089 & ~new_new_n12798__;
  assign new_new_n13027__ = ~pi089 & new_new_n12798__;
  assign new_new_n13028__ = ~new_new_n13026__ & ~new_new_n13027__;
  assign new_new_n13029__ = po017 & new_new_n13028__;
  assign new_new_n13030__ = new_new_n12515__ & new_new_n13029__;
  assign new_new_n13031__ = ~new_new_n12515__ & ~new_new_n13029__;
  assign new_new_n13032__ = ~new_new_n13030__ & ~new_new_n13031__;
  assign new_new_n13033__ = pi090 & ~new_new_n13032__;
  assign new_new_n13034__ = ~pi090 & new_new_n13032__;
  assign new_new_n13035__ = ~new_new_n12525__ & ~new_new_n12526__;
  assign new_new_n13036__ = pi088 & ~po017;
  assign new_new_n13037__ = ~new_new_n12796__ & po017;
  assign new_new_n13038__ = ~new_new_n13036__ & ~new_new_n13037__;
  assign new_new_n13039__ = new_new_n13035__ & ~new_new_n13038__;
  assign new_new_n13040__ = ~new_new_n13035__ & new_new_n13038__;
  assign new_new_n13041__ = ~new_new_n13039__ & ~new_new_n13040__;
  assign new_new_n13042__ = ~pi089 & ~new_new_n13041__;
  assign new_new_n13043__ = pi089 & new_new_n13041__;
  assign new_new_n13044__ = ~new_new_n12794__ & po017;
  assign new_new_n13045__ = pi087 & ~po017;
  assign new_new_n13046__ = ~new_new_n13044__ & ~new_new_n13045__;
  assign new_new_n13047__ = ~new_new_n12534__ & ~new_new_n12535__;
  assign new_new_n13048__ = ~new_new_n13046__ & new_new_n13047__;
  assign new_new_n13049__ = new_new_n13046__ & ~new_new_n13047__;
  assign new_new_n13050__ = ~new_new_n13048__ & ~new_new_n13049__;
  assign new_new_n13051__ = ~pi088 & ~new_new_n13050__;
  assign new_new_n13052__ = pi088 & new_new_n13050__;
  assign new_new_n13053__ = ~new_new_n12543__ & ~new_new_n12544__;
  assign new_new_n13054__ = pi086 & ~po017;
  assign new_new_n13055__ = ~new_new_n12792__ & po017;
  assign new_new_n13056__ = ~new_new_n13054__ & ~new_new_n13055__;
  assign new_new_n13057__ = new_new_n13053__ & new_new_n13056__;
  assign new_new_n13058__ = ~new_new_n13053__ & ~new_new_n13056__;
  assign new_new_n13059__ = ~new_new_n13057__ & ~new_new_n13058__;
  assign new_new_n13060__ = pi087 & ~new_new_n13059__;
  assign new_new_n13061__ = ~pi087 & new_new_n13059__;
  assign new_new_n13062__ = ~new_new_n12552__ & ~new_new_n12553__;
  assign new_new_n13063__ = pi085 & ~po017;
  assign new_new_n13064__ = ~new_new_n12790__ & po017;
  assign new_new_n13065__ = ~new_new_n13063__ & ~new_new_n13064__;
  assign new_new_n13066__ = new_new_n13062__ & new_new_n13065__;
  assign new_new_n13067__ = ~new_new_n13062__ & ~new_new_n13065__;
  assign new_new_n13068__ = ~new_new_n13066__ & ~new_new_n13067__;
  assign new_new_n13069__ = pi086 & ~new_new_n13068__;
  assign new_new_n13070__ = ~pi086 & new_new_n13068__;
  assign new_new_n13071__ = new_new_n12788__ & po017;
  assign new_new_n13072__ = ~pi084 & ~po017;
  assign new_new_n13073__ = ~new_new_n13071__ & ~new_new_n13072__;
  assign new_new_n13074__ = ~new_new_n12561__ & ~new_new_n12562__;
  assign new_new_n13075__ = ~new_new_n13073__ & ~new_new_n13074__;
  assign new_new_n13076__ = new_new_n13073__ & new_new_n13074__;
  assign new_new_n13077__ = ~new_new_n13075__ & ~new_new_n13076__;
  assign new_new_n13078__ = pi085 & new_new_n13077__;
  assign new_new_n13079__ = ~pi085 & ~new_new_n13077__;
  assign new_new_n13080__ = ~new_new_n12570__ & ~new_new_n12571__;
  assign new_new_n13081__ = pi083 & ~po017;
  assign new_new_n13082__ = ~new_new_n12786__ & po017;
  assign new_new_n13083__ = ~new_new_n13081__ & ~new_new_n13082__;
  assign new_new_n13084__ = new_new_n13080__ & ~new_new_n13083__;
  assign new_new_n13085__ = ~new_new_n13080__ & new_new_n13083__;
  assign new_new_n13086__ = ~new_new_n13084__ & ~new_new_n13085__;
  assign new_new_n13087__ = pi084 & new_new_n13086__;
  assign new_new_n13088__ = ~pi084 & ~new_new_n13086__;
  assign new_new_n13089__ = ~new_new_n12579__ & ~new_new_n12580__;
  assign new_new_n13090__ = ~new_new_n12784__ & po017;
  assign new_new_n13091__ = ~pi082 & ~po017;
  assign new_new_n13092__ = ~new_new_n13090__ & ~new_new_n13091__;
  assign new_new_n13093__ = new_new_n13089__ & ~new_new_n13092__;
  assign new_new_n13094__ = ~new_new_n13089__ & new_new_n13092__;
  assign new_new_n13095__ = ~new_new_n13093__ & ~new_new_n13094__;
  assign new_new_n13096__ = pi083 & ~new_new_n13095__;
  assign new_new_n13097__ = ~pi083 & new_new_n13095__;
  assign new_new_n13098__ = ~new_new_n12588__ & ~new_new_n12589__;
  assign new_new_n13099__ = ~new_new_n12782__ & po017;
  assign new_new_n13100__ = ~pi081 & ~po017;
  assign new_new_n13101__ = ~new_new_n13099__ & ~new_new_n13100__;
  assign new_new_n13102__ = new_new_n13098__ & ~new_new_n13101__;
  assign new_new_n13103__ = ~new_new_n13098__ & new_new_n13101__;
  assign new_new_n13104__ = ~new_new_n13102__ & ~new_new_n13103__;
  assign new_new_n13105__ = pi082 & ~new_new_n13104__;
  assign new_new_n13106__ = ~pi082 & new_new_n13104__;
  assign new_new_n13107__ = ~new_new_n12597__ & ~new_new_n12598__;
  assign new_new_n13108__ = ~new_new_n12780__ & po017;
  assign new_new_n13109__ = ~pi080 & ~po017;
  assign new_new_n13110__ = ~new_new_n13108__ & ~new_new_n13109__;
  assign new_new_n13111__ = new_new_n13107__ & ~new_new_n13110__;
  assign new_new_n13112__ = ~new_new_n13107__ & new_new_n13110__;
  assign new_new_n13113__ = ~new_new_n13111__ & ~new_new_n13112__;
  assign new_new_n13114__ = pi081 & ~new_new_n13113__;
  assign new_new_n13115__ = ~pi081 & new_new_n13113__;
  assign new_new_n13116__ = ~new_new_n12606__ & ~new_new_n12607__;
  assign new_new_n13117__ = pi079 & ~po017;
  assign new_new_n13118__ = ~new_new_n12778__ & po017;
  assign new_new_n13119__ = ~new_new_n13117__ & ~new_new_n13118__;
  assign new_new_n13120__ = new_new_n13116__ & ~new_new_n13119__;
  assign new_new_n13121__ = ~new_new_n13116__ & new_new_n13119__;
  assign new_new_n13122__ = ~new_new_n13120__ & ~new_new_n13121__;
  assign new_new_n13123__ = pi080 & new_new_n13122__;
  assign new_new_n13124__ = ~pi080 & ~new_new_n13122__;
  assign new_new_n13125__ = ~new_new_n12615__ & ~new_new_n12616__;
  assign new_new_n13126__ = ~new_new_n12776__ & po017;
  assign new_new_n13127__ = ~pi078 & ~po017;
  assign new_new_n13128__ = ~new_new_n13126__ & ~new_new_n13127__;
  assign new_new_n13129__ = new_new_n13125__ & ~new_new_n13128__;
  assign new_new_n13130__ = ~new_new_n13125__ & new_new_n13128__;
  assign new_new_n13131__ = ~new_new_n13129__ & ~new_new_n13130__;
  assign new_new_n13132__ = pi079 & ~new_new_n13131__;
  assign new_new_n13133__ = ~pi079 & new_new_n13131__;
  assign new_new_n13134__ = ~new_new_n12624__ & ~new_new_n12625__;
  assign new_new_n13135__ = ~new_new_n12774__ & po017;
  assign new_new_n13136__ = ~pi077 & ~po017;
  assign new_new_n13137__ = ~new_new_n13135__ & ~new_new_n13136__;
  assign new_new_n13138__ = new_new_n13134__ & ~new_new_n13137__;
  assign new_new_n13139__ = ~new_new_n13134__ & new_new_n13137__;
  assign new_new_n13140__ = ~new_new_n13138__ & ~new_new_n13139__;
  assign new_new_n13141__ = pi078 & ~new_new_n13140__;
  assign new_new_n13142__ = ~pi078 & new_new_n13140__;
  assign new_new_n13143__ = ~new_new_n12633__ & ~new_new_n12634__;
  assign new_new_n13144__ = ~new_new_n12772__ & po017;
  assign new_new_n13145__ = ~pi076 & ~po017;
  assign new_new_n13146__ = ~new_new_n13144__ & ~new_new_n13145__;
  assign new_new_n13147__ = new_new_n13143__ & ~new_new_n13146__;
  assign new_new_n13148__ = ~new_new_n13143__ & new_new_n13146__;
  assign new_new_n13149__ = ~new_new_n13147__ & ~new_new_n13148__;
  assign new_new_n13150__ = pi077 & ~new_new_n13149__;
  assign new_new_n13151__ = ~pi077 & new_new_n13149__;
  assign new_new_n13152__ = ~new_new_n12642__ & ~new_new_n12643__;
  assign new_new_n13153__ = ~new_new_n12770__ & po017;
  assign new_new_n13154__ = ~pi075 & ~po017;
  assign new_new_n13155__ = ~new_new_n13153__ & ~new_new_n13154__;
  assign new_new_n13156__ = new_new_n13152__ & ~new_new_n13155__;
  assign new_new_n13157__ = ~new_new_n13152__ & new_new_n13155__;
  assign new_new_n13158__ = ~new_new_n13156__ & ~new_new_n13157__;
  assign new_new_n13159__ = pi076 & ~new_new_n13158__;
  assign new_new_n13160__ = ~pi076 & new_new_n13158__;
  assign new_new_n13161__ = ~new_new_n12768__ & po017;
  assign new_new_n13162__ = pi074 & ~po017;
  assign new_new_n13163__ = ~new_new_n13161__ & ~new_new_n13162__;
  assign new_new_n13164__ = ~new_new_n12651__ & ~new_new_n12652__;
  assign new_new_n13165__ = ~new_new_n13163__ & new_new_n13164__;
  assign new_new_n13166__ = new_new_n13163__ & ~new_new_n13164__;
  assign new_new_n13167__ = ~new_new_n13165__ & ~new_new_n13166__;
  assign new_new_n13168__ = ~pi075 & ~new_new_n13167__;
  assign new_new_n13169__ = pi075 & new_new_n13167__;
  assign new_new_n13170__ = ~new_new_n12660__ & ~new_new_n12661__;
  assign new_new_n13171__ = pi073 & ~po017;
  assign new_new_n13172__ = ~new_new_n12766__ & po017;
  assign new_new_n13173__ = ~new_new_n13171__ & ~new_new_n13172__;
  assign new_new_n13174__ = new_new_n13170__ & ~new_new_n13173__;
  assign new_new_n13175__ = ~new_new_n13170__ & new_new_n13173__;
  assign new_new_n13176__ = ~new_new_n13174__ & ~new_new_n13175__;
  assign new_new_n13177__ = ~pi074 & ~new_new_n13176__;
  assign new_new_n13178__ = pi074 & new_new_n13176__;
  assign new_new_n13179__ = ~new_new_n12669__ & ~new_new_n12670__;
  assign new_new_n13180__ = ~new_new_n12764__ & po017;
  assign new_new_n13181__ = ~pi072 & ~po017;
  assign new_new_n13182__ = ~new_new_n13180__ & ~new_new_n13181__;
  assign new_new_n13183__ = new_new_n13179__ & new_new_n13182__;
  assign new_new_n13184__ = ~new_new_n13179__ & ~new_new_n13182__;
  assign new_new_n13185__ = ~new_new_n13183__ & ~new_new_n13184__;
  assign new_new_n13186__ = pi073 & new_new_n13185__;
  assign new_new_n13187__ = ~pi073 & ~new_new_n13185__;
  assign new_new_n13188__ = new_new_n12762__ & po017;
  assign new_new_n13189__ = pi071 & ~po017;
  assign new_new_n13190__ = ~new_new_n13188__ & ~new_new_n13189__;
  assign new_new_n13191__ = ~new_new_n12678__ & ~new_new_n12679__;
  assign new_new_n13192__ = ~new_new_n13190__ & ~new_new_n13191__;
  assign new_new_n13193__ = new_new_n13190__ & new_new_n13191__;
  assign new_new_n13194__ = ~new_new_n13192__ & ~new_new_n13193__;
  assign new_new_n13195__ = pi072 & ~new_new_n13194__;
  assign new_new_n13196__ = ~pi072 & new_new_n13194__;
  assign new_new_n13197__ = ~pi069 & ~new_new_n12758__;
  assign new_new_n13198__ = pi069 & new_new_n12758__;
  assign new_new_n13199__ = ~new_new_n13197__ & ~new_new_n13198__;
  assign new_new_n13200__ = po017 & new_new_n13199__;
  assign new_new_n13201__ = new_new_n12693__ & new_new_n13200__;
  assign new_new_n13202__ = ~new_new_n12693__ & ~new_new_n13200__;
  assign new_new_n13203__ = ~new_new_n13201__ & ~new_new_n13202__;
  assign new_new_n13204__ = pi070 & new_new_n13203__;
  assign new_new_n13205__ = ~pi070 & ~new_new_n13203__;
  assign new_new_n13206__ = ~new_new_n12710__ & ~new_new_n12711__;
  assign new_new_n13207__ = new_new_n12754__ & po017;
  assign new_new_n13208__ = ~pi067 & ~po017;
  assign new_new_n13209__ = ~new_new_n13207__ & ~new_new_n13208__;
  assign new_new_n13210__ = ~new_new_n13206__ & ~new_new_n13209__;
  assign new_new_n13211__ = new_new_n13206__ & new_new_n13209__;
  assign new_new_n13212__ = ~new_new_n13210__ & ~new_new_n13211__;
  assign new_new_n13213__ = ~pi068 & ~new_new_n13212__;
  assign new_new_n13214__ = pi068 & new_new_n13212__;
  assign new_new_n13215__ = pi065 & new_new_n12712__;
  assign new_new_n13216__ = pi018 & new_new_n12714__;
  assign new_new_n13217__ = ~new_new_n12715__ & ~new_new_n13216__;
  assign new_new_n13218__ = ~new_new_n12713__ & ~new_new_n13217__;
  assign new_new_n13219__ = ~new_new_n13215__ & ~new_new_n13218__;
  assign new_new_n13220__ = pi066 & ~new_new_n13219__;
  assign new_new_n13221__ = ~pi066 & new_new_n13219__;
  assign new_new_n13222__ = ~new_new_n13220__ & ~new_new_n13221__;
  assign new_new_n13223__ = po017 & new_new_n13222__;
  assign new_new_n13224__ = ~new_new_n12750__ & new_new_n13223__;
  assign new_new_n13225__ = new_new_n12750__ & ~new_new_n13223__;
  assign new_new_n13226__ = ~new_new_n13224__ & ~new_new_n13225__;
  assign new_new_n13227__ = ~pi067 & ~new_new_n13226__;
  assign new_new_n13228__ = pi067 & new_new_n13226__;
  assign new_new_n13229__ = pi016 & ~pi065;
  assign new_new_n13230__ = pi017 & po017;
  assign new_new_n13231__ = pi065 & new_new_n13217__;
  assign new_new_n13232__ = ~pi065 & ~new_new_n13217__;
  assign new_new_n13233__ = ~new_new_n13231__ & ~new_new_n13232__;
  assign new_new_n13234__ = ~new_new_n13229__ & ~new_new_n13233__;
  assign new_new_n13235__ = new_new_n13230__ & new_new_n13234__;
  assign new_new_n13236__ = ~new_new_n12717__ & po017;
  assign new_new_n13237__ = ~pi016 & ~new_new_n12718__;
  assign new_new_n13238__ = ~new_new_n13217__ & new_new_n13237__;
  assign new_new_n13239__ = ~new_new_n13236__ & new_new_n13238__;
  assign new_new_n13240__ = ~new_new_n13235__ & ~new_new_n13239__;
  assign new_new_n13241__ = pi064 & ~new_new_n13240__;
  assign new_new_n13242__ = ~po017 & new_new_n13217__;
  assign new_new_n13243__ = pi064 & po017;
  assign new_new_n13244__ = new_new_n12717__ & ~new_new_n13243__;
  assign new_new_n13245__ = po017 & ~new_new_n13217__;
  assign new_new_n13246__ = ~new_new_n13242__ & ~new_new_n13245__;
  assign new_new_n13247__ = new_new_n13244__ & new_new_n13246__;
  assign new_new_n13248__ = ~pi066 & ~new_new_n13247__;
  assign new_new_n13249__ = ~new_new_n13241__ & new_new_n13248__;
  assign new_new_n13250__ = ~pi016 & pi065;
  assign new_new_n13251__ = new_new_n12712__ & ~new_new_n13250__;
  assign new_new_n13252__ = ~new_new_n13233__ & new_new_n13251__;
  assign new_new_n13253__ = pi017 & new_new_n403__;
  assign new_new_n13254__ = ~new_new_n13217__ & new_new_n13253__;
  assign new_new_n13255__ = ~new_new_n13252__ & ~new_new_n13254__;
  assign new_new_n13256__ = po017 & ~new_new_n13255__;
  assign new_new_n13257__ = pi065 & po017;
  assign new_new_n13258__ = pi016 & ~new_new_n13257__;
  assign new_new_n13259__ = ~pi065 & ~po017;
  assign new_new_n13260__ = ~pi017 & ~new_new_n13259__;
  assign new_new_n13261__ = new_new_n13258__ & ~new_new_n13260__;
  assign new_new_n13262__ = pi017 & ~new_new_n426__;
  assign new_new_n13263__ = ~po017 & new_new_n13262__;
  assign new_new_n13264__ = ~new_new_n332__ & ~new_new_n13263__;
  assign new_new_n13265__ = ~new_new_n13261__ & new_new_n13264__;
  assign new_new_n13266__ = new_new_n13217__ & ~new_new_n13265__;
  assign new_new_n13267__ = ~new_new_n13249__ & ~new_new_n13256__;
  assign new_new_n13268__ = ~new_new_n13266__ & new_new_n13267__;
  assign new_new_n13269__ = ~new_new_n13228__ & ~new_new_n13268__;
  assign new_new_n13270__ = ~new_new_n13227__ & ~new_new_n13269__;
  assign new_new_n13271__ = ~new_new_n13214__ & ~new_new_n13270__;
  assign new_new_n13272__ = ~new_new_n13213__ & ~new_new_n13271__;
  assign new_new_n13273__ = pi069 & new_new_n13272__;
  assign new_new_n13274__ = ~pi069 & ~new_new_n13272__;
  assign new_new_n13275__ = ~new_new_n12703__ & ~new_new_n12704__;
  assign new_new_n13276__ = ~new_new_n12756__ & po017;
  assign new_new_n13277__ = ~pi068 & ~po017;
  assign new_new_n13278__ = ~new_new_n13276__ & ~new_new_n13277__;
  assign new_new_n13279__ = new_new_n13275__ & ~new_new_n13278__;
  assign new_new_n13280__ = ~new_new_n13275__ & new_new_n13278__;
  assign new_new_n13281__ = ~new_new_n13279__ & ~new_new_n13280__;
  assign new_new_n13282__ = ~new_new_n13274__ & ~new_new_n13281__;
  assign new_new_n13283__ = ~new_new_n13273__ & ~new_new_n13282__;
  assign new_new_n13284__ = ~new_new_n13205__ & ~new_new_n13283__;
  assign new_new_n13285__ = ~new_new_n13204__ & ~new_new_n13284__;
  assign new_new_n13286__ = pi071 & ~new_new_n13285__;
  assign new_new_n13287__ = ~pi071 & new_new_n13285__;
  assign new_new_n13288__ = new_new_n12760__ & po017;
  assign new_new_n13289__ = pi070 & ~po017;
  assign new_new_n13290__ = ~new_new_n13288__ & ~new_new_n13289__;
  assign new_new_n13291__ = ~new_new_n12687__ & ~new_new_n12688__;
  assign new_new_n13292__ = ~new_new_n13290__ & ~new_new_n13291__;
  assign new_new_n13293__ = new_new_n13290__ & new_new_n13291__;
  assign new_new_n13294__ = ~new_new_n13292__ & ~new_new_n13293__;
  assign new_new_n13295__ = ~new_new_n13287__ & ~new_new_n13294__;
  assign new_new_n13296__ = ~new_new_n13286__ & ~new_new_n13295__;
  assign new_new_n13297__ = ~new_new_n13196__ & ~new_new_n13296__;
  assign new_new_n13298__ = ~new_new_n13195__ & ~new_new_n13297__;
  assign new_new_n13299__ = ~new_new_n13187__ & ~new_new_n13298__;
  assign new_new_n13300__ = ~new_new_n13186__ & ~new_new_n13299__;
  assign new_new_n13301__ = ~new_new_n13178__ & new_new_n13300__;
  assign new_new_n13302__ = ~new_new_n13177__ & ~new_new_n13301__;
  assign new_new_n13303__ = ~new_new_n13169__ & ~new_new_n13302__;
  assign new_new_n13304__ = ~new_new_n13168__ & ~new_new_n13303__;
  assign new_new_n13305__ = ~new_new_n13160__ & new_new_n13304__;
  assign new_new_n13306__ = ~new_new_n13159__ & ~new_new_n13305__;
  assign new_new_n13307__ = ~new_new_n13151__ & ~new_new_n13306__;
  assign new_new_n13308__ = ~new_new_n13150__ & ~new_new_n13307__;
  assign new_new_n13309__ = ~new_new_n13142__ & ~new_new_n13308__;
  assign new_new_n13310__ = ~new_new_n13141__ & ~new_new_n13309__;
  assign new_new_n13311__ = ~new_new_n13133__ & ~new_new_n13310__;
  assign new_new_n13312__ = ~new_new_n13132__ & ~new_new_n13311__;
  assign new_new_n13313__ = ~new_new_n13124__ & ~new_new_n13312__;
  assign new_new_n13314__ = ~new_new_n13123__ & ~new_new_n13313__;
  assign new_new_n13315__ = ~new_new_n13115__ & ~new_new_n13314__;
  assign new_new_n13316__ = ~new_new_n13114__ & ~new_new_n13315__;
  assign new_new_n13317__ = ~new_new_n13106__ & ~new_new_n13316__;
  assign new_new_n13318__ = ~new_new_n13105__ & ~new_new_n13317__;
  assign new_new_n13319__ = ~new_new_n13097__ & ~new_new_n13318__;
  assign new_new_n13320__ = ~new_new_n13096__ & ~new_new_n13319__;
  assign new_new_n13321__ = ~new_new_n13088__ & ~new_new_n13320__;
  assign new_new_n13322__ = ~new_new_n13087__ & ~new_new_n13321__;
  assign new_new_n13323__ = ~new_new_n13079__ & ~new_new_n13322__;
  assign new_new_n13324__ = ~new_new_n13078__ & ~new_new_n13323__;
  assign new_new_n13325__ = ~new_new_n13070__ & ~new_new_n13324__;
  assign new_new_n13326__ = ~new_new_n13069__ & ~new_new_n13325__;
  assign new_new_n13327__ = ~new_new_n13061__ & ~new_new_n13326__;
  assign new_new_n13328__ = ~new_new_n13060__ & ~new_new_n13327__;
  assign new_new_n13329__ = ~new_new_n13052__ & new_new_n13328__;
  assign new_new_n13330__ = ~new_new_n13051__ & ~new_new_n13329__;
  assign new_new_n13331__ = ~new_new_n13043__ & ~new_new_n13330__;
  assign new_new_n13332__ = ~new_new_n13042__ & ~new_new_n13331__;
  assign new_new_n13333__ = ~new_new_n13034__ & new_new_n13332__;
  assign new_new_n13334__ = ~new_new_n13033__ & ~new_new_n13333__;
  assign new_new_n13335__ = ~new_new_n13025__ & new_new_n13334__;
  assign new_new_n13336__ = ~new_new_n13024__ & ~new_new_n13335__;
  assign new_new_n13337__ = ~new_new_n13016__ & ~new_new_n13336__;
  assign new_new_n13338__ = ~new_new_n13015__ & ~new_new_n13337__;
  assign new_new_n13339__ = ~new_new_n13007__ & ~new_new_n13338__;
  assign new_new_n13340__ = ~new_new_n13006__ & ~new_new_n13339__;
  assign new_new_n13341__ = ~new_new_n12998__ & ~new_new_n13340__;
  assign new_new_n13342__ = ~new_new_n12997__ & ~new_new_n13341__;
  assign new_new_n13343__ = ~new_new_n12989__ & ~new_new_n13342__;
  assign new_new_n13344__ = ~new_new_n12988__ & ~new_new_n13343__;
  assign new_new_n13345__ = ~new_new_n12980__ & new_new_n13344__;
  assign new_new_n13346__ = ~new_new_n12979__ & ~new_new_n13345__;
  assign new_new_n13347__ = ~new_new_n12971__ & new_new_n13346__;
  assign new_new_n13348__ = ~new_new_n12970__ & ~new_new_n13347__;
  assign new_new_n13349__ = ~new_new_n12962__ & ~new_new_n13348__;
  assign new_new_n13350__ = ~new_new_n12961__ & ~new_new_n13349__;
  assign new_new_n13351__ = ~new_new_n12953__ & ~new_new_n13350__;
  assign new_new_n13352__ = ~new_new_n12952__ & ~new_new_n13351__;
  assign new_new_n13353__ = ~new_new_n12944__ & ~new_new_n13352__;
  assign new_new_n13354__ = ~new_new_n12943__ & ~new_new_n13353__;
  assign new_new_n13355__ = ~new_new_n12935__ & ~new_new_n13354__;
  assign new_new_n13356__ = ~new_new_n12934__ & ~new_new_n13355__;
  assign new_new_n13357__ = ~new_new_n12926__ & ~new_new_n13356__;
  assign new_new_n13358__ = ~new_new_n12925__ & ~new_new_n13357__;
  assign new_new_n13359__ = ~new_new_n12917__ & ~new_new_n13358__;
  assign new_new_n13360__ = ~new_new_n12916__ & ~new_new_n13359__;
  assign new_new_n13361__ = pi104 & new_new_n13360__;
  assign new_new_n13362__ = ~pi104 & ~new_new_n13360__;
  assign new_new_n13363__ = ~new_new_n12390__ & ~new_new_n12391__;
  assign new_new_n13364__ = pi103 & ~po017;
  assign new_new_n13365__ = ~new_new_n12826__ & po017;
  assign new_new_n13366__ = ~new_new_n13364__ & ~new_new_n13365__;
  assign new_new_n13367__ = new_new_n13363__ & ~new_new_n13366__;
  assign new_new_n13368__ = ~new_new_n13363__ & new_new_n13366__;
  assign new_new_n13369__ = ~new_new_n13367__ & ~new_new_n13368__;
  assign new_new_n13370__ = ~new_new_n13362__ & new_new_n13369__;
  assign new_new_n13371__ = ~new_new_n13361__ & ~new_new_n13370__;
  assign new_new_n13372__ = ~new_new_n12908__ & ~new_new_n13371__;
  assign new_new_n13373__ = ~new_new_n12907__ & ~new_new_n13372__;
  assign new_new_n13374__ = ~new_new_n12899__ & ~new_new_n13373__;
  assign new_new_n13375__ = ~new_new_n12898__ & ~new_new_n13374__;
  assign new_new_n13376__ = ~new_new_n12890__ & ~new_new_n13375__;
  assign new_new_n13377__ = ~new_new_n12889__ & ~new_new_n13376__;
  assign new_new_n13378__ = ~new_new_n12881__ & ~new_new_n13377__;
  assign new_new_n13379__ = ~new_new_n12880__ & ~new_new_n13378__;
  assign new_new_n13380__ = ~new_new_n12872__ & ~new_new_n13379__;
  assign new_new_n13381__ = ~new_new_n12871__ & ~new_new_n13380__;
  assign new_new_n13382__ = ~new_new_n12870__ & new_new_n13381__;
  assign new_new_n13383__ = ~new_new_n12869__ & ~new_new_n13382__;
  assign new_new_n13384__ = ~new_new_n12861__ & new_new_n13383__;
  assign po016 = new_new_n12860__ & ~new_new_n13384__;
  assign new_new_n13386__ = pi109 & ~new_new_n13379__;
  assign new_new_n13387__ = ~pi109 & new_new_n13379__;
  assign new_new_n13388__ = ~new_new_n13386__ & ~new_new_n13387__;
  assign new_new_n13389__ = po016 & new_new_n13388__;
  assign new_new_n13390__ = new_new_n12858__ & new_new_n13389__;
  assign new_new_n13391__ = ~new_new_n12858__ & ~new_new_n13389__;
  assign new_new_n13392__ = ~new_new_n13390__ & ~new_new_n13391__;
  assign new_new_n13393__ = ~pi110 & new_new_n13392__;
  assign new_new_n13394__ = pi110 & ~new_new_n13392__;
  assign new_new_n13395__ = ~new_new_n12880__ & ~new_new_n12881__;
  assign new_new_n13396__ = ~new_new_n13377__ & po016;
  assign new_new_n13397__ = pi108 & ~po016;
  assign new_new_n13398__ = ~new_new_n13396__ & ~new_new_n13397__;
  assign new_new_n13399__ = new_new_n13395__ & ~new_new_n13398__;
  assign new_new_n13400__ = ~new_new_n13395__ & new_new_n13398__;
  assign new_new_n13401__ = ~new_new_n13399__ & ~new_new_n13400__;
  assign new_new_n13402__ = ~pi109 & ~new_new_n13401__;
  assign new_new_n13403__ = pi109 & new_new_n13401__;
  assign new_new_n13404__ = ~new_new_n12889__ & ~new_new_n12890__;
  assign new_new_n13405__ = ~new_new_n13375__ & po016;
  assign new_new_n13406__ = pi107 & ~po016;
  assign new_new_n13407__ = ~new_new_n13405__ & ~new_new_n13406__;
  assign new_new_n13408__ = new_new_n13404__ & ~new_new_n13407__;
  assign new_new_n13409__ = ~new_new_n13404__ & new_new_n13407__;
  assign new_new_n13410__ = ~new_new_n13408__ & ~new_new_n13409__;
  assign new_new_n13411__ = ~pi108 & ~new_new_n13410__;
  assign new_new_n13412__ = pi108 & new_new_n13410__;
  assign new_new_n13413__ = ~new_new_n13373__ & po016;
  assign new_new_n13414__ = pi106 & ~po016;
  assign new_new_n13415__ = ~new_new_n13413__ & ~new_new_n13414__;
  assign new_new_n13416__ = ~new_new_n12898__ & ~new_new_n12899__;
  assign new_new_n13417__ = ~new_new_n13415__ & new_new_n13416__;
  assign new_new_n13418__ = new_new_n13415__ & ~new_new_n13416__;
  assign new_new_n13419__ = ~new_new_n13417__ & ~new_new_n13418__;
  assign new_new_n13420__ = ~pi107 & ~new_new_n13419__;
  assign new_new_n13421__ = pi107 & new_new_n13419__;
  assign new_new_n13422__ = ~new_new_n12907__ & ~new_new_n12908__;
  assign new_new_n13423__ = ~new_new_n13371__ & po016;
  assign new_new_n13424__ = pi105 & ~po016;
  assign new_new_n13425__ = ~new_new_n13423__ & ~new_new_n13424__;
  assign new_new_n13426__ = new_new_n13422__ & ~new_new_n13425__;
  assign new_new_n13427__ = ~new_new_n13422__ & new_new_n13425__;
  assign new_new_n13428__ = ~new_new_n13426__ & ~new_new_n13427__;
  assign new_new_n13429__ = ~pi106 & ~new_new_n13428__;
  assign new_new_n13430__ = pi106 & new_new_n13428__;
  assign new_new_n13431__ = ~new_new_n13361__ & ~new_new_n13362__;
  assign new_new_n13432__ = po016 & new_new_n13431__;
  assign new_new_n13433__ = ~new_new_n13369__ & ~new_new_n13432__;
  assign new_new_n13434__ = new_new_n13369__ & new_new_n13432__;
  assign new_new_n13435__ = ~new_new_n13433__ & ~new_new_n13434__;
  assign new_new_n13436__ = pi105 & new_new_n13435__;
  assign new_new_n13437__ = ~pi105 & ~new_new_n13435__;
  assign new_new_n13438__ = ~new_new_n12916__ & ~new_new_n12917__;
  assign new_new_n13439__ = ~new_new_n13358__ & po016;
  assign new_new_n13440__ = ~pi103 & ~po016;
  assign new_new_n13441__ = ~new_new_n13439__ & ~new_new_n13440__;
  assign new_new_n13442__ = new_new_n13438__ & ~new_new_n13441__;
  assign new_new_n13443__ = ~new_new_n13438__ & new_new_n13441__;
  assign new_new_n13444__ = ~new_new_n13442__ & ~new_new_n13443__;
  assign new_new_n13445__ = pi104 & ~new_new_n13444__;
  assign new_new_n13446__ = ~pi104 & new_new_n13444__;
  assign new_new_n13447__ = ~pi102 & ~new_new_n13356__;
  assign new_new_n13448__ = pi102 & new_new_n13356__;
  assign new_new_n13449__ = ~new_new_n13447__ & ~new_new_n13448__;
  assign new_new_n13450__ = po016 & new_new_n13449__;
  assign new_new_n13451__ = new_new_n12924__ & new_new_n13450__;
  assign new_new_n13452__ = ~new_new_n12924__ & ~new_new_n13450__;
  assign new_new_n13453__ = ~new_new_n13451__ & ~new_new_n13452__;
  assign new_new_n13454__ = pi103 & new_new_n13453__;
  assign new_new_n13455__ = ~pi103 & ~new_new_n13453__;
  assign new_new_n13456__ = ~new_new_n12934__ & ~new_new_n12935__;
  assign new_new_n13457__ = ~new_new_n13354__ & po016;
  assign new_new_n13458__ = ~pi101 & ~po016;
  assign new_new_n13459__ = ~new_new_n13457__ & ~new_new_n13458__;
  assign new_new_n13460__ = new_new_n13456__ & ~new_new_n13459__;
  assign new_new_n13461__ = ~new_new_n13456__ & new_new_n13459__;
  assign new_new_n13462__ = ~new_new_n13460__ & ~new_new_n13461__;
  assign new_new_n13463__ = pi102 & ~new_new_n13462__;
  assign new_new_n13464__ = ~pi102 & new_new_n13462__;
  assign new_new_n13465__ = ~new_new_n12943__ & ~new_new_n12944__;
  assign new_new_n13466__ = ~new_new_n13352__ & po016;
  assign new_new_n13467__ = ~pi100 & ~po016;
  assign new_new_n13468__ = ~new_new_n13466__ & ~new_new_n13467__;
  assign new_new_n13469__ = new_new_n13465__ & ~new_new_n13468__;
  assign new_new_n13470__ = ~new_new_n13465__ & new_new_n13468__;
  assign new_new_n13471__ = ~new_new_n13469__ & ~new_new_n13470__;
  assign new_new_n13472__ = pi101 & ~new_new_n13471__;
  assign new_new_n13473__ = ~pi101 & new_new_n13471__;
  assign new_new_n13474__ = ~new_new_n12952__ & ~new_new_n12953__;
  assign new_new_n13475__ = ~new_new_n13350__ & po016;
  assign new_new_n13476__ = ~pi099 & ~po016;
  assign new_new_n13477__ = ~new_new_n13475__ & ~new_new_n13476__;
  assign new_new_n13478__ = new_new_n13474__ & ~new_new_n13477__;
  assign new_new_n13479__ = ~new_new_n13474__ & new_new_n13477__;
  assign new_new_n13480__ = ~new_new_n13478__ & ~new_new_n13479__;
  assign new_new_n13481__ = ~pi100 & new_new_n13480__;
  assign new_new_n13482__ = pi100 & ~new_new_n13480__;
  assign new_new_n13483__ = ~pi098 & ~new_new_n13348__;
  assign new_new_n13484__ = pi098 & new_new_n13348__;
  assign new_new_n13485__ = ~new_new_n13483__ & ~new_new_n13484__;
  assign new_new_n13486__ = po016 & new_new_n13485__;
  assign new_new_n13487__ = new_new_n12960__ & new_new_n13486__;
  assign new_new_n13488__ = ~new_new_n12960__ & ~new_new_n13486__;
  assign new_new_n13489__ = ~new_new_n13487__ & ~new_new_n13488__;
  assign new_new_n13490__ = ~pi099 & ~new_new_n13489__;
  assign new_new_n13491__ = pi099 & new_new_n13489__;
  assign new_new_n13492__ = ~new_new_n12970__ & ~new_new_n12971__;
  assign new_new_n13493__ = ~new_new_n13346__ & po016;
  assign new_new_n13494__ = pi097 & ~po016;
  assign new_new_n13495__ = ~new_new_n13493__ & ~new_new_n13494__;
  assign new_new_n13496__ = new_new_n13492__ & ~new_new_n13495__;
  assign new_new_n13497__ = ~new_new_n13492__ & new_new_n13495__;
  assign new_new_n13498__ = ~new_new_n13496__ & ~new_new_n13497__;
  assign new_new_n13499__ = ~pi098 & ~new_new_n13498__;
  assign new_new_n13500__ = pi098 & new_new_n13498__;
  assign new_new_n13501__ = new_new_n13344__ & po016;
  assign new_new_n13502__ = pi096 & ~po016;
  assign new_new_n13503__ = ~new_new_n13501__ & ~new_new_n13502__;
  assign new_new_n13504__ = ~new_new_n12979__ & ~new_new_n12980__;
  assign new_new_n13505__ = ~new_new_n13503__ & ~new_new_n13504__;
  assign new_new_n13506__ = new_new_n13503__ & new_new_n13504__;
  assign new_new_n13507__ = ~new_new_n13505__ & ~new_new_n13506__;
  assign new_new_n13508__ = pi097 & ~new_new_n13507__;
  assign new_new_n13509__ = ~pi097 & new_new_n13507__;
  assign new_new_n13510__ = ~pi095 & ~new_new_n13342__;
  assign new_new_n13511__ = pi095 & new_new_n13342__;
  assign new_new_n13512__ = ~new_new_n13510__ & ~new_new_n13511__;
  assign new_new_n13513__ = po016 & new_new_n13512__;
  assign new_new_n13514__ = new_new_n12987__ & new_new_n13513__;
  assign new_new_n13515__ = ~new_new_n12987__ & ~new_new_n13513__;
  assign new_new_n13516__ = ~new_new_n13514__ & ~new_new_n13515__;
  assign new_new_n13517__ = ~pi096 & ~new_new_n13516__;
  assign new_new_n13518__ = pi096 & new_new_n13516__;
  assign new_new_n13519__ = ~new_new_n12997__ & ~new_new_n12998__;
  assign new_new_n13520__ = ~new_new_n13340__ & po016;
  assign new_new_n13521__ = ~pi094 & ~po016;
  assign new_new_n13522__ = ~new_new_n13520__ & ~new_new_n13521__;
  assign new_new_n13523__ = new_new_n13519__ & ~new_new_n13522__;
  assign new_new_n13524__ = ~new_new_n13519__ & new_new_n13522__;
  assign new_new_n13525__ = ~new_new_n13523__ & ~new_new_n13524__;
  assign new_new_n13526__ = ~pi095 & new_new_n13525__;
  assign new_new_n13527__ = pi095 & ~new_new_n13525__;
  assign new_new_n13528__ = ~pi093 & ~new_new_n13338__;
  assign new_new_n13529__ = pi093 & new_new_n13338__;
  assign new_new_n13530__ = ~new_new_n13528__ & ~new_new_n13529__;
  assign new_new_n13531__ = po016 & new_new_n13530__;
  assign new_new_n13532__ = new_new_n13005__ & new_new_n13531__;
  assign new_new_n13533__ = ~new_new_n13005__ & ~new_new_n13531__;
  assign new_new_n13534__ = ~new_new_n13532__ & ~new_new_n13533__;
  assign new_new_n13535__ = ~pi094 & ~new_new_n13534__;
  assign new_new_n13536__ = pi094 & new_new_n13534__;
  assign new_new_n13537__ = ~new_new_n13015__ & ~new_new_n13016__;
  assign new_new_n13538__ = ~new_new_n13336__ & po016;
  assign new_new_n13539__ = ~pi092 & ~po016;
  assign new_new_n13540__ = ~new_new_n13538__ & ~new_new_n13539__;
  assign new_new_n13541__ = ~new_new_n13537__ & ~new_new_n13540__;
  assign new_new_n13542__ = new_new_n13537__ & new_new_n13540__;
  assign new_new_n13543__ = ~new_new_n13541__ & ~new_new_n13542__;
  assign new_new_n13544__ = ~pi093 & ~new_new_n13543__;
  assign new_new_n13545__ = pi093 & new_new_n13543__;
  assign new_new_n13546__ = new_new_n13334__ & po016;
  assign new_new_n13547__ = ~pi091 & ~po016;
  assign new_new_n13548__ = ~new_new_n13546__ & ~new_new_n13547__;
  assign new_new_n13549__ = ~new_new_n13024__ & ~new_new_n13025__;
  assign new_new_n13550__ = ~new_new_n13548__ & ~new_new_n13549__;
  assign new_new_n13551__ = new_new_n13548__ & new_new_n13549__;
  assign new_new_n13552__ = ~new_new_n13550__ & ~new_new_n13551__;
  assign new_new_n13553__ = ~pi092 & ~new_new_n13552__;
  assign new_new_n13554__ = pi092 & new_new_n13552__;
  assign new_new_n13555__ = ~new_new_n13033__ & ~new_new_n13034__;
  assign new_new_n13556__ = ~new_new_n13332__ & po016;
  assign new_new_n13557__ = ~pi090 & ~po016;
  assign new_new_n13558__ = ~new_new_n13556__ & ~new_new_n13557__;
  assign new_new_n13559__ = new_new_n13555__ & ~new_new_n13558__;
  assign new_new_n13560__ = ~new_new_n13555__ & new_new_n13558__;
  assign new_new_n13561__ = ~new_new_n13559__ & ~new_new_n13560__;
  assign new_new_n13562__ = pi091 & ~new_new_n13561__;
  assign new_new_n13563__ = ~pi091 & new_new_n13561__;
  assign new_new_n13564__ = ~pi089 & ~new_new_n13330__;
  assign new_new_n13565__ = pi089 & new_new_n13330__;
  assign new_new_n13566__ = ~new_new_n13564__ & ~new_new_n13565__;
  assign new_new_n13567__ = po016 & new_new_n13566__;
  assign new_new_n13568__ = new_new_n13041__ & new_new_n13567__;
  assign new_new_n13569__ = ~new_new_n13041__ & ~new_new_n13567__;
  assign new_new_n13570__ = ~new_new_n13568__ & ~new_new_n13569__;
  assign new_new_n13571__ = ~pi090 & ~new_new_n13570__;
  assign new_new_n13572__ = pi090 & new_new_n13570__;
  assign new_new_n13573__ = ~new_new_n13328__ & po016;
  assign new_new_n13574__ = pi088 & ~po016;
  assign new_new_n13575__ = ~new_new_n13573__ & ~new_new_n13574__;
  assign new_new_n13576__ = ~new_new_n13051__ & ~new_new_n13052__;
  assign new_new_n13577__ = new_new_n13575__ & new_new_n13576__;
  assign new_new_n13578__ = ~new_new_n13575__ & ~new_new_n13576__;
  assign new_new_n13579__ = ~new_new_n13577__ & ~new_new_n13578__;
  assign new_new_n13580__ = pi089 & ~new_new_n13579__;
  assign new_new_n13581__ = ~pi089 & new_new_n13579__;
  assign new_new_n13582__ = ~new_new_n13060__ & ~new_new_n13061__;
  assign new_new_n13583__ = pi087 & ~po016;
  assign new_new_n13584__ = ~new_new_n13326__ & po016;
  assign new_new_n13585__ = ~new_new_n13583__ & ~new_new_n13584__;
  assign new_new_n13586__ = new_new_n13582__ & new_new_n13585__;
  assign new_new_n13587__ = ~new_new_n13582__ & ~new_new_n13585__;
  assign new_new_n13588__ = ~new_new_n13586__ & ~new_new_n13587__;
  assign new_new_n13589__ = pi088 & ~new_new_n13588__;
  assign new_new_n13590__ = ~pi088 & new_new_n13588__;
  assign new_new_n13591__ = ~new_new_n13069__ & ~new_new_n13070__;
  assign new_new_n13592__ = ~new_new_n13324__ & po016;
  assign new_new_n13593__ = pi086 & ~po016;
  assign new_new_n13594__ = ~new_new_n13592__ & ~new_new_n13593__;
  assign new_new_n13595__ = new_new_n13591__ & new_new_n13594__;
  assign new_new_n13596__ = ~new_new_n13591__ & ~new_new_n13594__;
  assign new_new_n13597__ = ~new_new_n13595__ & ~new_new_n13596__;
  assign new_new_n13598__ = pi087 & ~new_new_n13597__;
  assign new_new_n13599__ = ~pi087 & new_new_n13597__;
  assign new_new_n13600__ = new_new_n13322__ & po016;
  assign new_new_n13601__ = ~pi085 & ~po016;
  assign new_new_n13602__ = ~new_new_n13600__ & ~new_new_n13601__;
  assign new_new_n13603__ = ~new_new_n13078__ & ~new_new_n13079__;
  assign new_new_n13604__ = ~new_new_n13602__ & ~new_new_n13603__;
  assign new_new_n13605__ = new_new_n13602__ & new_new_n13603__;
  assign new_new_n13606__ = ~new_new_n13604__ & ~new_new_n13605__;
  assign new_new_n13607__ = ~pi086 & ~new_new_n13606__;
  assign new_new_n13608__ = pi086 & new_new_n13606__;
  assign new_new_n13609__ = new_new_n13320__ & po016;
  assign new_new_n13610__ = ~pi084 & ~po016;
  assign new_new_n13611__ = ~new_new_n13609__ & ~new_new_n13610__;
  assign new_new_n13612__ = ~new_new_n13087__ & ~new_new_n13088__;
  assign new_new_n13613__ = ~new_new_n13611__ & ~new_new_n13612__;
  assign new_new_n13614__ = new_new_n13611__ & new_new_n13612__;
  assign new_new_n13615__ = ~new_new_n13613__ & ~new_new_n13614__;
  assign new_new_n13616__ = pi085 & new_new_n13615__;
  assign new_new_n13617__ = ~pi085 & ~new_new_n13615__;
  assign new_new_n13618__ = ~new_new_n13096__ & ~new_new_n13097__;
  assign new_new_n13619__ = ~new_new_n13318__ & po016;
  assign new_new_n13620__ = pi083 & ~po016;
  assign new_new_n13621__ = ~new_new_n13619__ & ~new_new_n13620__;
  assign new_new_n13622__ = new_new_n13618__ & new_new_n13621__;
  assign new_new_n13623__ = ~new_new_n13618__ & ~new_new_n13621__;
  assign new_new_n13624__ = ~new_new_n13622__ & ~new_new_n13623__;
  assign new_new_n13625__ = pi084 & ~new_new_n13624__;
  assign new_new_n13626__ = ~pi084 & new_new_n13624__;
  assign new_new_n13627__ = pi082 & ~new_new_n13316__;
  assign new_new_n13628__ = ~pi082 & new_new_n13316__;
  assign new_new_n13629__ = ~new_new_n13627__ & ~new_new_n13628__;
  assign new_new_n13630__ = po016 & new_new_n13629__;
  assign new_new_n13631__ = new_new_n13104__ & new_new_n13630__;
  assign new_new_n13632__ = ~new_new_n13104__ & ~new_new_n13630__;
  assign new_new_n13633__ = ~new_new_n13631__ & ~new_new_n13632__;
  assign new_new_n13634__ = pi083 & ~new_new_n13633__;
  assign new_new_n13635__ = pi081 & ~new_new_n13314__;
  assign new_new_n13636__ = ~pi081 & new_new_n13314__;
  assign new_new_n13637__ = ~new_new_n13635__ & ~new_new_n13636__;
  assign new_new_n13638__ = po016 & new_new_n13637__;
  assign new_new_n13639__ = new_new_n13113__ & new_new_n13638__;
  assign new_new_n13640__ = ~new_new_n13113__ & ~new_new_n13638__;
  assign new_new_n13641__ = ~new_new_n13639__ & ~new_new_n13640__;
  assign new_new_n13642__ = pi082 & ~new_new_n13641__;
  assign new_new_n13643__ = ~pi082 & new_new_n13641__;
  assign new_new_n13644__ = ~new_new_n13312__ & po016;
  assign new_new_n13645__ = pi080 & ~po016;
  assign new_new_n13646__ = ~new_new_n13644__ & ~new_new_n13645__;
  assign new_new_n13647__ = ~new_new_n13123__ & ~new_new_n13124__;
  assign new_new_n13648__ = ~new_new_n13646__ & new_new_n13647__;
  assign new_new_n13649__ = new_new_n13646__ & ~new_new_n13647__;
  assign new_new_n13650__ = ~new_new_n13648__ & ~new_new_n13649__;
  assign new_new_n13651__ = pi081 & new_new_n13650__;
  assign new_new_n13652__ = ~pi081 & ~new_new_n13650__;
  assign new_new_n13653__ = ~pi079 & ~new_new_n13310__;
  assign new_new_n13654__ = pi079 & new_new_n13310__;
  assign new_new_n13655__ = ~new_new_n13653__ & ~new_new_n13654__;
  assign new_new_n13656__ = po016 & ~new_new_n13655__;
  assign new_new_n13657__ = new_new_n13131__ & new_new_n13656__;
  assign new_new_n13658__ = ~new_new_n13131__ & ~new_new_n13656__;
  assign new_new_n13659__ = ~new_new_n13657__ & ~new_new_n13658__;
  assign new_new_n13660__ = pi080 & ~new_new_n13659__;
  assign new_new_n13661__ = ~pi080 & new_new_n13659__;
  assign new_new_n13662__ = ~new_new_n13141__ & ~new_new_n13142__;
  assign new_new_n13663__ = ~new_new_n13308__ & po016;
  assign new_new_n13664__ = pi078 & ~po016;
  assign new_new_n13665__ = ~new_new_n13663__ & ~new_new_n13664__;
  assign new_new_n13666__ = new_new_n13662__ & new_new_n13665__;
  assign new_new_n13667__ = ~new_new_n13662__ & ~new_new_n13665__;
  assign new_new_n13668__ = ~new_new_n13666__ & ~new_new_n13667__;
  assign new_new_n13669__ = pi079 & ~new_new_n13668__;
  assign new_new_n13670__ = ~pi079 & new_new_n13668__;
  assign new_new_n13671__ = pi077 & ~new_new_n13306__;
  assign new_new_n13672__ = ~pi077 & new_new_n13306__;
  assign new_new_n13673__ = ~new_new_n13671__ & ~new_new_n13672__;
  assign new_new_n13674__ = po016 & new_new_n13673__;
  assign new_new_n13675__ = ~new_new_n13149__ & ~new_new_n13674__;
  assign new_new_n13676__ = new_new_n13149__ & new_new_n13674__;
  assign new_new_n13677__ = ~new_new_n13675__ & ~new_new_n13676__;
  assign new_new_n13678__ = pi078 & ~new_new_n13677__;
  assign new_new_n13679__ = ~pi078 & new_new_n13677__;
  assign new_new_n13680__ = ~new_new_n13159__ & ~new_new_n13160__;
  assign new_new_n13681__ = ~new_new_n13304__ & po016;
  assign new_new_n13682__ = ~pi076 & ~po016;
  assign new_new_n13683__ = ~new_new_n13681__ & ~new_new_n13682__;
  assign new_new_n13684__ = new_new_n13680__ & ~new_new_n13683__;
  assign new_new_n13685__ = ~new_new_n13680__ & new_new_n13683__;
  assign new_new_n13686__ = ~new_new_n13684__ & ~new_new_n13685__;
  assign new_new_n13687__ = ~pi077 & new_new_n13686__;
  assign new_new_n13688__ = pi077 & ~new_new_n13686__;
  assign new_new_n13689__ = ~pi075 & ~new_new_n13302__;
  assign new_new_n13690__ = pi075 & new_new_n13302__;
  assign new_new_n13691__ = ~new_new_n13689__ & ~new_new_n13690__;
  assign new_new_n13692__ = po016 & new_new_n13691__;
  assign new_new_n13693__ = new_new_n13167__ & new_new_n13692__;
  assign new_new_n13694__ = ~new_new_n13167__ & ~new_new_n13692__;
  assign new_new_n13695__ = ~new_new_n13693__ & ~new_new_n13694__;
  assign new_new_n13696__ = ~pi076 & ~new_new_n13695__;
  assign new_new_n13697__ = pi076 & new_new_n13695__;
  assign new_new_n13698__ = ~new_new_n13177__ & ~new_new_n13178__;
  assign new_new_n13699__ = ~new_new_n13300__ & po016;
  assign new_new_n13700__ = pi074 & ~po016;
  assign new_new_n13701__ = ~new_new_n13699__ & ~new_new_n13700__;
  assign new_new_n13702__ = new_new_n13698__ & ~new_new_n13701__;
  assign new_new_n13703__ = ~new_new_n13698__ & new_new_n13701__;
  assign new_new_n13704__ = ~new_new_n13702__ & ~new_new_n13703__;
  assign new_new_n13705__ = ~pi075 & ~new_new_n13704__;
  assign new_new_n13706__ = pi075 & new_new_n13704__;
  assign new_new_n13707__ = ~new_new_n13298__ & po016;
  assign new_new_n13708__ = pi073 & ~po016;
  assign new_new_n13709__ = ~new_new_n13707__ & ~new_new_n13708__;
  assign new_new_n13710__ = ~new_new_n13186__ & ~new_new_n13187__;
  assign new_new_n13711__ = ~new_new_n13709__ & new_new_n13710__;
  assign new_new_n13712__ = new_new_n13709__ & ~new_new_n13710__;
  assign new_new_n13713__ = ~new_new_n13711__ & ~new_new_n13712__;
  assign new_new_n13714__ = ~pi074 & ~new_new_n13713__;
  assign new_new_n13715__ = pi074 & new_new_n13713__;
  assign new_new_n13716__ = ~new_new_n13195__ & ~new_new_n13196__;
  assign new_new_n13717__ = ~new_new_n13296__ & po016;
  assign new_new_n13718__ = pi072 & ~po016;
  assign new_new_n13719__ = ~new_new_n13717__ & ~new_new_n13718__;
  assign new_new_n13720__ = new_new_n13716__ & ~new_new_n13719__;
  assign new_new_n13721__ = ~new_new_n13716__ & new_new_n13719__;
  assign new_new_n13722__ = ~new_new_n13720__ & ~new_new_n13721__;
  assign new_new_n13723__ = ~pi073 & ~new_new_n13722__;
  assign new_new_n13724__ = pi073 & new_new_n13722__;
  assign new_new_n13725__ = ~new_new_n13286__ & ~new_new_n13287__;
  assign new_new_n13726__ = po016 & new_new_n13725__;
  assign new_new_n13727__ = ~new_new_n13294__ & ~new_new_n13726__;
  assign new_new_n13728__ = new_new_n13294__ & new_new_n13726__;
  assign new_new_n13729__ = ~new_new_n13727__ & ~new_new_n13728__;
  assign new_new_n13730__ = pi072 & ~new_new_n13729__;
  assign new_new_n13731__ = ~pi072 & new_new_n13729__;
  assign new_new_n13732__ = ~new_new_n13204__ & ~new_new_n13205__;
  assign new_new_n13733__ = new_new_n13283__ & po016;
  assign new_new_n13734__ = ~pi070 & ~po016;
  assign new_new_n13735__ = ~new_new_n13733__ & ~new_new_n13734__;
  assign new_new_n13736__ = ~new_new_n13732__ & ~new_new_n13735__;
  assign new_new_n13737__ = new_new_n13732__ & new_new_n13735__;
  assign new_new_n13738__ = ~new_new_n13736__ & ~new_new_n13737__;
  assign new_new_n13739__ = pi071 & new_new_n13738__;
  assign new_new_n13740__ = ~pi071 & ~new_new_n13738__;
  assign new_new_n13741__ = ~new_new_n13213__ & ~new_new_n13214__;
  assign new_new_n13742__ = ~new_new_n13270__ & po016;
  assign new_new_n13743__ = ~pi068 & ~po016;
  assign new_new_n13744__ = ~new_new_n13742__ & ~new_new_n13743__;
  assign new_new_n13745__ = new_new_n13741__ & ~new_new_n13744__;
  assign new_new_n13746__ = ~new_new_n13741__ & new_new_n13744__;
  assign new_new_n13747__ = ~new_new_n13745__ & ~new_new_n13746__;
  assign new_new_n13748__ = pi069 & ~new_new_n13747__;
  assign new_new_n13749__ = ~pi069 & new_new_n13747__;
  assign new_new_n13750__ = ~new_new_n13227__ & ~new_new_n13228__;
  assign new_new_n13751__ = ~new_new_n13268__ & po016;
  assign new_new_n13752__ = ~pi067 & ~po016;
  assign new_new_n13753__ = ~new_new_n13751__ & ~new_new_n13752__;
  assign new_new_n13754__ = new_new_n13750__ & ~new_new_n13753__;
  assign new_new_n13755__ = ~new_new_n13750__ & new_new_n13753__;
  assign new_new_n13756__ = ~new_new_n13754__ & ~new_new_n13755__;
  assign new_new_n13757__ = ~pi068 & new_new_n13756__;
  assign new_new_n13758__ = pi068 & ~new_new_n13756__;
  assign new_new_n13759__ = ~new_new_n13229__ & new_new_n13230__;
  assign new_new_n13760__ = ~pi017 & ~po017;
  assign new_new_n13761__ = ~pi065 & ~new_new_n13760__;
  assign new_new_n13762__ = ~pi016 & ~new_new_n13761__;
  assign new_new_n13763__ = ~new_new_n13759__ & ~new_new_n13762__;
  assign new_new_n13764__ = pi064 & ~new_new_n13763__;
  assign new_new_n13765__ = ~new_new_n13244__ & ~new_new_n13764__;
  assign new_new_n13766__ = pi066 & ~new_new_n13765__;
  assign new_new_n13767__ = ~pi066 & new_new_n13765__;
  assign new_new_n13768__ = ~new_new_n13766__ & ~new_new_n13767__;
  assign new_new_n13769__ = po016 & new_new_n13768__;
  assign new_new_n13770__ = ~new_new_n12713__ & ~new_new_n13215__;
  assign new_new_n13771__ = po017 & new_new_n13770__;
  assign new_new_n13772__ = new_new_n13217__ & ~new_new_n13771__;
  assign new_new_n13773__ = ~new_new_n13217__ & new_new_n13771__;
  assign new_new_n13774__ = ~new_new_n13772__ & ~new_new_n13773__;
  assign new_new_n13775__ = new_new_n13769__ & new_new_n13774__;
  assign new_new_n13776__ = ~new_new_n13769__ & ~new_new_n13774__;
  assign new_new_n13777__ = ~new_new_n13775__ & ~new_new_n13776__;
  assign new_new_n13778__ = ~pi067 & ~new_new_n13777__;
  assign new_new_n13779__ = pi067 & new_new_n13777__;
  assign new_new_n13780__ = pi016 & po016;
  assign new_new_n13781__ = pi015 & ~new_new_n13780__;
  assign new_new_n13782__ = pi065 & ~new_new_n13781__;
  assign new_new_n13783__ = ~pi016 & po016;
  assign new_new_n13784__ = pi016 & ~po016;
  assign new_new_n13785__ = ~pi015 & ~new_new_n13783__;
  assign new_new_n13786__ = ~new_new_n13784__ & new_new_n13785__;
  assign new_new_n13787__ = ~new_new_n13782__ & ~new_new_n13786__;
  assign new_new_n13788__ = pi064 & ~new_new_n13787__;
  assign new_new_n13789__ = pi064 & po016;
  assign new_new_n13790__ = new_new_n13250__ & ~new_new_n13789__;
  assign new_new_n13791__ = ~new_new_n13788__ & ~new_new_n13790__;
  assign new_new_n13792__ = pi066 & ~new_new_n13791__;
  assign new_new_n13793__ = ~pi066 & new_new_n13791__;
  assign new_new_n13794__ = ~new_new_n332__ & po016;
  assign new_new_n13795__ = ~new_new_n13243__ & ~new_new_n13794__;
  assign new_new_n13796__ = ~new_new_n13257__ & ~new_new_n13259__;
  assign new_new_n13797__ = ~pi065 & ~po016;
  assign new_new_n13798__ = ~pi016 & ~new_new_n403__;
  assign new_new_n13799__ = new_new_n13796__ & new_new_n13798__;
  assign new_new_n13800__ = ~new_new_n13797__ & new_new_n13799__;
  assign new_new_n13801__ = pi065 & ~new_new_n13789__;
  assign new_new_n13802__ = pi016 & ~new_new_n13796__;
  assign new_new_n13803__ = ~new_new_n13801__ & new_new_n13802__;
  assign new_new_n13804__ = ~new_new_n13795__ & ~new_new_n13800__;
  assign new_new_n13805__ = ~new_new_n13803__ & new_new_n13804__;
  assign new_new_n13806__ = ~pi017 & ~new_new_n13805__;
  assign new_new_n13807__ = pi065 & po016;
  assign new_new_n13808__ = ~new_new_n13243__ & ~new_new_n13807__;
  assign new_new_n13809__ = pi064 & ~new_new_n13258__;
  assign new_new_n13810__ = ~new_new_n13808__ & ~new_new_n13809__;
  assign new_new_n13811__ = ~new_new_n13250__ & po016;
  assign new_new_n13812__ = po017 & ~new_new_n13811__;
  assign new_new_n13813__ = new_new_n13259__ & new_new_n13783__;
  assign new_new_n13814__ = ~new_new_n13812__ & ~new_new_n13813__;
  assign new_new_n13815__ = pi064 & ~new_new_n13814__;
  assign new_new_n13816__ = ~new_new_n13810__ & ~new_new_n13815__;
  assign new_new_n13817__ = pi017 & ~new_new_n13816__;
  assign new_new_n13818__ = ~new_new_n13806__ & ~new_new_n13817__;
  assign new_new_n13819__ = ~new_new_n13793__ & ~new_new_n13818__;
  assign new_new_n13820__ = ~new_new_n13792__ & ~new_new_n13819__;
  assign new_new_n13821__ = ~new_new_n13779__ & new_new_n13820__;
  assign new_new_n13822__ = ~new_new_n13778__ & ~new_new_n13821__;
  assign new_new_n13823__ = ~new_new_n13758__ & ~new_new_n13822__;
  assign new_new_n13824__ = ~new_new_n13757__ & ~new_new_n13823__;
  assign new_new_n13825__ = ~new_new_n13749__ & new_new_n13824__;
  assign new_new_n13826__ = ~new_new_n13748__ & ~new_new_n13825__;
  assign new_new_n13827__ = pi070 & ~new_new_n13826__;
  assign new_new_n13828__ = ~pi070 & new_new_n13826__;
  assign new_new_n13829__ = ~new_new_n13273__ & ~new_new_n13274__;
  assign new_new_n13830__ = po016 & new_new_n13829__;
  assign new_new_n13831__ = ~new_new_n13281__ & ~new_new_n13830__;
  assign new_new_n13832__ = new_new_n13281__ & new_new_n13830__;
  assign new_new_n13833__ = ~new_new_n13831__ & ~new_new_n13832__;
  assign new_new_n13834__ = ~new_new_n13828__ & ~new_new_n13833__;
  assign new_new_n13835__ = ~new_new_n13827__ & ~new_new_n13834__;
  assign new_new_n13836__ = ~new_new_n13740__ & ~new_new_n13835__;
  assign new_new_n13837__ = ~new_new_n13739__ & ~new_new_n13836__;
  assign new_new_n13838__ = ~new_new_n13731__ & ~new_new_n13837__;
  assign new_new_n13839__ = ~new_new_n13730__ & ~new_new_n13838__;
  assign new_new_n13840__ = ~new_new_n13724__ & new_new_n13839__;
  assign new_new_n13841__ = ~new_new_n13723__ & ~new_new_n13840__;
  assign new_new_n13842__ = ~new_new_n13715__ & ~new_new_n13841__;
  assign new_new_n13843__ = ~new_new_n13714__ & ~new_new_n13842__;
  assign new_new_n13844__ = ~new_new_n13706__ & ~new_new_n13843__;
  assign new_new_n13845__ = ~new_new_n13705__ & ~new_new_n13844__;
  assign new_new_n13846__ = ~new_new_n13697__ & ~new_new_n13845__;
  assign new_new_n13847__ = ~new_new_n13696__ & ~new_new_n13846__;
  assign new_new_n13848__ = ~new_new_n13688__ & ~new_new_n13847__;
  assign new_new_n13849__ = ~new_new_n13687__ & ~new_new_n13848__;
  assign new_new_n13850__ = ~new_new_n13679__ & new_new_n13849__;
  assign new_new_n13851__ = ~new_new_n13678__ & ~new_new_n13850__;
  assign new_new_n13852__ = ~new_new_n13670__ & ~new_new_n13851__;
  assign new_new_n13853__ = ~new_new_n13669__ & ~new_new_n13852__;
  assign new_new_n13854__ = ~new_new_n13661__ & ~new_new_n13853__;
  assign new_new_n13855__ = ~new_new_n13660__ & ~new_new_n13854__;
  assign new_new_n13856__ = ~new_new_n13652__ & ~new_new_n13855__;
  assign new_new_n13857__ = ~new_new_n13651__ & ~new_new_n13856__;
  assign new_new_n13858__ = ~new_new_n13643__ & ~new_new_n13857__;
  assign new_new_n13859__ = ~new_new_n13642__ & ~new_new_n13858__;
  assign new_new_n13860__ = ~pi083 & new_new_n13633__;
  assign new_new_n13861__ = ~new_new_n13859__ & ~new_new_n13860__;
  assign new_new_n13862__ = ~new_new_n13634__ & ~new_new_n13861__;
  assign new_new_n13863__ = ~new_new_n13626__ & ~new_new_n13862__;
  assign new_new_n13864__ = ~new_new_n13625__ & ~new_new_n13863__;
  assign new_new_n13865__ = ~new_new_n13617__ & ~new_new_n13864__;
  assign new_new_n13866__ = ~new_new_n13616__ & ~new_new_n13865__;
  assign new_new_n13867__ = ~new_new_n13608__ & new_new_n13866__;
  assign new_new_n13868__ = ~new_new_n13607__ & ~new_new_n13867__;
  assign new_new_n13869__ = ~new_new_n13599__ & new_new_n13868__;
  assign new_new_n13870__ = ~new_new_n13598__ & ~new_new_n13869__;
  assign new_new_n13871__ = ~new_new_n13590__ & ~new_new_n13870__;
  assign new_new_n13872__ = ~new_new_n13589__ & ~new_new_n13871__;
  assign new_new_n13873__ = ~new_new_n13581__ & ~new_new_n13872__;
  assign new_new_n13874__ = ~new_new_n13580__ & ~new_new_n13873__;
  assign new_new_n13875__ = ~new_new_n13572__ & new_new_n13874__;
  assign new_new_n13876__ = ~new_new_n13571__ & ~new_new_n13875__;
  assign new_new_n13877__ = ~new_new_n13563__ & new_new_n13876__;
  assign new_new_n13878__ = ~new_new_n13562__ & ~new_new_n13877__;
  assign new_new_n13879__ = ~new_new_n13554__ & new_new_n13878__;
  assign new_new_n13880__ = ~new_new_n13553__ & ~new_new_n13879__;
  assign new_new_n13881__ = ~new_new_n13545__ & ~new_new_n13880__;
  assign new_new_n13882__ = ~new_new_n13544__ & ~new_new_n13881__;
  assign new_new_n13883__ = ~new_new_n13536__ & ~new_new_n13882__;
  assign new_new_n13884__ = ~new_new_n13535__ & ~new_new_n13883__;
  assign new_new_n13885__ = ~new_new_n13527__ & ~new_new_n13884__;
  assign new_new_n13886__ = ~new_new_n13526__ & ~new_new_n13885__;
  assign new_new_n13887__ = ~new_new_n13518__ & ~new_new_n13886__;
  assign new_new_n13888__ = ~new_new_n13517__ & ~new_new_n13887__;
  assign new_new_n13889__ = ~new_new_n13509__ & new_new_n13888__;
  assign new_new_n13890__ = ~new_new_n13508__ & ~new_new_n13889__;
  assign new_new_n13891__ = ~new_new_n13500__ & new_new_n13890__;
  assign new_new_n13892__ = ~new_new_n13499__ & ~new_new_n13891__;
  assign new_new_n13893__ = ~new_new_n13491__ & ~new_new_n13892__;
  assign new_new_n13894__ = ~new_new_n13490__ & ~new_new_n13893__;
  assign new_new_n13895__ = ~new_new_n13482__ & ~new_new_n13894__;
  assign new_new_n13896__ = ~new_new_n13481__ & ~new_new_n13895__;
  assign new_new_n13897__ = ~new_new_n13473__ & new_new_n13896__;
  assign new_new_n13898__ = ~new_new_n13472__ & ~new_new_n13897__;
  assign new_new_n13899__ = ~new_new_n13464__ & ~new_new_n13898__;
  assign new_new_n13900__ = ~new_new_n13463__ & ~new_new_n13899__;
  assign new_new_n13901__ = ~new_new_n13455__ & ~new_new_n13900__;
  assign new_new_n13902__ = ~new_new_n13454__ & ~new_new_n13901__;
  assign new_new_n13903__ = ~new_new_n13446__ & ~new_new_n13902__;
  assign new_new_n13904__ = ~new_new_n13445__ & ~new_new_n13903__;
  assign new_new_n13905__ = ~new_new_n13437__ & ~new_new_n13904__;
  assign new_new_n13906__ = ~new_new_n13436__ & ~new_new_n13905__;
  assign new_new_n13907__ = ~new_new_n13430__ & new_new_n13906__;
  assign new_new_n13908__ = ~new_new_n13429__ & ~new_new_n13907__;
  assign new_new_n13909__ = ~new_new_n13421__ & ~new_new_n13908__;
  assign new_new_n13910__ = ~new_new_n13420__ & ~new_new_n13909__;
  assign new_new_n13911__ = ~new_new_n13412__ & ~new_new_n13910__;
  assign new_new_n13912__ = ~new_new_n13411__ & ~new_new_n13911__;
  assign new_new_n13913__ = ~new_new_n13403__ & ~new_new_n13912__;
  assign new_new_n13914__ = ~new_new_n13402__ & ~new_new_n13913__;
  assign new_new_n13915__ = ~new_new_n13394__ & ~new_new_n13914__;
  assign new_new_n13916__ = ~new_new_n13393__ & ~new_new_n13915__;
  assign new_new_n13917__ = ~pi111 & ~new_new_n13916__;
  assign new_new_n13918__ = pi111 & new_new_n13916__;
  assign new_new_n13919__ = ~pi110 & ~new_new_n13381__;
  assign new_new_n13920__ = pi110 & new_new_n13381__;
  assign new_new_n13921__ = ~new_new_n13919__ & ~new_new_n13920__;
  assign new_new_n13922__ = new_new_n12860__ & ~new_new_n13921__;
  assign new_new_n13923__ = ~new_new_n12868__ & ~new_new_n13922__;
  assign new_new_n13924__ = new_new_n8065__ & new_new_n12845__;
  assign new_new_n13925__ = new_new_n12868__ & new_new_n13924__;
  assign new_new_n13926__ = ~new_new_n13921__ & new_new_n13925__;
  assign new_new_n13927__ = ~new_new_n13923__ & ~new_new_n13926__;
  assign new_new_n13928__ = ~new_new_n13918__ & ~new_new_n13927__;
  assign new_new_n13929__ = ~new_new_n13917__ & ~new_new_n13928__;
  assign new_new_n13930__ = pi112 & new_new_n13929__;
  assign new_new_n13931__ = ~pi111 & new_new_n13383__;
  assign new_new_n13932__ = pi111 & ~new_new_n13383__;
  assign new_new_n13933__ = ~new_new_n13931__ & ~new_new_n13932__;
  assign new_new_n13934__ = ~pi112 & new_new_n13933__;
  assign new_new_n13935__ = ~new_new_n13929__ & new_new_n13934__;
  assign new_new_n13936__ = new_new_n12849__ & ~new_new_n13930__;
  assign new_new_n13937__ = ~new_new_n13935__ & new_new_n13936__;
  assign new_new_n13938__ = new_new_n12845__ & ~new_new_n13937__;
  assign new_new_n13939__ = pi112 & ~new_new_n11785__;
  assign new_new_n13940__ = ~new_new_n13929__ & ~new_new_n13939__;
  assign new_new_n13941__ = new_new_n274__ & ~new_new_n13933__;
  assign new_new_n13942__ = ~pi112 & new_new_n12845__;
  assign new_new_n13943__ = ~new_new_n13941__ & new_new_n13942__;
  assign new_new_n13944__ = ~new_new_n13940__ & ~new_new_n13943__;
  assign po015 = new_new_n12849__ & ~new_new_n13944__;
  assign new_new_n13946__ = ~new_new_n13917__ & ~new_new_n13918__;
  assign new_new_n13947__ = po015 & new_new_n13946__;
  assign new_new_n13948__ = new_new_n13927__ & ~new_new_n13947__;
  assign new_new_n13949__ = ~new_new_n13927__ & new_new_n13947__;
  assign new_new_n13950__ = ~new_new_n13948__ & ~new_new_n13949__;
  assign new_new_n13951__ = pi112 & ~new_new_n13950__;
  assign new_new_n13952__ = ~pi112 & new_new_n13950__;
  assign new_new_n13953__ = ~new_new_n13393__ & ~new_new_n13394__;
  assign new_new_n13954__ = ~new_new_n13914__ & po015;
  assign new_new_n13955__ = ~pi110 & ~po015;
  assign new_new_n13956__ = ~new_new_n13954__ & ~new_new_n13955__;
  assign new_new_n13957__ = new_new_n13953__ & ~new_new_n13956__;
  assign new_new_n13958__ = ~new_new_n13953__ & new_new_n13956__;
  assign new_new_n13959__ = ~new_new_n13957__ & ~new_new_n13958__;
  assign new_new_n13960__ = pi111 & ~new_new_n13959__;
  assign new_new_n13961__ = ~pi111 & new_new_n13959__;
  assign new_new_n13962__ = ~new_new_n13402__ & ~new_new_n13403__;
  assign new_new_n13963__ = ~new_new_n13912__ & po015;
  assign new_new_n13964__ = ~pi109 & ~po015;
  assign new_new_n13965__ = ~new_new_n13963__ & ~new_new_n13964__;
  assign new_new_n13966__ = new_new_n13962__ & ~new_new_n13965__;
  assign new_new_n13967__ = ~new_new_n13962__ & new_new_n13965__;
  assign new_new_n13968__ = ~new_new_n13966__ & ~new_new_n13967__;
  assign new_new_n13969__ = pi110 & ~new_new_n13968__;
  assign new_new_n13970__ = ~pi110 & new_new_n13968__;
  assign new_new_n13971__ = ~pi108 & ~new_new_n13910__;
  assign new_new_n13972__ = pi108 & new_new_n13910__;
  assign new_new_n13973__ = ~new_new_n13971__ & ~new_new_n13972__;
  assign new_new_n13974__ = po015 & new_new_n13973__;
  assign new_new_n13975__ = new_new_n13410__ & new_new_n13974__;
  assign new_new_n13976__ = ~new_new_n13410__ & ~new_new_n13974__;
  assign new_new_n13977__ = ~new_new_n13975__ & ~new_new_n13976__;
  assign new_new_n13978__ = ~pi109 & ~new_new_n13977__;
  assign new_new_n13979__ = pi109 & new_new_n13977__;
  assign new_new_n13980__ = ~new_new_n13420__ & ~new_new_n13421__;
  assign new_new_n13981__ = ~new_new_n13908__ & po015;
  assign new_new_n13982__ = ~pi107 & ~po015;
  assign new_new_n13983__ = ~new_new_n13981__ & ~new_new_n13982__;
  assign new_new_n13984__ = ~new_new_n13980__ & ~new_new_n13983__;
  assign new_new_n13985__ = new_new_n13980__ & new_new_n13983__;
  assign new_new_n13986__ = ~new_new_n13984__ & ~new_new_n13985__;
  assign new_new_n13987__ = ~pi108 & ~new_new_n13986__;
  assign new_new_n13988__ = pi108 & new_new_n13986__;
  assign new_new_n13989__ = ~new_new_n13436__ & ~new_new_n13437__;
  assign new_new_n13990__ = new_new_n13904__ & po015;
  assign new_new_n13991__ = ~pi105 & ~po015;
  assign new_new_n13992__ = ~new_new_n13990__ & ~new_new_n13991__;
  assign new_new_n13993__ = ~new_new_n13989__ & ~new_new_n13992__;
  assign new_new_n13994__ = new_new_n13989__ & new_new_n13992__;
  assign new_new_n13995__ = ~new_new_n13993__ & ~new_new_n13994__;
  assign new_new_n13996__ = ~pi106 & ~new_new_n13995__;
  assign new_new_n13997__ = pi106 & new_new_n13995__;
  assign new_new_n13998__ = ~new_new_n13902__ & po015;
  assign new_new_n13999__ = pi104 & ~po015;
  assign new_new_n14000__ = ~new_new_n13998__ & ~new_new_n13999__;
  assign new_new_n14001__ = ~new_new_n13445__ & ~new_new_n13446__;
  assign new_new_n14002__ = ~new_new_n14000__ & new_new_n14001__;
  assign new_new_n14003__ = new_new_n14000__ & ~new_new_n14001__;
  assign new_new_n14004__ = ~new_new_n14002__ & ~new_new_n14003__;
  assign new_new_n14005__ = ~pi105 & ~new_new_n14004__;
  assign new_new_n14006__ = pi105 & new_new_n14004__;
  assign new_new_n14007__ = ~new_new_n13900__ & po015;
  assign new_new_n14008__ = pi103 & ~po015;
  assign new_new_n14009__ = ~new_new_n14007__ & ~new_new_n14008__;
  assign new_new_n14010__ = ~new_new_n13454__ & ~new_new_n13455__;
  assign new_new_n14011__ = ~new_new_n14009__ & new_new_n14010__;
  assign new_new_n14012__ = new_new_n14009__ & ~new_new_n14010__;
  assign new_new_n14013__ = ~new_new_n14011__ & ~new_new_n14012__;
  assign new_new_n14014__ = ~pi104 & ~new_new_n14013__;
  assign new_new_n14015__ = pi104 & new_new_n14013__;
  assign new_new_n14016__ = pi102 & ~new_new_n13898__;
  assign new_new_n14017__ = ~pi102 & new_new_n13898__;
  assign new_new_n14018__ = ~new_new_n14016__ & ~new_new_n14017__;
  assign new_new_n14019__ = po015 & new_new_n14018__;
  assign new_new_n14020__ = new_new_n13462__ & new_new_n14019__;
  assign new_new_n14021__ = ~new_new_n13462__ & ~new_new_n14019__;
  assign new_new_n14022__ = ~new_new_n14020__ & ~new_new_n14021__;
  assign new_new_n14023__ = pi103 & ~new_new_n14022__;
  assign new_new_n14024__ = ~pi103 & new_new_n14022__;
  assign new_new_n14025__ = ~new_new_n13472__ & ~new_new_n13473__;
  assign new_new_n14026__ = ~new_new_n13896__ & po015;
  assign new_new_n14027__ = ~pi101 & ~po015;
  assign new_new_n14028__ = ~new_new_n14026__ & ~new_new_n14027__;
  assign new_new_n14029__ = new_new_n14025__ & ~new_new_n14028__;
  assign new_new_n14030__ = ~new_new_n14025__ & new_new_n14028__;
  assign new_new_n14031__ = ~new_new_n14029__ & ~new_new_n14030__;
  assign new_new_n14032__ = pi102 & ~new_new_n14031__;
  assign new_new_n14033__ = ~pi102 & new_new_n14031__;
  assign new_new_n14034__ = ~new_new_n13481__ & ~new_new_n13482__;
  assign new_new_n14035__ = ~new_new_n13894__ & po015;
  assign new_new_n14036__ = ~pi100 & ~po015;
  assign new_new_n14037__ = ~new_new_n14035__ & ~new_new_n14036__;
  assign new_new_n14038__ = new_new_n14034__ & ~new_new_n14037__;
  assign new_new_n14039__ = ~new_new_n14034__ & new_new_n14037__;
  assign new_new_n14040__ = ~new_new_n14038__ & ~new_new_n14039__;
  assign new_new_n14041__ = pi101 & ~new_new_n14040__;
  assign new_new_n14042__ = ~pi101 & new_new_n14040__;
  assign new_new_n14043__ = ~pi099 & ~new_new_n13892__;
  assign new_new_n14044__ = pi099 & new_new_n13892__;
  assign new_new_n14045__ = ~new_new_n14043__ & ~new_new_n14044__;
  assign new_new_n14046__ = po015 & new_new_n14045__;
  assign new_new_n14047__ = new_new_n13489__ & ~new_new_n14046__;
  assign new_new_n14048__ = ~new_new_n13489__ & new_new_n14046__;
  assign new_new_n14049__ = ~new_new_n14047__ & ~new_new_n14048__;
  assign new_new_n14050__ = pi100 & ~new_new_n14049__;
  assign new_new_n14051__ = ~pi100 & new_new_n14049__;
  assign new_new_n14052__ = ~new_new_n13499__ & ~new_new_n13500__;
  assign new_new_n14053__ = ~new_new_n13890__ & po015;
  assign new_new_n14054__ = pi098 & ~po015;
  assign new_new_n14055__ = ~new_new_n14053__ & ~new_new_n14054__;
  assign new_new_n14056__ = new_new_n14052__ & ~new_new_n14055__;
  assign new_new_n14057__ = ~new_new_n14052__ & new_new_n14055__;
  assign new_new_n14058__ = ~new_new_n14056__ & ~new_new_n14057__;
  assign new_new_n14059__ = ~pi099 & ~new_new_n14058__;
  assign new_new_n14060__ = pi099 & new_new_n14058__;
  assign new_new_n14061__ = ~new_new_n13508__ & ~new_new_n13509__;
  assign new_new_n14062__ = ~new_new_n13888__ & po015;
  assign new_new_n14063__ = ~pi097 & ~po015;
  assign new_new_n14064__ = ~new_new_n14062__ & ~new_new_n14063__;
  assign new_new_n14065__ = new_new_n14061__ & new_new_n14064__;
  assign new_new_n14066__ = ~new_new_n14061__ & ~new_new_n14064__;
  assign new_new_n14067__ = ~new_new_n14065__ & ~new_new_n14066__;
  assign new_new_n14068__ = ~pi098 & ~new_new_n14067__;
  assign new_new_n14069__ = pi098 & new_new_n14067__;
  assign new_new_n14070__ = ~new_new_n13517__ & ~new_new_n13518__;
  assign new_new_n14071__ = ~new_new_n13886__ & po015;
  assign new_new_n14072__ = ~pi096 & ~po015;
  assign new_new_n14073__ = ~new_new_n14071__ & ~new_new_n14072__;
  assign new_new_n14074__ = ~new_new_n14070__ & ~new_new_n14073__;
  assign new_new_n14075__ = new_new_n14070__ & new_new_n14073__;
  assign new_new_n14076__ = ~new_new_n14074__ & ~new_new_n14075__;
  assign new_new_n14077__ = ~pi097 & ~new_new_n14076__;
  assign new_new_n14078__ = pi097 & new_new_n14076__;
  assign new_new_n14079__ = new_new_n13884__ & po015;
  assign new_new_n14080__ = pi095 & ~po015;
  assign new_new_n14081__ = ~new_new_n14079__ & ~new_new_n14080__;
  assign new_new_n14082__ = ~new_new_n13526__ & ~new_new_n13527__;
  assign new_new_n14083__ = ~new_new_n14081__ & ~new_new_n14082__;
  assign new_new_n14084__ = new_new_n14081__ & new_new_n14082__;
  assign new_new_n14085__ = ~new_new_n14083__ & ~new_new_n14084__;
  assign new_new_n14086__ = ~pi096 & new_new_n14085__;
  assign new_new_n14087__ = pi096 & ~new_new_n14085__;
  assign new_new_n14088__ = ~new_new_n13535__ & ~new_new_n13536__;
  assign new_new_n14089__ = ~new_new_n13882__ & po015;
  assign new_new_n14090__ = ~pi094 & ~po015;
  assign new_new_n14091__ = ~new_new_n14089__ & ~new_new_n14090__;
  assign new_new_n14092__ = ~new_new_n14088__ & ~new_new_n14091__;
  assign new_new_n14093__ = new_new_n14088__ & new_new_n14091__;
  assign new_new_n14094__ = ~new_new_n14092__ & ~new_new_n14093__;
  assign new_new_n14095__ = ~pi095 & ~new_new_n14094__;
  assign new_new_n14096__ = pi095 & new_new_n14094__;
  assign new_new_n14097__ = ~new_new_n13544__ & ~new_new_n13545__;
  assign new_new_n14098__ = ~new_new_n13880__ & po015;
  assign new_new_n14099__ = ~pi093 & ~po015;
  assign new_new_n14100__ = ~new_new_n14098__ & ~new_new_n14099__;
  assign new_new_n14101__ = ~new_new_n14097__ & ~new_new_n14100__;
  assign new_new_n14102__ = new_new_n14097__ & new_new_n14100__;
  assign new_new_n14103__ = ~new_new_n14101__ & ~new_new_n14102__;
  assign new_new_n14104__ = ~pi094 & ~new_new_n14103__;
  assign new_new_n14105__ = pi094 & new_new_n14103__;
  assign new_new_n14106__ = new_new_n13878__ & po015;
  assign new_new_n14107__ = ~pi092 & ~po015;
  assign new_new_n14108__ = ~new_new_n14106__ & ~new_new_n14107__;
  assign new_new_n14109__ = ~new_new_n13553__ & ~new_new_n13554__;
  assign new_new_n14110__ = ~new_new_n14108__ & ~new_new_n14109__;
  assign new_new_n14111__ = new_new_n14108__ & new_new_n14109__;
  assign new_new_n14112__ = ~new_new_n14110__ & ~new_new_n14111__;
  assign new_new_n14113__ = ~pi093 & ~new_new_n14112__;
  assign new_new_n14114__ = pi093 & new_new_n14112__;
  assign new_new_n14115__ = ~new_new_n13562__ & ~new_new_n13563__;
  assign new_new_n14116__ = ~new_new_n13876__ & po015;
  assign new_new_n14117__ = ~pi091 & ~po015;
  assign new_new_n14118__ = ~new_new_n14116__ & ~new_new_n14117__;
  assign new_new_n14119__ = new_new_n14115__ & ~new_new_n14118__;
  assign new_new_n14120__ = ~new_new_n14115__ & new_new_n14118__;
  assign new_new_n14121__ = ~new_new_n14119__ & ~new_new_n14120__;
  assign new_new_n14122__ = pi092 & ~new_new_n14121__;
  assign new_new_n14123__ = ~pi092 & new_new_n14121__;
  assign new_new_n14124__ = ~new_new_n13874__ & po015;
  assign new_new_n14125__ = pi090 & ~po015;
  assign new_new_n14126__ = ~new_new_n14124__ & ~new_new_n14125__;
  assign new_new_n14127__ = ~new_new_n13571__ & ~new_new_n13572__;
  assign new_new_n14128__ = ~new_new_n14126__ & new_new_n14127__;
  assign new_new_n14129__ = new_new_n14126__ & ~new_new_n14127__;
  assign new_new_n14130__ = ~new_new_n14128__ & ~new_new_n14129__;
  assign new_new_n14131__ = ~pi091 & ~new_new_n14130__;
  assign new_new_n14132__ = pi091 & new_new_n14130__;
  assign new_new_n14133__ = ~new_new_n13580__ & ~new_new_n13581__;
  assign new_new_n14134__ = ~new_new_n13872__ & po015;
  assign new_new_n14135__ = pi089 & ~po015;
  assign new_new_n14136__ = ~new_new_n14134__ & ~new_new_n14135__;
  assign new_new_n14137__ = new_new_n14133__ & new_new_n14136__;
  assign new_new_n14138__ = ~new_new_n14133__ & ~new_new_n14136__;
  assign new_new_n14139__ = ~new_new_n14137__ & ~new_new_n14138__;
  assign new_new_n14140__ = ~pi090 & new_new_n14139__;
  assign new_new_n14141__ = pi090 & ~new_new_n14139__;
  assign new_new_n14142__ = pi088 & ~new_new_n13870__;
  assign new_new_n14143__ = ~pi088 & new_new_n13870__;
  assign new_new_n14144__ = ~new_new_n14142__ & ~new_new_n14143__;
  assign new_new_n14145__ = po015 & new_new_n14144__;
  assign new_new_n14146__ = ~new_new_n13588__ & ~new_new_n14145__;
  assign new_new_n14147__ = new_new_n13588__ & new_new_n14145__;
  assign new_new_n14148__ = ~new_new_n14146__ & ~new_new_n14147__;
  assign new_new_n14149__ = ~pi089 & new_new_n14148__;
  assign new_new_n14150__ = pi089 & ~new_new_n14148__;
  assign new_new_n14151__ = ~new_new_n13598__ & ~new_new_n13599__;
  assign new_new_n14152__ = ~new_new_n13868__ & po015;
  assign new_new_n14153__ = ~pi087 & ~po015;
  assign new_new_n14154__ = ~new_new_n14152__ & ~new_new_n14153__;
  assign new_new_n14155__ = new_new_n14151__ & new_new_n14154__;
  assign new_new_n14156__ = ~new_new_n14151__ & ~new_new_n14154__;
  assign new_new_n14157__ = ~new_new_n14155__ & ~new_new_n14156__;
  assign new_new_n14158__ = ~pi088 & ~new_new_n14157__;
  assign new_new_n14159__ = pi088 & new_new_n14157__;
  assign new_new_n14160__ = new_new_n13866__ & po015;
  assign new_new_n14161__ = ~pi086 & ~po015;
  assign new_new_n14162__ = ~new_new_n14160__ & ~new_new_n14161__;
  assign new_new_n14163__ = ~new_new_n13607__ & ~new_new_n13608__;
  assign new_new_n14164__ = ~new_new_n14162__ & ~new_new_n14163__;
  assign new_new_n14165__ = new_new_n14162__ & new_new_n14163__;
  assign new_new_n14166__ = ~new_new_n14164__ & ~new_new_n14165__;
  assign new_new_n14167__ = ~pi087 & ~new_new_n14166__;
  assign new_new_n14168__ = pi087 & new_new_n14166__;
  assign new_new_n14169__ = ~new_new_n13864__ & po015;
  assign new_new_n14170__ = pi085 & ~po015;
  assign new_new_n14171__ = ~new_new_n14169__ & ~new_new_n14170__;
  assign new_new_n14172__ = ~new_new_n13616__ & ~new_new_n13617__;
  assign new_new_n14173__ = ~new_new_n14171__ & new_new_n14172__;
  assign new_new_n14174__ = new_new_n14171__ & ~new_new_n14172__;
  assign new_new_n14175__ = ~new_new_n14173__ & ~new_new_n14174__;
  assign new_new_n14176__ = pi086 & new_new_n14175__;
  assign new_new_n14177__ = ~pi086 & ~new_new_n14175__;
  assign new_new_n14178__ = ~pi084 & ~new_new_n13862__;
  assign new_new_n14179__ = pi084 & new_new_n13862__;
  assign new_new_n14180__ = ~new_new_n14178__ & ~new_new_n14179__;
  assign new_new_n14181__ = po015 & ~new_new_n14180__;
  assign new_new_n14182__ = ~new_new_n13624__ & ~new_new_n14181__;
  assign new_new_n14183__ = new_new_n13624__ & new_new_n14181__;
  assign new_new_n14184__ = ~new_new_n14182__ & ~new_new_n14183__;
  assign new_new_n14185__ = pi085 & ~new_new_n14184__;
  assign new_new_n14186__ = ~pi085 & new_new_n14184__;
  assign new_new_n14187__ = ~new_new_n13634__ & ~new_new_n13860__;
  assign new_new_n14188__ = pi083 & ~po015;
  assign new_new_n14189__ = ~new_new_n13859__ & po015;
  assign new_new_n14190__ = ~new_new_n14188__ & ~new_new_n14189__;
  assign new_new_n14191__ = new_new_n14187__ & new_new_n14190__;
  assign new_new_n14192__ = ~new_new_n14187__ & ~new_new_n14190__;
  assign new_new_n14193__ = ~new_new_n14191__ & ~new_new_n14192__;
  assign new_new_n14194__ = pi084 & ~new_new_n14193__;
  assign new_new_n14195__ = ~pi084 & new_new_n14193__;
  assign new_new_n14196__ = ~new_new_n13642__ & ~new_new_n13643__;
  assign new_new_n14197__ = ~new_new_n13857__ & po015;
  assign new_new_n14198__ = pi082 & ~po015;
  assign new_new_n14199__ = ~new_new_n14197__ & ~new_new_n14198__;
  assign new_new_n14200__ = new_new_n14196__ & new_new_n14199__;
  assign new_new_n14201__ = ~new_new_n14196__ & ~new_new_n14199__;
  assign new_new_n14202__ = ~new_new_n14200__ & ~new_new_n14201__;
  assign new_new_n14203__ = pi083 & ~new_new_n14202__;
  assign new_new_n14204__ = ~pi083 & new_new_n14202__;
  assign new_new_n14205__ = new_new_n13855__ & po015;
  assign new_new_n14206__ = ~pi081 & ~po015;
  assign new_new_n14207__ = ~new_new_n14205__ & ~new_new_n14206__;
  assign new_new_n14208__ = ~new_new_n13651__ & ~new_new_n13652__;
  assign new_new_n14209__ = ~new_new_n14207__ & ~new_new_n14208__;
  assign new_new_n14210__ = new_new_n14207__ & new_new_n14208__;
  assign new_new_n14211__ = ~new_new_n14209__ & ~new_new_n14210__;
  assign new_new_n14212__ = ~pi082 & ~new_new_n14211__;
  assign new_new_n14213__ = pi082 & new_new_n14211__;
  assign new_new_n14214__ = ~new_new_n13660__ & ~new_new_n13661__;
  assign new_new_n14215__ = pi080 & ~po015;
  assign new_new_n14216__ = ~new_new_n13853__ & po015;
  assign new_new_n14217__ = ~new_new_n14215__ & ~new_new_n14216__;
  assign new_new_n14218__ = new_new_n14214__ & new_new_n14217__;
  assign new_new_n14219__ = ~new_new_n14214__ & ~new_new_n14217__;
  assign new_new_n14220__ = ~new_new_n14218__ & ~new_new_n14219__;
  assign new_new_n14221__ = pi081 & ~new_new_n14220__;
  assign new_new_n14222__ = ~pi081 & new_new_n14220__;
  assign new_new_n14223__ = ~new_new_n13669__ & ~new_new_n13670__;
  assign new_new_n14224__ = ~new_new_n13851__ & po015;
  assign new_new_n14225__ = pi079 & ~po015;
  assign new_new_n14226__ = ~new_new_n14224__ & ~new_new_n14225__;
  assign new_new_n14227__ = new_new_n14223__ & new_new_n14226__;
  assign new_new_n14228__ = ~new_new_n14223__ & ~new_new_n14226__;
  assign new_new_n14229__ = ~new_new_n14227__ & ~new_new_n14228__;
  assign new_new_n14230__ = pi080 & ~new_new_n14229__;
  assign new_new_n14231__ = ~pi080 & new_new_n14229__;
  assign new_new_n14232__ = new_new_n13849__ & po015;
  assign new_new_n14233__ = pi078 & ~po015;
  assign new_new_n14234__ = ~new_new_n14232__ & ~new_new_n14233__;
  assign new_new_n14235__ = ~new_new_n13678__ & ~new_new_n13679__;
  assign new_new_n14236__ = ~new_new_n14234__ & ~new_new_n14235__;
  assign new_new_n14237__ = new_new_n14234__ & new_new_n14235__;
  assign new_new_n14238__ = ~new_new_n14236__ & ~new_new_n14237__;
  assign new_new_n14239__ = pi079 & ~new_new_n14238__;
  assign new_new_n14240__ = ~pi079 & new_new_n14238__;
  assign new_new_n14241__ = ~new_new_n13687__ & ~new_new_n13688__;
  assign new_new_n14242__ = ~new_new_n13847__ & po015;
  assign new_new_n14243__ = ~pi077 & ~po015;
  assign new_new_n14244__ = ~new_new_n14242__ & ~new_new_n14243__;
  assign new_new_n14245__ = new_new_n14241__ & ~new_new_n14244__;
  assign new_new_n14246__ = ~new_new_n14241__ & new_new_n14244__;
  assign new_new_n14247__ = ~new_new_n14245__ & ~new_new_n14246__;
  assign new_new_n14248__ = pi078 & ~new_new_n14247__;
  assign new_new_n14249__ = ~pi078 & new_new_n14247__;
  assign new_new_n14250__ = ~new_new_n13696__ & ~new_new_n13697__;
  assign new_new_n14251__ = ~new_new_n13845__ & po015;
  assign new_new_n14252__ = ~pi076 & ~po015;
  assign new_new_n14253__ = ~new_new_n14251__ & ~new_new_n14252__;
  assign new_new_n14254__ = new_new_n14250__ & ~new_new_n14253__;
  assign new_new_n14255__ = ~new_new_n14250__ & new_new_n14253__;
  assign new_new_n14256__ = ~new_new_n14254__ & ~new_new_n14255__;
  assign new_new_n14257__ = pi077 & ~new_new_n14256__;
  assign new_new_n14258__ = ~pi077 & new_new_n14256__;
  assign new_new_n14259__ = ~pi075 & ~new_new_n13843__;
  assign new_new_n14260__ = pi075 & new_new_n13843__;
  assign new_new_n14261__ = ~new_new_n14259__ & ~new_new_n14260__;
  assign new_new_n14262__ = po015 & new_new_n14261__;
  assign new_new_n14263__ = new_new_n13704__ & new_new_n14262__;
  assign new_new_n14264__ = ~new_new_n13704__ & ~new_new_n14262__;
  assign new_new_n14265__ = ~new_new_n14263__ & ~new_new_n14264__;
  assign new_new_n14266__ = pi076 & new_new_n14265__;
  assign new_new_n14267__ = ~pi076 & ~new_new_n14265__;
  assign new_new_n14268__ = ~new_new_n13714__ & ~new_new_n13715__;
  assign new_new_n14269__ = ~new_new_n13841__ & po015;
  assign new_new_n14270__ = ~pi074 & ~po015;
  assign new_new_n14271__ = ~new_new_n14269__ & ~new_new_n14270__;
  assign new_new_n14272__ = new_new_n14268__ & ~new_new_n14271__;
  assign new_new_n14273__ = ~new_new_n14268__ & new_new_n14271__;
  assign new_new_n14274__ = ~new_new_n14272__ & ~new_new_n14273__;
  assign new_new_n14275__ = pi075 & ~new_new_n14274__;
  assign new_new_n14276__ = ~pi075 & new_new_n14274__;
  assign new_new_n14277__ = ~new_new_n13839__ & po015;
  assign new_new_n14278__ = pi073 & ~po015;
  assign new_new_n14279__ = ~new_new_n14277__ & ~new_new_n14278__;
  assign new_new_n14280__ = ~new_new_n13723__ & ~new_new_n13724__;
  assign new_new_n14281__ = ~new_new_n14279__ & new_new_n14280__;
  assign new_new_n14282__ = new_new_n14279__ & ~new_new_n14280__;
  assign new_new_n14283__ = ~new_new_n14281__ & ~new_new_n14282__;
  assign new_new_n14284__ = ~pi074 & ~new_new_n14283__;
  assign new_new_n14285__ = pi074 & new_new_n14283__;
  assign new_new_n14286__ = ~new_new_n13837__ & po015;
  assign new_new_n14287__ = pi072 & ~po015;
  assign new_new_n14288__ = ~new_new_n14286__ & ~new_new_n14287__;
  assign new_new_n14289__ = ~new_new_n13730__ & ~new_new_n13731__;
  assign new_new_n14290__ = ~new_new_n14288__ & new_new_n14289__;
  assign new_new_n14291__ = new_new_n14288__ & ~new_new_n14289__;
  assign new_new_n14292__ = ~new_new_n14290__ & ~new_new_n14291__;
  assign new_new_n14293__ = ~pi073 & ~new_new_n14292__;
  assign new_new_n14294__ = pi073 & new_new_n14292__;
  assign new_new_n14295__ = ~new_new_n13739__ & ~new_new_n13740__;
  assign new_new_n14296__ = new_new_n13835__ & po015;
  assign new_new_n14297__ = ~pi071 & ~po015;
  assign new_new_n14298__ = ~new_new_n14296__ & ~new_new_n14297__;
  assign new_new_n14299__ = ~new_new_n14295__ & ~new_new_n14298__;
  assign new_new_n14300__ = new_new_n14295__ & new_new_n14298__;
  assign new_new_n14301__ = ~new_new_n14299__ & ~new_new_n14300__;
  assign new_new_n14302__ = ~pi072 & ~new_new_n14301__;
  assign new_new_n14303__ = pi072 & new_new_n14301__;
  assign new_new_n14304__ = ~new_new_n13827__ & po015;
  assign new_new_n14305__ = ~new_new_n13828__ & new_new_n14304__;
  assign new_new_n14306__ = new_new_n13833__ & ~new_new_n14305__;
  assign new_new_n14307__ = new_new_n13834__ & new_new_n14304__;
  assign new_new_n14308__ = ~new_new_n14306__ & ~new_new_n14307__;
  assign new_new_n14309__ = ~pi071 & ~new_new_n14308__;
  assign new_new_n14310__ = pi071 & new_new_n14308__;
  assign new_new_n14311__ = new_new_n13824__ & po015;
  assign new_new_n14312__ = pi069 & ~po015;
  assign new_new_n14313__ = ~new_new_n14311__ & ~new_new_n14312__;
  assign new_new_n14314__ = ~new_new_n13748__ & ~new_new_n13749__;
  assign new_new_n14315__ = ~new_new_n14313__ & ~new_new_n14314__;
  assign new_new_n14316__ = new_new_n14313__ & new_new_n14314__;
  assign new_new_n14317__ = ~new_new_n14315__ & ~new_new_n14316__;
  assign new_new_n14318__ = pi070 & ~new_new_n14317__;
  assign new_new_n14319__ = ~pi070 & new_new_n14317__;
  assign new_new_n14320__ = ~new_new_n13757__ & ~new_new_n13758__;
  assign new_new_n14321__ = ~new_new_n13822__ & po015;
  assign new_new_n14322__ = ~pi068 & ~po015;
  assign new_new_n14323__ = ~new_new_n14321__ & ~new_new_n14322__;
  assign new_new_n14324__ = new_new_n14320__ & ~new_new_n14323__;
  assign new_new_n14325__ = ~new_new_n14320__ & new_new_n14323__;
  assign new_new_n14326__ = ~new_new_n14324__ & ~new_new_n14325__;
  assign new_new_n14327__ = pi069 & ~new_new_n14326__;
  assign new_new_n14328__ = ~pi069 & new_new_n14326__;
  assign new_new_n14329__ = ~new_new_n13778__ & ~new_new_n13779__;
  assign new_new_n14330__ = new_new_n13820__ & po015;
  assign new_new_n14331__ = ~pi067 & ~po015;
  assign new_new_n14332__ = ~new_new_n14330__ & ~new_new_n14331__;
  assign new_new_n14333__ = ~new_new_n14329__ & ~new_new_n14332__;
  assign new_new_n14334__ = new_new_n14329__ & new_new_n14332__;
  assign new_new_n14335__ = ~new_new_n14333__ & ~new_new_n14334__;
  assign new_new_n14336__ = ~pi068 & ~new_new_n14335__;
  assign new_new_n14337__ = pi068 & new_new_n14335__;
  assign new_new_n14338__ = ~new_new_n13792__ & po015;
  assign new_new_n14339__ = ~new_new_n13793__ & new_new_n14338__;
  assign new_new_n14340__ = new_new_n13818__ & ~new_new_n14339__;
  assign new_new_n14341__ = new_new_n13819__ & new_new_n14338__;
  assign new_new_n14342__ = ~new_new_n14340__ & ~new_new_n14341__;
  assign new_new_n14343__ = ~pi067 & ~new_new_n14342__;
  assign new_new_n14344__ = pi067 & new_new_n14342__;
  assign new_new_n14345__ = ~pi014 & pi064;
  assign new_new_n14346__ = ~pi065 & ~new_new_n14345__;
  assign new_new_n14347__ = pi064 & po015;
  assign new_new_n14348__ = ~pi015 & ~new_new_n14347__;
  assign new_new_n14349__ = ~new_new_n14346__ & new_new_n14348__;
  assign new_new_n14350__ = ~pi014 & pi065;
  assign new_new_n14351__ = pi014 & ~pi065;
  assign new_new_n14352__ = pi015 & ~new_new_n14351__;
  assign new_new_n14353__ = po015 & new_new_n14352__;
  assign new_new_n14354__ = ~new_new_n14350__ & ~new_new_n14353__;
  assign new_new_n14355__ = pi064 & ~new_new_n14354__;
  assign new_new_n14356__ = ~new_new_n14349__ & ~new_new_n14355__;
  assign new_new_n14357__ = pi066 & ~new_new_n14356__;
  assign new_new_n14358__ = ~pi066 & new_new_n14356__;
  assign new_new_n14359__ = ~new_new_n332__ & po015;
  assign new_new_n14360__ = ~new_new_n13789__ & ~new_new_n14359__;
  assign new_new_n14361__ = po016 & ~po015;
  assign new_new_n14362__ = ~new_new_n426__ & ~po016;
  assign new_new_n14363__ = ~pi015 & ~new_new_n13807__;
  assign new_new_n14364__ = ~new_new_n14362__ & new_new_n14363__;
  assign new_new_n14365__ = ~new_new_n14361__ & new_new_n14364__;
  assign new_new_n14366__ = pi065 & po015;
  assign new_new_n14367__ = po016 & ~new_new_n14366__;
  assign new_new_n14368__ = pi015 & ~new_new_n13801__;
  assign new_new_n14369__ = ~new_new_n14367__ & new_new_n14368__;
  assign new_new_n14370__ = ~new_new_n14360__ & ~new_new_n14365__;
  assign new_new_n14371__ = ~new_new_n14369__ & new_new_n14370__;
  assign new_new_n14372__ = ~pi016 & ~new_new_n14371__;
  assign new_new_n14373__ = new_new_n13797__ & po015;
  assign new_new_n14374__ = ~new_new_n13807__ & ~new_new_n14373__;
  assign new_new_n14375__ = ~pi015 & ~new_new_n14374__;
  assign new_new_n14376__ = ~new_new_n14361__ & ~new_new_n14375__;
  assign new_new_n14377__ = pi064 & ~new_new_n14376__;
  assign new_new_n14378__ = ~new_new_n13789__ & ~new_new_n14366__;
  assign new_new_n14379__ = pi015 & ~new_new_n13807__;
  assign new_new_n14380__ = pi064 & ~new_new_n14379__;
  assign new_new_n14381__ = ~new_new_n14378__ & ~new_new_n14380__;
  assign new_new_n14382__ = ~new_new_n14377__ & ~new_new_n14381__;
  assign new_new_n14383__ = pi016 & ~new_new_n14382__;
  assign new_new_n14384__ = ~new_new_n14372__ & ~new_new_n14383__;
  assign new_new_n14385__ = ~new_new_n14358__ & ~new_new_n14384__;
  assign new_new_n14386__ = ~new_new_n14357__ & ~new_new_n14385__;
  assign new_new_n14387__ = ~new_new_n14344__ & new_new_n14386__;
  assign new_new_n14388__ = ~new_new_n14343__ & ~new_new_n14387__;
  assign new_new_n14389__ = ~new_new_n14337__ & ~new_new_n14388__;
  assign new_new_n14390__ = ~new_new_n14336__ & ~new_new_n14389__;
  assign new_new_n14391__ = ~new_new_n14328__ & new_new_n14390__;
  assign new_new_n14392__ = ~new_new_n14327__ & ~new_new_n14391__;
  assign new_new_n14393__ = ~new_new_n14319__ & ~new_new_n14392__;
  assign new_new_n14394__ = ~new_new_n14318__ & ~new_new_n14393__;
  assign new_new_n14395__ = ~new_new_n14310__ & new_new_n14394__;
  assign new_new_n14396__ = ~new_new_n14309__ & ~new_new_n14395__;
  assign new_new_n14397__ = ~new_new_n14303__ & ~new_new_n14396__;
  assign new_new_n14398__ = ~new_new_n14302__ & ~new_new_n14397__;
  assign new_new_n14399__ = ~new_new_n14294__ & ~new_new_n14398__;
  assign new_new_n14400__ = ~new_new_n14293__ & ~new_new_n14399__;
  assign new_new_n14401__ = ~new_new_n14285__ & ~new_new_n14400__;
  assign new_new_n14402__ = ~new_new_n14284__ & ~new_new_n14401__;
  assign new_new_n14403__ = ~new_new_n14276__ & new_new_n14402__;
  assign new_new_n14404__ = ~new_new_n14275__ & ~new_new_n14403__;
  assign new_new_n14405__ = ~new_new_n14267__ & ~new_new_n14404__;
  assign new_new_n14406__ = ~new_new_n14266__ & ~new_new_n14405__;
  assign new_new_n14407__ = ~new_new_n14258__ & ~new_new_n14406__;
  assign new_new_n14408__ = ~new_new_n14257__ & ~new_new_n14407__;
  assign new_new_n14409__ = ~new_new_n14249__ & ~new_new_n14408__;
  assign new_new_n14410__ = ~new_new_n14248__ & ~new_new_n14409__;
  assign new_new_n14411__ = ~new_new_n14240__ & ~new_new_n14410__;
  assign new_new_n14412__ = ~new_new_n14239__ & ~new_new_n14411__;
  assign new_new_n14413__ = ~new_new_n14231__ & ~new_new_n14412__;
  assign new_new_n14414__ = ~new_new_n14230__ & ~new_new_n14413__;
  assign new_new_n14415__ = ~new_new_n14222__ & ~new_new_n14414__;
  assign new_new_n14416__ = ~new_new_n14221__ & ~new_new_n14415__;
  assign new_new_n14417__ = ~new_new_n14213__ & new_new_n14416__;
  assign new_new_n14418__ = ~new_new_n14212__ & ~new_new_n14417__;
  assign new_new_n14419__ = ~new_new_n14204__ & new_new_n14418__;
  assign new_new_n14420__ = ~new_new_n14203__ & ~new_new_n14419__;
  assign new_new_n14421__ = ~new_new_n14195__ & ~new_new_n14420__;
  assign new_new_n14422__ = ~new_new_n14194__ & ~new_new_n14421__;
  assign new_new_n14423__ = ~new_new_n14186__ & ~new_new_n14422__;
  assign new_new_n14424__ = ~new_new_n14185__ & ~new_new_n14423__;
  assign new_new_n14425__ = ~new_new_n14177__ & ~new_new_n14424__;
  assign new_new_n14426__ = ~new_new_n14176__ & ~new_new_n14425__;
  assign new_new_n14427__ = ~new_new_n14168__ & new_new_n14426__;
  assign new_new_n14428__ = ~new_new_n14167__ & ~new_new_n14427__;
  assign new_new_n14429__ = ~new_new_n14159__ & ~new_new_n14428__;
  assign new_new_n14430__ = ~new_new_n14158__ & ~new_new_n14429__;
  assign new_new_n14431__ = ~new_new_n14150__ & ~new_new_n14430__;
  assign new_new_n14432__ = ~new_new_n14149__ & ~new_new_n14431__;
  assign new_new_n14433__ = ~new_new_n14141__ & ~new_new_n14432__;
  assign new_new_n14434__ = ~new_new_n14140__ & ~new_new_n14433__;
  assign new_new_n14435__ = ~new_new_n14132__ & ~new_new_n14434__;
  assign new_new_n14436__ = ~new_new_n14131__ & ~new_new_n14435__;
  assign new_new_n14437__ = ~new_new_n14123__ & new_new_n14436__;
  assign new_new_n14438__ = ~new_new_n14122__ & ~new_new_n14437__;
  assign new_new_n14439__ = ~new_new_n14114__ & new_new_n14438__;
  assign new_new_n14440__ = ~new_new_n14113__ & ~new_new_n14439__;
  assign new_new_n14441__ = ~new_new_n14105__ & ~new_new_n14440__;
  assign new_new_n14442__ = ~new_new_n14104__ & ~new_new_n14441__;
  assign new_new_n14443__ = ~new_new_n14096__ & ~new_new_n14442__;
  assign new_new_n14444__ = ~new_new_n14095__ & ~new_new_n14443__;
  assign new_new_n14445__ = ~new_new_n14087__ & ~new_new_n14444__;
  assign new_new_n14446__ = ~new_new_n14086__ & ~new_new_n14445__;
  assign new_new_n14447__ = ~new_new_n14078__ & ~new_new_n14446__;
  assign new_new_n14448__ = ~new_new_n14077__ & ~new_new_n14447__;
  assign new_new_n14449__ = ~new_new_n14069__ & ~new_new_n14448__;
  assign new_new_n14450__ = ~new_new_n14068__ & ~new_new_n14449__;
  assign new_new_n14451__ = ~new_new_n14060__ & ~new_new_n14450__;
  assign new_new_n14452__ = ~new_new_n14059__ & ~new_new_n14451__;
  assign new_new_n14453__ = ~new_new_n14051__ & new_new_n14452__;
  assign new_new_n14454__ = ~new_new_n14050__ & ~new_new_n14453__;
  assign new_new_n14455__ = ~new_new_n14042__ & ~new_new_n14454__;
  assign new_new_n14456__ = ~new_new_n14041__ & ~new_new_n14455__;
  assign new_new_n14457__ = ~new_new_n14033__ & ~new_new_n14456__;
  assign new_new_n14458__ = ~new_new_n14032__ & ~new_new_n14457__;
  assign new_new_n14459__ = ~new_new_n14024__ & ~new_new_n14458__;
  assign new_new_n14460__ = ~new_new_n14023__ & ~new_new_n14459__;
  assign new_new_n14461__ = ~new_new_n14015__ & new_new_n14460__;
  assign new_new_n14462__ = ~new_new_n14014__ & ~new_new_n14461__;
  assign new_new_n14463__ = ~new_new_n14006__ & ~new_new_n14462__;
  assign new_new_n14464__ = ~new_new_n14005__ & ~new_new_n14463__;
  assign new_new_n14465__ = ~new_new_n13997__ & ~new_new_n14464__;
  assign new_new_n14466__ = ~new_new_n13996__ & ~new_new_n14465__;
  assign new_new_n14467__ = pi107 & new_new_n14466__;
  assign new_new_n14468__ = ~pi107 & ~new_new_n14466__;
  assign new_new_n14469__ = pi106 & ~new_new_n13906__;
  assign new_new_n14470__ = ~pi106 & new_new_n13906__;
  assign new_new_n14471__ = ~new_new_n14469__ & ~new_new_n14470__;
  assign new_new_n14472__ = po015 & new_new_n14471__;
  assign new_new_n14473__ = new_new_n13428__ & ~new_new_n14472__;
  assign new_new_n14474__ = ~new_new_n13428__ & new_new_n14472__;
  assign new_new_n14475__ = ~new_new_n14473__ & ~new_new_n14474__;
  assign new_new_n14476__ = ~new_new_n14468__ & ~new_new_n14475__;
  assign new_new_n14477__ = ~new_new_n14467__ & ~new_new_n14476__;
  assign new_new_n14478__ = ~new_new_n13988__ & new_new_n14477__;
  assign new_new_n14479__ = ~new_new_n13987__ & ~new_new_n14478__;
  assign new_new_n14480__ = ~new_new_n13979__ & ~new_new_n14479__;
  assign new_new_n14481__ = ~new_new_n13978__ & ~new_new_n14480__;
  assign new_new_n14482__ = ~new_new_n13970__ & new_new_n14481__;
  assign new_new_n14483__ = ~new_new_n13969__ & ~new_new_n14482__;
  assign new_new_n14484__ = ~new_new_n13961__ & ~new_new_n14483__;
  assign new_new_n14485__ = ~new_new_n13960__ & ~new_new_n14484__;
  assign new_new_n14486__ = ~new_new_n13952__ & ~new_new_n14485__;
  assign new_new_n14487__ = ~new_new_n13951__ & ~new_new_n14486__;
  assign new_new_n14488__ = ~pi113 & new_new_n14487__;
  assign new_new_n14489__ = pi113 & ~new_new_n14487__;
  assign new_new_n14490__ = new_new_n12848__ & ~new_new_n14488__;
  assign new_new_n14491__ = ~new_new_n14489__ & new_new_n14490__;
  assign new_new_n14492__ = new_new_n13938__ & ~new_new_n14491__;
  assign new_new_n14493__ = ~pi113 & new_new_n13938__;
  assign new_new_n14494__ = ~new_new_n14487__ & ~new_new_n14493__;
  assign new_new_n14495__ = pi113 & ~new_new_n12845__;
  assign new_new_n14496__ = new_new_n12848__ & ~new_new_n14495__;
  assign po014 = ~new_new_n14494__ & new_new_n14496__;
  assign new_new_n14498__ = ~new_new_n14485__ & po014;
  assign new_new_n14499__ = pi112 & ~po014;
  assign new_new_n14500__ = ~new_new_n14498__ & ~new_new_n14499__;
  assign new_new_n14501__ = ~new_new_n13951__ & ~new_new_n13952__;
  assign new_new_n14502__ = ~new_new_n14500__ & new_new_n14501__;
  assign new_new_n14503__ = new_new_n14500__ & ~new_new_n14501__;
  assign new_new_n14504__ = ~new_new_n14502__ & ~new_new_n14503__;
  assign new_new_n14505__ = pi113 & new_new_n14504__;
  assign new_new_n14506__ = ~pi113 & ~new_new_n14504__;
  assign new_new_n14507__ = ~new_new_n13960__ & ~new_new_n13961__;
  assign new_new_n14508__ = ~new_new_n14483__ & po014;
  assign new_new_n14509__ = pi111 & ~po014;
  assign new_new_n14510__ = ~new_new_n14508__ & ~new_new_n14509__;
  assign new_new_n14511__ = new_new_n14507__ & new_new_n14510__;
  assign new_new_n14512__ = ~new_new_n14507__ & ~new_new_n14510__;
  assign new_new_n14513__ = ~new_new_n14511__ & ~new_new_n14512__;
  assign new_new_n14514__ = pi112 & ~new_new_n14513__;
  assign new_new_n14515__ = ~pi112 & new_new_n14513__;
  assign new_new_n14516__ = new_new_n14481__ & po014;
  assign new_new_n14517__ = pi110 & ~po014;
  assign new_new_n14518__ = ~new_new_n14516__ & ~new_new_n14517__;
  assign new_new_n14519__ = ~new_new_n13969__ & ~new_new_n13970__;
  assign new_new_n14520__ = ~new_new_n14518__ & ~new_new_n14519__;
  assign new_new_n14521__ = new_new_n14518__ & new_new_n14519__;
  assign new_new_n14522__ = ~new_new_n14520__ & ~new_new_n14521__;
  assign new_new_n14523__ = pi111 & ~new_new_n14522__;
  assign new_new_n14524__ = ~pi111 & new_new_n14522__;
  assign new_new_n14525__ = ~new_new_n14477__ & po014;
  assign new_new_n14526__ = pi108 & ~po014;
  assign new_new_n14527__ = ~new_new_n14525__ & ~new_new_n14526__;
  assign new_new_n14528__ = ~new_new_n13987__ & ~new_new_n13988__;
  assign new_new_n14529__ = ~new_new_n14527__ & new_new_n14528__;
  assign new_new_n14530__ = new_new_n14527__ & ~new_new_n14528__;
  assign new_new_n14531__ = ~new_new_n14529__ & ~new_new_n14530__;
  assign new_new_n14532__ = ~pi109 & ~new_new_n14531__;
  assign new_new_n14533__ = pi109 & new_new_n14531__;
  assign new_new_n14534__ = ~new_new_n14467__ & ~new_new_n14468__;
  assign new_new_n14535__ = po014 & new_new_n14534__;
  assign new_new_n14536__ = new_new_n14475__ & new_new_n14535__;
  assign new_new_n14537__ = ~new_new_n14475__ & ~new_new_n14535__;
  assign new_new_n14538__ = ~new_new_n14536__ & ~new_new_n14537__;
  assign new_new_n14539__ = pi108 & ~new_new_n14538__;
  assign new_new_n14540__ = ~pi108 & new_new_n14538__;
  assign new_new_n14541__ = ~new_new_n13996__ & ~new_new_n13997__;
  assign new_new_n14542__ = ~new_new_n14464__ & po014;
  assign new_new_n14543__ = ~pi106 & ~po014;
  assign new_new_n14544__ = ~new_new_n14542__ & ~new_new_n14543__;
  assign new_new_n14545__ = new_new_n14541__ & ~new_new_n14544__;
  assign new_new_n14546__ = ~new_new_n14541__ & new_new_n14544__;
  assign new_new_n14547__ = ~new_new_n14545__ & ~new_new_n14546__;
  assign new_new_n14548__ = ~pi107 & new_new_n14547__;
  assign new_new_n14549__ = pi107 & ~new_new_n14547__;
  assign new_new_n14550__ = ~pi105 & ~new_new_n14462__;
  assign new_new_n14551__ = pi105 & new_new_n14462__;
  assign new_new_n14552__ = ~new_new_n14550__ & ~new_new_n14551__;
  assign new_new_n14553__ = po014 & new_new_n14552__;
  assign new_new_n14554__ = new_new_n14004__ & new_new_n14553__;
  assign new_new_n14555__ = ~new_new_n14004__ & ~new_new_n14553__;
  assign new_new_n14556__ = ~new_new_n14554__ & ~new_new_n14555__;
  assign new_new_n14557__ = ~pi106 & ~new_new_n14556__;
  assign new_new_n14558__ = pi106 & new_new_n14556__;
  assign new_new_n14559__ = ~new_new_n14023__ & ~new_new_n14024__;
  assign new_new_n14560__ = ~new_new_n14458__ & po014;
  assign new_new_n14561__ = pi103 & ~po014;
  assign new_new_n14562__ = ~new_new_n14560__ & ~new_new_n14561__;
  assign new_new_n14563__ = new_new_n14559__ & new_new_n14562__;
  assign new_new_n14564__ = ~new_new_n14559__ & ~new_new_n14562__;
  assign new_new_n14565__ = ~new_new_n14563__ & ~new_new_n14564__;
  assign new_new_n14566__ = pi104 & ~new_new_n14565__;
  assign new_new_n14567__ = ~pi104 & new_new_n14565__;
  assign new_new_n14568__ = pi102 & ~new_new_n14456__;
  assign new_new_n14569__ = ~pi102 & new_new_n14456__;
  assign new_new_n14570__ = ~new_new_n14568__ & ~new_new_n14569__;
  assign new_new_n14571__ = po014 & new_new_n14570__;
  assign new_new_n14572__ = new_new_n14031__ & new_new_n14571__;
  assign new_new_n14573__ = ~new_new_n14031__ & ~new_new_n14571__;
  assign new_new_n14574__ = ~new_new_n14572__ & ~new_new_n14573__;
  assign new_new_n14575__ = pi103 & ~new_new_n14574__;
  assign new_new_n14576__ = ~pi103 & new_new_n14574__;
  assign new_new_n14577__ = ~new_new_n14041__ & ~new_new_n14042__;
  assign new_new_n14578__ = ~new_new_n14454__ & po014;
  assign new_new_n14579__ = pi101 & ~po014;
  assign new_new_n14580__ = ~new_new_n14578__ & ~new_new_n14579__;
  assign new_new_n14581__ = new_new_n14577__ & new_new_n14580__;
  assign new_new_n14582__ = ~new_new_n14577__ & ~new_new_n14580__;
  assign new_new_n14583__ = ~new_new_n14581__ & ~new_new_n14582__;
  assign new_new_n14584__ = pi102 & ~new_new_n14583__;
  assign new_new_n14585__ = ~pi102 & new_new_n14583__;
  assign new_new_n14586__ = new_new_n14452__ & po014;
  assign new_new_n14587__ = pi100 & ~po014;
  assign new_new_n14588__ = ~new_new_n14586__ & ~new_new_n14587__;
  assign new_new_n14589__ = ~new_new_n14050__ & ~new_new_n14051__;
  assign new_new_n14590__ = ~new_new_n14588__ & ~new_new_n14589__;
  assign new_new_n14591__ = new_new_n14588__ & new_new_n14589__;
  assign new_new_n14592__ = ~new_new_n14590__ & ~new_new_n14591__;
  assign new_new_n14593__ = pi101 & ~new_new_n14592__;
  assign new_new_n14594__ = ~pi101 & new_new_n14592__;
  assign new_new_n14595__ = ~new_new_n14059__ & ~new_new_n14060__;
  assign new_new_n14596__ = ~new_new_n14450__ & po014;
  assign new_new_n14597__ = ~pi099 & ~po014;
  assign new_new_n14598__ = ~new_new_n14596__ & ~new_new_n14597__;
  assign new_new_n14599__ = new_new_n14595__ & ~new_new_n14598__;
  assign new_new_n14600__ = ~new_new_n14595__ & new_new_n14598__;
  assign new_new_n14601__ = ~new_new_n14599__ & ~new_new_n14600__;
  assign new_new_n14602__ = pi100 & ~new_new_n14601__;
  assign new_new_n14603__ = ~pi100 & new_new_n14601__;
  assign new_new_n14604__ = ~pi098 & ~new_new_n14448__;
  assign new_new_n14605__ = pi098 & new_new_n14448__;
  assign new_new_n14606__ = ~new_new_n14604__ & ~new_new_n14605__;
  assign new_new_n14607__ = po014 & new_new_n14606__;
  assign new_new_n14608__ = new_new_n14067__ & new_new_n14607__;
  assign new_new_n14609__ = ~new_new_n14067__ & ~new_new_n14607__;
  assign new_new_n14610__ = ~new_new_n14608__ & ~new_new_n14609__;
  assign new_new_n14611__ = ~pi099 & ~new_new_n14610__;
  assign new_new_n14612__ = pi099 & new_new_n14610__;
  assign new_new_n14613__ = ~pi097 & ~new_new_n14446__;
  assign new_new_n14614__ = pi097 & new_new_n14446__;
  assign new_new_n14615__ = ~new_new_n14613__ & ~new_new_n14614__;
  assign new_new_n14616__ = po014 & new_new_n14615__;
  assign new_new_n14617__ = ~new_new_n14076__ & new_new_n14616__;
  assign new_new_n14618__ = new_new_n14076__ & ~new_new_n14616__;
  assign new_new_n14619__ = ~new_new_n14617__ & ~new_new_n14618__;
  assign new_new_n14620__ = pi098 & ~new_new_n14619__;
  assign new_new_n14621__ = ~pi098 & new_new_n14619__;
  assign new_new_n14622__ = ~new_new_n14086__ & ~new_new_n14087__;
  assign new_new_n14623__ = ~new_new_n14444__ & po014;
  assign new_new_n14624__ = ~pi096 & ~po014;
  assign new_new_n14625__ = ~new_new_n14623__ & ~new_new_n14624__;
  assign new_new_n14626__ = new_new_n14622__ & ~new_new_n14625__;
  assign new_new_n14627__ = ~new_new_n14622__ & new_new_n14625__;
  assign new_new_n14628__ = ~new_new_n14626__ & ~new_new_n14627__;
  assign new_new_n14629__ = pi097 & ~new_new_n14628__;
  assign new_new_n14630__ = ~pi097 & new_new_n14628__;
  assign new_new_n14631__ = ~pi095 & ~new_new_n14442__;
  assign new_new_n14632__ = pi095 & new_new_n14442__;
  assign new_new_n14633__ = ~new_new_n14631__ & ~new_new_n14632__;
  assign new_new_n14634__ = po014 & new_new_n14633__;
  assign new_new_n14635__ = ~new_new_n14094__ & new_new_n14634__;
  assign new_new_n14636__ = new_new_n14094__ & ~new_new_n14634__;
  assign new_new_n14637__ = ~new_new_n14635__ & ~new_new_n14636__;
  assign new_new_n14638__ = pi096 & ~new_new_n14637__;
  assign new_new_n14639__ = ~pi096 & new_new_n14637__;
  assign new_new_n14640__ = ~new_new_n14113__ & ~new_new_n14114__;
  assign new_new_n14641__ = ~new_new_n14438__ & po014;
  assign new_new_n14642__ = pi093 & ~po014;
  assign new_new_n14643__ = ~new_new_n14641__ & ~new_new_n14642__;
  assign new_new_n14644__ = new_new_n14640__ & ~new_new_n14643__;
  assign new_new_n14645__ = ~new_new_n14640__ & new_new_n14643__;
  assign new_new_n14646__ = ~new_new_n14644__ & ~new_new_n14645__;
  assign new_new_n14647__ = pi094 & new_new_n14646__;
  assign new_new_n14648__ = ~pi094 & ~new_new_n14646__;
  assign new_new_n14649__ = ~new_new_n14122__ & ~new_new_n14123__;
  assign new_new_n14650__ = ~new_new_n14436__ & po014;
  assign new_new_n14651__ = ~pi092 & ~po014;
  assign new_new_n14652__ = ~new_new_n14650__ & ~new_new_n14651__;
  assign new_new_n14653__ = new_new_n14649__ & ~new_new_n14652__;
  assign new_new_n14654__ = ~new_new_n14649__ & new_new_n14652__;
  assign new_new_n14655__ = ~new_new_n14653__ & ~new_new_n14654__;
  assign new_new_n14656__ = pi093 & ~new_new_n14655__;
  assign new_new_n14657__ = ~pi093 & new_new_n14655__;
  assign new_new_n14658__ = ~new_new_n14131__ & ~new_new_n14132__;
  assign new_new_n14659__ = ~new_new_n14434__ & po014;
  assign new_new_n14660__ = ~pi091 & ~po014;
  assign new_new_n14661__ = ~new_new_n14659__ & ~new_new_n14660__;
  assign new_new_n14662__ = new_new_n14658__ & ~new_new_n14661__;
  assign new_new_n14663__ = ~new_new_n14658__ & new_new_n14661__;
  assign new_new_n14664__ = ~new_new_n14662__ & ~new_new_n14663__;
  assign new_new_n14665__ = pi092 & ~new_new_n14664__;
  assign new_new_n14666__ = ~pi092 & new_new_n14664__;
  assign new_new_n14667__ = ~new_new_n14140__ & ~new_new_n14141__;
  assign new_new_n14668__ = ~new_new_n14432__ & po014;
  assign new_new_n14669__ = ~pi090 & ~po014;
  assign new_new_n14670__ = ~new_new_n14668__ & ~new_new_n14669__;
  assign new_new_n14671__ = new_new_n14667__ & ~new_new_n14670__;
  assign new_new_n14672__ = ~new_new_n14667__ & new_new_n14670__;
  assign new_new_n14673__ = ~new_new_n14671__ & ~new_new_n14672__;
  assign new_new_n14674__ = pi091 & ~new_new_n14673__;
  assign new_new_n14675__ = ~pi091 & new_new_n14673__;
  assign new_new_n14676__ = ~new_new_n14149__ & ~new_new_n14150__;
  assign new_new_n14677__ = ~new_new_n14430__ & po014;
  assign new_new_n14678__ = ~pi089 & ~po014;
  assign new_new_n14679__ = ~new_new_n14677__ & ~new_new_n14678__;
  assign new_new_n14680__ = new_new_n14676__ & ~new_new_n14679__;
  assign new_new_n14681__ = ~new_new_n14676__ & new_new_n14679__;
  assign new_new_n14682__ = ~new_new_n14680__ & ~new_new_n14681__;
  assign new_new_n14683__ = pi090 & ~new_new_n14682__;
  assign new_new_n14684__ = ~pi090 & new_new_n14682__;
  assign new_new_n14685__ = ~pi088 & ~new_new_n14428__;
  assign new_new_n14686__ = pi088 & new_new_n14428__;
  assign new_new_n14687__ = ~new_new_n14685__ & ~new_new_n14686__;
  assign new_new_n14688__ = po014 & new_new_n14687__;
  assign new_new_n14689__ = new_new_n14157__ & new_new_n14688__;
  assign new_new_n14690__ = ~new_new_n14157__ & ~new_new_n14688__;
  assign new_new_n14691__ = ~new_new_n14689__ & ~new_new_n14690__;
  assign new_new_n14692__ = ~pi089 & ~new_new_n14691__;
  assign new_new_n14693__ = pi089 & new_new_n14691__;
  assign new_new_n14694__ = ~new_new_n14167__ & ~new_new_n14168__;
  assign new_new_n14695__ = new_new_n14426__ & po014;
  assign new_new_n14696__ = ~pi087 & ~po014;
  assign new_new_n14697__ = ~new_new_n14695__ & ~new_new_n14696__;
  assign new_new_n14698__ = ~new_new_n14694__ & ~new_new_n14697__;
  assign new_new_n14699__ = new_new_n14694__ & new_new_n14697__;
  assign new_new_n14700__ = ~new_new_n14698__ & ~new_new_n14699__;
  assign new_new_n14701__ = ~pi088 & ~new_new_n14700__;
  assign new_new_n14702__ = pi088 & new_new_n14700__;
  assign new_new_n14703__ = new_new_n14424__ & po014;
  assign new_new_n14704__ = ~pi086 & ~po014;
  assign new_new_n14705__ = ~new_new_n14703__ & ~new_new_n14704__;
  assign new_new_n14706__ = ~new_new_n14176__ & ~new_new_n14177__;
  assign new_new_n14707__ = ~new_new_n14705__ & ~new_new_n14706__;
  assign new_new_n14708__ = new_new_n14705__ & new_new_n14706__;
  assign new_new_n14709__ = ~new_new_n14707__ & ~new_new_n14708__;
  assign new_new_n14710__ = ~pi087 & ~new_new_n14709__;
  assign new_new_n14711__ = pi087 & new_new_n14709__;
  assign new_new_n14712__ = ~new_new_n14422__ & po014;
  assign new_new_n14713__ = pi085 & ~po014;
  assign new_new_n14714__ = ~new_new_n14712__ & ~new_new_n14713__;
  assign new_new_n14715__ = ~new_new_n14185__ & ~new_new_n14186__;
  assign new_new_n14716__ = ~new_new_n14714__ & new_new_n14715__;
  assign new_new_n14717__ = new_new_n14714__ & ~new_new_n14715__;
  assign new_new_n14718__ = ~new_new_n14716__ & ~new_new_n14717__;
  assign new_new_n14719__ = pi086 & new_new_n14718__;
  assign new_new_n14720__ = ~pi086 & ~new_new_n14718__;
  assign new_new_n14721__ = pi084 & ~new_new_n14420__;
  assign new_new_n14722__ = ~pi084 & new_new_n14420__;
  assign new_new_n14723__ = ~new_new_n14721__ & ~new_new_n14722__;
  assign new_new_n14724__ = po014 & new_new_n14723__;
  assign new_new_n14725__ = new_new_n14193__ & new_new_n14724__;
  assign new_new_n14726__ = ~new_new_n14193__ & ~new_new_n14724__;
  assign new_new_n14727__ = ~new_new_n14725__ & ~new_new_n14726__;
  assign new_new_n14728__ = pi085 & ~new_new_n14727__;
  assign new_new_n14729__ = ~pi085 & new_new_n14727__;
  assign new_new_n14730__ = ~new_new_n14203__ & ~new_new_n14204__;
  assign new_new_n14731__ = ~new_new_n14418__ & po014;
  assign new_new_n14732__ = ~pi083 & ~po014;
  assign new_new_n14733__ = ~new_new_n14731__ & ~new_new_n14732__;
  assign new_new_n14734__ = new_new_n14730__ & ~new_new_n14733__;
  assign new_new_n14735__ = ~new_new_n14730__ & new_new_n14733__;
  assign new_new_n14736__ = ~new_new_n14734__ & ~new_new_n14735__;
  assign new_new_n14737__ = pi084 & ~new_new_n14736__;
  assign new_new_n14738__ = ~pi084 & new_new_n14736__;
  assign new_new_n14739__ = ~new_new_n14212__ & ~new_new_n14213__;
  assign new_new_n14740__ = ~new_new_n14416__ & po014;
  assign new_new_n14741__ = pi082 & ~po014;
  assign new_new_n14742__ = ~new_new_n14740__ & ~new_new_n14741__;
  assign new_new_n14743__ = new_new_n14739__ & ~new_new_n14742__;
  assign new_new_n14744__ = ~new_new_n14739__ & new_new_n14742__;
  assign new_new_n14745__ = ~new_new_n14743__ & ~new_new_n14744__;
  assign new_new_n14746__ = ~pi083 & ~new_new_n14745__;
  assign new_new_n14747__ = pi083 & new_new_n14745__;
  assign new_new_n14748__ = ~new_new_n14221__ & ~new_new_n14222__;
  assign new_new_n14749__ = ~new_new_n14414__ & po014;
  assign new_new_n14750__ = pi081 & ~po014;
  assign new_new_n14751__ = ~new_new_n14749__ & ~new_new_n14750__;
  assign new_new_n14752__ = new_new_n14748__ & ~new_new_n14751__;
  assign new_new_n14753__ = ~new_new_n14748__ & new_new_n14751__;
  assign new_new_n14754__ = ~new_new_n14752__ & ~new_new_n14753__;
  assign new_new_n14755__ = ~pi082 & ~new_new_n14754__;
  assign new_new_n14756__ = pi082 & new_new_n14754__;
  assign new_new_n14757__ = ~new_new_n14230__ & ~new_new_n14231__;
  assign new_new_n14758__ = pi080 & ~po014;
  assign new_new_n14759__ = ~new_new_n14412__ & po014;
  assign new_new_n14760__ = ~new_new_n14758__ & ~new_new_n14759__;
  assign new_new_n14761__ = new_new_n14757__ & new_new_n14760__;
  assign new_new_n14762__ = ~new_new_n14757__ & ~new_new_n14760__;
  assign new_new_n14763__ = ~new_new_n14761__ & ~new_new_n14762__;
  assign new_new_n14764__ = pi081 & ~new_new_n14763__;
  assign new_new_n14765__ = ~pi081 & new_new_n14763__;
  assign new_new_n14766__ = ~new_new_n14239__ & ~new_new_n14240__;
  assign new_new_n14767__ = ~new_new_n14410__ & po014;
  assign new_new_n14768__ = pi079 & ~po014;
  assign new_new_n14769__ = ~new_new_n14767__ & ~new_new_n14768__;
  assign new_new_n14770__ = new_new_n14766__ & ~new_new_n14769__;
  assign new_new_n14771__ = ~new_new_n14766__ & new_new_n14769__;
  assign new_new_n14772__ = ~new_new_n14770__ & ~new_new_n14771__;
  assign new_new_n14773__ = ~pi080 & ~new_new_n14772__;
  assign new_new_n14774__ = pi080 & new_new_n14772__;
  assign new_new_n14775__ = ~new_new_n14248__ & ~new_new_n14249__;
  assign new_new_n14776__ = pi078 & ~po014;
  assign new_new_n14777__ = ~new_new_n14408__ & po014;
  assign new_new_n14778__ = ~new_new_n14776__ & ~new_new_n14777__;
  assign new_new_n14779__ = new_new_n14775__ & new_new_n14778__;
  assign new_new_n14780__ = ~new_new_n14775__ & ~new_new_n14778__;
  assign new_new_n14781__ = ~new_new_n14779__ & ~new_new_n14780__;
  assign new_new_n14782__ = ~pi079 & new_new_n14781__;
  assign new_new_n14783__ = pi079 & ~new_new_n14781__;
  assign new_new_n14784__ = ~new_new_n14257__ & ~new_new_n14258__;
  assign new_new_n14785__ = ~new_new_n14406__ & po014;
  assign new_new_n14786__ = pi077 & ~po014;
  assign new_new_n14787__ = ~new_new_n14785__ & ~new_new_n14786__;
  assign new_new_n14788__ = new_new_n14784__ & ~new_new_n14787__;
  assign new_new_n14789__ = ~new_new_n14784__ & new_new_n14787__;
  assign new_new_n14790__ = ~new_new_n14788__ & ~new_new_n14789__;
  assign new_new_n14791__ = ~pi078 & ~new_new_n14790__;
  assign new_new_n14792__ = pi078 & new_new_n14790__;
  assign new_new_n14793__ = ~new_new_n14404__ & po014;
  assign new_new_n14794__ = pi076 & ~po014;
  assign new_new_n14795__ = ~new_new_n14793__ & ~new_new_n14794__;
  assign new_new_n14796__ = ~new_new_n14266__ & ~new_new_n14267__;
  assign new_new_n14797__ = ~new_new_n14795__ & new_new_n14796__;
  assign new_new_n14798__ = new_new_n14795__ & ~new_new_n14796__;
  assign new_new_n14799__ = ~new_new_n14797__ & ~new_new_n14798__;
  assign new_new_n14800__ = pi077 & new_new_n14799__;
  assign new_new_n14801__ = ~pi077 & ~new_new_n14799__;
  assign new_new_n14802__ = ~new_new_n14275__ & ~new_new_n14276__;
  assign new_new_n14803__ = ~new_new_n14402__ & po014;
  assign new_new_n14804__ = ~pi075 & ~po014;
  assign new_new_n14805__ = ~new_new_n14803__ & ~new_new_n14804__;
  assign new_new_n14806__ = new_new_n14802__ & ~new_new_n14805__;
  assign new_new_n14807__ = ~new_new_n14802__ & new_new_n14805__;
  assign new_new_n14808__ = ~new_new_n14806__ & ~new_new_n14807__;
  assign new_new_n14809__ = pi076 & ~new_new_n14808__;
  assign new_new_n14810__ = ~pi076 & new_new_n14808__;
  assign new_new_n14811__ = ~new_new_n14284__ & ~new_new_n14285__;
  assign new_new_n14812__ = ~new_new_n14400__ & po014;
  assign new_new_n14813__ = ~pi074 & ~po014;
  assign new_new_n14814__ = ~new_new_n14812__ & ~new_new_n14813__;
  assign new_new_n14815__ = new_new_n14811__ & ~new_new_n14814__;
  assign new_new_n14816__ = ~new_new_n14811__ & new_new_n14814__;
  assign new_new_n14817__ = ~new_new_n14815__ & ~new_new_n14816__;
  assign new_new_n14818__ = pi075 & ~new_new_n14817__;
  assign new_new_n14819__ = ~pi075 & new_new_n14817__;
  assign new_new_n14820__ = ~new_new_n14293__ & ~new_new_n14294__;
  assign new_new_n14821__ = ~new_new_n14398__ & po014;
  assign new_new_n14822__ = ~pi073 & ~po014;
  assign new_new_n14823__ = ~new_new_n14821__ & ~new_new_n14822__;
  assign new_new_n14824__ = ~new_new_n14820__ & ~new_new_n14823__;
  assign new_new_n14825__ = new_new_n14820__ & new_new_n14823__;
  assign new_new_n14826__ = ~new_new_n14824__ & ~new_new_n14825__;
  assign new_new_n14827__ = ~pi074 & ~new_new_n14826__;
  assign new_new_n14828__ = pi074 & new_new_n14826__;
  assign new_new_n14829__ = ~pi072 & ~new_new_n14396__;
  assign new_new_n14830__ = pi072 & new_new_n14396__;
  assign new_new_n14831__ = ~new_new_n14829__ & ~new_new_n14830__;
  assign new_new_n14832__ = po014 & new_new_n14831__;
  assign new_new_n14833__ = ~new_new_n14301__ & ~new_new_n14832__;
  assign new_new_n14834__ = new_new_n14301__ & new_new_n14832__;
  assign new_new_n14835__ = ~new_new_n14833__ & ~new_new_n14834__;
  assign new_new_n14836__ = ~pi073 & ~new_new_n14835__;
  assign new_new_n14837__ = pi073 & new_new_n14835__;
  assign new_new_n14838__ = new_new_n14394__ & po014;
  assign new_new_n14839__ = ~pi071 & ~po014;
  assign new_new_n14840__ = ~new_new_n14838__ & ~new_new_n14839__;
  assign new_new_n14841__ = ~new_new_n14309__ & ~new_new_n14310__;
  assign new_new_n14842__ = ~new_new_n14840__ & ~new_new_n14841__;
  assign new_new_n14843__ = new_new_n14840__ & new_new_n14841__;
  assign new_new_n14844__ = ~new_new_n14842__ & ~new_new_n14843__;
  assign new_new_n14845__ = ~pi072 & ~new_new_n14844__;
  assign new_new_n14846__ = pi072 & new_new_n14844__;
  assign new_new_n14847__ = ~new_new_n14318__ & ~new_new_n14319__;
  assign new_new_n14848__ = ~new_new_n14392__ & po014;
  assign new_new_n14849__ = pi070 & ~po014;
  assign new_new_n14850__ = ~new_new_n14848__ & ~new_new_n14849__;
  assign new_new_n14851__ = new_new_n14847__ & ~new_new_n14850__;
  assign new_new_n14852__ = ~new_new_n14847__ & new_new_n14850__;
  assign new_new_n14853__ = ~new_new_n14851__ & ~new_new_n14852__;
  assign new_new_n14854__ = ~pi071 & ~new_new_n14853__;
  assign new_new_n14855__ = pi071 & new_new_n14853__;
  assign new_new_n14856__ = ~new_new_n14336__ & ~new_new_n14337__;
  assign new_new_n14857__ = ~new_new_n14388__ & po014;
  assign new_new_n14858__ = ~pi068 & ~po014;
  assign new_new_n14859__ = ~new_new_n14857__ & ~new_new_n14858__;
  assign new_new_n14860__ = new_new_n14856__ & ~new_new_n14859__;
  assign new_new_n14861__ = ~new_new_n14856__ & new_new_n14859__;
  assign new_new_n14862__ = ~new_new_n14860__ & ~new_new_n14861__;
  assign new_new_n14863__ = pi069 & ~new_new_n14862__;
  assign new_new_n14864__ = ~pi069 & new_new_n14862__;
  assign new_new_n14865__ = pi065 & new_new_n14345__;
  assign new_new_n14866__ = pi015 & new_new_n14347__;
  assign new_new_n14867__ = ~new_new_n14348__ & ~new_new_n14866__;
  assign new_new_n14868__ = ~new_new_n14346__ & ~new_new_n14867__;
  assign new_new_n14869__ = ~new_new_n14865__ & ~new_new_n14868__;
  assign new_new_n14870__ = pi066 & ~new_new_n14869__;
  assign new_new_n14871__ = ~pi066 & new_new_n14869__;
  assign new_new_n14872__ = ~new_new_n14870__ & ~new_new_n14871__;
  assign new_new_n14873__ = po014 & new_new_n14872__;
  assign new_new_n14874__ = ~new_new_n14384__ & new_new_n14873__;
  assign new_new_n14875__ = new_new_n14384__ & ~new_new_n14873__;
  assign new_new_n14876__ = ~new_new_n14874__ & ~new_new_n14875__;
  assign new_new_n14877__ = ~pi067 & ~new_new_n14876__;
  assign new_new_n14878__ = pi067 & new_new_n14876__;
  assign new_new_n14879__ = pi013 & ~pi065;
  assign new_new_n14880__ = pi014 & po014;
  assign new_new_n14881__ = pi065 & new_new_n14867__;
  assign new_new_n14882__ = ~pi065 & ~new_new_n14867__;
  assign new_new_n14883__ = ~new_new_n14881__ & ~new_new_n14882__;
  assign new_new_n14884__ = ~new_new_n14879__ & ~new_new_n14883__;
  assign new_new_n14885__ = new_new_n14880__ & new_new_n14884__;
  assign new_new_n14886__ = ~new_new_n14350__ & po014;
  assign new_new_n14887__ = ~pi013 & ~new_new_n14351__;
  assign new_new_n14888__ = ~new_new_n14867__ & new_new_n14887__;
  assign new_new_n14889__ = ~new_new_n14886__ & new_new_n14888__;
  assign new_new_n14890__ = ~new_new_n14885__ & ~new_new_n14889__;
  assign new_new_n14891__ = pi064 & ~new_new_n14890__;
  assign new_new_n14892__ = pi064 & po014;
  assign new_new_n14893__ = new_new_n14350__ & ~new_new_n14892__;
  assign new_new_n14894__ = ~po014 & ~new_new_n14867__;
  assign new_new_n14895__ = po014 & new_new_n14867__;
  assign new_new_n14896__ = ~new_new_n14894__ & ~new_new_n14895__;
  assign new_new_n14897__ = new_new_n14893__ & ~new_new_n14896__;
  assign new_new_n14898__ = ~pi066 & ~new_new_n14897__;
  assign new_new_n14899__ = ~new_new_n14891__ & new_new_n14898__;
  assign new_new_n14900__ = ~pi013 & pi065;
  assign new_new_n14901__ = new_new_n14345__ & ~new_new_n14900__;
  assign new_new_n14902__ = ~new_new_n14883__ & new_new_n14901__;
  assign new_new_n14903__ = pi014 & new_new_n403__;
  assign new_new_n14904__ = ~new_new_n14867__ & new_new_n14903__;
  assign new_new_n14905__ = ~new_new_n14902__ & ~new_new_n14904__;
  assign new_new_n14906__ = po014 & ~new_new_n14905__;
  assign new_new_n14907__ = pi065 & po014;
  assign new_new_n14908__ = pi013 & ~new_new_n14907__;
  assign new_new_n14909__ = ~pi065 & ~po014;
  assign new_new_n14910__ = ~pi014 & ~new_new_n14909__;
  assign new_new_n14911__ = new_new_n14908__ & ~new_new_n14910__;
  assign new_new_n14912__ = pi014 & ~new_new_n426__;
  assign new_new_n14913__ = ~po014 & new_new_n14912__;
  assign new_new_n14914__ = ~new_new_n332__ & ~new_new_n14913__;
  assign new_new_n14915__ = ~new_new_n14911__ & new_new_n14914__;
  assign new_new_n14916__ = new_new_n14867__ & ~new_new_n14915__;
  assign new_new_n14917__ = ~new_new_n14899__ & ~new_new_n14906__;
  assign new_new_n14918__ = ~new_new_n14916__ & new_new_n14917__;
  assign new_new_n14919__ = ~new_new_n14878__ & ~new_new_n14918__;
  assign new_new_n14920__ = ~new_new_n14877__ & ~new_new_n14919__;
  assign new_new_n14921__ = pi068 & new_new_n14920__;
  assign new_new_n14922__ = ~pi068 & ~new_new_n14920__;
  assign new_new_n14923__ = ~new_new_n14343__ & ~new_new_n14344__;
  assign new_new_n14924__ = new_new_n14386__ & po014;
  assign new_new_n14925__ = ~pi067 & ~po014;
  assign new_new_n14926__ = ~new_new_n14924__ & ~new_new_n14925__;
  assign new_new_n14927__ = ~new_new_n14923__ & ~new_new_n14926__;
  assign new_new_n14928__ = new_new_n14923__ & new_new_n14926__;
  assign new_new_n14929__ = ~new_new_n14927__ & ~new_new_n14928__;
  assign new_new_n14930__ = ~new_new_n14922__ & new_new_n14929__;
  assign new_new_n14931__ = ~new_new_n14921__ & ~new_new_n14930__;
  assign new_new_n14932__ = ~new_new_n14864__ & ~new_new_n14931__;
  assign new_new_n14933__ = ~new_new_n14863__ & ~new_new_n14932__;
  assign new_new_n14934__ = ~pi070 & new_new_n14933__;
  assign new_new_n14935__ = pi070 & ~new_new_n14933__;
  assign new_new_n14936__ = ~new_new_n14327__ & ~new_new_n14328__;
  assign new_new_n14937__ = ~new_new_n14390__ & po014;
  assign new_new_n14938__ = ~pi069 & ~po014;
  assign new_new_n14939__ = ~new_new_n14937__ & ~new_new_n14938__;
  assign new_new_n14940__ = new_new_n14936__ & ~new_new_n14939__;
  assign new_new_n14941__ = ~new_new_n14936__ & new_new_n14939__;
  assign new_new_n14942__ = ~new_new_n14940__ & ~new_new_n14941__;
  assign new_new_n14943__ = ~new_new_n14935__ & new_new_n14942__;
  assign new_new_n14944__ = ~new_new_n14934__ & ~new_new_n14943__;
  assign new_new_n14945__ = ~new_new_n14855__ & ~new_new_n14944__;
  assign new_new_n14946__ = ~new_new_n14854__ & ~new_new_n14945__;
  assign new_new_n14947__ = ~new_new_n14846__ & ~new_new_n14946__;
  assign new_new_n14948__ = ~new_new_n14845__ & ~new_new_n14947__;
  assign new_new_n14949__ = ~new_new_n14837__ & ~new_new_n14948__;
  assign new_new_n14950__ = ~new_new_n14836__ & ~new_new_n14949__;
  assign new_new_n14951__ = ~new_new_n14828__ & ~new_new_n14950__;
  assign new_new_n14952__ = ~new_new_n14827__ & ~new_new_n14951__;
  assign new_new_n14953__ = ~new_new_n14819__ & new_new_n14952__;
  assign new_new_n14954__ = ~new_new_n14818__ & ~new_new_n14953__;
  assign new_new_n14955__ = ~new_new_n14810__ & ~new_new_n14954__;
  assign new_new_n14956__ = ~new_new_n14809__ & ~new_new_n14955__;
  assign new_new_n14957__ = ~new_new_n14801__ & ~new_new_n14956__;
  assign new_new_n14958__ = ~new_new_n14800__ & ~new_new_n14957__;
  assign new_new_n14959__ = ~new_new_n14792__ & new_new_n14958__;
  assign new_new_n14960__ = ~new_new_n14791__ & ~new_new_n14959__;
  assign new_new_n14961__ = ~new_new_n14783__ & ~new_new_n14960__;
  assign new_new_n14962__ = ~new_new_n14782__ & ~new_new_n14961__;
  assign new_new_n14963__ = ~new_new_n14774__ & ~new_new_n14962__;
  assign new_new_n14964__ = ~new_new_n14773__ & ~new_new_n14963__;
  assign new_new_n14965__ = ~new_new_n14765__ & new_new_n14964__;
  assign new_new_n14966__ = ~new_new_n14764__ & ~new_new_n14965__;
  assign new_new_n14967__ = ~new_new_n14756__ & new_new_n14966__;
  assign new_new_n14968__ = ~new_new_n14755__ & ~new_new_n14967__;
  assign new_new_n14969__ = ~new_new_n14747__ & ~new_new_n14968__;
  assign new_new_n14970__ = ~new_new_n14746__ & ~new_new_n14969__;
  assign new_new_n14971__ = ~new_new_n14738__ & new_new_n14970__;
  assign new_new_n14972__ = ~new_new_n14737__ & ~new_new_n14971__;
  assign new_new_n14973__ = ~new_new_n14729__ & ~new_new_n14972__;
  assign new_new_n14974__ = ~new_new_n14728__ & ~new_new_n14973__;
  assign new_new_n14975__ = ~new_new_n14720__ & ~new_new_n14974__;
  assign new_new_n14976__ = ~new_new_n14719__ & ~new_new_n14975__;
  assign new_new_n14977__ = ~new_new_n14711__ & new_new_n14976__;
  assign new_new_n14978__ = ~new_new_n14710__ & ~new_new_n14977__;
  assign new_new_n14979__ = ~new_new_n14702__ & ~new_new_n14978__;
  assign new_new_n14980__ = ~new_new_n14701__ & ~new_new_n14979__;
  assign new_new_n14981__ = ~new_new_n14693__ & ~new_new_n14980__;
  assign new_new_n14982__ = ~new_new_n14692__ & ~new_new_n14981__;
  assign new_new_n14983__ = ~new_new_n14684__ & new_new_n14982__;
  assign new_new_n14984__ = ~new_new_n14683__ & ~new_new_n14983__;
  assign new_new_n14985__ = ~new_new_n14675__ & ~new_new_n14984__;
  assign new_new_n14986__ = ~new_new_n14674__ & ~new_new_n14985__;
  assign new_new_n14987__ = ~new_new_n14666__ & ~new_new_n14986__;
  assign new_new_n14988__ = ~new_new_n14665__ & ~new_new_n14987__;
  assign new_new_n14989__ = ~new_new_n14657__ & ~new_new_n14988__;
  assign new_new_n14990__ = ~new_new_n14656__ & ~new_new_n14989__;
  assign new_new_n14991__ = ~new_new_n14648__ & ~new_new_n14990__;
  assign new_new_n14992__ = ~new_new_n14647__ & ~new_new_n14991__;
  assign new_new_n14993__ = ~pi095 & new_new_n14992__;
  assign new_new_n14994__ = pi095 & ~new_new_n14992__;
  assign new_new_n14995__ = ~pi094 & ~new_new_n14440__;
  assign new_new_n14996__ = pi094 & new_new_n14440__;
  assign new_new_n14997__ = ~new_new_n14995__ & ~new_new_n14996__;
  assign new_new_n14998__ = po014 & new_new_n14997__;
  assign new_new_n14999__ = ~new_new_n14103__ & new_new_n14998__;
  assign new_new_n15000__ = new_new_n14103__ & ~new_new_n14998__;
  assign new_new_n15001__ = ~new_new_n14999__ & ~new_new_n15000__;
  assign new_new_n15002__ = ~new_new_n14994__ & new_new_n15001__;
  assign new_new_n15003__ = ~new_new_n14993__ & ~new_new_n15002__;
  assign new_new_n15004__ = ~new_new_n14639__ & new_new_n15003__;
  assign new_new_n15005__ = ~new_new_n14638__ & ~new_new_n15004__;
  assign new_new_n15006__ = ~new_new_n14630__ & ~new_new_n15005__;
  assign new_new_n15007__ = ~new_new_n14629__ & ~new_new_n15006__;
  assign new_new_n15008__ = ~new_new_n14621__ & ~new_new_n15007__;
  assign new_new_n15009__ = ~new_new_n14620__ & ~new_new_n15008__;
  assign new_new_n15010__ = ~new_new_n14612__ & new_new_n15009__;
  assign new_new_n15011__ = ~new_new_n14611__ & ~new_new_n15010__;
  assign new_new_n15012__ = ~new_new_n14603__ & new_new_n15011__;
  assign new_new_n15013__ = ~new_new_n14602__ & ~new_new_n15012__;
  assign new_new_n15014__ = ~new_new_n14594__ & ~new_new_n15013__;
  assign new_new_n15015__ = ~new_new_n14593__ & ~new_new_n15014__;
  assign new_new_n15016__ = ~new_new_n14585__ & ~new_new_n15015__;
  assign new_new_n15017__ = ~new_new_n14584__ & ~new_new_n15016__;
  assign new_new_n15018__ = ~new_new_n14576__ & ~new_new_n15017__;
  assign new_new_n15019__ = ~new_new_n14575__ & ~new_new_n15018__;
  assign new_new_n15020__ = ~new_new_n14567__ & ~new_new_n15019__;
  assign new_new_n15021__ = ~new_new_n14566__ & ~new_new_n15020__;
  assign new_new_n15022__ = ~pi105 & new_new_n15021__;
  assign new_new_n15023__ = pi105 & ~new_new_n15021__;
  assign new_new_n15024__ = ~new_new_n14460__ & po014;
  assign new_new_n15025__ = pi104 & ~po014;
  assign new_new_n15026__ = ~new_new_n15024__ & ~new_new_n15025__;
  assign new_new_n15027__ = ~new_new_n14014__ & ~new_new_n14015__;
  assign new_new_n15028__ = ~new_new_n15026__ & new_new_n15027__;
  assign new_new_n15029__ = new_new_n15026__ & ~new_new_n15027__;
  assign new_new_n15030__ = ~new_new_n15028__ & ~new_new_n15029__;
  assign new_new_n15031__ = ~new_new_n15023__ & ~new_new_n15030__;
  assign new_new_n15032__ = ~new_new_n15022__ & ~new_new_n15031__;
  assign new_new_n15033__ = ~new_new_n14558__ & ~new_new_n15032__;
  assign new_new_n15034__ = ~new_new_n14557__ & ~new_new_n15033__;
  assign new_new_n15035__ = ~new_new_n14549__ & ~new_new_n15034__;
  assign new_new_n15036__ = ~new_new_n14548__ & ~new_new_n15035__;
  assign new_new_n15037__ = ~new_new_n14540__ & new_new_n15036__;
  assign new_new_n15038__ = ~new_new_n14539__ & ~new_new_n15037__;
  assign new_new_n15039__ = ~new_new_n14533__ & new_new_n15038__;
  assign new_new_n15040__ = ~new_new_n14532__ & ~new_new_n15039__;
  assign new_new_n15041__ = ~pi110 & ~new_new_n15040__;
  assign new_new_n15042__ = pi110 & new_new_n15040__;
  assign new_new_n15043__ = ~new_new_n13978__ & ~new_new_n13979__;
  assign new_new_n15044__ = ~new_new_n14479__ & po014;
  assign new_new_n15045__ = ~pi109 & ~po014;
  assign new_new_n15046__ = ~new_new_n15044__ & ~new_new_n15045__;
  assign new_new_n15047__ = new_new_n15043__ & ~new_new_n15046__;
  assign new_new_n15048__ = ~new_new_n15043__ & new_new_n15046__;
  assign new_new_n15049__ = ~new_new_n15047__ & ~new_new_n15048__;
  assign new_new_n15050__ = ~new_new_n15042__ & new_new_n15049__;
  assign new_new_n15051__ = ~new_new_n15041__ & ~new_new_n15050__;
  assign new_new_n15052__ = ~new_new_n14524__ & new_new_n15051__;
  assign new_new_n15053__ = ~new_new_n14523__ & ~new_new_n15052__;
  assign new_new_n15054__ = ~new_new_n14515__ & ~new_new_n15053__;
  assign new_new_n15055__ = ~new_new_n14514__ & ~new_new_n15054__;
  assign new_new_n15056__ = ~new_new_n14506__ & ~new_new_n15055__;
  assign new_new_n15057__ = ~new_new_n14505__ & ~new_new_n15056__;
  assign new_new_n15058__ = ~pi114 & new_new_n15057__;
  assign new_new_n15059__ = pi114 & ~new_new_n15057__;
  assign new_new_n15060__ = new_new_n12847__ & ~new_new_n15058__;
  assign new_new_n15061__ = ~new_new_n15059__ & new_new_n15060__;
  assign new_new_n15062__ = new_new_n14492__ & ~new_new_n15061__;
  assign new_new_n15063__ = pi114 & ~new_new_n14492__;
  assign new_new_n15064__ = new_new_n12847__ & ~new_new_n15063__;
  assign new_new_n15065__ = ~pi113 & new_new_n15055__;
  assign new_new_n15066__ = pi113 & ~new_new_n15055__;
  assign new_new_n15067__ = ~new_new_n15065__ & ~new_new_n15066__;
  assign new_new_n15068__ = new_new_n15064__ & new_new_n15067__;
  assign new_new_n15069__ = ~new_new_n14504__ & ~new_new_n15068__;
  assign new_new_n15070__ = ~pi114 & new_new_n14492__;
  assign new_new_n15071__ = new_new_n12847__ & new_new_n15070__;
  assign new_new_n15072__ = new_new_n14504__ & new_new_n15071__;
  assign new_new_n15073__ = new_new_n15067__ & new_new_n15072__;
  assign new_new_n15074__ = ~new_new_n15069__ & ~new_new_n15073__;
  assign new_new_n15075__ = ~pi114 & ~new_new_n15074__;
  assign new_new_n15076__ = pi114 & ~new_new_n15069__;
  assign new_new_n15077__ = ~new_new_n14514__ & ~new_new_n14515__;
  assign new_new_n15078__ = ~new_new_n15057__ & ~new_new_n15070__;
  assign po013 = new_new_n15064__ & ~new_new_n15078__;
  assign new_new_n15080__ = ~new_new_n15053__ & po013;
  assign new_new_n15081__ = pi112 & ~po013;
  assign new_new_n15082__ = ~new_new_n15080__ & ~new_new_n15081__;
  assign new_new_n15083__ = new_new_n15077__ & new_new_n15082__;
  assign new_new_n15084__ = ~new_new_n15077__ & ~new_new_n15082__;
  assign new_new_n15085__ = ~new_new_n15083__ & ~new_new_n15084__;
  assign new_new_n15086__ = pi113 & ~new_new_n15085__;
  assign new_new_n15087__ = ~pi113 & new_new_n15085__;
  assign new_new_n15088__ = new_new_n15051__ & po013;
  assign new_new_n15089__ = pi111 & ~po013;
  assign new_new_n15090__ = ~new_new_n15088__ & ~new_new_n15089__;
  assign new_new_n15091__ = ~new_new_n14523__ & ~new_new_n14524__;
  assign new_new_n15092__ = ~new_new_n15090__ & ~new_new_n15091__;
  assign new_new_n15093__ = new_new_n15090__ & new_new_n15091__;
  assign new_new_n15094__ = ~new_new_n15092__ & ~new_new_n15093__;
  assign new_new_n15095__ = pi112 & ~new_new_n15094__;
  assign new_new_n15096__ = ~pi112 & new_new_n15094__;
  assign new_new_n15097__ = ~new_new_n15041__ & ~new_new_n15042__;
  assign new_new_n15098__ = po013 & new_new_n15097__;
  assign new_new_n15099__ = new_new_n15049__ & new_new_n15098__;
  assign new_new_n15100__ = ~new_new_n15049__ & ~new_new_n15098__;
  assign new_new_n15101__ = ~new_new_n15099__ & ~new_new_n15100__;
  assign new_new_n15102__ = pi111 & ~new_new_n15101__;
  assign new_new_n15103__ = ~pi111 & new_new_n15101__;
  assign new_new_n15104__ = new_new_n15038__ & po013;
  assign new_new_n15105__ = ~pi109 & ~po013;
  assign new_new_n15106__ = ~new_new_n15104__ & ~new_new_n15105__;
  assign new_new_n15107__ = ~new_new_n14532__ & ~new_new_n14533__;
  assign new_new_n15108__ = ~new_new_n15106__ & ~new_new_n15107__;
  assign new_new_n15109__ = new_new_n15106__ & new_new_n15107__;
  assign new_new_n15110__ = ~new_new_n15108__ & ~new_new_n15109__;
  assign new_new_n15111__ = pi110 & new_new_n15110__;
  assign new_new_n15112__ = ~pi110 & ~new_new_n15110__;
  assign new_new_n15113__ = new_new_n15036__ & po013;
  assign new_new_n15114__ = pi108 & ~po013;
  assign new_new_n15115__ = ~new_new_n15113__ & ~new_new_n15114__;
  assign new_new_n15116__ = ~new_new_n14539__ & ~new_new_n14540__;
  assign new_new_n15117__ = ~new_new_n15115__ & ~new_new_n15116__;
  assign new_new_n15118__ = new_new_n15115__ & new_new_n15116__;
  assign new_new_n15119__ = ~new_new_n15117__ & ~new_new_n15118__;
  assign new_new_n15120__ = pi109 & ~new_new_n15119__;
  assign new_new_n15121__ = ~pi109 & new_new_n15119__;
  assign new_new_n15122__ = ~new_new_n14548__ & ~new_new_n14549__;
  assign new_new_n15123__ = ~new_new_n15034__ & po013;
  assign new_new_n15124__ = ~pi107 & ~po013;
  assign new_new_n15125__ = ~new_new_n15123__ & ~new_new_n15124__;
  assign new_new_n15126__ = new_new_n15122__ & ~new_new_n15125__;
  assign new_new_n15127__ = ~new_new_n15122__ & new_new_n15125__;
  assign new_new_n15128__ = ~new_new_n15126__ & ~new_new_n15127__;
  assign new_new_n15129__ = pi108 & ~new_new_n15128__;
  assign new_new_n15130__ = ~pi108 & new_new_n15128__;
  assign new_new_n15131__ = ~pi106 & ~new_new_n15032__;
  assign new_new_n15132__ = pi106 & new_new_n15032__;
  assign new_new_n15133__ = ~new_new_n15131__ & ~new_new_n15132__;
  assign new_new_n15134__ = po013 & new_new_n15133__;
  assign new_new_n15135__ = new_new_n14556__ & new_new_n15134__;
  assign new_new_n15136__ = ~new_new_n14556__ & ~new_new_n15134__;
  assign new_new_n15137__ = ~new_new_n15135__ & ~new_new_n15136__;
  assign new_new_n15138__ = ~pi107 & ~new_new_n15137__;
  assign new_new_n15139__ = pi107 & new_new_n15137__;
  assign new_new_n15140__ = ~new_new_n15022__ & ~new_new_n15023__;
  assign new_new_n15141__ = po013 & new_new_n15140__;
  assign new_new_n15142__ = new_new_n15030__ & new_new_n15141__;
  assign new_new_n15143__ = ~new_new_n15030__ & ~new_new_n15141__;
  assign new_new_n15144__ = ~new_new_n15142__ & ~new_new_n15143__;
  assign new_new_n15145__ = ~pi106 & ~new_new_n15144__;
  assign new_new_n15146__ = pi106 & new_new_n15144__;
  assign new_new_n15147__ = ~new_new_n15019__ & po013;
  assign new_new_n15148__ = pi104 & ~po013;
  assign new_new_n15149__ = ~new_new_n15147__ & ~new_new_n15148__;
  assign new_new_n15150__ = ~new_new_n14566__ & ~new_new_n14567__;
  assign new_new_n15151__ = new_new_n15149__ & new_new_n15150__;
  assign new_new_n15152__ = ~new_new_n15149__ & ~new_new_n15150__;
  assign new_new_n15153__ = ~new_new_n15151__ & ~new_new_n15152__;
  assign new_new_n15154__ = pi105 & ~new_new_n15153__;
  assign new_new_n15155__ = ~pi105 & new_new_n15153__;
  assign new_new_n15156__ = ~new_new_n14575__ & ~new_new_n14576__;
  assign new_new_n15157__ = pi103 & ~po013;
  assign new_new_n15158__ = ~new_new_n15017__ & po013;
  assign new_new_n15159__ = ~new_new_n15157__ & ~new_new_n15158__;
  assign new_new_n15160__ = new_new_n15156__ & new_new_n15159__;
  assign new_new_n15161__ = ~new_new_n15156__ & ~new_new_n15159__;
  assign new_new_n15162__ = ~new_new_n15160__ & ~new_new_n15161__;
  assign new_new_n15163__ = pi104 & ~new_new_n15162__;
  assign new_new_n15164__ = ~pi104 & new_new_n15162__;
  assign new_new_n15165__ = ~new_new_n14584__ & ~new_new_n14585__;
  assign new_new_n15166__ = pi102 & ~po013;
  assign new_new_n15167__ = ~new_new_n15015__ & po013;
  assign new_new_n15168__ = ~new_new_n15166__ & ~new_new_n15167__;
  assign new_new_n15169__ = new_new_n15165__ & new_new_n15168__;
  assign new_new_n15170__ = ~new_new_n15165__ & ~new_new_n15168__;
  assign new_new_n15171__ = ~new_new_n15169__ & ~new_new_n15170__;
  assign new_new_n15172__ = pi103 & ~new_new_n15171__;
  assign new_new_n15173__ = ~pi103 & new_new_n15171__;
  assign new_new_n15174__ = ~new_new_n14593__ & ~new_new_n14594__;
  assign new_new_n15175__ = ~new_new_n15013__ & po013;
  assign new_new_n15176__ = pi101 & ~po013;
  assign new_new_n15177__ = ~new_new_n15175__ & ~new_new_n15176__;
  assign new_new_n15178__ = new_new_n15174__ & new_new_n15177__;
  assign new_new_n15179__ = ~new_new_n15174__ & ~new_new_n15177__;
  assign new_new_n15180__ = ~new_new_n15178__ & ~new_new_n15179__;
  assign new_new_n15181__ = pi102 & ~new_new_n15180__;
  assign new_new_n15182__ = ~pi102 & new_new_n15180__;
  assign new_new_n15183__ = new_new_n15011__ & po013;
  assign new_new_n15184__ = pi100 & ~po013;
  assign new_new_n15185__ = ~new_new_n15183__ & ~new_new_n15184__;
  assign new_new_n15186__ = ~new_new_n14602__ & ~new_new_n14603__;
  assign new_new_n15187__ = ~new_new_n15185__ & ~new_new_n15186__;
  assign new_new_n15188__ = new_new_n15185__ & new_new_n15186__;
  assign new_new_n15189__ = ~new_new_n15187__ & ~new_new_n15188__;
  assign new_new_n15190__ = pi101 & ~new_new_n15189__;
  assign new_new_n15191__ = ~pi101 & new_new_n15189__;
  assign new_new_n15192__ = ~new_new_n14611__ & ~new_new_n14612__;
  assign new_new_n15193__ = new_new_n15009__ & po013;
  assign new_new_n15194__ = ~pi099 & ~po013;
  assign new_new_n15195__ = ~new_new_n15193__ & ~new_new_n15194__;
  assign new_new_n15196__ = ~new_new_n15192__ & ~new_new_n15195__;
  assign new_new_n15197__ = new_new_n15192__ & new_new_n15195__;
  assign new_new_n15198__ = ~new_new_n15196__ & ~new_new_n15197__;
  assign new_new_n15199__ = pi100 & new_new_n15198__;
  assign new_new_n15200__ = ~pi100 & ~new_new_n15198__;
  assign new_new_n15201__ = pi098 & ~new_new_n15007__;
  assign new_new_n15202__ = ~pi098 & new_new_n15007__;
  assign new_new_n15203__ = ~new_new_n15201__ & ~new_new_n15202__;
  assign new_new_n15204__ = po013 & new_new_n15203__;
  assign new_new_n15205__ = new_new_n14619__ & new_new_n15204__;
  assign new_new_n15206__ = ~new_new_n14619__ & ~new_new_n15204__;
  assign new_new_n15207__ = ~new_new_n15205__ & ~new_new_n15206__;
  assign new_new_n15208__ = pi099 & ~new_new_n15207__;
  assign new_new_n15209__ = ~pi099 & new_new_n15207__;
  assign new_new_n15210__ = ~new_new_n14629__ & ~new_new_n14630__;
  assign new_new_n15211__ = ~new_new_n15005__ & po013;
  assign new_new_n15212__ = pi097 & ~po013;
  assign new_new_n15213__ = ~new_new_n15211__ & ~new_new_n15212__;
  assign new_new_n15214__ = new_new_n15210__ & new_new_n15213__;
  assign new_new_n15215__ = ~new_new_n15210__ & ~new_new_n15213__;
  assign new_new_n15216__ = ~new_new_n15214__ & ~new_new_n15215__;
  assign new_new_n15217__ = pi098 & ~new_new_n15216__;
  assign new_new_n15218__ = ~pi098 & new_new_n15216__;
  assign new_new_n15219__ = new_new_n15003__ & po013;
  assign new_new_n15220__ = pi096 & ~po013;
  assign new_new_n15221__ = ~new_new_n15219__ & ~new_new_n15220__;
  assign new_new_n15222__ = ~new_new_n14638__ & ~new_new_n14639__;
  assign new_new_n15223__ = ~new_new_n15221__ & ~new_new_n15222__;
  assign new_new_n15224__ = new_new_n15221__ & new_new_n15222__;
  assign new_new_n15225__ = ~new_new_n15223__ & ~new_new_n15224__;
  assign new_new_n15226__ = pi097 & ~new_new_n15225__;
  assign new_new_n15227__ = ~pi097 & new_new_n15225__;
  assign new_new_n15228__ = ~new_new_n14993__ & ~new_new_n14994__;
  assign new_new_n15229__ = po013 & new_new_n15228__;
  assign new_new_n15230__ = new_new_n15001__ & new_new_n15229__;
  assign new_new_n15231__ = ~new_new_n15001__ & ~new_new_n15229__;
  assign new_new_n15232__ = ~new_new_n15230__ & ~new_new_n15231__;
  assign new_new_n15233__ = pi096 & ~new_new_n15232__;
  assign new_new_n15234__ = ~pi096 & new_new_n15232__;
  assign new_new_n15235__ = new_new_n14990__ & po013;
  assign new_new_n15236__ = ~pi094 & ~po013;
  assign new_new_n15237__ = ~new_new_n15235__ & ~new_new_n15236__;
  assign new_new_n15238__ = ~new_new_n14647__ & ~new_new_n14648__;
  assign new_new_n15239__ = ~new_new_n15237__ & ~new_new_n15238__;
  assign new_new_n15240__ = new_new_n15237__ & new_new_n15238__;
  assign new_new_n15241__ = ~new_new_n15239__ & ~new_new_n15240__;
  assign new_new_n15242__ = pi095 & new_new_n15241__;
  assign new_new_n15243__ = ~pi095 & ~new_new_n15241__;
  assign new_new_n15244__ = pi093 & ~new_new_n14988__;
  assign new_new_n15245__ = ~pi093 & new_new_n14988__;
  assign new_new_n15246__ = ~new_new_n15244__ & ~new_new_n15245__;
  assign new_new_n15247__ = po013 & new_new_n15246__;
  assign new_new_n15248__ = new_new_n14655__ & new_new_n15247__;
  assign new_new_n15249__ = ~new_new_n14655__ & ~new_new_n15247__;
  assign new_new_n15250__ = ~new_new_n15248__ & ~new_new_n15249__;
  assign new_new_n15251__ = pi094 & ~new_new_n15250__;
  assign new_new_n15252__ = ~pi094 & new_new_n15250__;
  assign new_new_n15253__ = pi092 & ~new_new_n14986__;
  assign new_new_n15254__ = ~pi092 & new_new_n14986__;
  assign new_new_n15255__ = ~new_new_n15253__ & ~new_new_n15254__;
  assign new_new_n15256__ = po013 & new_new_n15255__;
  assign new_new_n15257__ = new_new_n14664__ & new_new_n15256__;
  assign new_new_n15258__ = ~new_new_n14664__ & ~new_new_n15256__;
  assign new_new_n15259__ = ~new_new_n15257__ & ~new_new_n15258__;
  assign new_new_n15260__ = pi093 & ~new_new_n15259__;
  assign new_new_n15261__ = ~pi093 & new_new_n15259__;
  assign new_new_n15262__ = ~new_new_n14674__ & ~new_new_n14675__;
  assign new_new_n15263__ = ~new_new_n14984__ & po013;
  assign new_new_n15264__ = pi091 & ~po013;
  assign new_new_n15265__ = ~new_new_n15263__ & ~new_new_n15264__;
  assign new_new_n15266__ = new_new_n15262__ & ~new_new_n15265__;
  assign new_new_n15267__ = ~new_new_n15262__ & new_new_n15265__;
  assign new_new_n15268__ = ~new_new_n15266__ & ~new_new_n15267__;
  assign new_new_n15269__ = pi092 & new_new_n15268__;
  assign new_new_n15270__ = ~pi092 & ~new_new_n15268__;
  assign new_new_n15271__ = ~new_new_n14683__ & ~new_new_n14684__;
  assign new_new_n15272__ = ~new_new_n14982__ & po013;
  assign new_new_n15273__ = ~pi090 & ~po013;
  assign new_new_n15274__ = ~new_new_n15272__ & ~new_new_n15273__;
  assign new_new_n15275__ = new_new_n15271__ & ~new_new_n15274__;
  assign new_new_n15276__ = ~new_new_n15271__ & new_new_n15274__;
  assign new_new_n15277__ = ~new_new_n15275__ & ~new_new_n15276__;
  assign new_new_n15278__ = pi091 & ~new_new_n15277__;
  assign new_new_n15279__ = ~pi091 & new_new_n15277__;
  assign new_new_n15280__ = ~new_new_n14692__ & ~new_new_n14693__;
  assign new_new_n15281__ = ~new_new_n14980__ & po013;
  assign new_new_n15282__ = ~pi089 & ~po013;
  assign new_new_n15283__ = ~new_new_n15281__ & ~new_new_n15282__;
  assign new_new_n15284__ = new_new_n15280__ & ~new_new_n15283__;
  assign new_new_n15285__ = ~new_new_n15280__ & new_new_n15283__;
  assign new_new_n15286__ = ~new_new_n15284__ & ~new_new_n15285__;
  assign new_new_n15287__ = pi090 & ~new_new_n15286__;
  assign new_new_n15288__ = ~pi090 & new_new_n15286__;
  assign new_new_n15289__ = ~new_new_n14701__ & ~new_new_n14702__;
  assign new_new_n15290__ = ~new_new_n14978__ & po013;
  assign new_new_n15291__ = ~pi088 & ~po013;
  assign new_new_n15292__ = ~new_new_n15290__ & ~new_new_n15291__;
  assign new_new_n15293__ = new_new_n15289__ & ~new_new_n15292__;
  assign new_new_n15294__ = ~new_new_n15289__ & new_new_n15292__;
  assign new_new_n15295__ = ~new_new_n15293__ & ~new_new_n15294__;
  assign new_new_n15296__ = ~pi089 & new_new_n15295__;
  assign new_new_n15297__ = pi089 & ~new_new_n15295__;
  assign new_new_n15298__ = ~new_new_n14710__ & ~new_new_n14711__;
  assign new_new_n15299__ = ~new_new_n14976__ & po013;
  assign new_new_n15300__ = pi087 & ~po013;
  assign new_new_n15301__ = ~new_new_n15299__ & ~new_new_n15300__;
  assign new_new_n15302__ = new_new_n15298__ & ~new_new_n15301__;
  assign new_new_n15303__ = ~new_new_n15298__ & new_new_n15301__;
  assign new_new_n15304__ = ~new_new_n15302__ & ~new_new_n15303__;
  assign new_new_n15305__ = ~pi088 & ~new_new_n15304__;
  assign new_new_n15306__ = pi088 & new_new_n15304__;
  assign new_new_n15307__ = ~new_new_n14974__ & po013;
  assign new_new_n15308__ = pi086 & ~po013;
  assign new_new_n15309__ = ~new_new_n15307__ & ~new_new_n15308__;
  assign new_new_n15310__ = ~new_new_n14719__ & ~new_new_n14720__;
  assign new_new_n15311__ = ~new_new_n15309__ & new_new_n15310__;
  assign new_new_n15312__ = new_new_n15309__ & ~new_new_n15310__;
  assign new_new_n15313__ = ~new_new_n15311__ & ~new_new_n15312__;
  assign new_new_n15314__ = ~pi087 & ~new_new_n15313__;
  assign new_new_n15315__ = pi087 & new_new_n15313__;
  assign new_new_n15316__ = ~new_new_n14972__ & po013;
  assign new_new_n15317__ = pi085 & ~po013;
  assign new_new_n15318__ = ~new_new_n15316__ & ~new_new_n15317__;
  assign new_new_n15319__ = ~new_new_n14728__ & ~new_new_n14729__;
  assign new_new_n15320__ = ~new_new_n15318__ & new_new_n15319__;
  assign new_new_n15321__ = new_new_n15318__ & ~new_new_n15319__;
  assign new_new_n15322__ = ~new_new_n15320__ & ~new_new_n15321__;
  assign new_new_n15323__ = ~pi086 & ~new_new_n15322__;
  assign new_new_n15324__ = pi086 & new_new_n15322__;
  assign new_new_n15325__ = ~new_new_n14737__ & ~new_new_n14738__;
  assign new_new_n15326__ = ~new_new_n14970__ & po013;
  assign new_new_n15327__ = ~pi084 & ~po013;
  assign new_new_n15328__ = ~new_new_n15326__ & ~new_new_n15327__;
  assign new_new_n15329__ = new_new_n15325__ & ~new_new_n15328__;
  assign new_new_n15330__ = ~new_new_n15325__ & new_new_n15328__;
  assign new_new_n15331__ = ~new_new_n15329__ & ~new_new_n15330__;
  assign new_new_n15332__ = pi085 & ~new_new_n15331__;
  assign new_new_n15333__ = ~pi085 & new_new_n15331__;
  assign new_new_n15334__ = ~pi083 & ~new_new_n14968__;
  assign new_new_n15335__ = pi083 & new_new_n14968__;
  assign new_new_n15336__ = ~new_new_n15334__ & ~new_new_n15335__;
  assign new_new_n15337__ = po013 & new_new_n15336__;
  assign new_new_n15338__ = new_new_n14745__ & new_new_n15337__;
  assign new_new_n15339__ = ~new_new_n14745__ & ~new_new_n15337__;
  assign new_new_n15340__ = ~new_new_n15338__ & ~new_new_n15339__;
  assign new_new_n15341__ = ~pi084 & ~new_new_n15340__;
  assign new_new_n15342__ = pi084 & new_new_n15340__;
  assign new_new_n15343__ = ~new_new_n14755__ & ~new_new_n14756__;
  assign new_new_n15344__ = ~new_new_n14966__ & po013;
  assign new_new_n15345__ = pi082 & ~po013;
  assign new_new_n15346__ = ~new_new_n15344__ & ~new_new_n15345__;
  assign new_new_n15347__ = new_new_n15343__ & ~new_new_n15346__;
  assign new_new_n15348__ = ~new_new_n15343__ & new_new_n15346__;
  assign new_new_n15349__ = ~new_new_n15347__ & ~new_new_n15348__;
  assign new_new_n15350__ = ~pi083 & ~new_new_n15349__;
  assign new_new_n15351__ = pi083 & new_new_n15349__;
  assign new_new_n15352__ = ~new_new_n14764__ & ~new_new_n14765__;
  assign new_new_n15353__ = ~new_new_n14964__ & po013;
  assign new_new_n15354__ = ~pi081 & ~po013;
  assign new_new_n15355__ = ~new_new_n15353__ & ~new_new_n15354__;
  assign new_new_n15356__ = new_new_n15352__ & ~new_new_n15355__;
  assign new_new_n15357__ = ~new_new_n15352__ & new_new_n15355__;
  assign new_new_n15358__ = ~new_new_n15356__ & ~new_new_n15357__;
  assign new_new_n15359__ = ~pi082 & new_new_n15358__;
  assign new_new_n15360__ = pi082 & ~new_new_n15358__;
  assign new_new_n15361__ = ~pi080 & ~new_new_n14962__;
  assign new_new_n15362__ = pi080 & new_new_n14962__;
  assign new_new_n15363__ = ~new_new_n15361__ & ~new_new_n15362__;
  assign new_new_n15364__ = po013 & new_new_n15363__;
  assign new_new_n15365__ = new_new_n14772__ & new_new_n15364__;
  assign new_new_n15366__ = ~new_new_n14772__ & ~new_new_n15364__;
  assign new_new_n15367__ = ~new_new_n15365__ & ~new_new_n15366__;
  assign new_new_n15368__ = ~pi081 & ~new_new_n15367__;
  assign new_new_n15369__ = pi081 & new_new_n15367__;
  assign new_new_n15370__ = ~new_new_n14782__ & ~new_new_n14783__;
  assign new_new_n15371__ = ~new_new_n14960__ & po013;
  assign new_new_n15372__ = ~pi079 & ~po013;
  assign new_new_n15373__ = ~new_new_n15371__ & ~new_new_n15372__;
  assign new_new_n15374__ = new_new_n15370__ & ~new_new_n15373__;
  assign new_new_n15375__ = ~new_new_n15370__ & new_new_n15373__;
  assign new_new_n15376__ = ~new_new_n15374__ & ~new_new_n15375__;
  assign new_new_n15377__ = pi080 & ~new_new_n15376__;
  assign new_new_n15378__ = ~pi080 & new_new_n15376__;
  assign new_new_n15379__ = ~new_new_n14791__ & ~new_new_n14792__;
  assign new_new_n15380__ = ~new_new_n14958__ & po013;
  assign new_new_n15381__ = pi078 & ~po013;
  assign new_new_n15382__ = ~new_new_n15380__ & ~new_new_n15381__;
  assign new_new_n15383__ = new_new_n15379__ & ~new_new_n15382__;
  assign new_new_n15384__ = ~new_new_n15379__ & new_new_n15382__;
  assign new_new_n15385__ = ~new_new_n15383__ & ~new_new_n15384__;
  assign new_new_n15386__ = pi079 & new_new_n15385__;
  assign new_new_n15387__ = ~pi079 & ~new_new_n15385__;
  assign new_new_n15388__ = ~new_new_n14956__ & po013;
  assign new_new_n15389__ = pi077 & ~po013;
  assign new_new_n15390__ = ~new_new_n15388__ & ~new_new_n15389__;
  assign new_new_n15391__ = ~new_new_n14800__ & ~new_new_n14801__;
  assign new_new_n15392__ = ~new_new_n15390__ & new_new_n15391__;
  assign new_new_n15393__ = new_new_n15390__ & ~new_new_n15391__;
  assign new_new_n15394__ = ~new_new_n15392__ & ~new_new_n15393__;
  assign new_new_n15395__ = pi078 & new_new_n15394__;
  assign new_new_n15396__ = ~pi078 & ~new_new_n15394__;
  assign new_new_n15397__ = ~new_new_n14809__ & ~new_new_n14810__;
  assign new_new_n15398__ = ~new_new_n14954__ & po013;
  assign new_new_n15399__ = pi076 & ~po013;
  assign new_new_n15400__ = ~new_new_n15398__ & ~new_new_n15399__;
  assign new_new_n15401__ = new_new_n15397__ & new_new_n15400__;
  assign new_new_n15402__ = ~new_new_n15397__ & ~new_new_n15400__;
  assign new_new_n15403__ = ~new_new_n15401__ & ~new_new_n15402__;
  assign new_new_n15404__ = pi077 & ~new_new_n15403__;
  assign new_new_n15405__ = ~pi077 & new_new_n15403__;
  assign new_new_n15406__ = new_new_n14952__ & po013;
  assign new_new_n15407__ = pi075 & ~po013;
  assign new_new_n15408__ = ~new_new_n15406__ & ~new_new_n15407__;
  assign new_new_n15409__ = ~new_new_n14818__ & ~new_new_n14819__;
  assign new_new_n15410__ = ~new_new_n15408__ & ~new_new_n15409__;
  assign new_new_n15411__ = new_new_n15408__ & new_new_n15409__;
  assign new_new_n15412__ = ~new_new_n15410__ & ~new_new_n15411__;
  assign new_new_n15413__ = pi076 & ~new_new_n15412__;
  assign new_new_n15414__ = ~pi076 & new_new_n15412__;
  assign new_new_n15415__ = ~new_new_n14827__ & ~new_new_n14828__;
  assign new_new_n15416__ = ~new_new_n14950__ & po013;
  assign new_new_n15417__ = ~pi074 & ~po013;
  assign new_new_n15418__ = ~new_new_n15416__ & ~new_new_n15417__;
  assign new_new_n15419__ = new_new_n15415__ & ~new_new_n15418__;
  assign new_new_n15420__ = ~new_new_n15415__ & new_new_n15418__;
  assign new_new_n15421__ = ~new_new_n15419__ & ~new_new_n15420__;
  assign new_new_n15422__ = pi075 & ~new_new_n15421__;
  assign new_new_n15423__ = ~pi075 & new_new_n15421__;
  assign new_new_n15424__ = ~new_new_n14836__ & ~new_new_n14837__;
  assign new_new_n15425__ = ~new_new_n14948__ & po013;
  assign new_new_n15426__ = ~pi073 & ~po013;
  assign new_new_n15427__ = ~new_new_n15425__ & ~new_new_n15426__;
  assign new_new_n15428__ = new_new_n15424__ & ~new_new_n15427__;
  assign new_new_n15429__ = ~new_new_n15424__ & new_new_n15427__;
  assign new_new_n15430__ = ~new_new_n15428__ & ~new_new_n15429__;
  assign new_new_n15431__ = pi074 & ~new_new_n15430__;
  assign new_new_n15432__ = ~pi074 & new_new_n15430__;
  assign new_new_n15433__ = ~new_new_n14845__ & ~new_new_n14846__;
  assign new_new_n15434__ = ~new_new_n14946__ & po013;
  assign new_new_n15435__ = ~pi072 & ~po013;
  assign new_new_n15436__ = ~new_new_n15434__ & ~new_new_n15435__;
  assign new_new_n15437__ = new_new_n15433__ & ~new_new_n15436__;
  assign new_new_n15438__ = ~new_new_n15433__ & new_new_n15436__;
  assign new_new_n15439__ = ~new_new_n15437__ & ~new_new_n15438__;
  assign new_new_n15440__ = pi073 & ~new_new_n15439__;
  assign new_new_n15441__ = ~pi073 & new_new_n15439__;
  assign new_new_n15442__ = ~new_new_n14854__ & ~new_new_n14855__;
  assign new_new_n15443__ = ~new_new_n14944__ & po013;
  assign new_new_n15444__ = ~pi071 & ~po013;
  assign new_new_n15445__ = ~new_new_n15443__ & ~new_new_n15444__;
  assign new_new_n15446__ = ~new_new_n15442__ & ~new_new_n15445__;
  assign new_new_n15447__ = new_new_n15442__ & new_new_n15445__;
  assign new_new_n15448__ = ~new_new_n15446__ & ~new_new_n15447__;
  assign new_new_n15449__ = pi072 & new_new_n15448__;
  assign new_new_n15450__ = ~pi072 & ~new_new_n15448__;
  assign new_new_n15451__ = ~new_new_n14934__ & ~new_new_n14935__;
  assign new_new_n15452__ = po013 & new_new_n15451__;
  assign new_new_n15453__ = ~new_new_n14942__ & ~new_new_n15452__;
  assign new_new_n15454__ = new_new_n14942__ & new_new_n15452__;
  assign new_new_n15455__ = ~new_new_n15453__ & ~new_new_n15454__;
  assign new_new_n15456__ = ~pi071 & new_new_n15455__;
  assign new_new_n15457__ = pi069 & ~new_new_n14931__;
  assign new_new_n15458__ = ~pi069 & new_new_n14931__;
  assign new_new_n15459__ = ~new_new_n15457__ & ~new_new_n15458__;
  assign new_new_n15460__ = po013 & new_new_n15459__;
  assign new_new_n15461__ = new_new_n14862__ & new_new_n15460__;
  assign new_new_n15462__ = ~new_new_n14862__ & ~new_new_n15460__;
  assign new_new_n15463__ = ~new_new_n15461__ & ~new_new_n15462__;
  assign new_new_n15464__ = pi070 & ~new_new_n15463__;
  assign new_new_n15465__ = ~pi070 & new_new_n15463__;
  assign new_new_n15466__ = ~new_new_n14921__ & ~new_new_n14922__;
  assign new_new_n15467__ = po013 & new_new_n15466__;
  assign new_new_n15468__ = new_new_n14929__ & ~new_new_n15467__;
  assign new_new_n15469__ = ~new_new_n14929__ & new_new_n15467__;
  assign new_new_n15470__ = ~new_new_n15468__ & ~new_new_n15469__;
  assign new_new_n15471__ = pi069 & ~new_new_n15470__;
  assign new_new_n15472__ = ~pi069 & new_new_n15470__;
  assign new_new_n15473__ = ~new_new_n14877__ & ~new_new_n14878__;
  assign new_new_n15474__ = ~new_new_n14918__ & po013;
  assign new_new_n15475__ = ~pi067 & ~po013;
  assign new_new_n15476__ = ~new_new_n15474__ & ~new_new_n15475__;
  assign new_new_n15477__ = new_new_n15473__ & ~new_new_n15476__;
  assign new_new_n15478__ = ~new_new_n15473__ & new_new_n15476__;
  assign new_new_n15479__ = ~new_new_n15477__ & ~new_new_n15478__;
  assign new_new_n15480__ = pi068 & ~new_new_n15479__;
  assign new_new_n15481__ = ~pi068 & new_new_n15479__;
  assign new_new_n15482__ = ~new_new_n14879__ & new_new_n14880__;
  assign new_new_n15483__ = ~pi014 & ~po014;
  assign new_new_n15484__ = ~pi065 & ~new_new_n15483__;
  assign new_new_n15485__ = ~pi013 & ~new_new_n15484__;
  assign new_new_n15486__ = ~new_new_n15482__ & ~new_new_n15485__;
  assign new_new_n15487__ = pi064 & ~new_new_n15486__;
  assign new_new_n15488__ = ~new_new_n14893__ & ~new_new_n15487__;
  assign new_new_n15489__ = ~pi066 & ~new_new_n15488__;
  assign new_new_n15490__ = pi066 & new_new_n15488__;
  assign new_new_n15491__ = ~new_new_n15489__ & ~new_new_n15490__;
  assign new_new_n15492__ = po013 & ~new_new_n15491__;
  assign new_new_n15493__ = ~new_new_n14346__ & ~new_new_n14865__;
  assign new_new_n15494__ = ~new_new_n14867__ & ~new_new_n15493__;
  assign new_new_n15495__ = ~new_new_n14896__ & new_new_n15493__;
  assign new_new_n15496__ = ~new_new_n15494__ & ~new_new_n15495__;
  assign new_new_n15497__ = new_new_n15492__ & ~new_new_n15496__;
  assign new_new_n15498__ = ~new_new_n15492__ & new_new_n15496__;
  assign new_new_n15499__ = ~new_new_n15497__ & ~new_new_n15498__;
  assign new_new_n15500__ = pi067 & new_new_n15499__;
  assign new_new_n15501__ = ~pi067 & ~new_new_n15499__;
  assign new_new_n15502__ = pi013 & po013;
  assign new_new_n15503__ = ~pi013 & ~po013;
  assign new_new_n15504__ = ~pi065 & ~new_new_n15502__;
  assign new_new_n15505__ = ~new_new_n15503__ & new_new_n15504__;
  assign new_new_n15506__ = ~pi012 & ~new_new_n15505__;
  assign new_new_n15507__ = pi065 & new_new_n15502__;
  assign new_new_n15508__ = ~new_new_n15506__ & ~new_new_n15507__;
  assign new_new_n15509__ = pi064 & ~new_new_n15508__;
  assign new_new_n15510__ = pi064 & po013;
  assign new_new_n15511__ = new_new_n14900__ & ~new_new_n15510__;
  assign new_new_n15512__ = ~new_new_n15509__ & ~new_new_n15511__;
  assign new_new_n15513__ = pi066 & ~new_new_n15512__;
  assign new_new_n15514__ = ~pi066 & new_new_n15512__;
  assign new_new_n15515__ = pi065 & po013;
  assign new_new_n15516__ = ~new_new_n14892__ & ~new_new_n15515__;
  assign new_new_n15517__ = pi064 & ~new_new_n14908__;
  assign new_new_n15518__ = ~new_new_n15516__ & ~new_new_n15517__;
  assign new_new_n15519__ = ~pi065 & po013;
  assign new_new_n15520__ = po014 & new_new_n15519__;
  assign new_new_n15521__ = ~po014 & ~new_new_n15519__;
  assign new_new_n15522__ = pi064 & ~new_new_n15502__;
  assign new_new_n15523__ = ~new_new_n15520__ & new_new_n15522__;
  assign new_new_n15524__ = ~new_new_n15521__ & new_new_n15523__;
  assign new_new_n15525__ = ~new_new_n15518__ & ~new_new_n15524__;
  assign new_new_n15526__ = pi014 & ~new_new_n15525__;
  assign new_new_n15527__ = ~new_new_n332__ & po013;
  assign new_new_n15528__ = ~new_new_n14892__ & ~new_new_n15527__;
  assign new_new_n15529__ = ~new_new_n14907__ & ~new_new_n14909__;
  assign new_new_n15530__ = pi065 & ~new_new_n15510__;
  assign new_new_n15531__ = pi013 & ~new_new_n15529__;
  assign new_new_n15532__ = ~new_new_n15530__ & new_new_n15531__;
  assign new_new_n15533__ = ~pi065 & ~po013;
  assign new_new_n15534__ = ~pi013 & ~new_new_n403__;
  assign new_new_n15535__ = new_new_n15529__ & new_new_n15534__;
  assign new_new_n15536__ = ~new_new_n15533__ & new_new_n15535__;
  assign new_new_n15537__ = ~new_new_n15528__ & ~new_new_n15536__;
  assign new_new_n15538__ = ~new_new_n15532__ & new_new_n15537__;
  assign new_new_n15539__ = ~pi014 & ~new_new_n15538__;
  assign new_new_n15540__ = ~new_new_n15526__ & ~new_new_n15539__;
  assign new_new_n15541__ = ~new_new_n15514__ & ~new_new_n15540__;
  assign new_new_n15542__ = ~new_new_n15513__ & ~new_new_n15541__;
  assign new_new_n15543__ = ~new_new_n15501__ & ~new_new_n15542__;
  assign new_new_n15544__ = ~new_new_n15500__ & ~new_new_n15543__;
  assign new_new_n15545__ = ~new_new_n15481__ & ~new_new_n15544__;
  assign new_new_n15546__ = ~new_new_n15480__ & ~new_new_n15545__;
  assign new_new_n15547__ = ~new_new_n15472__ & ~new_new_n15546__;
  assign new_new_n15548__ = ~new_new_n15471__ & ~new_new_n15547__;
  assign new_new_n15549__ = ~new_new_n15465__ & ~new_new_n15548__;
  assign new_new_n15550__ = ~new_new_n15464__ & ~new_new_n15549__;
  assign new_new_n15551__ = ~new_new_n15456__ & ~new_new_n15550__;
  assign new_new_n15552__ = pi071 & ~new_new_n15455__;
  assign new_new_n15553__ = ~new_new_n15551__ & ~new_new_n15552__;
  assign new_new_n15554__ = ~new_new_n15450__ & ~new_new_n15553__;
  assign new_new_n15555__ = ~new_new_n15449__ & ~new_new_n15554__;
  assign new_new_n15556__ = ~new_new_n15441__ & ~new_new_n15555__;
  assign new_new_n15557__ = ~new_new_n15440__ & ~new_new_n15556__;
  assign new_new_n15558__ = ~new_new_n15432__ & ~new_new_n15557__;
  assign new_new_n15559__ = ~new_new_n15431__ & ~new_new_n15558__;
  assign new_new_n15560__ = ~new_new_n15423__ & ~new_new_n15559__;
  assign new_new_n15561__ = ~new_new_n15422__ & ~new_new_n15560__;
  assign new_new_n15562__ = ~new_new_n15414__ & ~new_new_n15561__;
  assign new_new_n15563__ = ~new_new_n15413__ & ~new_new_n15562__;
  assign new_new_n15564__ = ~new_new_n15405__ & ~new_new_n15563__;
  assign new_new_n15565__ = ~new_new_n15404__ & ~new_new_n15564__;
  assign new_new_n15566__ = ~new_new_n15396__ & ~new_new_n15565__;
  assign new_new_n15567__ = ~new_new_n15395__ & ~new_new_n15566__;
  assign new_new_n15568__ = ~new_new_n15387__ & ~new_new_n15567__;
  assign new_new_n15569__ = ~new_new_n15386__ & ~new_new_n15568__;
  assign new_new_n15570__ = ~new_new_n15378__ & ~new_new_n15569__;
  assign new_new_n15571__ = ~new_new_n15377__ & ~new_new_n15570__;
  assign new_new_n15572__ = ~new_new_n15369__ & new_new_n15571__;
  assign new_new_n15573__ = ~new_new_n15368__ & ~new_new_n15572__;
  assign new_new_n15574__ = ~new_new_n15360__ & ~new_new_n15573__;
  assign new_new_n15575__ = ~new_new_n15359__ & ~new_new_n15574__;
  assign new_new_n15576__ = ~new_new_n15351__ & ~new_new_n15575__;
  assign new_new_n15577__ = ~new_new_n15350__ & ~new_new_n15576__;
  assign new_new_n15578__ = ~new_new_n15342__ & ~new_new_n15577__;
  assign new_new_n15579__ = ~new_new_n15341__ & ~new_new_n15578__;
  assign new_new_n15580__ = ~new_new_n15333__ & new_new_n15579__;
  assign new_new_n15581__ = ~new_new_n15332__ & ~new_new_n15580__;
  assign new_new_n15582__ = ~new_new_n15324__ & new_new_n15581__;
  assign new_new_n15583__ = ~new_new_n15323__ & ~new_new_n15582__;
  assign new_new_n15584__ = ~new_new_n15315__ & ~new_new_n15583__;
  assign new_new_n15585__ = ~new_new_n15314__ & ~new_new_n15584__;
  assign new_new_n15586__ = ~new_new_n15306__ & ~new_new_n15585__;
  assign new_new_n15587__ = ~new_new_n15305__ & ~new_new_n15586__;
  assign new_new_n15588__ = ~new_new_n15297__ & ~new_new_n15587__;
  assign new_new_n15589__ = ~new_new_n15296__ & ~new_new_n15588__;
  assign new_new_n15590__ = ~new_new_n15288__ & new_new_n15589__;
  assign new_new_n15591__ = ~new_new_n15287__ & ~new_new_n15590__;
  assign new_new_n15592__ = ~new_new_n15279__ & ~new_new_n15591__;
  assign new_new_n15593__ = ~new_new_n15278__ & ~new_new_n15592__;
  assign new_new_n15594__ = ~new_new_n15270__ & ~new_new_n15593__;
  assign new_new_n15595__ = ~new_new_n15269__ & ~new_new_n15594__;
  assign new_new_n15596__ = ~new_new_n15261__ & ~new_new_n15595__;
  assign new_new_n15597__ = ~new_new_n15260__ & ~new_new_n15596__;
  assign new_new_n15598__ = ~new_new_n15252__ & ~new_new_n15597__;
  assign new_new_n15599__ = ~new_new_n15251__ & ~new_new_n15598__;
  assign new_new_n15600__ = ~new_new_n15243__ & ~new_new_n15599__;
  assign new_new_n15601__ = ~new_new_n15242__ & ~new_new_n15600__;
  assign new_new_n15602__ = ~new_new_n15234__ & ~new_new_n15601__;
  assign new_new_n15603__ = ~new_new_n15233__ & ~new_new_n15602__;
  assign new_new_n15604__ = ~new_new_n15227__ & ~new_new_n15603__;
  assign new_new_n15605__ = ~new_new_n15226__ & ~new_new_n15604__;
  assign new_new_n15606__ = ~new_new_n15218__ & ~new_new_n15605__;
  assign new_new_n15607__ = ~new_new_n15217__ & ~new_new_n15606__;
  assign new_new_n15608__ = ~new_new_n15209__ & ~new_new_n15607__;
  assign new_new_n15609__ = ~new_new_n15208__ & ~new_new_n15608__;
  assign new_new_n15610__ = ~new_new_n15200__ & ~new_new_n15609__;
  assign new_new_n15611__ = ~new_new_n15199__ & ~new_new_n15610__;
  assign new_new_n15612__ = ~new_new_n15191__ & ~new_new_n15611__;
  assign new_new_n15613__ = ~new_new_n15190__ & ~new_new_n15612__;
  assign new_new_n15614__ = ~new_new_n15182__ & ~new_new_n15613__;
  assign new_new_n15615__ = ~new_new_n15181__ & ~new_new_n15614__;
  assign new_new_n15616__ = ~new_new_n15173__ & ~new_new_n15615__;
  assign new_new_n15617__ = ~new_new_n15172__ & ~new_new_n15616__;
  assign new_new_n15618__ = ~new_new_n15164__ & ~new_new_n15617__;
  assign new_new_n15619__ = ~new_new_n15163__ & ~new_new_n15618__;
  assign new_new_n15620__ = ~new_new_n15155__ & ~new_new_n15619__;
  assign new_new_n15621__ = ~new_new_n15154__ & ~new_new_n15620__;
  assign new_new_n15622__ = ~new_new_n15146__ & new_new_n15621__;
  assign new_new_n15623__ = ~new_new_n15145__ & ~new_new_n15622__;
  assign new_new_n15624__ = ~new_new_n15139__ & ~new_new_n15623__;
  assign new_new_n15625__ = ~new_new_n15138__ & ~new_new_n15624__;
  assign new_new_n15626__ = ~new_new_n15130__ & new_new_n15625__;
  assign new_new_n15627__ = ~new_new_n15129__ & ~new_new_n15626__;
  assign new_new_n15628__ = ~new_new_n15121__ & ~new_new_n15627__;
  assign new_new_n15629__ = ~new_new_n15120__ & ~new_new_n15628__;
  assign new_new_n15630__ = ~new_new_n15112__ & ~new_new_n15629__;
  assign new_new_n15631__ = ~new_new_n15111__ & ~new_new_n15630__;
  assign new_new_n15632__ = ~new_new_n15103__ & ~new_new_n15631__;
  assign new_new_n15633__ = ~new_new_n15102__ & ~new_new_n15632__;
  assign new_new_n15634__ = ~new_new_n15096__ & ~new_new_n15633__;
  assign new_new_n15635__ = ~new_new_n15095__ & ~new_new_n15634__;
  assign new_new_n15636__ = ~new_new_n15087__ & ~new_new_n15635__;
  assign new_new_n15637__ = ~new_new_n15086__ & ~new_new_n15636__;
  assign new_new_n15638__ = ~new_new_n15076__ & new_new_n15637__;
  assign new_new_n15639__ = ~new_new_n15075__ & ~new_new_n15638__;
  assign new_new_n15640__ = ~pi115 & ~new_new_n15639__;
  assign new_new_n15641__ = pi115 & new_new_n15639__;
  assign new_new_n15642__ = ~new_new_n15640__ & ~new_new_n15641__;
  assign new_new_n15643__ = ~pi116 & ~new_new_n15642__;
  assign new_new_n15644__ = ~new_new_n15062__ & ~new_new_n15640__;
  assign new_new_n15645__ = new_new_n12846__ & ~new_new_n15641__;
  assign po012 = ~new_new_n15644__ & new_new_n15645__;
  assign new_new_n15647__ = pi114 & ~new_new_n15637__;
  assign new_new_n15648__ = ~pi114 & new_new_n15637__;
  assign new_new_n15649__ = ~new_new_n15647__ & ~new_new_n15648__;
  assign new_new_n15650__ = po012 & new_new_n15649__;
  assign new_new_n15651__ = ~new_new_n15074__ & new_new_n15650__;
  assign new_new_n15652__ = new_new_n15074__ & ~new_new_n15650__;
  assign new_new_n15653__ = ~new_new_n15651__ & ~new_new_n15652__;
  assign new_new_n15654__ = pi115 & ~new_new_n15653__;
  assign new_new_n15655__ = ~pi115 & new_new_n15653__;
  assign new_new_n15656__ = ~new_new_n15086__ & ~new_new_n15087__;
  assign new_new_n15657__ = ~new_new_n15635__ & po012;
  assign new_new_n15658__ = pi113 & ~po012;
  assign new_new_n15659__ = ~new_new_n15657__ & ~new_new_n15658__;
  assign new_new_n15660__ = new_new_n15656__ & new_new_n15659__;
  assign new_new_n15661__ = ~new_new_n15656__ & ~new_new_n15659__;
  assign new_new_n15662__ = ~new_new_n15660__ & ~new_new_n15661__;
  assign new_new_n15663__ = pi114 & ~new_new_n15662__;
  assign new_new_n15664__ = ~pi114 & new_new_n15662__;
  assign new_new_n15665__ = pi112 & ~new_new_n15633__;
  assign new_new_n15666__ = ~pi112 & new_new_n15633__;
  assign new_new_n15667__ = ~new_new_n15665__ & ~new_new_n15666__;
  assign new_new_n15668__ = po012 & new_new_n15667__;
  assign new_new_n15669__ = ~new_new_n15094__ & ~new_new_n15668__;
  assign new_new_n15670__ = new_new_n15094__ & new_new_n15668__;
  assign new_new_n15671__ = ~new_new_n15669__ & ~new_new_n15670__;
  assign new_new_n15672__ = pi113 & ~new_new_n15671__;
  assign new_new_n15673__ = ~pi113 & new_new_n15671__;
  assign new_new_n15674__ = ~new_new_n15102__ & ~new_new_n15103__;
  assign new_new_n15675__ = ~new_new_n15631__ & po012;
  assign new_new_n15676__ = pi111 & ~po012;
  assign new_new_n15677__ = ~new_new_n15675__ & ~new_new_n15676__;
  assign new_new_n15678__ = new_new_n15674__ & new_new_n15677__;
  assign new_new_n15679__ = ~new_new_n15674__ & ~new_new_n15677__;
  assign new_new_n15680__ = ~new_new_n15678__ & ~new_new_n15679__;
  assign new_new_n15681__ = pi112 & ~new_new_n15680__;
  assign new_new_n15682__ = ~pi112 & new_new_n15680__;
  assign new_new_n15683__ = new_new_n15629__ & po012;
  assign new_new_n15684__ = ~pi110 & ~po012;
  assign new_new_n15685__ = ~new_new_n15683__ & ~new_new_n15684__;
  assign new_new_n15686__ = ~new_new_n15111__ & ~new_new_n15112__;
  assign new_new_n15687__ = ~new_new_n15685__ & ~new_new_n15686__;
  assign new_new_n15688__ = new_new_n15685__ & new_new_n15686__;
  assign new_new_n15689__ = ~new_new_n15687__ & ~new_new_n15688__;
  assign new_new_n15690__ = ~pi111 & ~new_new_n15689__;
  assign new_new_n15691__ = pi111 & new_new_n15689__;
  assign new_new_n15692__ = ~new_new_n15120__ & ~new_new_n15121__;
  assign new_new_n15693__ = ~new_new_n15627__ & po012;
  assign new_new_n15694__ = pi109 & ~po012;
  assign new_new_n15695__ = ~new_new_n15693__ & ~new_new_n15694__;
  assign new_new_n15696__ = new_new_n15692__ & ~new_new_n15695__;
  assign new_new_n15697__ = ~new_new_n15692__ & new_new_n15695__;
  assign new_new_n15698__ = ~new_new_n15696__ & ~new_new_n15697__;
  assign new_new_n15699__ = ~pi110 & ~new_new_n15698__;
  assign new_new_n15700__ = pi110 & new_new_n15698__;
  assign new_new_n15701__ = ~new_new_n15129__ & ~new_new_n15130__;
  assign new_new_n15702__ = ~new_new_n15625__ & po012;
  assign new_new_n15703__ = ~pi108 & ~po012;
  assign new_new_n15704__ = ~new_new_n15702__ & ~new_new_n15703__;
  assign new_new_n15705__ = new_new_n15701__ & ~new_new_n15704__;
  assign new_new_n15706__ = ~new_new_n15701__ & new_new_n15704__;
  assign new_new_n15707__ = ~new_new_n15705__ & ~new_new_n15706__;
  assign new_new_n15708__ = pi109 & ~new_new_n15707__;
  assign new_new_n15709__ = ~pi109 & new_new_n15707__;
  assign new_new_n15710__ = ~new_new_n15138__ & ~new_new_n15139__;
  assign new_new_n15711__ = ~new_new_n15623__ & po012;
  assign new_new_n15712__ = ~pi107 & ~po012;
  assign new_new_n15713__ = ~new_new_n15711__ & ~new_new_n15712__;
  assign new_new_n15714__ = new_new_n15710__ & ~new_new_n15713__;
  assign new_new_n15715__ = ~new_new_n15710__ & new_new_n15713__;
  assign new_new_n15716__ = ~new_new_n15714__ & ~new_new_n15715__;
  assign new_new_n15717__ = pi108 & ~new_new_n15716__;
  assign new_new_n15718__ = ~pi108 & new_new_n15716__;
  assign new_new_n15719__ = ~new_new_n15621__ & po012;
  assign new_new_n15720__ = pi106 & ~po012;
  assign new_new_n15721__ = ~new_new_n15719__ & ~new_new_n15720__;
  assign new_new_n15722__ = ~new_new_n15145__ & ~new_new_n15146__;
  assign new_new_n15723__ = ~new_new_n15721__ & new_new_n15722__;
  assign new_new_n15724__ = new_new_n15721__ & ~new_new_n15722__;
  assign new_new_n15725__ = ~new_new_n15723__ & ~new_new_n15724__;
  assign new_new_n15726__ = ~pi107 & ~new_new_n15725__;
  assign new_new_n15727__ = pi107 & new_new_n15725__;
  assign new_new_n15728__ = ~new_new_n15154__ & ~new_new_n15155__;
  assign new_new_n15729__ = ~new_new_n15619__ & po012;
  assign new_new_n15730__ = pi105 & ~po012;
  assign new_new_n15731__ = ~new_new_n15729__ & ~new_new_n15730__;
  assign new_new_n15732__ = new_new_n15728__ & new_new_n15731__;
  assign new_new_n15733__ = ~new_new_n15728__ & ~new_new_n15731__;
  assign new_new_n15734__ = ~new_new_n15732__ & ~new_new_n15733__;
  assign new_new_n15735__ = pi106 & ~new_new_n15734__;
  assign new_new_n15736__ = ~pi106 & new_new_n15734__;
  assign new_new_n15737__ = pi104 & ~new_new_n15617__;
  assign new_new_n15738__ = ~pi104 & new_new_n15617__;
  assign new_new_n15739__ = ~new_new_n15737__ & ~new_new_n15738__;
  assign new_new_n15740__ = po012 & new_new_n15739__;
  assign new_new_n15741__ = new_new_n15162__ & new_new_n15740__;
  assign new_new_n15742__ = ~new_new_n15162__ & ~new_new_n15740__;
  assign new_new_n15743__ = ~new_new_n15741__ & ~new_new_n15742__;
  assign new_new_n15744__ = pi105 & ~new_new_n15743__;
  assign new_new_n15745__ = ~pi105 & new_new_n15743__;
  assign new_new_n15746__ = ~pi103 & ~new_new_n15615__;
  assign new_new_n15747__ = pi103 & new_new_n15615__;
  assign new_new_n15748__ = ~new_new_n15746__ & ~new_new_n15747__;
  assign new_new_n15749__ = po012 & ~new_new_n15748__;
  assign new_new_n15750__ = new_new_n15171__ & new_new_n15749__;
  assign new_new_n15751__ = ~new_new_n15171__ & ~new_new_n15749__;
  assign new_new_n15752__ = ~new_new_n15750__ & ~new_new_n15751__;
  assign new_new_n15753__ = pi104 & ~new_new_n15752__;
  assign new_new_n15754__ = ~pi104 & new_new_n15752__;
  assign new_new_n15755__ = ~new_new_n15181__ & ~new_new_n15182__;
  assign new_new_n15756__ = pi102 & ~po012;
  assign new_new_n15757__ = ~new_new_n15613__ & po012;
  assign new_new_n15758__ = ~new_new_n15756__ & ~new_new_n15757__;
  assign new_new_n15759__ = new_new_n15755__ & new_new_n15758__;
  assign new_new_n15760__ = ~new_new_n15755__ & ~new_new_n15758__;
  assign new_new_n15761__ = ~new_new_n15759__ & ~new_new_n15760__;
  assign new_new_n15762__ = pi103 & ~new_new_n15761__;
  assign new_new_n15763__ = ~pi103 & new_new_n15761__;
  assign new_new_n15764__ = ~new_new_n15190__ & ~new_new_n15191__;
  assign new_new_n15765__ = ~new_new_n15611__ & po012;
  assign new_new_n15766__ = pi101 & ~po012;
  assign new_new_n15767__ = ~new_new_n15765__ & ~new_new_n15766__;
  assign new_new_n15768__ = new_new_n15764__ & ~new_new_n15767__;
  assign new_new_n15769__ = ~new_new_n15764__ & new_new_n15767__;
  assign new_new_n15770__ = ~new_new_n15768__ & ~new_new_n15769__;
  assign new_new_n15771__ = ~pi102 & ~new_new_n15770__;
  assign new_new_n15772__ = pi102 & new_new_n15770__;
  assign new_new_n15773__ = ~new_new_n15199__ & ~new_new_n15200__;
  assign new_new_n15774__ = new_new_n15609__ & po012;
  assign new_new_n15775__ = ~pi100 & ~po012;
  assign new_new_n15776__ = ~new_new_n15774__ & ~new_new_n15775__;
  assign new_new_n15777__ = ~new_new_n15773__ & ~new_new_n15776__;
  assign new_new_n15778__ = new_new_n15773__ & new_new_n15776__;
  assign new_new_n15779__ = ~new_new_n15777__ & ~new_new_n15778__;
  assign new_new_n15780__ = ~pi101 & ~new_new_n15779__;
  assign new_new_n15781__ = pi101 & new_new_n15779__;
  assign new_new_n15782__ = ~new_new_n15208__ & ~new_new_n15209__;
  assign new_new_n15783__ = ~new_new_n15607__ & po012;
  assign new_new_n15784__ = pi099 & ~po012;
  assign new_new_n15785__ = ~new_new_n15783__ & ~new_new_n15784__;
  assign new_new_n15786__ = new_new_n15782__ & ~new_new_n15785__;
  assign new_new_n15787__ = ~new_new_n15782__ & new_new_n15785__;
  assign new_new_n15788__ = ~new_new_n15786__ & ~new_new_n15787__;
  assign new_new_n15789__ = pi100 & new_new_n15788__;
  assign new_new_n15790__ = ~pi100 & ~new_new_n15788__;
  assign new_new_n15791__ = pi098 & ~new_new_n15605__;
  assign new_new_n15792__ = ~pi098 & new_new_n15605__;
  assign new_new_n15793__ = ~new_new_n15791__ & ~new_new_n15792__;
  assign new_new_n15794__ = po012 & new_new_n15793__;
  assign new_new_n15795__ = ~new_new_n15216__ & ~new_new_n15794__;
  assign new_new_n15796__ = new_new_n15216__ & new_new_n15794__;
  assign new_new_n15797__ = ~new_new_n15795__ & ~new_new_n15796__;
  assign new_new_n15798__ = pi099 & ~new_new_n15797__;
  assign new_new_n15799__ = ~pi099 & new_new_n15797__;
  assign new_new_n15800__ = pi097 & ~new_new_n15603__;
  assign new_new_n15801__ = ~pi097 & new_new_n15603__;
  assign new_new_n15802__ = ~new_new_n15800__ & ~new_new_n15801__;
  assign new_new_n15803__ = po012 & new_new_n15802__;
  assign new_new_n15804__ = new_new_n15225__ & new_new_n15803__;
  assign new_new_n15805__ = ~new_new_n15225__ & ~new_new_n15803__;
  assign new_new_n15806__ = ~new_new_n15804__ & ~new_new_n15805__;
  assign new_new_n15807__ = pi098 & ~new_new_n15806__;
  assign new_new_n15808__ = ~pi098 & new_new_n15806__;
  assign new_new_n15809__ = ~new_new_n15233__ & ~new_new_n15234__;
  assign new_new_n15810__ = ~new_new_n15601__ & po012;
  assign new_new_n15811__ = pi096 & ~po012;
  assign new_new_n15812__ = ~new_new_n15810__ & ~new_new_n15811__;
  assign new_new_n15813__ = new_new_n15809__ & ~new_new_n15812__;
  assign new_new_n15814__ = ~new_new_n15809__ & new_new_n15812__;
  assign new_new_n15815__ = ~new_new_n15813__ & ~new_new_n15814__;
  assign new_new_n15816__ = ~pi097 & ~new_new_n15815__;
  assign new_new_n15817__ = pi097 & new_new_n15815__;
  assign new_new_n15818__ = ~new_new_n15599__ & po012;
  assign new_new_n15819__ = pi095 & ~po012;
  assign new_new_n15820__ = ~new_new_n15818__ & ~new_new_n15819__;
  assign new_new_n15821__ = ~new_new_n15242__ & ~new_new_n15243__;
  assign new_new_n15822__ = ~new_new_n15820__ & new_new_n15821__;
  assign new_new_n15823__ = new_new_n15820__ & ~new_new_n15821__;
  assign new_new_n15824__ = ~new_new_n15822__ & ~new_new_n15823__;
  assign new_new_n15825__ = pi096 & new_new_n15824__;
  assign new_new_n15826__ = ~pi096 & ~new_new_n15824__;
  assign new_new_n15827__ = ~new_new_n15251__ & ~new_new_n15252__;
  assign new_new_n15828__ = ~new_new_n15597__ & po012;
  assign new_new_n15829__ = pi094 & ~po012;
  assign new_new_n15830__ = ~new_new_n15828__ & ~new_new_n15829__;
  assign new_new_n15831__ = new_new_n15827__ & ~new_new_n15830__;
  assign new_new_n15832__ = ~new_new_n15827__ & new_new_n15830__;
  assign new_new_n15833__ = ~new_new_n15831__ & ~new_new_n15832__;
  assign new_new_n15834__ = pi095 & new_new_n15833__;
  assign new_new_n15835__ = ~pi095 & ~new_new_n15833__;
  assign new_new_n15836__ = pi093 & ~new_new_n15595__;
  assign new_new_n15837__ = ~pi093 & new_new_n15595__;
  assign new_new_n15838__ = ~new_new_n15836__ & ~new_new_n15837__;
  assign new_new_n15839__ = po012 & new_new_n15838__;
  assign new_new_n15840__ = new_new_n15259__ & new_new_n15839__;
  assign new_new_n15841__ = ~new_new_n15259__ & ~new_new_n15839__;
  assign new_new_n15842__ = ~new_new_n15840__ & ~new_new_n15841__;
  assign new_new_n15843__ = pi094 & ~new_new_n15842__;
  assign new_new_n15844__ = ~pi094 & new_new_n15842__;
  assign new_new_n15845__ = ~new_new_n15269__ & ~new_new_n15270__;
  assign new_new_n15846__ = ~new_new_n15593__ & po012;
  assign new_new_n15847__ = pi092 & ~po012;
  assign new_new_n15848__ = ~new_new_n15846__ & ~new_new_n15847__;
  assign new_new_n15849__ = new_new_n15845__ & ~new_new_n15848__;
  assign new_new_n15850__ = ~new_new_n15845__ & new_new_n15848__;
  assign new_new_n15851__ = ~new_new_n15849__ & ~new_new_n15850__;
  assign new_new_n15852__ = ~pi093 & ~new_new_n15851__;
  assign new_new_n15853__ = pi093 & new_new_n15851__;
  assign new_new_n15854__ = pi091 & ~new_new_n15591__;
  assign new_new_n15855__ = ~pi091 & new_new_n15591__;
  assign new_new_n15856__ = ~new_new_n15854__ & ~new_new_n15855__;
  assign new_new_n15857__ = po012 & new_new_n15856__;
  assign new_new_n15858__ = new_new_n15277__ & new_new_n15857__;
  assign new_new_n15859__ = ~new_new_n15277__ & ~new_new_n15857__;
  assign new_new_n15860__ = ~new_new_n15858__ & ~new_new_n15859__;
  assign new_new_n15861__ = pi092 & ~new_new_n15860__;
  assign new_new_n15862__ = ~new_new_n15287__ & ~new_new_n15288__;
  assign new_new_n15863__ = ~new_new_n15589__ & po012;
  assign new_new_n15864__ = ~pi090 & ~po012;
  assign new_new_n15865__ = ~new_new_n15863__ & ~new_new_n15864__;
  assign new_new_n15866__ = new_new_n15862__ & ~new_new_n15865__;
  assign new_new_n15867__ = ~new_new_n15862__ & new_new_n15865__;
  assign new_new_n15868__ = ~new_new_n15866__ & ~new_new_n15867__;
  assign new_new_n15869__ = pi091 & ~new_new_n15868__;
  assign new_new_n15870__ = ~pi091 & new_new_n15868__;
  assign new_new_n15871__ = ~new_new_n15296__ & ~new_new_n15297__;
  assign new_new_n15872__ = ~new_new_n15587__ & po012;
  assign new_new_n15873__ = ~pi089 & ~po012;
  assign new_new_n15874__ = ~new_new_n15872__ & ~new_new_n15873__;
  assign new_new_n15875__ = new_new_n15871__ & ~new_new_n15874__;
  assign new_new_n15876__ = ~new_new_n15871__ & new_new_n15874__;
  assign new_new_n15877__ = ~new_new_n15875__ & ~new_new_n15876__;
  assign new_new_n15878__ = pi090 & ~new_new_n15877__;
  assign new_new_n15879__ = ~pi090 & new_new_n15877__;
  assign new_new_n15880__ = ~pi088 & ~new_new_n15585__;
  assign new_new_n15881__ = pi088 & new_new_n15585__;
  assign new_new_n15882__ = ~new_new_n15880__ & ~new_new_n15881__;
  assign new_new_n15883__ = po012 & new_new_n15882__;
  assign new_new_n15884__ = new_new_n15304__ & new_new_n15883__;
  assign new_new_n15885__ = ~new_new_n15304__ & ~new_new_n15883__;
  assign new_new_n15886__ = ~new_new_n15884__ & ~new_new_n15885__;
  assign new_new_n15887__ = ~pi089 & ~new_new_n15886__;
  assign new_new_n15888__ = pi089 & new_new_n15886__;
  assign new_new_n15889__ = ~pi087 & ~new_new_n15583__;
  assign new_new_n15890__ = pi087 & new_new_n15583__;
  assign new_new_n15891__ = ~new_new_n15889__ & ~new_new_n15890__;
  assign new_new_n15892__ = po012 & new_new_n15891__;
  assign new_new_n15893__ = new_new_n15313__ & new_new_n15892__;
  assign new_new_n15894__ = ~new_new_n15313__ & ~new_new_n15892__;
  assign new_new_n15895__ = ~new_new_n15893__ & ~new_new_n15894__;
  assign new_new_n15896__ = ~pi088 & ~new_new_n15895__;
  assign new_new_n15897__ = pi088 & new_new_n15895__;
  assign new_new_n15898__ = ~new_new_n15581__ & po012;
  assign new_new_n15899__ = pi086 & ~po012;
  assign new_new_n15900__ = ~new_new_n15898__ & ~new_new_n15899__;
  assign new_new_n15901__ = ~new_new_n15323__ & ~new_new_n15324__;
  assign new_new_n15902__ = ~new_new_n15900__ & new_new_n15901__;
  assign new_new_n15903__ = new_new_n15900__ & ~new_new_n15901__;
  assign new_new_n15904__ = ~new_new_n15902__ & ~new_new_n15903__;
  assign new_new_n15905__ = pi087 & new_new_n15904__;
  assign new_new_n15906__ = ~pi087 & ~new_new_n15904__;
  assign new_new_n15907__ = ~new_new_n15332__ & ~new_new_n15333__;
  assign new_new_n15908__ = ~new_new_n15579__ & po012;
  assign new_new_n15909__ = ~pi085 & ~po012;
  assign new_new_n15910__ = ~new_new_n15908__ & ~new_new_n15909__;
  assign new_new_n15911__ = new_new_n15907__ & ~new_new_n15910__;
  assign new_new_n15912__ = ~new_new_n15907__ & new_new_n15910__;
  assign new_new_n15913__ = ~new_new_n15911__ & ~new_new_n15912__;
  assign new_new_n15914__ = pi086 & ~new_new_n15913__;
  assign new_new_n15915__ = ~pi086 & new_new_n15913__;
  assign new_new_n15916__ = ~pi084 & ~new_new_n15577__;
  assign new_new_n15917__ = pi084 & new_new_n15577__;
  assign new_new_n15918__ = ~new_new_n15916__ & ~new_new_n15917__;
  assign new_new_n15919__ = po012 & new_new_n15918__;
  assign new_new_n15920__ = new_new_n15340__ & new_new_n15919__;
  assign new_new_n15921__ = ~new_new_n15340__ & ~new_new_n15919__;
  assign new_new_n15922__ = ~new_new_n15920__ & ~new_new_n15921__;
  assign new_new_n15923__ = ~pi085 & ~new_new_n15922__;
  assign new_new_n15924__ = pi085 & new_new_n15922__;
  assign new_new_n15925__ = ~pi083 & ~new_new_n15575__;
  assign new_new_n15926__ = pi083 & new_new_n15575__;
  assign new_new_n15927__ = ~new_new_n15925__ & ~new_new_n15926__;
  assign new_new_n15928__ = po012 & new_new_n15927__;
  assign new_new_n15929__ = new_new_n15349__ & new_new_n15928__;
  assign new_new_n15930__ = ~new_new_n15349__ & ~new_new_n15928__;
  assign new_new_n15931__ = ~new_new_n15929__ & ~new_new_n15930__;
  assign new_new_n15932__ = ~pi084 & ~new_new_n15931__;
  assign new_new_n15933__ = pi084 & new_new_n15931__;
  assign new_new_n15934__ = ~new_new_n15359__ & ~new_new_n15360__;
  assign new_new_n15935__ = ~new_new_n15573__ & po012;
  assign new_new_n15936__ = ~pi082 & ~po012;
  assign new_new_n15937__ = ~new_new_n15935__ & ~new_new_n15936__;
  assign new_new_n15938__ = new_new_n15934__ & ~new_new_n15937__;
  assign new_new_n15939__ = ~new_new_n15934__ & new_new_n15937__;
  assign new_new_n15940__ = ~new_new_n15938__ & ~new_new_n15939__;
  assign new_new_n15941__ = ~pi083 & new_new_n15940__;
  assign new_new_n15942__ = pi083 & ~new_new_n15940__;
  assign new_new_n15943__ = ~new_new_n15571__ & po012;
  assign new_new_n15944__ = pi081 & ~po012;
  assign new_new_n15945__ = ~new_new_n15943__ & ~new_new_n15944__;
  assign new_new_n15946__ = ~new_new_n15368__ & ~new_new_n15369__;
  assign new_new_n15947__ = ~new_new_n15945__ & new_new_n15946__;
  assign new_new_n15948__ = new_new_n15945__ & ~new_new_n15946__;
  assign new_new_n15949__ = ~new_new_n15947__ & ~new_new_n15948__;
  assign new_new_n15950__ = ~pi082 & ~new_new_n15949__;
  assign new_new_n15951__ = pi082 & new_new_n15949__;
  assign new_new_n15952__ = pi080 & ~new_new_n15569__;
  assign new_new_n15953__ = ~pi080 & new_new_n15569__;
  assign new_new_n15954__ = ~new_new_n15952__ & ~new_new_n15953__;
  assign new_new_n15955__ = po012 & new_new_n15954__;
  assign new_new_n15956__ = new_new_n15376__ & new_new_n15955__;
  assign new_new_n15957__ = ~new_new_n15376__ & ~new_new_n15955__;
  assign new_new_n15958__ = ~new_new_n15956__ & ~new_new_n15957__;
  assign new_new_n15959__ = ~pi081 & new_new_n15958__;
  assign new_new_n15960__ = pi081 & ~new_new_n15958__;
  assign new_new_n15961__ = ~new_new_n15386__ & ~new_new_n15387__;
  assign new_new_n15962__ = ~new_new_n15567__ & po012;
  assign new_new_n15963__ = pi079 & ~po012;
  assign new_new_n15964__ = ~new_new_n15962__ & ~new_new_n15963__;
  assign new_new_n15965__ = new_new_n15961__ & ~new_new_n15964__;
  assign new_new_n15966__ = ~new_new_n15961__ & new_new_n15964__;
  assign new_new_n15967__ = ~new_new_n15965__ & ~new_new_n15966__;
  assign new_new_n15968__ = ~pi080 & ~new_new_n15967__;
  assign new_new_n15969__ = pi080 & new_new_n15967__;
  assign new_new_n15970__ = ~new_new_n15565__ & po012;
  assign new_new_n15971__ = pi078 & ~po012;
  assign new_new_n15972__ = ~new_new_n15970__ & ~new_new_n15971__;
  assign new_new_n15973__ = ~new_new_n15395__ & ~new_new_n15396__;
  assign new_new_n15974__ = ~new_new_n15972__ & new_new_n15973__;
  assign new_new_n15975__ = new_new_n15972__ & ~new_new_n15973__;
  assign new_new_n15976__ = ~new_new_n15974__ & ~new_new_n15975__;
  assign new_new_n15977__ = ~pi079 & ~new_new_n15976__;
  assign new_new_n15978__ = pi079 & new_new_n15976__;
  assign new_new_n15979__ = ~new_new_n15404__ & ~new_new_n15405__;
  assign new_new_n15980__ = pi077 & ~po012;
  assign new_new_n15981__ = ~new_new_n15563__ & po012;
  assign new_new_n15982__ = ~new_new_n15980__ & ~new_new_n15981__;
  assign new_new_n15983__ = new_new_n15979__ & new_new_n15982__;
  assign new_new_n15984__ = ~new_new_n15979__ & ~new_new_n15982__;
  assign new_new_n15985__ = ~new_new_n15983__ & ~new_new_n15984__;
  assign new_new_n15986__ = pi078 & ~new_new_n15985__;
  assign new_new_n15987__ = ~pi078 & new_new_n15985__;
  assign new_new_n15988__ = ~new_new_n15413__ & ~new_new_n15414__;
  assign new_new_n15989__ = pi076 & ~po012;
  assign new_new_n15990__ = ~new_new_n15561__ & po012;
  assign new_new_n15991__ = ~new_new_n15989__ & ~new_new_n15990__;
  assign new_new_n15992__ = new_new_n15988__ & new_new_n15991__;
  assign new_new_n15993__ = ~new_new_n15988__ & ~new_new_n15991__;
  assign new_new_n15994__ = ~new_new_n15992__ & ~new_new_n15993__;
  assign new_new_n15995__ = pi077 & ~new_new_n15994__;
  assign new_new_n15996__ = ~pi077 & new_new_n15994__;
  assign new_new_n15997__ = ~new_new_n15559__ & po012;
  assign new_new_n15998__ = pi075 & ~po012;
  assign new_new_n15999__ = ~new_new_n15997__ & ~new_new_n15998__;
  assign new_new_n16000__ = ~new_new_n15422__ & ~new_new_n15423__;
  assign new_new_n16001__ = ~new_new_n15999__ & new_new_n16000__;
  assign new_new_n16002__ = new_new_n15999__ & ~new_new_n16000__;
  assign new_new_n16003__ = ~new_new_n16001__ & ~new_new_n16002__;
  assign new_new_n16004__ = pi076 & new_new_n16003__;
  assign new_new_n16005__ = ~pi076 & ~new_new_n16003__;
  assign new_new_n16006__ = ~new_new_n15431__ & ~new_new_n15432__;
  assign new_new_n16007__ = pi074 & ~po012;
  assign new_new_n16008__ = ~new_new_n15557__ & po012;
  assign new_new_n16009__ = ~new_new_n16007__ & ~new_new_n16008__;
  assign new_new_n16010__ = new_new_n16006__ & new_new_n16009__;
  assign new_new_n16011__ = ~new_new_n16006__ & ~new_new_n16009__;
  assign new_new_n16012__ = ~new_new_n16010__ & ~new_new_n16011__;
  assign new_new_n16013__ = pi075 & ~new_new_n16012__;
  assign new_new_n16014__ = ~pi075 & new_new_n16012__;
  assign new_new_n16015__ = ~new_new_n15440__ & ~new_new_n15441__;
  assign new_new_n16016__ = ~new_new_n15555__ & po012;
  assign new_new_n16017__ = pi073 & ~po012;
  assign new_new_n16018__ = ~new_new_n16016__ & ~new_new_n16017__;
  assign new_new_n16019__ = new_new_n16015__ & new_new_n16018__;
  assign new_new_n16020__ = ~new_new_n16015__ & ~new_new_n16018__;
  assign new_new_n16021__ = ~new_new_n16019__ & ~new_new_n16020__;
  assign new_new_n16022__ = pi074 & ~new_new_n16021__;
  assign new_new_n16023__ = ~pi074 & new_new_n16021__;
  assign new_new_n16024__ = new_new_n15553__ & po012;
  assign new_new_n16025__ = ~pi072 & ~po012;
  assign new_new_n16026__ = ~new_new_n16024__ & ~new_new_n16025__;
  assign new_new_n16027__ = ~new_new_n15449__ & ~new_new_n15450__;
  assign new_new_n16028__ = ~new_new_n16026__ & ~new_new_n16027__;
  assign new_new_n16029__ = new_new_n16026__ & new_new_n16027__;
  assign new_new_n16030__ = ~new_new_n16028__ & ~new_new_n16029__;
  assign new_new_n16031__ = pi073 & new_new_n16030__;
  assign new_new_n16032__ = ~pi073 & ~new_new_n16030__;
  assign new_new_n16033__ = ~new_new_n15550__ & po012;
  assign new_new_n16034__ = pi071 & ~po012;
  assign new_new_n16035__ = ~new_new_n16033__ & ~new_new_n16034__;
  assign new_new_n16036__ = ~new_new_n15456__ & ~new_new_n15552__;
  assign new_new_n16037__ = new_new_n16035__ & new_new_n16036__;
  assign new_new_n16038__ = ~new_new_n16035__ & ~new_new_n16036__;
  assign new_new_n16039__ = ~new_new_n16037__ & ~new_new_n16038__;
  assign new_new_n16040__ = pi072 & ~new_new_n16039__;
  assign new_new_n16041__ = ~pi072 & new_new_n16039__;
  assign new_new_n16042__ = ~new_new_n15464__ & ~new_new_n15465__;
  assign new_new_n16043__ = pi070 & ~po012;
  assign new_new_n16044__ = ~new_new_n15548__ & po012;
  assign new_new_n16045__ = ~new_new_n16043__ & ~new_new_n16044__;
  assign new_new_n16046__ = new_new_n16042__ & new_new_n16045__;
  assign new_new_n16047__ = ~new_new_n16042__ & ~new_new_n16045__;
  assign new_new_n16048__ = ~new_new_n16046__ & ~new_new_n16047__;
  assign new_new_n16049__ = pi071 & ~new_new_n16048__;
  assign new_new_n16050__ = ~pi071 & new_new_n16048__;
  assign new_new_n16051__ = ~new_new_n15546__ & po012;
  assign new_new_n16052__ = pi069 & ~po012;
  assign new_new_n16053__ = ~new_new_n16051__ & ~new_new_n16052__;
  assign new_new_n16054__ = ~new_new_n15471__ & ~new_new_n15472__;
  assign new_new_n16055__ = ~new_new_n16053__ & new_new_n16054__;
  assign new_new_n16056__ = new_new_n16053__ & ~new_new_n16054__;
  assign new_new_n16057__ = ~new_new_n16055__ & ~new_new_n16056__;
  assign new_new_n16058__ = pi070 & new_new_n16057__;
  assign new_new_n16059__ = ~pi070 & ~new_new_n16057__;
  assign new_new_n16060__ = new_new_n15542__ & po012;
  assign new_new_n16061__ = ~pi067 & ~po012;
  assign new_new_n16062__ = ~new_new_n16060__ & ~new_new_n16061__;
  assign new_new_n16063__ = ~new_new_n15500__ & ~new_new_n15501__;
  assign new_new_n16064__ = ~new_new_n16062__ & ~new_new_n16063__;
  assign new_new_n16065__ = new_new_n16062__ & new_new_n16063__;
  assign new_new_n16066__ = ~new_new_n16064__ & ~new_new_n16065__;
  assign new_new_n16067__ = ~pi068 & ~new_new_n16066__;
  assign new_new_n16068__ = pi068 & new_new_n16066__;
  assign new_new_n16069__ = ~new_new_n15513__ & po012;
  assign new_new_n16070__ = ~new_new_n15514__ & new_new_n16069__;
  assign new_new_n16071__ = new_new_n15540__ & ~new_new_n16070__;
  assign new_new_n16072__ = new_new_n15541__ & new_new_n16069__;
  assign new_new_n16073__ = ~new_new_n16071__ & ~new_new_n16072__;
  assign new_new_n16074__ = pi067 & new_new_n16073__;
  assign new_new_n16075__ = ~pi067 & ~new_new_n16073__;
  assign new_new_n16076__ = pi012 & po012;
  assign new_new_n16077__ = pi011 & ~pi065;
  assign new_new_n16078__ = new_new_n16076__ & ~new_new_n16077__;
  assign new_new_n16079__ = ~pi012 & ~po012;
  assign new_new_n16080__ = ~pi065 & ~new_new_n16079__;
  assign new_new_n16081__ = ~pi011 & ~new_new_n16080__;
  assign new_new_n16082__ = ~new_new_n16078__ & ~new_new_n16081__;
  assign new_new_n16083__ = pi064 & ~new_new_n16082__;
  assign new_new_n16084__ = pi064 & po012;
  assign new_new_n16085__ = ~pi012 & pi065;
  assign new_new_n16086__ = ~new_new_n16084__ & new_new_n16085__;
  assign new_new_n16087__ = ~new_new_n16083__ & ~new_new_n16086__;
  assign new_new_n16088__ = pi066 & ~new_new_n16087__;
  assign new_new_n16089__ = new_new_n15519__ & po012;
  assign new_new_n16090__ = new_new_n426__ & ~po013;
  assign new_new_n16091__ = ~new_new_n16089__ & ~new_new_n16090__;
  assign new_new_n16092__ = ~pi012 & ~new_new_n16091__;
  assign new_new_n16093__ = ~new_new_n332__ & po012;
  assign new_new_n16094__ = ~new_new_n15510__ & ~new_new_n16093__;
  assign new_new_n16095__ = pi065 & po012;
  assign new_new_n16096__ = po013 & ~new_new_n16095__;
  assign new_new_n16097__ = pi012 & ~new_new_n15530__;
  assign new_new_n16098__ = ~new_new_n16096__ & new_new_n16097__;
  assign new_new_n16099__ = ~new_new_n16092__ & ~new_new_n16094__;
  assign new_new_n16100__ = ~new_new_n16098__ & new_new_n16099__;
  assign new_new_n16101__ = ~pi013 & ~new_new_n16100__;
  assign new_new_n16102__ = ~new_new_n15510__ & ~new_new_n16095__;
  assign new_new_n16103__ = pi012 & ~new_new_n15515__;
  assign new_new_n16104__ = pi064 & ~new_new_n16103__;
  assign new_new_n16105__ = ~new_new_n16102__ & ~new_new_n16104__;
  assign new_new_n16106__ = ~pi065 & po012;
  assign new_new_n16107__ = ~po013 & ~new_new_n16106__;
  assign new_new_n16108__ = pi064 & ~new_new_n16076__;
  assign new_new_n16109__ = ~new_new_n16089__ & new_new_n16108__;
  assign new_new_n16110__ = ~new_new_n16107__ & new_new_n16109__;
  assign new_new_n16111__ = ~new_new_n16105__ & ~new_new_n16110__;
  assign new_new_n16112__ = pi013 & ~new_new_n16111__;
  assign new_new_n16113__ = ~new_new_n16101__ & ~new_new_n16112__;
  assign new_new_n16114__ = ~pi066 & new_new_n16087__;
  assign new_new_n16115__ = ~new_new_n16113__ & ~new_new_n16114__;
  assign new_new_n16116__ = ~new_new_n16088__ & ~new_new_n16115__;
  assign new_new_n16117__ = ~new_new_n16075__ & ~new_new_n16116__;
  assign new_new_n16118__ = ~new_new_n16074__ & ~new_new_n16117__;
  assign new_new_n16119__ = ~new_new_n16068__ & new_new_n16118__;
  assign new_new_n16120__ = ~new_new_n16067__ & ~new_new_n16119__;
  assign new_new_n16121__ = pi069 & new_new_n16120__;
  assign new_new_n16122__ = ~pi069 & ~new_new_n16120__;
  assign new_new_n16123__ = ~new_new_n15480__ & ~new_new_n15481__;
  assign new_new_n16124__ = ~new_new_n15544__ & po012;
  assign new_new_n16125__ = pi068 & ~po012;
  assign new_new_n16126__ = ~new_new_n16124__ & ~new_new_n16125__;
  assign new_new_n16127__ = new_new_n16123__ & new_new_n16126__;
  assign new_new_n16128__ = ~new_new_n16123__ & ~new_new_n16126__;
  assign new_new_n16129__ = ~new_new_n16127__ & ~new_new_n16128__;
  assign new_new_n16130__ = ~new_new_n16122__ & ~new_new_n16129__;
  assign new_new_n16131__ = ~new_new_n16121__ & ~new_new_n16130__;
  assign new_new_n16132__ = ~new_new_n16059__ & ~new_new_n16131__;
  assign new_new_n16133__ = ~new_new_n16058__ & ~new_new_n16132__;
  assign new_new_n16134__ = ~new_new_n16050__ & ~new_new_n16133__;
  assign new_new_n16135__ = ~new_new_n16049__ & ~new_new_n16134__;
  assign new_new_n16136__ = ~new_new_n16041__ & ~new_new_n16135__;
  assign new_new_n16137__ = ~new_new_n16040__ & ~new_new_n16136__;
  assign new_new_n16138__ = ~new_new_n16032__ & ~new_new_n16137__;
  assign new_new_n16139__ = ~new_new_n16031__ & ~new_new_n16138__;
  assign new_new_n16140__ = ~new_new_n16023__ & ~new_new_n16139__;
  assign new_new_n16141__ = ~new_new_n16022__ & ~new_new_n16140__;
  assign new_new_n16142__ = ~new_new_n16014__ & ~new_new_n16141__;
  assign new_new_n16143__ = ~new_new_n16013__ & ~new_new_n16142__;
  assign new_new_n16144__ = ~new_new_n16005__ & ~new_new_n16143__;
  assign new_new_n16145__ = ~new_new_n16004__ & ~new_new_n16144__;
  assign new_new_n16146__ = ~new_new_n15996__ & ~new_new_n16145__;
  assign new_new_n16147__ = ~new_new_n15995__ & ~new_new_n16146__;
  assign new_new_n16148__ = ~new_new_n15987__ & ~new_new_n16147__;
  assign new_new_n16149__ = ~new_new_n15986__ & ~new_new_n16148__;
  assign new_new_n16150__ = ~new_new_n15978__ & new_new_n16149__;
  assign new_new_n16151__ = ~new_new_n15977__ & ~new_new_n16150__;
  assign new_new_n16152__ = ~new_new_n15969__ & ~new_new_n16151__;
  assign new_new_n16153__ = ~new_new_n15968__ & ~new_new_n16152__;
  assign new_new_n16154__ = ~new_new_n15960__ & ~new_new_n16153__;
  assign new_new_n16155__ = ~new_new_n15959__ & ~new_new_n16154__;
  assign new_new_n16156__ = ~new_new_n15951__ & ~new_new_n16155__;
  assign new_new_n16157__ = ~new_new_n15950__ & ~new_new_n16156__;
  assign new_new_n16158__ = ~new_new_n15942__ & ~new_new_n16157__;
  assign new_new_n16159__ = ~new_new_n15941__ & ~new_new_n16158__;
  assign new_new_n16160__ = ~new_new_n15933__ & ~new_new_n16159__;
  assign new_new_n16161__ = ~new_new_n15932__ & ~new_new_n16160__;
  assign new_new_n16162__ = ~new_new_n15924__ & ~new_new_n16161__;
  assign new_new_n16163__ = ~new_new_n15923__ & ~new_new_n16162__;
  assign new_new_n16164__ = ~new_new_n15915__ & new_new_n16163__;
  assign new_new_n16165__ = ~new_new_n15914__ & ~new_new_n16164__;
  assign new_new_n16166__ = ~new_new_n15906__ & ~new_new_n16165__;
  assign new_new_n16167__ = ~new_new_n15905__ & ~new_new_n16166__;
  assign new_new_n16168__ = ~new_new_n15897__ & new_new_n16167__;
  assign new_new_n16169__ = ~new_new_n15896__ & ~new_new_n16168__;
  assign new_new_n16170__ = ~new_new_n15888__ & ~new_new_n16169__;
  assign new_new_n16171__ = ~new_new_n15887__ & ~new_new_n16170__;
  assign new_new_n16172__ = ~new_new_n15879__ & new_new_n16171__;
  assign new_new_n16173__ = ~new_new_n15878__ & ~new_new_n16172__;
  assign new_new_n16174__ = ~new_new_n15870__ & ~new_new_n16173__;
  assign new_new_n16175__ = ~new_new_n15869__ & ~new_new_n16174__;
  assign new_new_n16176__ = ~pi092 & new_new_n15860__;
  assign new_new_n16177__ = ~new_new_n16175__ & ~new_new_n16176__;
  assign new_new_n16178__ = ~new_new_n15861__ & ~new_new_n16177__;
  assign new_new_n16179__ = ~new_new_n15853__ & new_new_n16178__;
  assign new_new_n16180__ = ~new_new_n15852__ & ~new_new_n16179__;
  assign new_new_n16181__ = ~new_new_n15844__ & new_new_n16180__;
  assign new_new_n16182__ = ~new_new_n15843__ & ~new_new_n16181__;
  assign new_new_n16183__ = ~new_new_n15835__ & ~new_new_n16182__;
  assign new_new_n16184__ = ~new_new_n15834__ & ~new_new_n16183__;
  assign new_new_n16185__ = ~new_new_n15826__ & ~new_new_n16184__;
  assign new_new_n16186__ = ~new_new_n15825__ & ~new_new_n16185__;
  assign new_new_n16187__ = ~new_new_n15817__ & new_new_n16186__;
  assign new_new_n16188__ = ~new_new_n15816__ & ~new_new_n16187__;
  assign new_new_n16189__ = ~new_new_n15808__ & new_new_n16188__;
  assign new_new_n16190__ = ~new_new_n15807__ & ~new_new_n16189__;
  assign new_new_n16191__ = ~new_new_n15799__ & ~new_new_n16190__;
  assign new_new_n16192__ = ~new_new_n15798__ & ~new_new_n16191__;
  assign new_new_n16193__ = ~new_new_n15790__ & ~new_new_n16192__;
  assign new_new_n16194__ = ~new_new_n15789__ & ~new_new_n16193__;
  assign new_new_n16195__ = ~new_new_n15781__ & new_new_n16194__;
  assign new_new_n16196__ = ~new_new_n15780__ & ~new_new_n16195__;
  assign new_new_n16197__ = ~new_new_n15772__ & ~new_new_n16196__;
  assign new_new_n16198__ = ~new_new_n15771__ & ~new_new_n16197__;
  assign new_new_n16199__ = ~new_new_n15763__ & new_new_n16198__;
  assign new_new_n16200__ = ~new_new_n15762__ & ~new_new_n16199__;
  assign new_new_n16201__ = ~new_new_n15754__ & ~new_new_n16200__;
  assign new_new_n16202__ = ~new_new_n15753__ & ~new_new_n16201__;
  assign new_new_n16203__ = ~new_new_n15745__ & ~new_new_n16202__;
  assign new_new_n16204__ = ~new_new_n15744__ & ~new_new_n16203__;
  assign new_new_n16205__ = ~new_new_n15736__ & ~new_new_n16204__;
  assign new_new_n16206__ = ~new_new_n15735__ & ~new_new_n16205__;
  assign new_new_n16207__ = ~new_new_n15727__ & new_new_n16206__;
  assign new_new_n16208__ = ~new_new_n15726__ & ~new_new_n16207__;
  assign new_new_n16209__ = ~new_new_n15718__ & new_new_n16208__;
  assign new_new_n16210__ = ~new_new_n15717__ & ~new_new_n16209__;
  assign new_new_n16211__ = ~new_new_n15709__ & ~new_new_n16210__;
  assign new_new_n16212__ = ~new_new_n15708__ & ~new_new_n16211__;
  assign new_new_n16213__ = ~new_new_n15700__ & new_new_n16212__;
  assign new_new_n16214__ = ~new_new_n15699__ & ~new_new_n16213__;
  assign new_new_n16215__ = ~new_new_n15691__ & ~new_new_n16214__;
  assign new_new_n16216__ = ~new_new_n15690__ & ~new_new_n16215__;
  assign new_new_n16217__ = ~new_new_n15682__ & new_new_n16216__;
  assign new_new_n16218__ = ~new_new_n15681__ & ~new_new_n16217__;
  assign new_new_n16219__ = ~new_new_n15673__ & ~new_new_n16218__;
  assign new_new_n16220__ = ~new_new_n15672__ & ~new_new_n16219__;
  assign new_new_n16221__ = ~new_new_n15664__ & ~new_new_n16220__;
  assign new_new_n16222__ = ~new_new_n15663__ & ~new_new_n16221__;
  assign new_new_n16223__ = ~new_new_n15655__ & ~new_new_n16222__;
  assign new_new_n16224__ = ~new_new_n15654__ & ~new_new_n16223__;
  assign new_new_n16225__ = new_new_n15643__ & new_new_n16224__;
  assign new_new_n16226__ = pi116 & ~new_new_n16224__;
  assign new_new_n16227__ = new_new_n269__ & ~new_new_n16225__;
  assign new_new_n16228__ = ~new_new_n16226__ & new_new_n16227__;
  assign new_new_n16229__ = new_new_n15062__ & ~new_new_n16228__;
  assign new_new_n16230__ = ~new_new_n15654__ & ~new_new_n15655__;
  assign new_new_n16231__ = pi116 & ~new_new_n15062__;
  assign new_new_n16232__ = new_new_n16224__ & ~new_new_n16231__;
  assign new_new_n16233__ = new_new_n15062__ & new_new_n15643__;
  assign new_new_n16234__ = ~new_new_n16232__ & ~new_new_n16233__;
  assign po011 = new_new_n269__ & ~new_new_n16234__;
  assign new_new_n16236__ = ~new_new_n16222__ & po011;
  assign new_new_n16237__ = pi115 & ~po011;
  assign new_new_n16238__ = ~new_new_n16236__ & ~new_new_n16237__;
  assign new_new_n16239__ = new_new_n16230__ & ~new_new_n16238__;
  assign new_new_n16240__ = ~new_new_n16230__ & new_new_n16238__;
  assign new_new_n16241__ = ~new_new_n16239__ & ~new_new_n16240__;
  assign new_new_n16242__ = ~pi116 & ~new_new_n16241__;
  assign new_new_n16243__ = pi116 & new_new_n16241__;
  assign new_new_n16244__ = ~new_new_n15663__ & ~new_new_n15664__;
  assign new_new_n16245__ = pi114 & ~po011;
  assign new_new_n16246__ = ~new_new_n16220__ & po011;
  assign new_new_n16247__ = ~new_new_n16245__ & ~new_new_n16246__;
  assign new_new_n16248__ = new_new_n16244__ & new_new_n16247__;
  assign new_new_n16249__ = ~new_new_n16244__ & ~new_new_n16247__;
  assign new_new_n16250__ = ~new_new_n16248__ & ~new_new_n16249__;
  assign new_new_n16251__ = pi115 & ~new_new_n16250__;
  assign new_new_n16252__ = ~pi115 & new_new_n16250__;
  assign new_new_n16253__ = ~new_new_n16218__ & po011;
  assign new_new_n16254__ = pi113 & ~po011;
  assign new_new_n16255__ = ~new_new_n16253__ & ~new_new_n16254__;
  assign new_new_n16256__ = ~new_new_n15672__ & ~new_new_n15673__;
  assign new_new_n16257__ = ~new_new_n16255__ & new_new_n16256__;
  assign new_new_n16258__ = new_new_n16255__ & ~new_new_n16256__;
  assign new_new_n16259__ = ~new_new_n16257__ & ~new_new_n16258__;
  assign new_new_n16260__ = pi114 & new_new_n16259__;
  assign new_new_n16261__ = ~pi114 & ~new_new_n16259__;
  assign new_new_n16262__ = ~new_new_n15681__ & ~new_new_n15682__;
  assign new_new_n16263__ = ~new_new_n16216__ & po011;
  assign new_new_n16264__ = ~pi112 & ~po011;
  assign new_new_n16265__ = ~new_new_n16263__ & ~new_new_n16264__;
  assign new_new_n16266__ = new_new_n16262__ & ~new_new_n16265__;
  assign new_new_n16267__ = ~new_new_n16262__ & new_new_n16265__;
  assign new_new_n16268__ = ~new_new_n16266__ & ~new_new_n16267__;
  assign new_new_n16269__ = pi113 & ~new_new_n16268__;
  assign new_new_n16270__ = ~pi113 & new_new_n16268__;
  assign new_new_n16271__ = ~pi111 & ~new_new_n16214__;
  assign new_new_n16272__ = pi111 & new_new_n16214__;
  assign new_new_n16273__ = ~new_new_n16271__ & ~new_new_n16272__;
  assign new_new_n16274__ = po011 & new_new_n16273__;
  assign new_new_n16275__ = ~new_new_n15689__ & new_new_n16274__;
  assign new_new_n16276__ = new_new_n15689__ & ~new_new_n16274__;
  assign new_new_n16277__ = ~new_new_n16275__ & ~new_new_n16276__;
  assign new_new_n16278__ = pi112 & ~new_new_n16277__;
  assign new_new_n16279__ = ~pi112 & new_new_n16277__;
  assign new_new_n16280__ = ~new_new_n16212__ & po011;
  assign new_new_n16281__ = pi110 & ~po011;
  assign new_new_n16282__ = ~new_new_n16280__ & ~new_new_n16281__;
  assign new_new_n16283__ = ~new_new_n15699__ & ~new_new_n15700__;
  assign new_new_n16284__ = ~new_new_n16282__ & new_new_n16283__;
  assign new_new_n16285__ = new_new_n16282__ & ~new_new_n16283__;
  assign new_new_n16286__ = ~new_new_n16284__ & ~new_new_n16285__;
  assign new_new_n16287__ = pi111 & new_new_n16286__;
  assign new_new_n16288__ = ~pi111 & ~new_new_n16286__;
  assign new_new_n16289__ = pi109 & ~new_new_n16210__;
  assign new_new_n16290__ = ~pi109 & new_new_n16210__;
  assign new_new_n16291__ = ~new_new_n16289__ & ~new_new_n16290__;
  assign new_new_n16292__ = po011 & new_new_n16291__;
  assign new_new_n16293__ = new_new_n15707__ & new_new_n16292__;
  assign new_new_n16294__ = ~new_new_n15707__ & ~new_new_n16292__;
  assign new_new_n16295__ = ~new_new_n16293__ & ~new_new_n16294__;
  assign new_new_n16296__ = pi110 & ~new_new_n16295__;
  assign new_new_n16297__ = ~pi110 & new_new_n16295__;
  assign new_new_n16298__ = ~new_new_n15717__ & ~new_new_n15718__;
  assign new_new_n16299__ = ~new_new_n16208__ & po011;
  assign new_new_n16300__ = ~pi108 & ~po011;
  assign new_new_n16301__ = ~new_new_n16299__ & ~new_new_n16300__;
  assign new_new_n16302__ = new_new_n16298__ & ~new_new_n16301__;
  assign new_new_n16303__ = ~new_new_n16298__ & new_new_n16301__;
  assign new_new_n16304__ = ~new_new_n16302__ & ~new_new_n16303__;
  assign new_new_n16305__ = pi109 & ~new_new_n16304__;
  assign new_new_n16306__ = ~pi109 & new_new_n16304__;
  assign new_new_n16307__ = ~new_new_n16206__ & po011;
  assign new_new_n16308__ = pi107 & ~po011;
  assign new_new_n16309__ = ~new_new_n16307__ & ~new_new_n16308__;
  assign new_new_n16310__ = ~new_new_n15726__ & ~new_new_n15727__;
  assign new_new_n16311__ = ~new_new_n16309__ & new_new_n16310__;
  assign new_new_n16312__ = new_new_n16309__ & ~new_new_n16310__;
  assign new_new_n16313__ = ~new_new_n16311__ & ~new_new_n16312__;
  assign new_new_n16314__ = ~pi108 & ~new_new_n16313__;
  assign new_new_n16315__ = pi108 & new_new_n16313__;
  assign new_new_n16316__ = ~new_new_n15735__ & ~new_new_n15736__;
  assign new_new_n16317__ = ~new_new_n16204__ & po011;
  assign new_new_n16318__ = pi106 & ~po011;
  assign new_new_n16319__ = ~new_new_n16317__ & ~new_new_n16318__;
  assign new_new_n16320__ = new_new_n16316__ & new_new_n16319__;
  assign new_new_n16321__ = ~new_new_n16316__ & ~new_new_n16319__;
  assign new_new_n16322__ = ~new_new_n16320__ & ~new_new_n16321__;
  assign new_new_n16323__ = ~pi107 & new_new_n16322__;
  assign new_new_n16324__ = pi107 & ~new_new_n16322__;
  assign new_new_n16325__ = ~new_new_n15744__ & ~new_new_n15745__;
  assign new_new_n16326__ = ~new_new_n16202__ & po011;
  assign new_new_n16327__ = pi105 & ~po011;
  assign new_new_n16328__ = ~new_new_n16326__ & ~new_new_n16327__;
  assign new_new_n16329__ = new_new_n16325__ & ~new_new_n16328__;
  assign new_new_n16330__ = ~new_new_n16325__ & new_new_n16328__;
  assign new_new_n16331__ = ~new_new_n16329__ & ~new_new_n16330__;
  assign new_new_n16332__ = ~pi106 & ~new_new_n16331__;
  assign new_new_n16333__ = pi106 & new_new_n16331__;
  assign new_new_n16334__ = pi104 & ~new_new_n16200__;
  assign new_new_n16335__ = ~pi104 & new_new_n16200__;
  assign new_new_n16336__ = ~new_new_n16334__ & ~new_new_n16335__;
  assign new_new_n16337__ = po011 & new_new_n16336__;
  assign new_new_n16338__ = ~new_new_n15752__ & new_new_n16337__;
  assign new_new_n16339__ = new_new_n15752__ & ~new_new_n16337__;
  assign new_new_n16340__ = ~new_new_n16338__ & ~new_new_n16339__;
  assign new_new_n16341__ = ~pi105 & ~new_new_n16340__;
  assign new_new_n16342__ = pi105 & new_new_n16340__;
  assign new_new_n16343__ = ~new_new_n15762__ & ~new_new_n15763__;
  assign new_new_n16344__ = ~new_new_n16198__ & po011;
  assign new_new_n16345__ = ~pi103 & ~po011;
  assign new_new_n16346__ = ~new_new_n16344__ & ~new_new_n16345__;
  assign new_new_n16347__ = new_new_n16343__ & ~new_new_n16346__;
  assign new_new_n16348__ = ~new_new_n16343__ & new_new_n16346__;
  assign new_new_n16349__ = ~new_new_n16347__ & ~new_new_n16348__;
  assign new_new_n16350__ = pi104 & ~new_new_n16349__;
  assign new_new_n16351__ = ~pi104 & new_new_n16349__;
  assign new_new_n16352__ = ~pi102 & ~new_new_n16196__;
  assign new_new_n16353__ = pi102 & new_new_n16196__;
  assign new_new_n16354__ = ~new_new_n16352__ & ~new_new_n16353__;
  assign new_new_n16355__ = po011 & new_new_n16354__;
  assign new_new_n16356__ = new_new_n15770__ & new_new_n16355__;
  assign new_new_n16357__ = ~new_new_n15770__ & ~new_new_n16355__;
  assign new_new_n16358__ = ~new_new_n16356__ & ~new_new_n16357__;
  assign new_new_n16359__ = ~pi103 & ~new_new_n16358__;
  assign new_new_n16360__ = pi103 & new_new_n16358__;
  assign new_new_n16361__ = ~new_new_n15780__ & ~new_new_n15781__;
  assign new_new_n16362__ = new_new_n16194__ & po011;
  assign new_new_n16363__ = ~pi101 & ~po011;
  assign new_new_n16364__ = ~new_new_n16362__ & ~new_new_n16363__;
  assign new_new_n16365__ = ~new_new_n16361__ & ~new_new_n16364__;
  assign new_new_n16366__ = new_new_n16361__ & new_new_n16364__;
  assign new_new_n16367__ = ~new_new_n16365__ & ~new_new_n16366__;
  assign new_new_n16368__ = ~pi102 & ~new_new_n16367__;
  assign new_new_n16369__ = pi102 & new_new_n16367__;
  assign new_new_n16370__ = new_new_n16192__ & po011;
  assign new_new_n16371__ = ~pi100 & ~po011;
  assign new_new_n16372__ = ~new_new_n16370__ & ~new_new_n16371__;
  assign new_new_n16373__ = ~new_new_n15789__ & ~new_new_n15790__;
  assign new_new_n16374__ = ~new_new_n16372__ & ~new_new_n16373__;
  assign new_new_n16375__ = new_new_n16372__ & new_new_n16373__;
  assign new_new_n16376__ = ~new_new_n16374__ & ~new_new_n16375__;
  assign new_new_n16377__ = ~pi101 & ~new_new_n16376__;
  assign new_new_n16378__ = pi101 & new_new_n16376__;
  assign new_new_n16379__ = ~new_new_n16190__ & po011;
  assign new_new_n16380__ = pi099 & ~po011;
  assign new_new_n16381__ = ~new_new_n16379__ & ~new_new_n16380__;
  assign new_new_n16382__ = ~new_new_n15798__ & ~new_new_n15799__;
  assign new_new_n16383__ = ~new_new_n16381__ & new_new_n16382__;
  assign new_new_n16384__ = new_new_n16381__ & ~new_new_n16382__;
  assign new_new_n16385__ = ~new_new_n16383__ & ~new_new_n16384__;
  assign new_new_n16386__ = ~pi100 & ~new_new_n16385__;
  assign new_new_n16387__ = pi100 & new_new_n16385__;
  assign new_new_n16388__ = ~new_new_n15807__ & ~new_new_n15808__;
  assign new_new_n16389__ = ~new_new_n16188__ & po011;
  assign new_new_n16390__ = ~pi098 & ~po011;
  assign new_new_n16391__ = ~new_new_n16389__ & ~new_new_n16390__;
  assign new_new_n16392__ = new_new_n16388__ & ~new_new_n16391__;
  assign new_new_n16393__ = ~new_new_n16388__ & new_new_n16391__;
  assign new_new_n16394__ = ~new_new_n16392__ & ~new_new_n16393__;
  assign new_new_n16395__ = pi099 & ~new_new_n16394__;
  assign new_new_n16396__ = ~pi099 & new_new_n16394__;
  assign new_new_n16397__ = ~new_new_n15816__ & ~new_new_n15817__;
  assign new_new_n16398__ = ~new_new_n16186__ & po011;
  assign new_new_n16399__ = pi097 & ~po011;
  assign new_new_n16400__ = ~new_new_n16398__ & ~new_new_n16399__;
  assign new_new_n16401__ = new_new_n16397__ & ~new_new_n16400__;
  assign new_new_n16402__ = ~new_new_n16397__ & new_new_n16400__;
  assign new_new_n16403__ = ~new_new_n16401__ & ~new_new_n16402__;
  assign new_new_n16404__ = ~pi098 & ~new_new_n16403__;
  assign new_new_n16405__ = pi098 & new_new_n16403__;
  assign new_new_n16406__ = ~new_new_n16184__ & po011;
  assign new_new_n16407__ = pi096 & ~po011;
  assign new_new_n16408__ = ~new_new_n16406__ & ~new_new_n16407__;
  assign new_new_n16409__ = ~new_new_n15825__ & ~new_new_n15826__;
  assign new_new_n16410__ = ~new_new_n16408__ & new_new_n16409__;
  assign new_new_n16411__ = new_new_n16408__ & ~new_new_n16409__;
  assign new_new_n16412__ = ~new_new_n16410__ & ~new_new_n16411__;
  assign new_new_n16413__ = ~pi097 & ~new_new_n16412__;
  assign new_new_n16414__ = pi097 & new_new_n16412__;
  assign new_new_n16415__ = ~new_new_n16182__ & po011;
  assign new_new_n16416__ = pi095 & ~po011;
  assign new_new_n16417__ = ~new_new_n16415__ & ~new_new_n16416__;
  assign new_new_n16418__ = ~new_new_n15834__ & ~new_new_n15835__;
  assign new_new_n16419__ = ~new_new_n16417__ & new_new_n16418__;
  assign new_new_n16420__ = new_new_n16417__ & ~new_new_n16418__;
  assign new_new_n16421__ = ~new_new_n16419__ & ~new_new_n16420__;
  assign new_new_n16422__ = ~pi096 & ~new_new_n16421__;
  assign new_new_n16423__ = pi096 & new_new_n16421__;
  assign new_new_n16424__ = ~new_new_n15843__ & ~new_new_n15844__;
  assign new_new_n16425__ = ~new_new_n16180__ & po011;
  assign new_new_n16426__ = ~pi094 & ~po011;
  assign new_new_n16427__ = ~new_new_n16425__ & ~new_new_n16426__;
  assign new_new_n16428__ = new_new_n16424__ & ~new_new_n16427__;
  assign new_new_n16429__ = ~new_new_n16424__ & new_new_n16427__;
  assign new_new_n16430__ = ~new_new_n16428__ & ~new_new_n16429__;
  assign new_new_n16431__ = pi095 & ~new_new_n16430__;
  assign new_new_n16432__ = ~pi095 & new_new_n16430__;
  assign new_new_n16433__ = ~new_new_n16178__ & po011;
  assign new_new_n16434__ = pi093 & ~po011;
  assign new_new_n16435__ = ~new_new_n16433__ & ~new_new_n16434__;
  assign new_new_n16436__ = ~new_new_n15852__ & ~new_new_n15853__;
  assign new_new_n16437__ = ~new_new_n16435__ & new_new_n16436__;
  assign new_new_n16438__ = new_new_n16435__ & ~new_new_n16436__;
  assign new_new_n16439__ = ~new_new_n16437__ & ~new_new_n16438__;
  assign new_new_n16440__ = ~pi094 & ~new_new_n16439__;
  assign new_new_n16441__ = pi094 & new_new_n16439__;
  assign new_new_n16442__ = ~new_new_n15861__ & ~new_new_n16176__;
  assign new_new_n16443__ = ~new_new_n16175__ & po011;
  assign new_new_n16444__ = pi092 & ~po011;
  assign new_new_n16445__ = ~new_new_n16443__ & ~new_new_n16444__;
  assign new_new_n16446__ = new_new_n16442__ & ~new_new_n16445__;
  assign new_new_n16447__ = ~new_new_n16442__ & new_new_n16445__;
  assign new_new_n16448__ = ~new_new_n16446__ & ~new_new_n16447__;
  assign new_new_n16449__ = pi093 & new_new_n16448__;
  assign new_new_n16450__ = ~pi093 & ~new_new_n16448__;
  assign new_new_n16451__ = pi091 & ~new_new_n16173__;
  assign new_new_n16452__ = ~pi091 & new_new_n16173__;
  assign new_new_n16453__ = ~new_new_n16451__ & ~new_new_n16452__;
  assign new_new_n16454__ = po011 & new_new_n16453__;
  assign new_new_n16455__ = new_new_n15868__ & new_new_n16454__;
  assign new_new_n16456__ = ~new_new_n15868__ & ~new_new_n16454__;
  assign new_new_n16457__ = ~new_new_n16455__ & ~new_new_n16456__;
  assign new_new_n16458__ = pi092 & ~new_new_n16457__;
  assign new_new_n16459__ = ~pi092 & new_new_n16457__;
  assign new_new_n16460__ = ~new_new_n15878__ & ~new_new_n15879__;
  assign new_new_n16461__ = ~new_new_n16171__ & po011;
  assign new_new_n16462__ = ~pi090 & ~po011;
  assign new_new_n16463__ = ~new_new_n16461__ & ~new_new_n16462__;
  assign new_new_n16464__ = new_new_n16460__ & ~new_new_n16463__;
  assign new_new_n16465__ = ~new_new_n16460__ & new_new_n16463__;
  assign new_new_n16466__ = ~new_new_n16464__ & ~new_new_n16465__;
  assign new_new_n16467__ = ~pi091 & new_new_n16466__;
  assign new_new_n16468__ = pi091 & ~new_new_n16466__;
  assign new_new_n16469__ = ~pi089 & ~new_new_n16169__;
  assign new_new_n16470__ = pi089 & new_new_n16169__;
  assign new_new_n16471__ = ~new_new_n16469__ & ~new_new_n16470__;
  assign new_new_n16472__ = po011 & new_new_n16471__;
  assign new_new_n16473__ = new_new_n15886__ & new_new_n16472__;
  assign new_new_n16474__ = ~new_new_n15886__ & ~new_new_n16472__;
  assign new_new_n16475__ = ~new_new_n16473__ & ~new_new_n16474__;
  assign new_new_n16476__ = ~pi090 & ~new_new_n16475__;
  assign new_new_n16477__ = pi090 & new_new_n16475__;
  assign new_new_n16478__ = ~new_new_n16167__ & po011;
  assign new_new_n16479__ = pi088 & ~po011;
  assign new_new_n16480__ = ~new_new_n16478__ & ~new_new_n16479__;
  assign new_new_n16481__ = ~new_new_n15896__ & ~new_new_n15897__;
  assign new_new_n16482__ = ~new_new_n16480__ & new_new_n16481__;
  assign new_new_n16483__ = new_new_n16480__ & ~new_new_n16481__;
  assign new_new_n16484__ = ~new_new_n16482__ & ~new_new_n16483__;
  assign new_new_n16485__ = ~pi089 & ~new_new_n16484__;
  assign new_new_n16486__ = pi089 & new_new_n16484__;
  assign new_new_n16487__ = ~new_new_n16165__ & po011;
  assign new_new_n16488__ = pi087 & ~po011;
  assign new_new_n16489__ = ~new_new_n16487__ & ~new_new_n16488__;
  assign new_new_n16490__ = ~new_new_n15905__ & ~new_new_n15906__;
  assign new_new_n16491__ = ~new_new_n16489__ & new_new_n16490__;
  assign new_new_n16492__ = new_new_n16489__ & ~new_new_n16490__;
  assign new_new_n16493__ = ~new_new_n16491__ & ~new_new_n16492__;
  assign new_new_n16494__ = pi088 & new_new_n16493__;
  assign new_new_n16495__ = ~pi088 & ~new_new_n16493__;
  assign new_new_n16496__ = ~new_new_n15914__ & ~new_new_n15915__;
  assign new_new_n16497__ = ~new_new_n16163__ & po011;
  assign new_new_n16498__ = ~pi086 & ~po011;
  assign new_new_n16499__ = ~new_new_n16497__ & ~new_new_n16498__;
  assign new_new_n16500__ = new_new_n16496__ & ~new_new_n16499__;
  assign new_new_n16501__ = ~new_new_n16496__ & new_new_n16499__;
  assign new_new_n16502__ = ~new_new_n16500__ & ~new_new_n16501__;
  assign new_new_n16503__ = pi087 & ~new_new_n16502__;
  assign new_new_n16504__ = ~pi087 & new_new_n16502__;
  assign new_new_n16505__ = ~pi085 & ~new_new_n16161__;
  assign new_new_n16506__ = pi085 & new_new_n16161__;
  assign new_new_n16507__ = ~new_new_n16505__ & ~new_new_n16506__;
  assign new_new_n16508__ = po011 & new_new_n16507__;
  assign new_new_n16509__ = new_new_n15922__ & new_new_n16508__;
  assign new_new_n16510__ = ~new_new_n15922__ & ~new_new_n16508__;
  assign new_new_n16511__ = ~new_new_n16509__ & ~new_new_n16510__;
  assign new_new_n16512__ = ~pi086 & ~new_new_n16511__;
  assign new_new_n16513__ = pi086 & new_new_n16511__;
  assign new_new_n16514__ = ~pi084 & ~new_new_n16159__;
  assign new_new_n16515__ = pi084 & new_new_n16159__;
  assign new_new_n16516__ = ~new_new_n16514__ & ~new_new_n16515__;
  assign new_new_n16517__ = po011 & new_new_n16516__;
  assign new_new_n16518__ = new_new_n15931__ & new_new_n16517__;
  assign new_new_n16519__ = ~new_new_n15931__ & ~new_new_n16517__;
  assign new_new_n16520__ = ~new_new_n16518__ & ~new_new_n16519__;
  assign new_new_n16521__ = ~pi085 & ~new_new_n16520__;
  assign new_new_n16522__ = pi085 & new_new_n16520__;
  assign new_new_n16523__ = ~new_new_n15941__ & ~new_new_n15942__;
  assign new_new_n16524__ = ~new_new_n16157__ & po011;
  assign new_new_n16525__ = ~pi083 & ~po011;
  assign new_new_n16526__ = ~new_new_n16524__ & ~new_new_n16525__;
  assign new_new_n16527__ = new_new_n16523__ & ~new_new_n16526__;
  assign new_new_n16528__ = ~new_new_n16523__ & new_new_n16526__;
  assign new_new_n16529__ = ~new_new_n16527__ & ~new_new_n16528__;
  assign new_new_n16530__ = ~pi084 & new_new_n16529__;
  assign new_new_n16531__ = pi084 & ~new_new_n16529__;
  assign new_new_n16532__ = ~pi082 & ~new_new_n16155__;
  assign new_new_n16533__ = pi082 & new_new_n16155__;
  assign new_new_n16534__ = ~new_new_n16532__ & ~new_new_n16533__;
  assign new_new_n16535__ = po011 & new_new_n16534__;
  assign new_new_n16536__ = new_new_n15949__ & new_new_n16535__;
  assign new_new_n16537__ = ~new_new_n15949__ & ~new_new_n16535__;
  assign new_new_n16538__ = ~new_new_n16536__ & ~new_new_n16537__;
  assign new_new_n16539__ = ~pi083 & ~new_new_n16538__;
  assign new_new_n16540__ = pi083 & new_new_n16538__;
  assign new_new_n16541__ = ~new_new_n15959__ & ~new_new_n15960__;
  assign new_new_n16542__ = ~new_new_n16153__ & po011;
  assign new_new_n16543__ = ~pi081 & ~po011;
  assign new_new_n16544__ = ~new_new_n16542__ & ~new_new_n16543__;
  assign new_new_n16545__ = new_new_n16541__ & ~new_new_n16544__;
  assign new_new_n16546__ = ~new_new_n16541__ & new_new_n16544__;
  assign new_new_n16547__ = ~new_new_n16545__ & ~new_new_n16546__;
  assign new_new_n16548__ = pi082 & ~new_new_n16547__;
  assign new_new_n16549__ = ~pi082 & new_new_n16547__;
  assign new_new_n16550__ = ~pi080 & ~new_new_n16151__;
  assign new_new_n16551__ = pi080 & new_new_n16151__;
  assign new_new_n16552__ = ~new_new_n16550__ & ~new_new_n16551__;
  assign new_new_n16553__ = po011 & new_new_n16552__;
  assign new_new_n16554__ = new_new_n15967__ & new_new_n16553__;
  assign new_new_n16555__ = ~new_new_n15967__ & ~new_new_n16553__;
  assign new_new_n16556__ = ~new_new_n16554__ & ~new_new_n16555__;
  assign new_new_n16557__ = pi081 & new_new_n16556__;
  assign new_new_n16558__ = ~pi081 & ~new_new_n16556__;
  assign new_new_n16559__ = ~new_new_n16149__ & po011;
  assign new_new_n16560__ = pi079 & ~po011;
  assign new_new_n16561__ = ~new_new_n16559__ & ~new_new_n16560__;
  assign new_new_n16562__ = ~new_new_n15977__ & ~new_new_n15978__;
  assign new_new_n16563__ = ~new_new_n16561__ & new_new_n16562__;
  assign new_new_n16564__ = new_new_n16561__ & ~new_new_n16562__;
  assign new_new_n16565__ = ~new_new_n16563__ & ~new_new_n16564__;
  assign new_new_n16566__ = pi080 & new_new_n16565__;
  assign new_new_n16567__ = ~pi080 & ~new_new_n16565__;
  assign new_new_n16568__ = pi078 & ~new_new_n16147__;
  assign new_new_n16569__ = ~pi078 & new_new_n16147__;
  assign new_new_n16570__ = ~new_new_n16568__ & ~new_new_n16569__;
  assign new_new_n16571__ = po011 & new_new_n16570__;
  assign new_new_n16572__ = new_new_n15985__ & new_new_n16571__;
  assign new_new_n16573__ = ~new_new_n15985__ & ~new_new_n16571__;
  assign new_new_n16574__ = ~new_new_n16572__ & ~new_new_n16573__;
  assign new_new_n16575__ = pi079 & ~new_new_n16574__;
  assign new_new_n16576__ = ~pi079 & new_new_n16574__;
  assign new_new_n16577__ = pi077 & ~new_new_n16145__;
  assign new_new_n16578__ = ~pi077 & new_new_n16145__;
  assign new_new_n16579__ = ~new_new_n16577__ & ~new_new_n16578__;
  assign new_new_n16580__ = po011 & new_new_n16579__;
  assign new_new_n16581__ = new_new_n15994__ & new_new_n16580__;
  assign new_new_n16582__ = ~new_new_n15994__ & ~new_new_n16580__;
  assign new_new_n16583__ = ~new_new_n16581__ & ~new_new_n16582__;
  assign new_new_n16584__ = pi078 & ~new_new_n16583__;
  assign new_new_n16585__ = ~pi078 & new_new_n16583__;
  assign new_new_n16586__ = ~new_new_n16004__ & ~new_new_n16005__;
  assign new_new_n16587__ = ~new_new_n16143__ & po011;
  assign new_new_n16588__ = pi076 & ~po011;
  assign new_new_n16589__ = ~new_new_n16587__ & ~new_new_n16588__;
  assign new_new_n16590__ = new_new_n16586__ & ~new_new_n16589__;
  assign new_new_n16591__ = ~new_new_n16586__ & new_new_n16589__;
  assign new_new_n16592__ = ~new_new_n16590__ & ~new_new_n16591__;
  assign new_new_n16593__ = ~pi077 & ~new_new_n16592__;
  assign new_new_n16594__ = pi077 & new_new_n16592__;
  assign new_new_n16595__ = pi075 & ~new_new_n16141__;
  assign new_new_n16596__ = ~pi075 & new_new_n16141__;
  assign new_new_n16597__ = ~new_new_n16595__ & ~new_new_n16596__;
  assign new_new_n16598__ = po011 & new_new_n16597__;
  assign new_new_n16599__ = new_new_n16012__ & new_new_n16598__;
  assign new_new_n16600__ = ~new_new_n16012__ & ~new_new_n16598__;
  assign new_new_n16601__ = ~new_new_n16599__ & ~new_new_n16600__;
  assign new_new_n16602__ = pi076 & ~new_new_n16601__;
  assign new_new_n16603__ = ~pi076 & new_new_n16601__;
  assign new_new_n16604__ = pi074 & ~new_new_n16139__;
  assign new_new_n16605__ = ~pi074 & new_new_n16139__;
  assign new_new_n16606__ = ~new_new_n16604__ & ~new_new_n16605__;
  assign new_new_n16607__ = po011 & new_new_n16606__;
  assign new_new_n16608__ = ~new_new_n16021__ & ~new_new_n16607__;
  assign new_new_n16609__ = new_new_n16021__ & new_new_n16607__;
  assign new_new_n16610__ = ~new_new_n16608__ & ~new_new_n16609__;
  assign new_new_n16611__ = pi075 & ~new_new_n16610__;
  assign new_new_n16612__ = ~pi075 & new_new_n16610__;
  assign new_new_n16613__ = ~new_new_n16137__ & po011;
  assign new_new_n16614__ = pi073 & ~po011;
  assign new_new_n16615__ = ~new_new_n16613__ & ~new_new_n16614__;
  assign new_new_n16616__ = ~new_new_n16031__ & ~new_new_n16032__;
  assign new_new_n16617__ = ~new_new_n16615__ & new_new_n16616__;
  assign new_new_n16618__ = new_new_n16615__ & ~new_new_n16616__;
  assign new_new_n16619__ = ~new_new_n16617__ & ~new_new_n16618__;
  assign new_new_n16620__ = ~pi074 & ~new_new_n16619__;
  assign new_new_n16621__ = pi074 & new_new_n16619__;
  assign new_new_n16622__ = pi072 & ~new_new_n16135__;
  assign new_new_n16623__ = ~pi072 & new_new_n16135__;
  assign new_new_n16624__ = ~new_new_n16622__ & ~new_new_n16623__;
  assign new_new_n16625__ = po011 & new_new_n16624__;
  assign new_new_n16626__ = new_new_n16039__ & new_new_n16625__;
  assign new_new_n16627__ = ~new_new_n16039__ & ~new_new_n16625__;
  assign new_new_n16628__ = ~new_new_n16626__ & ~new_new_n16627__;
  assign new_new_n16629__ = ~pi073 & new_new_n16628__;
  assign new_new_n16630__ = pi073 & ~new_new_n16628__;
  assign new_new_n16631__ = pi071 & ~new_new_n16133__;
  assign new_new_n16632__ = ~pi071 & new_new_n16133__;
  assign new_new_n16633__ = ~new_new_n16631__ & ~new_new_n16632__;
  assign new_new_n16634__ = po011 & new_new_n16633__;
  assign new_new_n16635__ = new_new_n16048__ & new_new_n16634__;
  assign new_new_n16636__ = ~new_new_n16048__ & ~new_new_n16634__;
  assign new_new_n16637__ = ~new_new_n16635__ & ~new_new_n16636__;
  assign new_new_n16638__ = ~pi072 & new_new_n16637__;
  assign new_new_n16639__ = pi072 & ~new_new_n16637__;
  assign new_new_n16640__ = ~new_new_n16058__ & ~new_new_n16059__;
  assign new_new_n16641__ = new_new_n16131__ & po011;
  assign new_new_n16642__ = ~pi070 & ~po011;
  assign new_new_n16643__ = ~new_new_n16641__ & ~new_new_n16642__;
  assign new_new_n16644__ = ~new_new_n16640__ & ~new_new_n16643__;
  assign new_new_n16645__ = new_new_n16640__ & new_new_n16643__;
  assign new_new_n16646__ = ~new_new_n16644__ & ~new_new_n16645__;
  assign new_new_n16647__ = ~pi071 & ~new_new_n16646__;
  assign new_new_n16648__ = pi071 & new_new_n16646__;
  assign new_new_n16649__ = ~new_new_n16121__ & ~new_new_n16122__;
  assign new_new_n16650__ = po011 & new_new_n16649__;
  assign new_new_n16651__ = new_new_n16129__ & new_new_n16650__;
  assign new_new_n16652__ = ~new_new_n16129__ & ~new_new_n16650__;
  assign new_new_n16653__ = ~new_new_n16651__ & ~new_new_n16652__;
  assign new_new_n16654__ = pi070 & ~new_new_n16653__;
  assign new_new_n16655__ = ~pi070 & new_new_n16653__;
  assign new_new_n16656__ = ~new_new_n16118__ & po011;
  assign new_new_n16657__ = pi068 & ~po011;
  assign new_new_n16658__ = ~new_new_n16656__ & ~new_new_n16657__;
  assign new_new_n16659__ = ~new_new_n16067__ & ~new_new_n16068__;
  assign new_new_n16660__ = ~new_new_n16658__ & new_new_n16659__;
  assign new_new_n16661__ = new_new_n16658__ & ~new_new_n16659__;
  assign new_new_n16662__ = ~new_new_n16660__ & ~new_new_n16661__;
  assign new_new_n16663__ = ~pi069 & ~new_new_n16662__;
  assign new_new_n16664__ = pi069 & new_new_n16662__;
  assign new_new_n16665__ = ~new_new_n16088__ & po011;
  assign new_new_n16666__ = ~new_new_n16114__ & new_new_n16665__;
  assign new_new_n16667__ = new_new_n16113__ & ~new_new_n16666__;
  assign new_new_n16668__ = new_new_n16115__ & new_new_n16665__;
  assign new_new_n16669__ = ~new_new_n16667__ & ~new_new_n16668__;
  assign new_new_n16670__ = ~pi067 & ~new_new_n16669__;
  assign new_new_n16671__ = pi067 & new_new_n16669__;
  assign new_new_n16672__ = ~pi010 & pi064;
  assign new_new_n16673__ = pi064 & po011;
  assign new_new_n16674__ = pi011 & ~new_new_n16673__;
  assign new_new_n16675__ = ~pi011 & new_new_n16673__;
  assign new_new_n16676__ = ~new_new_n16674__ & ~new_new_n16675__;
  assign new_new_n16677__ = pi065 & new_new_n16676__;
  assign new_new_n16678__ = ~new_new_n16672__ & ~new_new_n16677__;
  assign new_new_n16679__ = ~pi065 & ~new_new_n16676__;
  assign new_new_n16680__ = ~new_new_n16678__ & ~new_new_n16679__;
  assign new_new_n16681__ = ~pi066 & ~new_new_n16680__;
  assign new_new_n16682__ = pi066 & new_new_n16680__;
  assign new_new_n16683__ = ~new_new_n332__ & po011;
  assign new_new_n16684__ = ~new_new_n16084__ & ~new_new_n16683__;
  assign new_new_n16685__ = ~pi065 & ~po012;
  assign new_new_n16686__ = ~new_new_n16095__ & ~new_new_n16685__;
  assign new_new_n16687__ = po012 & ~po011;
  assign new_new_n16688__ = ~pi011 & ~new_new_n403__;
  assign new_new_n16689__ = new_new_n16686__ & new_new_n16688__;
  assign new_new_n16690__ = ~new_new_n16687__ & new_new_n16689__;
  assign new_new_n16691__ = pi065 & ~new_new_n16673__;
  assign new_new_n16692__ = pi011 & ~new_new_n16686__;
  assign new_new_n16693__ = ~new_new_n16691__ & new_new_n16692__;
  assign new_new_n16694__ = ~new_new_n16684__ & ~new_new_n16690__;
  assign new_new_n16695__ = ~new_new_n16693__ & new_new_n16694__;
  assign new_new_n16696__ = ~pi012 & ~new_new_n16695__;
  assign new_new_n16697__ = ~pi065 & ~po011;
  assign new_new_n16698__ = ~pi011 & ~new_new_n16686__;
  assign new_new_n16699__ = ~new_new_n16697__ & new_new_n16698__;
  assign new_new_n16700__ = ~new_new_n16687__ & ~new_new_n16699__;
  assign new_new_n16701__ = pi064 & ~new_new_n16700__;
  assign new_new_n16702__ = pi065 & po011;
  assign new_new_n16703__ = ~new_new_n16084__ & ~new_new_n16702__;
  assign new_new_n16704__ = pi011 & ~new_new_n16095__;
  assign new_new_n16705__ = pi064 & ~new_new_n16704__;
  assign new_new_n16706__ = ~new_new_n16703__ & ~new_new_n16705__;
  assign new_new_n16707__ = ~new_new_n16701__ & ~new_new_n16706__;
  assign new_new_n16708__ = pi012 & ~new_new_n16707__;
  assign new_new_n16709__ = ~new_new_n16696__ & ~new_new_n16708__;
  assign new_new_n16710__ = ~new_new_n16682__ & new_new_n16709__;
  assign new_new_n16711__ = ~new_new_n16681__ & ~new_new_n16710__;
  assign new_new_n16712__ = ~new_new_n16671__ & ~new_new_n16711__;
  assign new_new_n16713__ = ~new_new_n16670__ & ~new_new_n16712__;
  assign new_new_n16714__ = pi068 & new_new_n16713__;
  assign new_new_n16715__ = ~pi068 & ~new_new_n16713__;
  assign new_new_n16716__ = ~new_new_n16074__ & ~new_new_n16075__;
  assign new_new_n16717__ = ~new_new_n16116__ & po011;
  assign new_new_n16718__ = pi067 & ~po011;
  assign new_new_n16719__ = ~new_new_n16717__ & ~new_new_n16718__;
  assign new_new_n16720__ = new_new_n16716__ & ~new_new_n16719__;
  assign new_new_n16721__ = ~new_new_n16716__ & new_new_n16719__;
  assign new_new_n16722__ = ~new_new_n16720__ & ~new_new_n16721__;
  assign new_new_n16723__ = ~new_new_n16715__ & new_new_n16722__;
  assign new_new_n16724__ = ~new_new_n16714__ & ~new_new_n16723__;
  assign new_new_n16725__ = ~new_new_n16664__ & new_new_n16724__;
  assign new_new_n16726__ = ~new_new_n16663__ & ~new_new_n16725__;
  assign new_new_n16727__ = ~new_new_n16655__ & new_new_n16726__;
  assign new_new_n16728__ = ~new_new_n16654__ & ~new_new_n16727__;
  assign new_new_n16729__ = ~new_new_n16648__ & new_new_n16728__;
  assign new_new_n16730__ = ~new_new_n16647__ & ~new_new_n16729__;
  assign new_new_n16731__ = ~new_new_n16639__ & ~new_new_n16730__;
  assign new_new_n16732__ = ~new_new_n16638__ & ~new_new_n16731__;
  assign new_new_n16733__ = ~new_new_n16630__ & ~new_new_n16732__;
  assign new_new_n16734__ = ~new_new_n16629__ & ~new_new_n16733__;
  assign new_new_n16735__ = ~new_new_n16621__ & ~new_new_n16734__;
  assign new_new_n16736__ = ~new_new_n16620__ & ~new_new_n16735__;
  assign new_new_n16737__ = ~new_new_n16612__ & new_new_n16736__;
  assign new_new_n16738__ = ~new_new_n16611__ & ~new_new_n16737__;
  assign new_new_n16739__ = ~new_new_n16603__ & ~new_new_n16738__;
  assign new_new_n16740__ = ~new_new_n16602__ & ~new_new_n16739__;
  assign new_new_n16741__ = ~new_new_n16594__ & new_new_n16740__;
  assign new_new_n16742__ = ~new_new_n16593__ & ~new_new_n16741__;
  assign new_new_n16743__ = ~new_new_n16585__ & new_new_n16742__;
  assign new_new_n16744__ = ~new_new_n16584__ & ~new_new_n16743__;
  assign new_new_n16745__ = ~new_new_n16576__ & ~new_new_n16744__;
  assign new_new_n16746__ = ~new_new_n16575__ & ~new_new_n16745__;
  assign new_new_n16747__ = ~new_new_n16567__ & ~new_new_n16746__;
  assign new_new_n16748__ = ~new_new_n16566__ & ~new_new_n16747__;
  assign new_new_n16749__ = ~new_new_n16558__ & ~new_new_n16748__;
  assign new_new_n16750__ = ~new_new_n16557__ & ~new_new_n16749__;
  assign new_new_n16751__ = ~new_new_n16549__ & ~new_new_n16750__;
  assign new_new_n16752__ = ~new_new_n16548__ & ~new_new_n16751__;
  assign new_new_n16753__ = ~new_new_n16540__ & new_new_n16752__;
  assign new_new_n16754__ = ~new_new_n16539__ & ~new_new_n16753__;
  assign new_new_n16755__ = ~new_new_n16531__ & ~new_new_n16754__;
  assign new_new_n16756__ = ~new_new_n16530__ & ~new_new_n16755__;
  assign new_new_n16757__ = ~new_new_n16522__ & ~new_new_n16756__;
  assign new_new_n16758__ = ~new_new_n16521__ & ~new_new_n16757__;
  assign new_new_n16759__ = ~new_new_n16513__ & ~new_new_n16758__;
  assign new_new_n16760__ = ~new_new_n16512__ & ~new_new_n16759__;
  assign new_new_n16761__ = ~new_new_n16504__ & new_new_n16760__;
  assign new_new_n16762__ = ~new_new_n16503__ & ~new_new_n16761__;
  assign new_new_n16763__ = ~new_new_n16495__ & ~new_new_n16762__;
  assign new_new_n16764__ = ~new_new_n16494__ & ~new_new_n16763__;
  assign new_new_n16765__ = ~new_new_n16486__ & new_new_n16764__;
  assign new_new_n16766__ = ~new_new_n16485__ & ~new_new_n16765__;
  assign new_new_n16767__ = ~new_new_n16477__ & ~new_new_n16766__;
  assign new_new_n16768__ = ~new_new_n16476__ & ~new_new_n16767__;
  assign new_new_n16769__ = ~new_new_n16468__ & ~new_new_n16768__;
  assign new_new_n16770__ = ~new_new_n16467__ & ~new_new_n16769__;
  assign new_new_n16771__ = ~new_new_n16459__ & new_new_n16770__;
  assign new_new_n16772__ = ~new_new_n16458__ & ~new_new_n16771__;
  assign new_new_n16773__ = ~new_new_n16450__ & ~new_new_n16772__;
  assign new_new_n16774__ = ~new_new_n16449__ & ~new_new_n16773__;
  assign new_new_n16775__ = ~new_new_n16441__ & new_new_n16774__;
  assign new_new_n16776__ = ~new_new_n16440__ & ~new_new_n16775__;
  assign new_new_n16777__ = ~new_new_n16432__ & new_new_n16776__;
  assign new_new_n16778__ = ~new_new_n16431__ & ~new_new_n16777__;
  assign new_new_n16779__ = ~new_new_n16423__ & new_new_n16778__;
  assign new_new_n16780__ = ~new_new_n16422__ & ~new_new_n16779__;
  assign new_new_n16781__ = ~new_new_n16414__ & ~new_new_n16780__;
  assign new_new_n16782__ = ~new_new_n16413__ & ~new_new_n16781__;
  assign new_new_n16783__ = ~new_new_n16405__ & ~new_new_n16782__;
  assign new_new_n16784__ = ~new_new_n16404__ & ~new_new_n16783__;
  assign new_new_n16785__ = ~new_new_n16396__ & new_new_n16784__;
  assign new_new_n16786__ = ~new_new_n16395__ & ~new_new_n16785__;
  assign new_new_n16787__ = ~new_new_n16387__ & new_new_n16786__;
  assign new_new_n16788__ = ~new_new_n16386__ & ~new_new_n16787__;
  assign new_new_n16789__ = ~new_new_n16378__ & ~new_new_n16788__;
  assign new_new_n16790__ = ~new_new_n16377__ & ~new_new_n16789__;
  assign new_new_n16791__ = ~new_new_n16369__ & ~new_new_n16790__;
  assign new_new_n16792__ = ~new_new_n16368__ & ~new_new_n16791__;
  assign new_new_n16793__ = ~new_new_n16360__ & ~new_new_n16792__;
  assign new_new_n16794__ = ~new_new_n16359__ & ~new_new_n16793__;
  assign new_new_n16795__ = ~new_new_n16351__ & new_new_n16794__;
  assign new_new_n16796__ = ~new_new_n16350__ & ~new_new_n16795__;
  assign new_new_n16797__ = ~new_new_n16342__ & new_new_n16796__;
  assign new_new_n16798__ = ~new_new_n16341__ & ~new_new_n16797__;
  assign new_new_n16799__ = ~new_new_n16333__ & ~new_new_n16798__;
  assign new_new_n16800__ = ~new_new_n16332__ & ~new_new_n16799__;
  assign new_new_n16801__ = ~new_new_n16324__ & ~new_new_n16800__;
  assign new_new_n16802__ = ~new_new_n16323__ & ~new_new_n16801__;
  assign new_new_n16803__ = ~new_new_n16315__ & ~new_new_n16802__;
  assign new_new_n16804__ = ~new_new_n16314__ & ~new_new_n16803__;
  assign new_new_n16805__ = ~new_new_n16306__ & new_new_n16804__;
  assign new_new_n16806__ = ~new_new_n16305__ & ~new_new_n16805__;
  assign new_new_n16807__ = ~new_new_n16297__ & ~new_new_n16806__;
  assign new_new_n16808__ = ~new_new_n16296__ & ~new_new_n16807__;
  assign new_new_n16809__ = ~new_new_n16288__ & ~new_new_n16808__;
  assign new_new_n16810__ = ~new_new_n16287__ & ~new_new_n16809__;
  assign new_new_n16811__ = ~new_new_n16279__ & ~new_new_n16810__;
  assign new_new_n16812__ = ~new_new_n16278__ & ~new_new_n16811__;
  assign new_new_n16813__ = ~new_new_n16270__ & ~new_new_n16812__;
  assign new_new_n16814__ = ~new_new_n16269__ & ~new_new_n16813__;
  assign new_new_n16815__ = ~new_new_n16261__ & ~new_new_n16814__;
  assign new_new_n16816__ = ~new_new_n16260__ & ~new_new_n16815__;
  assign new_new_n16817__ = ~new_new_n16252__ & ~new_new_n16816__;
  assign new_new_n16818__ = ~new_new_n16251__ & ~new_new_n16817__;
  assign new_new_n16819__ = ~new_new_n16243__ & new_new_n16818__;
  assign new_new_n16820__ = ~new_new_n16242__ & ~new_new_n16819__;
  assign new_new_n16821__ = ~pi117 & ~new_new_n16820__;
  assign new_new_n16822__ = new_new_n269__ & new_new_n16229__;
  assign new_new_n16823__ = ~pi117 & new_new_n16229__;
  assign new_new_n16824__ = pi117 & ~new_new_n16229__;
  assign new_new_n16825__ = ~pi121 & new_new_n264__;
  assign new_new_n16826__ = ~pi120 & new_new_n16825__;
  assign new_new_n16827__ = ~pi119 & new_new_n16826__;
  assign new_new_n16828__ = ~pi118 & new_new_n16827__;
  assign new_new_n16829__ = ~new_new_n16823__ & new_new_n16828__;
  assign new_new_n16830__ = ~new_new_n16824__ & new_new_n16829__;
  assign new_new_n16831__ = ~new_new_n16822__ & ~new_new_n16830__;
  assign new_new_n16832__ = new_new_n16820__ & ~new_new_n16822__;
  assign po010 = ~new_new_n16831__ & ~new_new_n16832__;
  assign new_new_n16834__ = pi117 & new_new_n16820__;
  assign new_new_n16835__ = ~new_new_n16821__ & ~new_new_n16834__;
  assign new_new_n16836__ = po010 & new_new_n16835__;
  assign new_new_n16837__ = new_new_n16229__ & ~new_new_n16836__;
  assign new_new_n16838__ = pi116 & new_new_n16818__;
  assign new_new_n16839__ = ~pi116 & ~new_new_n16818__;
  assign new_new_n16840__ = ~new_new_n16838__ & ~new_new_n16839__;
  assign new_new_n16841__ = ~new_new_n16831__ & ~new_new_n16840__;
  assign new_new_n16842__ = ~new_new_n16241__ & ~new_new_n16841__;
  assign new_new_n16843__ = new_new_n16241__ & new_new_n16822__;
  assign new_new_n16844__ = ~new_new_n16840__ & new_new_n16843__;
  assign new_new_n16845__ = ~new_new_n16842__ & ~new_new_n16844__;
  assign new_new_n16846__ = ~pi117 & ~new_new_n16845__;
  assign new_new_n16847__ = pi117 & new_new_n16845__;
  assign new_new_n16848__ = ~new_new_n16251__ & ~new_new_n16252__;
  assign new_new_n16849__ = pi115 & ~po010;
  assign new_new_n16850__ = ~new_new_n16816__ & po010;
  assign new_new_n16851__ = ~new_new_n16849__ & ~new_new_n16850__;
  assign new_new_n16852__ = new_new_n16848__ & new_new_n16851__;
  assign new_new_n16853__ = ~new_new_n16848__ & ~new_new_n16851__;
  assign new_new_n16854__ = ~new_new_n16852__ & ~new_new_n16853__;
  assign new_new_n16855__ = ~pi116 & new_new_n16854__;
  assign new_new_n16856__ = pi116 & ~new_new_n16854__;
  assign new_new_n16857__ = new_new_n16814__ & po010;
  assign new_new_n16858__ = ~pi114 & ~po010;
  assign new_new_n16859__ = ~new_new_n16857__ & ~new_new_n16858__;
  assign new_new_n16860__ = ~new_new_n16260__ & ~new_new_n16261__;
  assign new_new_n16861__ = ~new_new_n16859__ & ~new_new_n16860__;
  assign new_new_n16862__ = new_new_n16859__ & new_new_n16860__;
  assign new_new_n16863__ = ~new_new_n16861__ & ~new_new_n16862__;
  assign new_new_n16864__ = ~pi115 & ~new_new_n16863__;
  assign new_new_n16865__ = pi115 & new_new_n16863__;
  assign new_new_n16866__ = ~new_new_n16269__ & ~new_new_n16270__;
  assign new_new_n16867__ = pi113 & ~po010;
  assign new_new_n16868__ = ~new_new_n16812__ & po010;
  assign new_new_n16869__ = ~new_new_n16867__ & ~new_new_n16868__;
  assign new_new_n16870__ = new_new_n16866__ & new_new_n16869__;
  assign new_new_n16871__ = ~new_new_n16866__ & ~new_new_n16869__;
  assign new_new_n16872__ = ~new_new_n16870__ & ~new_new_n16871__;
  assign new_new_n16873__ = pi114 & ~new_new_n16872__;
  assign new_new_n16874__ = ~pi114 & new_new_n16872__;
  assign new_new_n16875__ = pi112 & ~new_new_n16810__;
  assign new_new_n16876__ = ~pi112 & new_new_n16810__;
  assign new_new_n16877__ = ~new_new_n16875__ & ~new_new_n16876__;
  assign new_new_n16878__ = po010 & new_new_n16877__;
  assign new_new_n16879__ = new_new_n16277__ & new_new_n16878__;
  assign new_new_n16880__ = ~new_new_n16277__ & ~new_new_n16878__;
  assign new_new_n16881__ = ~new_new_n16879__ & ~new_new_n16880__;
  assign new_new_n16882__ = ~pi113 & new_new_n16881__;
  assign new_new_n16883__ = pi113 & ~new_new_n16881__;
  assign new_new_n16884__ = new_new_n16808__ & po010;
  assign new_new_n16885__ = ~pi111 & ~po010;
  assign new_new_n16886__ = ~new_new_n16884__ & ~new_new_n16885__;
  assign new_new_n16887__ = ~new_new_n16287__ & ~new_new_n16288__;
  assign new_new_n16888__ = ~new_new_n16886__ & ~new_new_n16887__;
  assign new_new_n16889__ = new_new_n16886__ & new_new_n16887__;
  assign new_new_n16890__ = ~new_new_n16888__ & ~new_new_n16889__;
  assign new_new_n16891__ = ~pi112 & ~new_new_n16890__;
  assign new_new_n16892__ = pi112 & new_new_n16890__;
  assign new_new_n16893__ = ~new_new_n16296__ & ~new_new_n16297__;
  assign new_new_n16894__ = pi110 & ~po010;
  assign new_new_n16895__ = ~new_new_n16806__ & po010;
  assign new_new_n16896__ = ~new_new_n16894__ & ~new_new_n16895__;
  assign new_new_n16897__ = new_new_n16893__ & ~new_new_n16896__;
  assign new_new_n16898__ = ~new_new_n16893__ & new_new_n16896__;
  assign new_new_n16899__ = ~new_new_n16897__ & ~new_new_n16898__;
  assign new_new_n16900__ = pi111 & new_new_n16899__;
  assign new_new_n16901__ = ~pi111 & ~new_new_n16899__;
  assign new_new_n16902__ = ~new_new_n16305__ & ~new_new_n16306__;
  assign new_new_n16903__ = ~new_new_n16804__ & po010;
  assign new_new_n16904__ = ~pi109 & ~po010;
  assign new_new_n16905__ = ~new_new_n16903__ & ~new_new_n16904__;
  assign new_new_n16906__ = new_new_n16902__ & ~new_new_n16905__;
  assign new_new_n16907__ = ~new_new_n16902__ & new_new_n16905__;
  assign new_new_n16908__ = ~new_new_n16906__ & ~new_new_n16907__;
  assign new_new_n16909__ = pi110 & ~new_new_n16908__;
  assign new_new_n16910__ = ~pi110 & new_new_n16908__;
  assign new_new_n16911__ = ~new_new_n16323__ & ~new_new_n16324__;
  assign new_new_n16912__ = ~new_new_n16800__ & po010;
  assign new_new_n16913__ = ~pi107 & ~po010;
  assign new_new_n16914__ = ~new_new_n16912__ & ~new_new_n16913__;
  assign new_new_n16915__ = new_new_n16911__ & ~new_new_n16914__;
  assign new_new_n16916__ = ~new_new_n16911__ & new_new_n16914__;
  assign new_new_n16917__ = ~new_new_n16915__ & ~new_new_n16916__;
  assign new_new_n16918__ = pi108 & ~new_new_n16917__;
  assign new_new_n16919__ = ~pi108 & new_new_n16917__;
  assign new_new_n16920__ = ~new_new_n16332__ & ~new_new_n16333__;
  assign new_new_n16921__ = ~new_new_n16798__ & po010;
  assign new_new_n16922__ = ~pi106 & ~po010;
  assign new_new_n16923__ = ~new_new_n16921__ & ~new_new_n16922__;
  assign new_new_n16924__ = ~new_new_n16920__ & ~new_new_n16923__;
  assign new_new_n16925__ = new_new_n16920__ & new_new_n16923__;
  assign new_new_n16926__ = ~new_new_n16924__ & ~new_new_n16925__;
  assign new_new_n16927__ = ~pi107 & ~new_new_n16926__;
  assign new_new_n16928__ = pi107 & new_new_n16926__;
  assign new_new_n16929__ = new_new_n16796__ & po010;
  assign new_new_n16930__ = ~pi105 & ~po010;
  assign new_new_n16931__ = ~new_new_n16929__ & ~new_new_n16930__;
  assign new_new_n16932__ = ~new_new_n16341__ & ~new_new_n16342__;
  assign new_new_n16933__ = ~new_new_n16931__ & ~new_new_n16932__;
  assign new_new_n16934__ = new_new_n16931__ & new_new_n16932__;
  assign new_new_n16935__ = ~new_new_n16933__ & ~new_new_n16934__;
  assign new_new_n16936__ = ~pi106 & ~new_new_n16935__;
  assign new_new_n16937__ = pi106 & new_new_n16935__;
  assign new_new_n16938__ = ~new_new_n16350__ & ~new_new_n16351__;
  assign new_new_n16939__ = ~new_new_n16794__ & po010;
  assign new_new_n16940__ = ~pi104 & ~po010;
  assign new_new_n16941__ = ~new_new_n16939__ & ~new_new_n16940__;
  assign new_new_n16942__ = new_new_n16938__ & ~new_new_n16941__;
  assign new_new_n16943__ = ~new_new_n16938__ & new_new_n16941__;
  assign new_new_n16944__ = ~new_new_n16942__ & ~new_new_n16943__;
  assign new_new_n16945__ = pi105 & ~new_new_n16944__;
  assign new_new_n16946__ = ~pi105 & new_new_n16944__;
  assign new_new_n16947__ = ~pi103 & ~new_new_n16792__;
  assign new_new_n16948__ = pi103 & new_new_n16792__;
  assign new_new_n16949__ = ~new_new_n16947__ & ~new_new_n16948__;
  assign new_new_n16950__ = po010 & new_new_n16949__;
  assign new_new_n16951__ = new_new_n16358__ & new_new_n16950__;
  assign new_new_n16952__ = ~new_new_n16358__ & ~new_new_n16950__;
  assign new_new_n16953__ = ~new_new_n16951__ & ~new_new_n16952__;
  assign new_new_n16954__ = ~pi104 & ~new_new_n16953__;
  assign new_new_n16955__ = pi104 & new_new_n16953__;
  assign new_new_n16956__ = ~new_new_n16368__ & ~new_new_n16369__;
  assign new_new_n16957__ = ~new_new_n16790__ & po010;
  assign new_new_n16958__ = ~pi102 & ~po010;
  assign new_new_n16959__ = ~new_new_n16957__ & ~new_new_n16958__;
  assign new_new_n16960__ = new_new_n16956__ & ~new_new_n16959__;
  assign new_new_n16961__ = ~new_new_n16956__ & new_new_n16959__;
  assign new_new_n16962__ = ~new_new_n16960__ & ~new_new_n16961__;
  assign new_new_n16963__ = pi103 & ~new_new_n16962__;
  assign new_new_n16964__ = ~pi103 & new_new_n16962__;
  assign new_new_n16965__ = ~pi101 & ~new_new_n16788__;
  assign new_new_n16966__ = pi101 & new_new_n16788__;
  assign new_new_n16967__ = ~new_new_n16965__ & ~new_new_n16966__;
  assign new_new_n16968__ = po010 & new_new_n16967__;
  assign new_new_n16969__ = ~new_new_n16376__ & new_new_n16968__;
  assign new_new_n16970__ = new_new_n16376__ & ~new_new_n16968__;
  assign new_new_n16971__ = ~new_new_n16969__ & ~new_new_n16970__;
  assign new_new_n16972__ = pi102 & ~new_new_n16971__;
  assign new_new_n16973__ = ~pi102 & new_new_n16971__;
  assign new_new_n16974__ = ~new_new_n16786__ & po010;
  assign new_new_n16975__ = pi100 & ~po010;
  assign new_new_n16976__ = ~new_new_n16974__ & ~new_new_n16975__;
  assign new_new_n16977__ = ~new_new_n16386__ & ~new_new_n16387__;
  assign new_new_n16978__ = ~new_new_n16976__ & new_new_n16977__;
  assign new_new_n16979__ = new_new_n16976__ & ~new_new_n16977__;
  assign new_new_n16980__ = ~new_new_n16978__ & ~new_new_n16979__;
  assign new_new_n16981__ = ~pi101 & ~new_new_n16980__;
  assign new_new_n16982__ = pi101 & new_new_n16980__;
  assign new_new_n16983__ = ~new_new_n16395__ & ~new_new_n16396__;
  assign new_new_n16984__ = ~new_new_n16784__ & po010;
  assign new_new_n16985__ = ~pi099 & ~po010;
  assign new_new_n16986__ = ~new_new_n16984__ & ~new_new_n16985__;
  assign new_new_n16987__ = new_new_n16983__ & ~new_new_n16986__;
  assign new_new_n16988__ = ~new_new_n16983__ & new_new_n16986__;
  assign new_new_n16989__ = ~new_new_n16987__ & ~new_new_n16988__;
  assign new_new_n16990__ = ~pi100 & new_new_n16989__;
  assign new_new_n16991__ = pi100 & ~new_new_n16989__;
  assign new_new_n16992__ = ~pi098 & ~new_new_n16782__;
  assign new_new_n16993__ = pi098 & new_new_n16782__;
  assign new_new_n16994__ = ~new_new_n16992__ & ~new_new_n16993__;
  assign new_new_n16995__ = po010 & new_new_n16994__;
  assign new_new_n16996__ = new_new_n16403__ & new_new_n16995__;
  assign new_new_n16997__ = ~new_new_n16403__ & ~new_new_n16995__;
  assign new_new_n16998__ = ~new_new_n16996__ & ~new_new_n16997__;
  assign new_new_n16999__ = ~pi099 & ~new_new_n16998__;
  assign new_new_n17000__ = pi099 & new_new_n16998__;
  assign new_new_n17001__ = ~pi097 & ~new_new_n16780__;
  assign new_new_n17002__ = pi097 & new_new_n16780__;
  assign new_new_n17003__ = ~new_new_n17001__ & ~new_new_n17002__;
  assign new_new_n17004__ = po010 & new_new_n17003__;
  assign new_new_n17005__ = new_new_n16412__ & new_new_n17004__;
  assign new_new_n17006__ = ~new_new_n16412__ & ~new_new_n17004__;
  assign new_new_n17007__ = ~new_new_n17005__ & ~new_new_n17006__;
  assign new_new_n17008__ = ~pi098 & ~new_new_n17007__;
  assign new_new_n17009__ = pi098 & new_new_n17007__;
  assign new_new_n17010__ = ~new_new_n16422__ & ~new_new_n16423__;
  assign new_new_n17011__ = pi096 & ~po010;
  assign new_new_n17012__ = ~new_new_n16778__ & po010;
  assign new_new_n17013__ = ~new_new_n17011__ & ~new_new_n17012__;
  assign new_new_n17014__ = new_new_n17010__ & ~new_new_n17013__;
  assign new_new_n17015__ = ~new_new_n17010__ & new_new_n17013__;
  assign new_new_n17016__ = ~new_new_n17014__ & ~new_new_n17015__;
  assign new_new_n17017__ = ~pi097 & ~new_new_n17016__;
  assign new_new_n17018__ = pi097 & new_new_n17016__;
  assign new_new_n17019__ = ~new_new_n16431__ & ~new_new_n16432__;
  assign new_new_n17020__ = ~new_new_n16776__ & po010;
  assign new_new_n17021__ = ~pi095 & ~po010;
  assign new_new_n17022__ = ~new_new_n17020__ & ~new_new_n17021__;
  assign new_new_n17023__ = new_new_n17019__ & ~new_new_n17022__;
  assign new_new_n17024__ = ~new_new_n17019__ & new_new_n17022__;
  assign new_new_n17025__ = ~new_new_n17023__ & ~new_new_n17024__;
  assign new_new_n17026__ = ~pi096 & new_new_n17025__;
  assign new_new_n17027__ = pi096 & ~new_new_n17025__;
  assign new_new_n17028__ = ~new_new_n16774__ & po010;
  assign new_new_n17029__ = pi094 & ~po010;
  assign new_new_n17030__ = ~new_new_n17028__ & ~new_new_n17029__;
  assign new_new_n17031__ = ~new_new_n16440__ & ~new_new_n16441__;
  assign new_new_n17032__ = ~new_new_n17030__ & new_new_n17031__;
  assign new_new_n17033__ = new_new_n17030__ & ~new_new_n17031__;
  assign new_new_n17034__ = ~new_new_n17032__ & ~new_new_n17033__;
  assign new_new_n17035__ = ~pi095 & ~new_new_n17034__;
  assign new_new_n17036__ = pi095 & new_new_n17034__;
  assign new_new_n17037__ = ~new_new_n16772__ & po010;
  assign new_new_n17038__ = pi093 & ~po010;
  assign new_new_n17039__ = ~new_new_n17037__ & ~new_new_n17038__;
  assign new_new_n17040__ = ~new_new_n16449__ & ~new_new_n16450__;
  assign new_new_n17041__ = ~new_new_n17039__ & new_new_n17040__;
  assign new_new_n17042__ = new_new_n17039__ & ~new_new_n17040__;
  assign new_new_n17043__ = ~new_new_n17041__ & ~new_new_n17042__;
  assign new_new_n17044__ = pi094 & new_new_n17043__;
  assign new_new_n17045__ = ~pi094 & ~new_new_n17043__;
  assign new_new_n17046__ = ~new_new_n16458__ & ~new_new_n16459__;
  assign new_new_n17047__ = ~new_new_n16770__ & po010;
  assign new_new_n17048__ = ~pi092 & ~po010;
  assign new_new_n17049__ = ~new_new_n17047__ & ~new_new_n17048__;
  assign new_new_n17050__ = new_new_n17046__ & ~new_new_n17049__;
  assign new_new_n17051__ = ~new_new_n17046__ & new_new_n17049__;
  assign new_new_n17052__ = ~new_new_n17050__ & ~new_new_n17051__;
  assign new_new_n17053__ = pi093 & ~new_new_n17052__;
  assign new_new_n17054__ = ~pi093 & new_new_n17052__;
  assign new_new_n17055__ = ~new_new_n16467__ & ~new_new_n16468__;
  assign new_new_n17056__ = ~new_new_n16768__ & po010;
  assign new_new_n17057__ = ~pi091 & ~po010;
  assign new_new_n17058__ = ~new_new_n17056__ & ~new_new_n17057__;
  assign new_new_n17059__ = new_new_n17055__ & ~new_new_n17058__;
  assign new_new_n17060__ = ~new_new_n17055__ & new_new_n17058__;
  assign new_new_n17061__ = ~new_new_n17059__ & ~new_new_n17060__;
  assign new_new_n17062__ = pi092 & ~new_new_n17061__;
  assign new_new_n17063__ = ~pi092 & new_new_n17061__;
  assign new_new_n17064__ = ~pi090 & ~new_new_n16766__;
  assign new_new_n17065__ = pi090 & new_new_n16766__;
  assign new_new_n17066__ = ~new_new_n17064__ & ~new_new_n17065__;
  assign new_new_n17067__ = po010 & new_new_n17066__;
  assign new_new_n17068__ = ~new_new_n16475__ & ~new_new_n17067__;
  assign new_new_n17069__ = new_new_n16475__ & new_new_n17067__;
  assign new_new_n17070__ = ~new_new_n17068__ & ~new_new_n17069__;
  assign new_new_n17071__ = ~pi091 & ~new_new_n17070__;
  assign new_new_n17072__ = pi091 & new_new_n17070__;
  assign new_new_n17073__ = ~new_new_n16764__ & po010;
  assign new_new_n17074__ = pi089 & ~po010;
  assign new_new_n17075__ = ~new_new_n17073__ & ~new_new_n17074__;
  assign new_new_n17076__ = ~new_new_n16485__ & ~new_new_n16486__;
  assign new_new_n17077__ = ~new_new_n17075__ & new_new_n17076__;
  assign new_new_n17078__ = new_new_n17075__ & ~new_new_n17076__;
  assign new_new_n17079__ = ~new_new_n17077__ & ~new_new_n17078__;
  assign new_new_n17080__ = ~pi090 & ~new_new_n17079__;
  assign new_new_n17081__ = pi090 & new_new_n17079__;
  assign new_new_n17082__ = ~new_new_n16762__ & po010;
  assign new_new_n17083__ = pi088 & ~po010;
  assign new_new_n17084__ = ~new_new_n17082__ & ~new_new_n17083__;
  assign new_new_n17085__ = ~new_new_n16494__ & ~new_new_n16495__;
  assign new_new_n17086__ = ~new_new_n17084__ & new_new_n17085__;
  assign new_new_n17087__ = new_new_n17084__ & ~new_new_n17085__;
  assign new_new_n17088__ = ~new_new_n17086__ & ~new_new_n17087__;
  assign new_new_n17089__ = ~pi089 & ~new_new_n17088__;
  assign new_new_n17090__ = pi089 & new_new_n17088__;
  assign new_new_n17091__ = ~new_new_n16503__ & ~new_new_n16504__;
  assign new_new_n17092__ = ~new_new_n16760__ & po010;
  assign new_new_n17093__ = ~pi087 & ~po010;
  assign new_new_n17094__ = ~new_new_n17092__ & ~new_new_n17093__;
  assign new_new_n17095__ = new_new_n17091__ & ~new_new_n17094__;
  assign new_new_n17096__ = ~new_new_n17091__ & new_new_n17094__;
  assign new_new_n17097__ = ~new_new_n17095__ & ~new_new_n17096__;
  assign new_new_n17098__ = ~pi088 & new_new_n17097__;
  assign new_new_n17099__ = pi088 & ~new_new_n17097__;
  assign new_new_n17100__ = ~new_new_n16512__ & ~new_new_n16513__;
  assign new_new_n17101__ = ~new_new_n16758__ & po010;
  assign new_new_n17102__ = ~pi086 & ~po010;
  assign new_new_n17103__ = ~new_new_n17101__ & ~new_new_n17102__;
  assign new_new_n17104__ = new_new_n17100__ & ~new_new_n17103__;
  assign new_new_n17105__ = ~new_new_n17100__ & new_new_n17103__;
  assign new_new_n17106__ = ~new_new_n17104__ & ~new_new_n17105__;
  assign new_new_n17107__ = ~pi087 & new_new_n17106__;
  assign new_new_n17108__ = pi087 & ~new_new_n17106__;
  assign new_new_n17109__ = ~pi085 & ~new_new_n16756__;
  assign new_new_n17110__ = pi085 & new_new_n16756__;
  assign new_new_n17111__ = ~new_new_n17109__ & ~new_new_n17110__;
  assign new_new_n17112__ = po010 & new_new_n17111__;
  assign new_new_n17113__ = ~new_new_n16520__ & ~new_new_n17112__;
  assign new_new_n17114__ = new_new_n16520__ & new_new_n17112__;
  assign new_new_n17115__ = ~new_new_n17113__ & ~new_new_n17114__;
  assign new_new_n17116__ = ~pi086 & ~new_new_n17115__;
  assign new_new_n17117__ = pi086 & new_new_n17115__;
  assign new_new_n17118__ = ~new_new_n16530__ & ~new_new_n16531__;
  assign new_new_n17119__ = ~new_new_n16754__ & po010;
  assign new_new_n17120__ = ~pi084 & ~po010;
  assign new_new_n17121__ = ~new_new_n17119__ & ~new_new_n17120__;
  assign new_new_n17122__ = new_new_n17118__ & ~new_new_n17121__;
  assign new_new_n17123__ = ~new_new_n17118__ & new_new_n17121__;
  assign new_new_n17124__ = ~new_new_n17122__ & ~new_new_n17123__;
  assign new_new_n17125__ = ~pi085 & new_new_n17124__;
  assign new_new_n17126__ = pi085 & ~new_new_n17124__;
  assign new_new_n17127__ = ~new_new_n16752__ & po010;
  assign new_new_n17128__ = pi083 & ~po010;
  assign new_new_n17129__ = ~new_new_n17127__ & ~new_new_n17128__;
  assign new_new_n17130__ = ~new_new_n16539__ & ~new_new_n16540__;
  assign new_new_n17131__ = ~new_new_n17129__ & new_new_n17130__;
  assign new_new_n17132__ = new_new_n17129__ & ~new_new_n17130__;
  assign new_new_n17133__ = ~new_new_n17131__ & ~new_new_n17132__;
  assign new_new_n17134__ = ~pi084 & ~new_new_n17133__;
  assign new_new_n17135__ = pi084 & new_new_n17133__;
  assign new_new_n17136__ = pi082 & ~new_new_n16750__;
  assign new_new_n17137__ = ~pi082 & new_new_n16750__;
  assign new_new_n17138__ = ~new_new_n17136__ & ~new_new_n17137__;
  assign new_new_n17139__ = po010 & new_new_n17138__;
  assign new_new_n17140__ = new_new_n16547__ & new_new_n17139__;
  assign new_new_n17141__ = ~new_new_n16547__ & ~new_new_n17139__;
  assign new_new_n17142__ = ~new_new_n17140__ & ~new_new_n17141__;
  assign new_new_n17143__ = ~pi083 & new_new_n17142__;
  assign new_new_n17144__ = pi083 & ~new_new_n17142__;
  assign new_new_n17145__ = ~new_new_n16557__ & ~new_new_n16558__;
  assign new_new_n17146__ = pi081 & ~po010;
  assign new_new_n17147__ = ~new_new_n16748__ & po010;
  assign new_new_n17148__ = ~new_new_n17146__ & ~new_new_n17147__;
  assign new_new_n17149__ = new_new_n17145__ & ~new_new_n17148__;
  assign new_new_n17150__ = ~new_new_n17145__ & new_new_n17148__;
  assign new_new_n17151__ = ~new_new_n17149__ & ~new_new_n17150__;
  assign new_new_n17152__ = ~pi082 & ~new_new_n17151__;
  assign new_new_n17153__ = pi082 & new_new_n17151__;
  assign new_new_n17154__ = ~new_new_n16566__ & ~new_new_n16567__;
  assign new_new_n17155__ = pi080 & ~po010;
  assign new_new_n17156__ = ~new_new_n16746__ & po010;
  assign new_new_n17157__ = ~new_new_n17155__ & ~new_new_n17156__;
  assign new_new_n17158__ = new_new_n17154__ & ~new_new_n17157__;
  assign new_new_n17159__ = ~new_new_n17154__ & new_new_n17157__;
  assign new_new_n17160__ = ~new_new_n17158__ & ~new_new_n17159__;
  assign new_new_n17161__ = ~pi081 & ~new_new_n17160__;
  assign new_new_n17162__ = pi081 & new_new_n17160__;
  assign new_new_n17163__ = ~new_new_n16575__ & ~new_new_n16576__;
  assign new_new_n17164__ = pi079 & ~po010;
  assign new_new_n17165__ = ~new_new_n16744__ & po010;
  assign new_new_n17166__ = ~new_new_n17164__ & ~new_new_n17165__;
  assign new_new_n17167__ = new_new_n17163__ & ~new_new_n17166__;
  assign new_new_n17168__ = ~new_new_n17163__ & new_new_n17166__;
  assign new_new_n17169__ = ~new_new_n17167__ & ~new_new_n17168__;
  assign new_new_n17170__ = pi080 & new_new_n17169__;
  assign new_new_n17171__ = ~pi080 & ~new_new_n17169__;
  assign new_new_n17172__ = ~new_new_n16584__ & ~new_new_n16585__;
  assign new_new_n17173__ = ~new_new_n16742__ & po010;
  assign new_new_n17174__ = ~pi078 & ~po010;
  assign new_new_n17175__ = ~new_new_n17173__ & ~new_new_n17174__;
  assign new_new_n17176__ = new_new_n17172__ & ~new_new_n17175__;
  assign new_new_n17177__ = ~new_new_n17172__ & new_new_n17175__;
  assign new_new_n17178__ = ~new_new_n17176__ & ~new_new_n17177__;
  assign new_new_n17179__ = pi079 & ~new_new_n17178__;
  assign new_new_n17180__ = ~pi079 & new_new_n17178__;
  assign new_new_n17181__ = ~new_new_n16740__ & po010;
  assign new_new_n17182__ = pi077 & ~po010;
  assign new_new_n17183__ = ~new_new_n17181__ & ~new_new_n17182__;
  assign new_new_n17184__ = ~new_new_n16593__ & ~new_new_n16594__;
  assign new_new_n17185__ = ~new_new_n17183__ & new_new_n17184__;
  assign new_new_n17186__ = new_new_n17183__ & ~new_new_n17184__;
  assign new_new_n17187__ = ~new_new_n17185__ & ~new_new_n17186__;
  assign new_new_n17188__ = pi078 & new_new_n17187__;
  assign new_new_n17189__ = ~pi078 & ~new_new_n17187__;
  assign new_new_n17190__ = pi076 & ~new_new_n16738__;
  assign new_new_n17191__ = ~pi076 & new_new_n16738__;
  assign new_new_n17192__ = ~new_new_n17190__ & ~new_new_n17191__;
  assign new_new_n17193__ = po010 & new_new_n17192__;
  assign new_new_n17194__ = new_new_n16601__ & new_new_n17193__;
  assign new_new_n17195__ = ~new_new_n16601__ & ~new_new_n17193__;
  assign new_new_n17196__ = ~new_new_n17194__ & ~new_new_n17195__;
  assign new_new_n17197__ = pi077 & ~new_new_n17196__;
  assign new_new_n17198__ = ~pi077 & new_new_n17196__;
  assign new_new_n17199__ = new_new_n16736__ & po010;
  assign new_new_n17200__ = pi075 & ~po010;
  assign new_new_n17201__ = ~new_new_n17199__ & ~new_new_n17200__;
  assign new_new_n17202__ = ~new_new_n16611__ & ~new_new_n16612__;
  assign new_new_n17203__ = ~new_new_n17201__ & ~new_new_n17202__;
  assign new_new_n17204__ = new_new_n17201__ & new_new_n17202__;
  assign new_new_n17205__ = ~new_new_n17203__ & ~new_new_n17204__;
  assign new_new_n17206__ = pi076 & ~new_new_n17205__;
  assign new_new_n17207__ = ~pi076 & new_new_n17205__;
  assign new_new_n17208__ = ~new_new_n16620__ & ~new_new_n16621__;
  assign new_new_n17209__ = ~new_new_n16734__ & po010;
  assign new_new_n17210__ = ~pi074 & ~po010;
  assign new_new_n17211__ = ~new_new_n17209__ & ~new_new_n17210__;
  assign new_new_n17212__ = ~new_new_n17208__ & ~new_new_n17211__;
  assign new_new_n17213__ = new_new_n17208__ & new_new_n17211__;
  assign new_new_n17214__ = ~new_new_n17212__ & ~new_new_n17213__;
  assign new_new_n17215__ = pi075 & new_new_n17214__;
  assign new_new_n17216__ = ~pi075 & ~new_new_n17214__;
  assign new_new_n17217__ = new_new_n16732__ & po010;
  assign new_new_n17218__ = pi073 & ~po010;
  assign new_new_n17219__ = ~new_new_n17217__ & ~new_new_n17218__;
  assign new_new_n17220__ = ~new_new_n16629__ & ~new_new_n16630__;
  assign new_new_n17221__ = ~new_new_n17219__ & ~new_new_n17220__;
  assign new_new_n17222__ = new_new_n17219__ & new_new_n17220__;
  assign new_new_n17223__ = ~new_new_n17221__ & ~new_new_n17222__;
  assign new_new_n17224__ = pi074 & ~new_new_n17223__;
  assign new_new_n17225__ = ~pi074 & new_new_n17223__;
  assign new_new_n17226__ = new_new_n16730__ & po010;
  assign new_new_n17227__ = pi072 & ~po010;
  assign new_new_n17228__ = ~new_new_n17226__ & ~new_new_n17227__;
  assign new_new_n17229__ = ~new_new_n16638__ & ~new_new_n16639__;
  assign new_new_n17230__ = ~new_new_n17228__ & ~new_new_n17229__;
  assign new_new_n17231__ = new_new_n17228__ & new_new_n17229__;
  assign new_new_n17232__ = ~new_new_n17230__ & ~new_new_n17231__;
  assign new_new_n17233__ = pi073 & ~new_new_n17232__;
  assign new_new_n17234__ = ~pi073 & new_new_n17232__;
  assign new_new_n17235__ = new_new_n16728__ & po010;
  assign new_new_n17236__ = ~pi071 & ~po010;
  assign new_new_n17237__ = ~new_new_n17235__ & ~new_new_n17236__;
  assign new_new_n17238__ = ~new_new_n16647__ & ~new_new_n16648__;
  assign new_new_n17239__ = ~new_new_n17237__ & ~new_new_n17238__;
  assign new_new_n17240__ = new_new_n17237__ & new_new_n17238__;
  assign new_new_n17241__ = ~new_new_n17239__ & ~new_new_n17240__;
  assign new_new_n17242__ = ~pi072 & ~new_new_n17241__;
  assign new_new_n17243__ = pi072 & new_new_n17241__;
  assign new_new_n17244__ = ~new_new_n16654__ & ~new_new_n16655__;
  assign new_new_n17245__ = ~new_new_n16726__ & po010;
  assign new_new_n17246__ = ~pi070 & ~po010;
  assign new_new_n17247__ = ~new_new_n17245__ & ~new_new_n17246__;
  assign new_new_n17248__ = new_new_n17244__ & ~new_new_n17247__;
  assign new_new_n17249__ = ~new_new_n17244__ & new_new_n17247__;
  assign new_new_n17250__ = ~new_new_n17248__ & ~new_new_n17249__;
  assign new_new_n17251__ = pi071 & ~new_new_n17250__;
  assign new_new_n17252__ = ~pi071 & new_new_n17250__;
  assign new_new_n17253__ = ~new_new_n16724__ & po010;
  assign new_new_n17254__ = pi069 & ~po010;
  assign new_new_n17255__ = ~new_new_n17253__ & ~new_new_n17254__;
  assign new_new_n17256__ = ~new_new_n16663__ & ~new_new_n16664__;
  assign new_new_n17257__ = ~new_new_n17255__ & new_new_n17256__;
  assign new_new_n17258__ = new_new_n17255__ & ~new_new_n17256__;
  assign new_new_n17259__ = ~new_new_n17257__ & ~new_new_n17258__;
  assign new_new_n17260__ = pi070 & new_new_n17259__;
  assign new_new_n17261__ = ~pi070 & ~new_new_n17259__;
  assign new_new_n17262__ = ~new_new_n16670__ & ~new_new_n16671__;
  assign new_new_n17263__ = ~new_new_n16711__ & po010;
  assign new_new_n17264__ = ~pi067 & ~po010;
  assign new_new_n17265__ = ~new_new_n17263__ & ~new_new_n17264__;
  assign new_new_n17266__ = new_new_n17262__ & ~new_new_n17265__;
  assign new_new_n17267__ = ~new_new_n17262__ & new_new_n17265__;
  assign new_new_n17268__ = ~new_new_n17266__ & ~new_new_n17267__;
  assign new_new_n17269__ = ~pi068 & new_new_n17268__;
  assign new_new_n17270__ = pi068 & ~new_new_n17268__;
  assign new_new_n17271__ = ~new_new_n16681__ & ~new_new_n16682__;
  assign new_new_n17272__ = po010 & new_new_n17271__;
  assign new_new_n17273__ = new_new_n16709__ & ~new_new_n17272__;
  assign new_new_n17274__ = ~new_new_n16709__ & new_new_n17272__;
  assign new_new_n17275__ = ~new_new_n17273__ & ~new_new_n17274__;
  assign new_new_n17276__ = ~pi067 & ~new_new_n17275__;
  assign new_new_n17277__ = pi067 & new_new_n17275__;
  assign new_new_n17278__ = ~pi009 & pi065;
  assign new_new_n17279__ = new_new_n16672__ & ~new_new_n17278__;
  assign new_new_n17280__ = ~new_new_n16677__ & new_new_n17279__;
  assign new_new_n17281__ = ~new_new_n16679__ & new_new_n17280__;
  assign new_new_n17282__ = pi010 & ~pi064;
  assign new_new_n17283__ = new_new_n16677__ & new_new_n17282__;
  assign new_new_n17284__ = ~new_new_n17281__ & ~new_new_n17283__;
  assign new_new_n17285__ = po010 & ~new_new_n17284__;
  assign new_new_n17286__ = pi065 & po010;
  assign new_new_n17287__ = pi009 & ~new_new_n17286__;
  assign new_new_n17288__ = ~pi065 & ~po010;
  assign new_new_n17289__ = ~pi010 & ~new_new_n17288__;
  assign new_new_n17290__ = new_new_n17287__ & ~new_new_n17289__;
  assign new_new_n17291__ = ~new_new_n332__ & po010;
  assign new_new_n17292__ = ~pi010 & ~new_new_n332__;
  assign new_new_n17293__ = ~new_new_n426__ & ~new_new_n17292__;
  assign new_new_n17294__ = ~new_new_n17291__ & new_new_n17293__;
  assign new_new_n17295__ = ~new_new_n17290__ & ~new_new_n17294__;
  assign new_new_n17296__ = ~new_new_n16676__ & ~new_new_n17295__;
  assign new_new_n17297__ = pi064 & po010;
  assign new_new_n17298__ = pi065 & ~new_new_n17297__;
  assign new_new_n17299__ = ~pi010 & new_new_n17298__;
  assign new_new_n17300__ = new_new_n16676__ & po010;
  assign new_new_n17301__ = ~new_new_n16676__ & ~po010;
  assign new_new_n17302__ = ~new_new_n17300__ & ~new_new_n17301__;
  assign new_new_n17303__ = new_new_n17299__ & new_new_n17302__;
  assign new_new_n17304__ = ~pi010 & ~po010;
  assign new_new_n17305__ = ~pi065 & ~new_new_n17304__;
  assign new_new_n17306__ = pi010 & po010;
  assign new_new_n17307__ = ~pi009 & new_new_n16676__;
  assign new_new_n17308__ = ~new_new_n17306__ & new_new_n17307__;
  assign new_new_n17309__ = ~new_new_n17305__ & new_new_n17308__;
  assign new_new_n17310__ = pi009 & ~pi065;
  assign new_new_n17311__ = new_new_n17306__ & ~new_new_n17310__;
  assign new_new_n17312__ = ~new_new_n16677__ & ~new_new_n16679__;
  assign new_new_n17313__ = new_new_n17311__ & new_new_n17312__;
  assign new_new_n17314__ = ~new_new_n17309__ & ~new_new_n17313__;
  assign new_new_n17315__ = pi064 & ~new_new_n17314__;
  assign new_new_n17316__ = ~pi066 & ~new_new_n17303__;
  assign new_new_n17317__ = ~new_new_n17315__ & new_new_n17316__;
  assign new_new_n17318__ = ~new_new_n17285__ & ~new_new_n17296__;
  assign new_new_n17319__ = ~new_new_n17317__ & new_new_n17318__;
  assign new_new_n17320__ = ~new_new_n17277__ & ~new_new_n17319__;
  assign new_new_n17321__ = ~new_new_n17276__ & ~new_new_n17320__;
  assign new_new_n17322__ = ~new_new_n17270__ & ~new_new_n17321__;
  assign new_new_n17323__ = ~new_new_n17269__ & ~new_new_n17322__;
  assign new_new_n17324__ = pi069 & new_new_n17323__;
  assign new_new_n17325__ = ~pi069 & ~new_new_n17323__;
  assign new_new_n17326__ = ~new_new_n16714__ & ~new_new_n16715__;
  assign new_new_n17327__ = po010 & new_new_n17326__;
  assign new_new_n17328__ = new_new_n16722__ & new_new_n17327__;
  assign new_new_n17329__ = ~new_new_n16722__ & ~new_new_n17327__;
  assign new_new_n17330__ = ~new_new_n17328__ & ~new_new_n17329__;
  assign new_new_n17331__ = ~new_new_n17325__ & new_new_n17330__;
  assign new_new_n17332__ = ~new_new_n17324__ & ~new_new_n17331__;
  assign new_new_n17333__ = ~new_new_n17261__ & ~new_new_n17332__;
  assign new_new_n17334__ = ~new_new_n17260__ & ~new_new_n17333__;
  assign new_new_n17335__ = ~new_new_n17252__ & ~new_new_n17334__;
  assign new_new_n17336__ = ~new_new_n17251__ & ~new_new_n17335__;
  assign new_new_n17337__ = ~new_new_n17243__ & new_new_n17336__;
  assign new_new_n17338__ = ~new_new_n17242__ & ~new_new_n17337__;
  assign new_new_n17339__ = ~new_new_n17234__ & new_new_n17338__;
  assign new_new_n17340__ = ~new_new_n17233__ & ~new_new_n17339__;
  assign new_new_n17341__ = ~new_new_n17225__ & ~new_new_n17340__;
  assign new_new_n17342__ = ~new_new_n17224__ & ~new_new_n17341__;
  assign new_new_n17343__ = ~new_new_n17216__ & ~new_new_n17342__;
  assign new_new_n17344__ = ~new_new_n17215__ & ~new_new_n17343__;
  assign new_new_n17345__ = ~new_new_n17207__ & ~new_new_n17344__;
  assign new_new_n17346__ = ~new_new_n17206__ & ~new_new_n17345__;
  assign new_new_n17347__ = ~new_new_n17198__ & ~new_new_n17346__;
  assign new_new_n17348__ = ~new_new_n17197__ & ~new_new_n17347__;
  assign new_new_n17349__ = ~new_new_n17189__ & ~new_new_n17348__;
  assign new_new_n17350__ = ~new_new_n17188__ & ~new_new_n17349__;
  assign new_new_n17351__ = ~new_new_n17180__ & ~new_new_n17350__;
  assign new_new_n17352__ = ~new_new_n17179__ & ~new_new_n17351__;
  assign new_new_n17353__ = ~new_new_n17171__ & ~new_new_n17352__;
  assign new_new_n17354__ = ~new_new_n17170__ & ~new_new_n17353__;
  assign new_new_n17355__ = ~new_new_n17162__ & new_new_n17354__;
  assign new_new_n17356__ = ~new_new_n17161__ & ~new_new_n17355__;
  assign new_new_n17357__ = ~new_new_n17153__ & ~new_new_n17356__;
  assign new_new_n17358__ = ~new_new_n17152__ & ~new_new_n17357__;
  assign new_new_n17359__ = ~new_new_n17144__ & ~new_new_n17358__;
  assign new_new_n17360__ = ~new_new_n17143__ & ~new_new_n17359__;
  assign new_new_n17361__ = ~new_new_n17135__ & ~new_new_n17360__;
  assign new_new_n17362__ = ~new_new_n17134__ & ~new_new_n17361__;
  assign new_new_n17363__ = ~new_new_n17126__ & ~new_new_n17362__;
  assign new_new_n17364__ = ~new_new_n17125__ & ~new_new_n17363__;
  assign new_new_n17365__ = ~new_new_n17117__ & ~new_new_n17364__;
  assign new_new_n17366__ = ~new_new_n17116__ & ~new_new_n17365__;
  assign new_new_n17367__ = ~new_new_n17108__ & ~new_new_n17366__;
  assign new_new_n17368__ = ~new_new_n17107__ & ~new_new_n17367__;
  assign new_new_n17369__ = ~new_new_n17099__ & ~new_new_n17368__;
  assign new_new_n17370__ = ~new_new_n17098__ & ~new_new_n17369__;
  assign new_new_n17371__ = ~new_new_n17090__ & ~new_new_n17370__;
  assign new_new_n17372__ = ~new_new_n17089__ & ~new_new_n17371__;
  assign new_new_n17373__ = ~new_new_n17081__ & ~new_new_n17372__;
  assign new_new_n17374__ = ~new_new_n17080__ & ~new_new_n17373__;
  assign new_new_n17375__ = ~new_new_n17072__ & ~new_new_n17374__;
  assign new_new_n17376__ = ~new_new_n17071__ & ~new_new_n17375__;
  assign new_new_n17377__ = ~new_new_n17063__ & new_new_n17376__;
  assign new_new_n17378__ = ~new_new_n17062__ & ~new_new_n17377__;
  assign new_new_n17379__ = ~new_new_n17054__ & ~new_new_n17378__;
  assign new_new_n17380__ = ~new_new_n17053__ & ~new_new_n17379__;
  assign new_new_n17381__ = ~new_new_n17045__ & ~new_new_n17380__;
  assign new_new_n17382__ = ~new_new_n17044__ & ~new_new_n17381__;
  assign new_new_n17383__ = ~new_new_n17036__ & new_new_n17382__;
  assign new_new_n17384__ = ~new_new_n17035__ & ~new_new_n17383__;
  assign new_new_n17385__ = ~new_new_n17027__ & ~new_new_n17384__;
  assign new_new_n17386__ = ~new_new_n17026__ & ~new_new_n17385__;
  assign new_new_n17387__ = ~new_new_n17018__ & ~new_new_n17386__;
  assign new_new_n17388__ = ~new_new_n17017__ & ~new_new_n17387__;
  assign new_new_n17389__ = ~new_new_n17009__ & ~new_new_n17388__;
  assign new_new_n17390__ = ~new_new_n17008__ & ~new_new_n17389__;
  assign new_new_n17391__ = ~new_new_n17000__ & ~new_new_n17390__;
  assign new_new_n17392__ = ~new_new_n16999__ & ~new_new_n17391__;
  assign new_new_n17393__ = ~new_new_n16991__ & ~new_new_n17392__;
  assign new_new_n17394__ = ~new_new_n16990__ & ~new_new_n17393__;
  assign new_new_n17395__ = ~new_new_n16982__ & ~new_new_n17394__;
  assign new_new_n17396__ = ~new_new_n16981__ & ~new_new_n17395__;
  assign new_new_n17397__ = ~new_new_n16973__ & new_new_n17396__;
  assign new_new_n17398__ = ~new_new_n16972__ & ~new_new_n17397__;
  assign new_new_n17399__ = ~new_new_n16964__ & ~new_new_n17398__;
  assign new_new_n17400__ = ~new_new_n16963__ & ~new_new_n17399__;
  assign new_new_n17401__ = ~new_new_n16955__ & new_new_n17400__;
  assign new_new_n17402__ = ~new_new_n16954__ & ~new_new_n17401__;
  assign new_new_n17403__ = ~new_new_n16946__ & new_new_n17402__;
  assign new_new_n17404__ = ~new_new_n16945__ & ~new_new_n17403__;
  assign new_new_n17405__ = ~new_new_n16937__ & new_new_n17404__;
  assign new_new_n17406__ = ~new_new_n16936__ & ~new_new_n17405__;
  assign new_new_n17407__ = ~new_new_n16928__ & ~new_new_n17406__;
  assign new_new_n17408__ = ~new_new_n16927__ & ~new_new_n17407__;
  assign new_new_n17409__ = ~new_new_n16919__ & new_new_n17408__;
  assign new_new_n17410__ = ~new_new_n16918__ & ~new_new_n17409__;
  assign new_new_n17411__ = pi109 & ~new_new_n17410__;
  assign new_new_n17412__ = ~pi109 & new_new_n17410__;
  assign new_new_n17413__ = ~new_new_n16314__ & ~new_new_n16315__;
  assign new_new_n17414__ = ~new_new_n16802__ & po010;
  assign new_new_n17415__ = ~pi108 & ~po010;
  assign new_new_n17416__ = ~new_new_n17414__ & ~new_new_n17415__;
  assign new_new_n17417__ = new_new_n17413__ & ~new_new_n17416__;
  assign new_new_n17418__ = ~new_new_n17413__ & new_new_n17416__;
  assign new_new_n17419__ = ~new_new_n17417__ & ~new_new_n17418__;
  assign new_new_n17420__ = ~new_new_n17412__ & ~new_new_n17419__;
  assign new_new_n17421__ = ~new_new_n17411__ & ~new_new_n17420__;
  assign new_new_n17422__ = ~new_new_n16910__ & ~new_new_n17421__;
  assign new_new_n17423__ = ~new_new_n16909__ & ~new_new_n17422__;
  assign new_new_n17424__ = ~new_new_n16901__ & ~new_new_n17423__;
  assign new_new_n17425__ = ~new_new_n16900__ & ~new_new_n17424__;
  assign new_new_n17426__ = ~new_new_n16892__ & new_new_n17425__;
  assign new_new_n17427__ = ~new_new_n16891__ & ~new_new_n17426__;
  assign new_new_n17428__ = ~new_new_n16883__ & ~new_new_n17427__;
  assign new_new_n17429__ = ~new_new_n16882__ & ~new_new_n17428__;
  assign new_new_n17430__ = ~new_new_n16874__ & new_new_n17429__;
  assign new_new_n17431__ = ~new_new_n16873__ & ~new_new_n17430__;
  assign new_new_n17432__ = ~new_new_n16865__ & new_new_n17431__;
  assign new_new_n17433__ = ~new_new_n16864__ & ~new_new_n17432__;
  assign new_new_n17434__ = ~new_new_n16856__ & ~new_new_n17433__;
  assign new_new_n17435__ = ~new_new_n16855__ & ~new_new_n17434__;
  assign new_new_n17436__ = ~new_new_n16847__ & ~new_new_n17435__;
  assign new_new_n17437__ = ~new_new_n16846__ & ~new_new_n17436__;
  assign new_new_n17438__ = pi118 & new_new_n17437__;
  assign new_new_n17439__ = ~pi118 & ~new_new_n17437__;
  assign new_new_n17440__ = new_new_n16827__ & ~new_new_n17438__;
  assign new_new_n17441__ = ~new_new_n17439__ & new_new_n17440__;
  assign new_new_n17442__ = new_new_n16837__ & ~new_new_n17441__;
  assign new_new_n17443__ = pi118 & ~new_new_n16837__;
  assign new_new_n17444__ = new_new_n16827__ & ~new_new_n17443__;
  assign new_new_n17445__ = ~pi117 & new_new_n17435__;
  assign new_new_n17446__ = pi117 & ~new_new_n17435__;
  assign new_new_n17447__ = ~new_new_n17445__ & ~new_new_n17446__;
  assign new_new_n17448__ = new_new_n17444__ & ~new_new_n17447__;
  assign new_new_n17449__ = ~new_new_n16845__ & ~new_new_n17448__;
  assign new_new_n17450__ = ~pi118 & new_new_n16837__;
  assign new_new_n17451__ = new_new_n16827__ & new_new_n16845__;
  assign new_new_n17452__ = new_new_n17450__ & new_new_n17451__;
  assign new_new_n17453__ = ~new_new_n17447__ & new_new_n17452__;
  assign new_new_n17454__ = ~new_new_n17449__ & ~new_new_n17453__;
  assign new_new_n17455__ = pi118 & new_new_n17454__;
  assign new_new_n17456__ = ~pi118 & ~new_new_n17454__;
  assign new_new_n17457__ = ~new_new_n17455__ & ~new_new_n17456__;
  assign new_new_n17458__ = ~new_new_n16855__ & ~new_new_n16856__;
  assign new_new_n17459__ = new_new_n17437__ & ~new_new_n17450__;
  assign po009 = new_new_n17444__ & ~new_new_n17459__;
  assign new_new_n17461__ = ~new_new_n17433__ & po009;
  assign new_new_n17462__ = ~pi116 & ~po009;
  assign new_new_n17463__ = ~new_new_n17461__ & ~new_new_n17462__;
  assign new_new_n17464__ = new_new_n17458__ & ~new_new_n17463__;
  assign new_new_n17465__ = ~new_new_n17458__ & new_new_n17463__;
  assign new_new_n17466__ = ~new_new_n17464__ & ~new_new_n17465__;
  assign new_new_n17467__ = ~pi117 & new_new_n17466__;
  assign new_new_n17468__ = pi117 & ~new_new_n17466__;
  assign new_new_n17469__ = ~new_new_n17431__ & po009;
  assign new_new_n17470__ = pi115 & ~po009;
  assign new_new_n17471__ = ~new_new_n17469__ & ~new_new_n17470__;
  assign new_new_n17472__ = ~new_new_n16864__ & ~new_new_n16865__;
  assign new_new_n17473__ = ~new_new_n17471__ & new_new_n17472__;
  assign new_new_n17474__ = new_new_n17471__ & ~new_new_n17472__;
  assign new_new_n17475__ = ~new_new_n17473__ & ~new_new_n17474__;
  assign new_new_n17476__ = ~pi116 & ~new_new_n17475__;
  assign new_new_n17477__ = pi116 & new_new_n17475__;
  assign new_new_n17478__ = ~new_new_n16873__ & ~new_new_n16874__;
  assign new_new_n17479__ = ~new_new_n17429__ & po009;
  assign new_new_n17480__ = ~pi114 & ~po009;
  assign new_new_n17481__ = ~new_new_n17479__ & ~new_new_n17480__;
  assign new_new_n17482__ = new_new_n17478__ & ~new_new_n17481__;
  assign new_new_n17483__ = ~new_new_n17478__ & new_new_n17481__;
  assign new_new_n17484__ = ~new_new_n17482__ & ~new_new_n17483__;
  assign new_new_n17485__ = pi115 & ~new_new_n17484__;
  assign new_new_n17486__ = ~pi115 & new_new_n17484__;
  assign new_new_n17487__ = ~new_new_n16882__ & ~new_new_n16883__;
  assign new_new_n17488__ = ~new_new_n17427__ & po009;
  assign new_new_n17489__ = ~pi113 & ~po009;
  assign new_new_n17490__ = ~new_new_n17488__ & ~new_new_n17489__;
  assign new_new_n17491__ = new_new_n17487__ & ~new_new_n17490__;
  assign new_new_n17492__ = ~new_new_n17487__ & new_new_n17490__;
  assign new_new_n17493__ = ~new_new_n17491__ & ~new_new_n17492__;
  assign new_new_n17494__ = pi114 & ~new_new_n17493__;
  assign new_new_n17495__ = ~pi114 & new_new_n17493__;
  assign new_new_n17496__ = ~new_new_n17425__ & po009;
  assign new_new_n17497__ = pi112 & ~po009;
  assign new_new_n17498__ = ~new_new_n17496__ & ~new_new_n17497__;
  assign new_new_n17499__ = ~new_new_n16891__ & ~new_new_n16892__;
  assign new_new_n17500__ = ~new_new_n17498__ & new_new_n17499__;
  assign new_new_n17501__ = new_new_n17498__ & ~new_new_n17499__;
  assign new_new_n17502__ = ~new_new_n17500__ & ~new_new_n17501__;
  assign new_new_n17503__ = ~pi113 & ~new_new_n17502__;
  assign new_new_n17504__ = pi113 & new_new_n17502__;
  assign new_new_n17505__ = ~new_new_n16900__ & ~new_new_n16901__;
  assign new_new_n17506__ = ~new_new_n17423__ & po009;
  assign new_new_n17507__ = pi111 & ~po009;
  assign new_new_n17508__ = ~new_new_n17506__ & ~new_new_n17507__;
  assign new_new_n17509__ = new_new_n17505__ & ~new_new_n17508__;
  assign new_new_n17510__ = ~new_new_n17505__ & new_new_n17508__;
  assign new_new_n17511__ = ~new_new_n17509__ & ~new_new_n17510__;
  assign new_new_n17512__ = pi112 & new_new_n17511__;
  assign new_new_n17513__ = ~pi112 & ~new_new_n17511__;
  assign new_new_n17514__ = pi110 & ~new_new_n17421__;
  assign new_new_n17515__ = ~pi110 & new_new_n17421__;
  assign new_new_n17516__ = ~new_new_n17514__ & ~new_new_n17515__;
  assign new_new_n17517__ = po009 & new_new_n17516__;
  assign new_new_n17518__ = new_new_n16908__ & new_new_n17517__;
  assign new_new_n17519__ = ~new_new_n16908__ & ~new_new_n17517__;
  assign new_new_n17520__ = ~new_new_n17518__ & ~new_new_n17519__;
  assign new_new_n17521__ = pi111 & ~new_new_n17520__;
  assign new_new_n17522__ = ~pi111 & new_new_n17520__;
  assign new_new_n17523__ = ~new_new_n17411__ & ~new_new_n17412__;
  assign new_new_n17524__ = po009 & new_new_n17523__;
  assign new_new_n17525__ = new_new_n17419__ & new_new_n17524__;
  assign new_new_n17526__ = ~new_new_n17419__ & ~new_new_n17524__;
  assign new_new_n17527__ = ~new_new_n17525__ & ~new_new_n17526__;
  assign new_new_n17528__ = pi110 & ~new_new_n17527__;
  assign new_new_n17529__ = ~pi110 & new_new_n17527__;
  assign new_new_n17530__ = ~new_new_n16918__ & ~new_new_n16919__;
  assign new_new_n17531__ = ~new_new_n17408__ & po009;
  assign new_new_n17532__ = ~pi108 & ~po009;
  assign new_new_n17533__ = ~new_new_n17531__ & ~new_new_n17532__;
  assign new_new_n17534__ = new_new_n17530__ & ~new_new_n17533__;
  assign new_new_n17535__ = ~new_new_n17530__ & new_new_n17533__;
  assign new_new_n17536__ = ~new_new_n17534__ & ~new_new_n17535__;
  assign new_new_n17537__ = pi109 & ~new_new_n17536__;
  assign new_new_n17538__ = ~pi109 & new_new_n17536__;
  assign new_new_n17539__ = ~new_new_n16927__ & ~new_new_n16928__;
  assign new_new_n17540__ = ~new_new_n17406__ & po009;
  assign new_new_n17541__ = ~pi107 & ~po009;
  assign new_new_n17542__ = ~new_new_n17540__ & ~new_new_n17541__;
  assign new_new_n17543__ = ~new_new_n17539__ & ~new_new_n17542__;
  assign new_new_n17544__ = new_new_n17539__ & new_new_n17542__;
  assign new_new_n17545__ = ~new_new_n17543__ & ~new_new_n17544__;
  assign new_new_n17546__ = ~pi108 & ~new_new_n17545__;
  assign new_new_n17547__ = pi108 & new_new_n17545__;
  assign new_new_n17548__ = new_new_n17404__ & po009;
  assign new_new_n17549__ = ~pi106 & ~po009;
  assign new_new_n17550__ = ~new_new_n17548__ & ~new_new_n17549__;
  assign new_new_n17551__ = ~new_new_n16936__ & ~new_new_n16937__;
  assign new_new_n17552__ = ~new_new_n17550__ & ~new_new_n17551__;
  assign new_new_n17553__ = new_new_n17550__ & new_new_n17551__;
  assign new_new_n17554__ = ~new_new_n17552__ & ~new_new_n17553__;
  assign new_new_n17555__ = ~pi107 & ~new_new_n17554__;
  assign new_new_n17556__ = pi107 & new_new_n17554__;
  assign new_new_n17557__ = ~new_new_n16945__ & ~new_new_n16946__;
  assign new_new_n17558__ = ~new_new_n17402__ & po009;
  assign new_new_n17559__ = ~pi105 & ~po009;
  assign new_new_n17560__ = ~new_new_n17558__ & ~new_new_n17559__;
  assign new_new_n17561__ = new_new_n17557__ & ~new_new_n17560__;
  assign new_new_n17562__ = ~new_new_n17557__ & new_new_n17560__;
  assign new_new_n17563__ = ~new_new_n17561__ & ~new_new_n17562__;
  assign new_new_n17564__ = ~pi106 & new_new_n17563__;
  assign new_new_n17565__ = pi106 & ~new_new_n17563__;
  assign new_new_n17566__ = ~new_new_n17400__ & po009;
  assign new_new_n17567__ = pi104 & ~po009;
  assign new_new_n17568__ = ~new_new_n17566__ & ~new_new_n17567__;
  assign new_new_n17569__ = ~new_new_n16954__ & ~new_new_n16955__;
  assign new_new_n17570__ = ~new_new_n17568__ & new_new_n17569__;
  assign new_new_n17571__ = new_new_n17568__ & ~new_new_n17569__;
  assign new_new_n17572__ = ~new_new_n17570__ & ~new_new_n17571__;
  assign new_new_n17573__ = ~pi105 & ~new_new_n17572__;
  assign new_new_n17574__ = pi105 & new_new_n17572__;
  assign new_new_n17575__ = ~new_new_n16963__ & ~new_new_n16964__;
  assign new_new_n17576__ = ~new_new_n17398__ & po009;
  assign new_new_n17577__ = pi103 & ~po009;
  assign new_new_n17578__ = ~new_new_n17576__ & ~new_new_n17577__;
  assign new_new_n17579__ = new_new_n17575__ & new_new_n17578__;
  assign new_new_n17580__ = ~new_new_n17575__ & ~new_new_n17578__;
  assign new_new_n17581__ = ~new_new_n17579__ & ~new_new_n17580__;
  assign new_new_n17582__ = ~pi104 & new_new_n17581__;
  assign new_new_n17583__ = pi104 & ~new_new_n17581__;
  assign new_new_n17584__ = new_new_n17396__ & po009;
  assign new_new_n17585__ = pi102 & ~po009;
  assign new_new_n17586__ = ~new_new_n17584__ & ~new_new_n17585__;
  assign new_new_n17587__ = ~new_new_n16972__ & ~new_new_n16973__;
  assign new_new_n17588__ = ~new_new_n17586__ & ~new_new_n17587__;
  assign new_new_n17589__ = new_new_n17586__ & new_new_n17587__;
  assign new_new_n17590__ = ~new_new_n17588__ & ~new_new_n17589__;
  assign new_new_n17591__ = ~pi103 & new_new_n17590__;
  assign new_new_n17592__ = pi103 & ~new_new_n17590__;
  assign new_new_n17593__ = ~pi101 & ~new_new_n17394__;
  assign new_new_n17594__ = pi101 & new_new_n17394__;
  assign new_new_n17595__ = ~new_new_n17593__ & ~new_new_n17594__;
  assign new_new_n17596__ = po009 & new_new_n17595__;
  assign new_new_n17597__ = new_new_n16980__ & new_new_n17596__;
  assign new_new_n17598__ = ~new_new_n16980__ & ~new_new_n17596__;
  assign new_new_n17599__ = ~new_new_n17597__ & ~new_new_n17598__;
  assign new_new_n17600__ = ~pi102 & ~new_new_n17599__;
  assign new_new_n17601__ = pi102 & new_new_n17599__;
  assign new_new_n17602__ = ~new_new_n16990__ & ~new_new_n16991__;
  assign new_new_n17603__ = ~new_new_n17392__ & po009;
  assign new_new_n17604__ = ~pi100 & ~po009;
  assign new_new_n17605__ = ~new_new_n17603__ & ~new_new_n17604__;
  assign new_new_n17606__ = new_new_n17602__ & ~new_new_n17605__;
  assign new_new_n17607__ = ~new_new_n17602__ & new_new_n17605__;
  assign new_new_n17608__ = ~new_new_n17606__ & ~new_new_n17607__;
  assign new_new_n17609__ = pi101 & ~new_new_n17608__;
  assign new_new_n17610__ = ~pi101 & new_new_n17608__;
  assign new_new_n17611__ = ~new_new_n16999__ & ~new_new_n17000__;
  assign new_new_n17612__ = ~new_new_n17390__ & po009;
  assign new_new_n17613__ = ~pi099 & ~po009;
  assign new_new_n17614__ = ~new_new_n17612__ & ~new_new_n17613__;
  assign new_new_n17615__ = new_new_n17611__ & ~new_new_n17614__;
  assign new_new_n17616__ = ~new_new_n17611__ & new_new_n17614__;
  assign new_new_n17617__ = ~new_new_n17615__ & ~new_new_n17616__;
  assign new_new_n17618__ = pi100 & ~new_new_n17617__;
  assign new_new_n17619__ = ~pi100 & new_new_n17617__;
  assign new_new_n17620__ = ~pi098 & ~new_new_n17388__;
  assign new_new_n17621__ = pi098 & new_new_n17388__;
  assign new_new_n17622__ = ~new_new_n17620__ & ~new_new_n17621__;
  assign new_new_n17623__ = po009 & new_new_n17622__;
  assign new_new_n17624__ = ~new_new_n17007__ & ~new_new_n17623__;
  assign new_new_n17625__ = new_new_n17007__ & new_new_n17623__;
  assign new_new_n17626__ = ~new_new_n17624__ & ~new_new_n17625__;
  assign new_new_n17627__ = ~pi099 & ~new_new_n17626__;
  assign new_new_n17628__ = pi099 & new_new_n17626__;
  assign new_new_n17629__ = ~pi097 & ~new_new_n17386__;
  assign new_new_n17630__ = pi097 & new_new_n17386__;
  assign new_new_n17631__ = ~new_new_n17629__ & ~new_new_n17630__;
  assign new_new_n17632__ = po009 & new_new_n17631__;
  assign new_new_n17633__ = new_new_n17016__ & new_new_n17632__;
  assign new_new_n17634__ = ~new_new_n17016__ & ~new_new_n17632__;
  assign new_new_n17635__ = ~new_new_n17633__ & ~new_new_n17634__;
  assign new_new_n17636__ = ~pi098 & ~new_new_n17635__;
  assign new_new_n17637__ = pi098 & new_new_n17635__;
  assign new_new_n17638__ = ~new_new_n17026__ & ~new_new_n17027__;
  assign new_new_n17639__ = ~new_new_n17384__ & po009;
  assign new_new_n17640__ = ~pi096 & ~po009;
  assign new_new_n17641__ = ~new_new_n17639__ & ~new_new_n17640__;
  assign new_new_n17642__ = new_new_n17638__ & ~new_new_n17641__;
  assign new_new_n17643__ = ~new_new_n17638__ & new_new_n17641__;
  assign new_new_n17644__ = ~new_new_n17642__ & ~new_new_n17643__;
  assign new_new_n17645__ = pi097 & ~new_new_n17644__;
  assign new_new_n17646__ = ~pi097 & new_new_n17644__;
  assign new_new_n17647__ = ~new_new_n17382__ & po009;
  assign new_new_n17648__ = pi095 & ~po009;
  assign new_new_n17649__ = ~new_new_n17647__ & ~new_new_n17648__;
  assign new_new_n17650__ = ~new_new_n17035__ & ~new_new_n17036__;
  assign new_new_n17651__ = ~new_new_n17649__ & new_new_n17650__;
  assign new_new_n17652__ = new_new_n17649__ & ~new_new_n17650__;
  assign new_new_n17653__ = ~new_new_n17651__ & ~new_new_n17652__;
  assign new_new_n17654__ = ~pi096 & ~new_new_n17653__;
  assign new_new_n17655__ = pi096 & new_new_n17653__;
  assign new_new_n17656__ = ~new_new_n17044__ & ~new_new_n17045__;
  assign new_new_n17657__ = new_new_n17380__ & po009;
  assign new_new_n17658__ = ~pi094 & ~po009;
  assign new_new_n17659__ = ~new_new_n17657__ & ~new_new_n17658__;
  assign new_new_n17660__ = ~new_new_n17656__ & ~new_new_n17659__;
  assign new_new_n17661__ = new_new_n17656__ & new_new_n17659__;
  assign new_new_n17662__ = ~new_new_n17660__ & ~new_new_n17661__;
  assign new_new_n17663__ = ~pi095 & ~new_new_n17662__;
  assign new_new_n17664__ = pi095 & new_new_n17662__;
  assign new_new_n17665__ = pi093 & ~new_new_n17378__;
  assign new_new_n17666__ = ~pi093 & new_new_n17378__;
  assign new_new_n17667__ = ~new_new_n17665__ & ~new_new_n17666__;
  assign new_new_n17668__ = po009 & new_new_n17667__;
  assign new_new_n17669__ = new_new_n17052__ & new_new_n17668__;
  assign new_new_n17670__ = ~new_new_n17052__ & ~new_new_n17668__;
  assign new_new_n17671__ = ~new_new_n17669__ & ~new_new_n17670__;
  assign new_new_n17672__ = pi094 & ~new_new_n17671__;
  assign new_new_n17673__ = ~pi094 & new_new_n17671__;
  assign new_new_n17674__ = ~new_new_n17062__ & ~new_new_n17063__;
  assign new_new_n17675__ = ~new_new_n17376__ & po009;
  assign new_new_n17676__ = ~pi092 & ~po009;
  assign new_new_n17677__ = ~new_new_n17675__ & ~new_new_n17676__;
  assign new_new_n17678__ = new_new_n17674__ & ~new_new_n17677__;
  assign new_new_n17679__ = ~new_new_n17674__ & new_new_n17677__;
  assign new_new_n17680__ = ~new_new_n17678__ & ~new_new_n17679__;
  assign new_new_n17681__ = pi093 & ~new_new_n17680__;
  assign new_new_n17682__ = ~pi093 & new_new_n17680__;
  assign new_new_n17683__ = ~new_new_n17071__ & ~new_new_n17072__;
  assign new_new_n17684__ = ~new_new_n17374__ & po009;
  assign new_new_n17685__ = ~pi091 & ~po009;
  assign new_new_n17686__ = ~new_new_n17684__ & ~new_new_n17685__;
  assign new_new_n17687__ = new_new_n17683__ & ~new_new_n17686__;
  assign new_new_n17688__ = ~new_new_n17683__ & new_new_n17686__;
  assign new_new_n17689__ = ~new_new_n17687__ & ~new_new_n17688__;
  assign new_new_n17690__ = pi092 & ~new_new_n17689__;
  assign new_new_n17691__ = ~pi092 & new_new_n17689__;
  assign new_new_n17692__ = ~new_new_n17080__ & ~new_new_n17081__;
  assign new_new_n17693__ = ~new_new_n17372__ & po009;
  assign new_new_n17694__ = ~pi090 & ~po009;
  assign new_new_n17695__ = ~new_new_n17693__ & ~new_new_n17694__;
  assign new_new_n17696__ = new_new_n17692__ & ~new_new_n17695__;
  assign new_new_n17697__ = ~new_new_n17692__ & new_new_n17695__;
  assign new_new_n17698__ = ~new_new_n17696__ & ~new_new_n17697__;
  assign new_new_n17699__ = ~pi091 & new_new_n17698__;
  assign new_new_n17700__ = pi091 & ~new_new_n17698__;
  assign new_new_n17701__ = ~new_new_n17089__ & ~new_new_n17090__;
  assign new_new_n17702__ = ~new_new_n17370__ & po009;
  assign new_new_n17703__ = ~pi089 & ~po009;
  assign new_new_n17704__ = ~new_new_n17702__ & ~new_new_n17703__;
  assign new_new_n17705__ = ~new_new_n17701__ & ~new_new_n17704__;
  assign new_new_n17706__ = new_new_n17701__ & new_new_n17704__;
  assign new_new_n17707__ = ~new_new_n17705__ & ~new_new_n17706__;
  assign new_new_n17708__ = ~pi090 & ~new_new_n17707__;
  assign new_new_n17709__ = pi090 & new_new_n17707__;
  assign new_new_n17710__ = new_new_n17368__ & po009;
  assign new_new_n17711__ = pi088 & ~po009;
  assign new_new_n17712__ = ~new_new_n17710__ & ~new_new_n17711__;
  assign new_new_n17713__ = ~new_new_n17098__ & ~new_new_n17099__;
  assign new_new_n17714__ = ~new_new_n17712__ & ~new_new_n17713__;
  assign new_new_n17715__ = new_new_n17712__ & new_new_n17713__;
  assign new_new_n17716__ = ~new_new_n17714__ & ~new_new_n17715__;
  assign new_new_n17717__ = pi089 & ~new_new_n17716__;
  assign new_new_n17718__ = ~pi089 & new_new_n17716__;
  assign new_new_n17719__ = new_new_n17366__ & po009;
  assign new_new_n17720__ = pi087 & ~po009;
  assign new_new_n17721__ = ~new_new_n17719__ & ~new_new_n17720__;
  assign new_new_n17722__ = ~new_new_n17107__ & ~new_new_n17108__;
  assign new_new_n17723__ = ~new_new_n17721__ & ~new_new_n17722__;
  assign new_new_n17724__ = new_new_n17721__ & new_new_n17722__;
  assign new_new_n17725__ = ~new_new_n17723__ & ~new_new_n17724__;
  assign new_new_n17726__ = pi088 & ~new_new_n17725__;
  assign new_new_n17727__ = ~pi088 & new_new_n17725__;
  assign new_new_n17728__ = ~new_new_n17116__ & ~new_new_n17117__;
  assign new_new_n17729__ = ~new_new_n17364__ & po009;
  assign new_new_n17730__ = ~pi086 & ~po009;
  assign new_new_n17731__ = ~new_new_n17729__ & ~new_new_n17730__;
  assign new_new_n17732__ = new_new_n17728__ & ~new_new_n17731__;
  assign new_new_n17733__ = ~new_new_n17728__ & new_new_n17731__;
  assign new_new_n17734__ = ~new_new_n17732__ & ~new_new_n17733__;
  assign new_new_n17735__ = pi087 & ~new_new_n17734__;
  assign new_new_n17736__ = ~pi087 & new_new_n17734__;
  assign new_new_n17737__ = ~new_new_n17125__ & ~new_new_n17126__;
  assign new_new_n17738__ = ~new_new_n17362__ & po009;
  assign new_new_n17739__ = ~pi085 & ~po009;
  assign new_new_n17740__ = ~new_new_n17738__ & ~new_new_n17739__;
  assign new_new_n17741__ = new_new_n17737__ & ~new_new_n17740__;
  assign new_new_n17742__ = ~new_new_n17737__ & new_new_n17740__;
  assign new_new_n17743__ = ~new_new_n17741__ & ~new_new_n17742__;
  assign new_new_n17744__ = ~pi086 & new_new_n17743__;
  assign new_new_n17745__ = pi086 & ~new_new_n17743__;
  assign new_new_n17746__ = ~pi084 & ~new_new_n17360__;
  assign new_new_n17747__ = pi084 & new_new_n17360__;
  assign new_new_n17748__ = ~new_new_n17746__ & ~new_new_n17747__;
  assign new_new_n17749__ = po009 & new_new_n17748__;
  assign new_new_n17750__ = new_new_n17133__ & new_new_n17749__;
  assign new_new_n17751__ = ~new_new_n17133__ & ~new_new_n17749__;
  assign new_new_n17752__ = ~new_new_n17750__ & ~new_new_n17751__;
  assign new_new_n17753__ = ~pi085 & ~new_new_n17752__;
  assign new_new_n17754__ = pi085 & new_new_n17752__;
  assign new_new_n17755__ = ~new_new_n17143__ & ~new_new_n17144__;
  assign new_new_n17756__ = ~new_new_n17358__ & po009;
  assign new_new_n17757__ = ~pi083 & ~po009;
  assign new_new_n17758__ = ~new_new_n17756__ & ~new_new_n17757__;
  assign new_new_n17759__ = new_new_n17755__ & ~new_new_n17758__;
  assign new_new_n17760__ = ~new_new_n17755__ & new_new_n17758__;
  assign new_new_n17761__ = ~new_new_n17759__ & ~new_new_n17760__;
  assign new_new_n17762__ = pi084 & ~new_new_n17761__;
  assign new_new_n17763__ = ~pi084 & new_new_n17761__;
  assign new_new_n17764__ = ~pi082 & ~new_new_n17356__;
  assign new_new_n17765__ = pi082 & new_new_n17356__;
  assign new_new_n17766__ = ~new_new_n17764__ & ~new_new_n17765__;
  assign new_new_n17767__ = po009 & new_new_n17766__;
  assign new_new_n17768__ = new_new_n17151__ & new_new_n17767__;
  assign new_new_n17769__ = ~new_new_n17151__ & ~new_new_n17767__;
  assign new_new_n17770__ = ~new_new_n17768__ & ~new_new_n17769__;
  assign new_new_n17771__ = ~pi083 & ~new_new_n17770__;
  assign new_new_n17772__ = pi083 & new_new_n17770__;
  assign new_new_n17773__ = ~new_new_n17161__ & ~new_new_n17162__;
  assign new_new_n17774__ = ~new_new_n17354__ & po009;
  assign new_new_n17775__ = pi081 & ~po009;
  assign new_new_n17776__ = ~new_new_n17774__ & ~new_new_n17775__;
  assign new_new_n17777__ = new_new_n17773__ & ~new_new_n17776__;
  assign new_new_n17778__ = ~new_new_n17773__ & new_new_n17776__;
  assign new_new_n17779__ = ~new_new_n17777__ & ~new_new_n17778__;
  assign new_new_n17780__ = ~pi082 & ~new_new_n17779__;
  assign new_new_n17781__ = pi082 & new_new_n17779__;
  assign new_new_n17782__ = new_new_n17352__ & po009;
  assign new_new_n17783__ = ~pi080 & ~po009;
  assign new_new_n17784__ = ~new_new_n17782__ & ~new_new_n17783__;
  assign new_new_n17785__ = ~new_new_n17170__ & ~new_new_n17171__;
  assign new_new_n17786__ = ~new_new_n17784__ & ~new_new_n17785__;
  assign new_new_n17787__ = new_new_n17784__ & new_new_n17785__;
  assign new_new_n17788__ = ~new_new_n17786__ & ~new_new_n17787__;
  assign new_new_n17789__ = pi081 & new_new_n17788__;
  assign new_new_n17790__ = ~pi081 & ~new_new_n17788__;
  assign new_new_n17791__ = ~new_new_n17179__ & ~new_new_n17180__;
  assign new_new_n17792__ = ~new_new_n17350__ & po009;
  assign new_new_n17793__ = pi079 & ~po009;
  assign new_new_n17794__ = ~new_new_n17792__ & ~new_new_n17793__;
  assign new_new_n17795__ = new_new_n17791__ & new_new_n17794__;
  assign new_new_n17796__ = ~new_new_n17791__ & ~new_new_n17794__;
  assign new_new_n17797__ = ~new_new_n17795__ & ~new_new_n17796__;
  assign new_new_n17798__ = pi080 & ~new_new_n17797__;
  assign new_new_n17799__ = ~pi080 & new_new_n17797__;
  assign new_new_n17800__ = new_new_n17348__ & po009;
  assign new_new_n17801__ = ~pi078 & ~po009;
  assign new_new_n17802__ = ~new_new_n17800__ & ~new_new_n17801__;
  assign new_new_n17803__ = ~new_new_n17188__ & ~new_new_n17189__;
  assign new_new_n17804__ = ~new_new_n17802__ & ~new_new_n17803__;
  assign new_new_n17805__ = new_new_n17802__ & new_new_n17803__;
  assign new_new_n17806__ = ~new_new_n17804__ & ~new_new_n17805__;
  assign new_new_n17807__ = ~pi079 & ~new_new_n17806__;
  assign new_new_n17808__ = pi079 & new_new_n17806__;
  assign new_new_n17809__ = ~new_new_n17346__ & po009;
  assign new_new_n17810__ = pi077 & ~po009;
  assign new_new_n17811__ = ~new_new_n17809__ & ~new_new_n17810__;
  assign new_new_n17812__ = ~new_new_n17197__ & ~new_new_n17198__;
  assign new_new_n17813__ = ~new_new_n17811__ & new_new_n17812__;
  assign new_new_n17814__ = new_new_n17811__ & ~new_new_n17812__;
  assign new_new_n17815__ = ~new_new_n17813__ & ~new_new_n17814__;
  assign new_new_n17816__ = ~pi078 & ~new_new_n17815__;
  assign new_new_n17817__ = pi078 & new_new_n17815__;
  assign new_new_n17818__ = ~new_new_n17344__ & po009;
  assign new_new_n17819__ = pi076 & ~po009;
  assign new_new_n17820__ = ~new_new_n17818__ & ~new_new_n17819__;
  assign new_new_n17821__ = ~new_new_n17206__ & ~new_new_n17207__;
  assign new_new_n17822__ = ~new_new_n17820__ & new_new_n17821__;
  assign new_new_n17823__ = new_new_n17820__ & ~new_new_n17821__;
  assign new_new_n17824__ = ~new_new_n17822__ & ~new_new_n17823__;
  assign new_new_n17825__ = ~pi077 & ~new_new_n17824__;
  assign new_new_n17826__ = pi077 & new_new_n17824__;
  assign new_new_n17827__ = ~new_new_n17342__ & po009;
  assign new_new_n17828__ = pi075 & ~po009;
  assign new_new_n17829__ = ~new_new_n17827__ & ~new_new_n17828__;
  assign new_new_n17830__ = ~new_new_n17215__ & ~new_new_n17216__;
  assign new_new_n17831__ = ~new_new_n17829__ & new_new_n17830__;
  assign new_new_n17832__ = new_new_n17829__ & ~new_new_n17830__;
  assign new_new_n17833__ = ~new_new_n17831__ & ~new_new_n17832__;
  assign new_new_n17834__ = ~pi076 & ~new_new_n17833__;
  assign new_new_n17835__ = pi076 & new_new_n17833__;
  assign new_new_n17836__ = pi074 & ~new_new_n17340__;
  assign new_new_n17837__ = ~pi074 & new_new_n17340__;
  assign new_new_n17838__ = ~new_new_n17836__ & ~new_new_n17837__;
  assign new_new_n17839__ = po009 & new_new_n17838__;
  assign new_new_n17840__ = ~new_new_n17223__ & ~new_new_n17839__;
  assign new_new_n17841__ = new_new_n17223__ & new_new_n17839__;
  assign new_new_n17842__ = ~new_new_n17840__ & ~new_new_n17841__;
  assign new_new_n17843__ = ~pi075 & new_new_n17842__;
  assign new_new_n17844__ = pi075 & ~new_new_n17842__;
  assign new_new_n17845__ = ~new_new_n17233__ & ~new_new_n17234__;
  assign new_new_n17846__ = ~new_new_n17338__ & po009;
  assign new_new_n17847__ = ~pi073 & ~po009;
  assign new_new_n17848__ = ~new_new_n17846__ & ~new_new_n17847__;
  assign new_new_n17849__ = new_new_n17845__ & new_new_n17848__;
  assign new_new_n17850__ = ~new_new_n17845__ & ~new_new_n17848__;
  assign new_new_n17851__ = ~new_new_n17849__ & ~new_new_n17850__;
  assign new_new_n17852__ = ~pi074 & ~new_new_n17851__;
  assign new_new_n17853__ = pi074 & new_new_n17851__;
  assign new_new_n17854__ = new_new_n17336__ & po009;
  assign new_new_n17855__ = ~pi072 & ~po009;
  assign new_new_n17856__ = ~new_new_n17854__ & ~new_new_n17855__;
  assign new_new_n17857__ = ~new_new_n17242__ & ~new_new_n17243__;
  assign new_new_n17858__ = ~new_new_n17856__ & ~new_new_n17857__;
  assign new_new_n17859__ = new_new_n17856__ & new_new_n17857__;
  assign new_new_n17860__ = ~new_new_n17858__ & ~new_new_n17859__;
  assign new_new_n17861__ = pi073 & new_new_n17860__;
  assign new_new_n17862__ = ~pi073 & ~new_new_n17860__;
  assign new_new_n17863__ = pi071 & ~new_new_n17334__;
  assign new_new_n17864__ = ~pi071 & new_new_n17334__;
  assign new_new_n17865__ = ~new_new_n17863__ & ~new_new_n17864__;
  assign new_new_n17866__ = po009 & new_new_n17865__;
  assign new_new_n17867__ = new_new_n17250__ & new_new_n17866__;
  assign new_new_n17868__ = ~new_new_n17250__ & ~new_new_n17866__;
  assign new_new_n17869__ = ~new_new_n17867__ & ~new_new_n17868__;
  assign new_new_n17870__ = pi072 & ~new_new_n17869__;
  assign new_new_n17871__ = ~pi072 & new_new_n17869__;
  assign new_new_n17872__ = ~new_new_n17332__ & po009;
  assign new_new_n17873__ = pi070 & ~po009;
  assign new_new_n17874__ = ~new_new_n17872__ & ~new_new_n17873__;
  assign new_new_n17875__ = ~new_new_n17260__ & ~new_new_n17261__;
  assign new_new_n17876__ = ~new_new_n17874__ & new_new_n17875__;
  assign new_new_n17877__ = new_new_n17874__ & ~new_new_n17875__;
  assign new_new_n17878__ = ~new_new_n17876__ & ~new_new_n17877__;
  assign new_new_n17879__ = ~pi071 & ~new_new_n17878__;
  assign new_new_n17880__ = pi071 & new_new_n17878__;
  assign new_new_n17881__ = ~new_new_n17324__ & ~new_new_n17325__;
  assign new_new_n17882__ = po009 & new_new_n17881__;
  assign new_new_n17883__ = new_new_n17330__ & new_new_n17882__;
  assign new_new_n17884__ = ~new_new_n17330__ & ~new_new_n17882__;
  assign new_new_n17885__ = ~new_new_n17883__ & ~new_new_n17884__;
  assign new_new_n17886__ = ~pi070 & ~new_new_n17885__;
  assign new_new_n17887__ = pi070 & new_new_n17885__;
  assign new_new_n17888__ = new_new_n17321__ & po009;
  assign new_new_n17889__ = pi068 & ~po009;
  assign new_new_n17890__ = ~new_new_n17888__ & ~new_new_n17889__;
  assign new_new_n17891__ = ~new_new_n17269__ & ~new_new_n17270__;
  assign new_new_n17892__ = ~new_new_n17890__ & ~new_new_n17891__;
  assign new_new_n17893__ = new_new_n17890__ & new_new_n17891__;
  assign new_new_n17894__ = ~new_new_n17892__ & ~new_new_n17893__;
  assign new_new_n17895__ = ~pi069 & new_new_n17894__;
  assign new_new_n17896__ = pi069 & ~new_new_n17894__;
  assign new_new_n17897__ = ~new_new_n16673__ & ~new_new_n17291__;
  assign new_new_n17898__ = ~new_new_n16697__ & ~new_new_n16702__;
  assign new_new_n17899__ = ~new_new_n403__ & new_new_n17898__;
  assign new_new_n17900__ = new_new_n17289__ & new_new_n17899__;
  assign new_new_n17901__ = pi010 & ~new_new_n17898__;
  assign new_new_n17902__ = ~new_new_n17298__ & new_new_n17901__;
  assign new_new_n17903__ = ~new_new_n17897__ & ~new_new_n17900__;
  assign new_new_n17904__ = ~new_new_n17902__ & new_new_n17903__;
  assign new_new_n17905__ = pi011 & ~new_new_n17904__;
  assign new_new_n17906__ = ~new_new_n16673__ & ~new_new_n17286__;
  assign new_new_n17907__ = pi010 & ~new_new_n16702__;
  assign new_new_n17908__ = pi064 & ~new_new_n17907__;
  assign new_new_n17909__ = ~new_new_n17906__ & ~new_new_n17908__;
  assign new_new_n17910__ = ~pi065 & po010;
  assign new_new_n17911__ = po011 & new_new_n17910__;
  assign new_new_n17912__ = ~po011 & ~new_new_n17910__;
  assign new_new_n17913__ = pi064 & ~new_new_n17306__;
  assign new_new_n17914__ = ~new_new_n17911__ & new_new_n17913__;
  assign new_new_n17915__ = ~new_new_n17912__ & new_new_n17914__;
  assign new_new_n17916__ = ~new_new_n17909__ & ~new_new_n17915__;
  assign new_new_n17917__ = ~pi011 & ~new_new_n17916__;
  assign new_new_n17918__ = ~new_new_n17905__ & ~new_new_n17917__;
  assign new_new_n17919__ = ~pi009 & ~new_new_n17305__;
  assign new_new_n17920__ = ~new_new_n17311__ & ~new_new_n17919__;
  assign new_new_n17921__ = pi064 & ~new_new_n17920__;
  assign new_new_n17922__ = ~new_new_n17299__ & ~new_new_n17921__;
  assign new_new_n17923__ = ~pi066 & ~new_new_n17922__;
  assign new_new_n17924__ = pi066 & new_new_n17922__;
  assign new_new_n17925__ = ~new_new_n17923__ & ~new_new_n17924__;
  assign new_new_n17926__ = po009 & ~new_new_n17925__;
  assign new_new_n17927__ = ~new_new_n17918__ & new_new_n17926__;
  assign new_new_n17928__ = new_new_n17918__ & ~new_new_n17926__;
  assign new_new_n17929__ = ~new_new_n17927__ & ~new_new_n17928__;
  assign new_new_n17930__ = pi067 & ~new_new_n17929__;
  assign new_new_n17931__ = pi009 & po009;
  assign new_new_n17932__ = pi008 & ~pi065;
  assign new_new_n17933__ = new_new_n17931__ & ~new_new_n17932__;
  assign new_new_n17934__ = ~pi009 & ~po009;
  assign new_new_n17935__ = ~pi065 & ~new_new_n17934__;
  assign new_new_n17936__ = ~pi008 & ~new_new_n17935__;
  assign new_new_n17937__ = ~new_new_n17933__ & ~new_new_n17936__;
  assign new_new_n17938__ = pi064 & ~new_new_n17937__;
  assign new_new_n17939__ = pi064 & po009;
  assign new_new_n17940__ = new_new_n17278__ & ~new_new_n17939__;
  assign new_new_n17941__ = ~new_new_n17938__ & ~new_new_n17940__;
  assign new_new_n17942__ = pi066 & ~new_new_n17941__;
  assign new_new_n17943__ = po009 & new_new_n17910__;
  assign new_new_n17944__ = new_new_n426__ & ~po010;
  assign new_new_n17945__ = ~new_new_n17943__ & ~new_new_n17944__;
  assign new_new_n17946__ = ~pi009 & ~new_new_n17945__;
  assign new_new_n17947__ = ~new_new_n332__ & po009;
  assign new_new_n17948__ = ~new_new_n17297__ & ~new_new_n17947__;
  assign new_new_n17949__ = pi065 & po009;
  assign new_new_n17950__ = po010 & ~new_new_n17949__;
  assign new_new_n17951__ = pi009 & ~new_new_n17298__;
  assign new_new_n17952__ = ~new_new_n17950__ & new_new_n17951__;
  assign new_new_n17953__ = ~new_new_n17946__ & ~new_new_n17948__;
  assign new_new_n17954__ = ~new_new_n17952__ & new_new_n17953__;
  assign new_new_n17955__ = ~pi010 & ~new_new_n17954__;
  assign new_new_n17956__ = ~new_new_n17297__ & ~new_new_n17949__;
  assign new_new_n17957__ = pi064 & ~new_new_n17287__;
  assign new_new_n17958__ = ~new_new_n17956__ & ~new_new_n17957__;
  assign new_new_n17959__ = ~pi065 & po009;
  assign new_new_n17960__ = ~po010 & ~new_new_n17959__;
  assign new_new_n17961__ = pi064 & ~new_new_n17931__;
  assign new_new_n17962__ = ~new_new_n17943__ & new_new_n17961__;
  assign new_new_n17963__ = ~new_new_n17960__ & new_new_n17962__;
  assign new_new_n17964__ = ~new_new_n17958__ & ~new_new_n17963__;
  assign new_new_n17965__ = pi010 & ~new_new_n17964__;
  assign new_new_n17966__ = ~new_new_n17955__ & ~new_new_n17965__;
  assign new_new_n17967__ = ~pi066 & new_new_n17941__;
  assign new_new_n17968__ = ~new_new_n17966__ & ~new_new_n17967__;
  assign new_new_n17969__ = ~new_new_n17942__ & ~new_new_n17968__;
  assign new_new_n17970__ = ~pi067 & new_new_n17929__;
  assign new_new_n17971__ = ~new_new_n17969__ & ~new_new_n17970__;
  assign new_new_n17972__ = ~new_new_n17930__ & ~new_new_n17971__;
  assign new_new_n17973__ = ~pi068 & new_new_n17972__;
  assign new_new_n17974__ = pi068 & ~new_new_n17972__;
  assign new_new_n17975__ = ~pi067 & ~new_new_n17319__;
  assign new_new_n17976__ = pi067 & new_new_n17319__;
  assign new_new_n17977__ = ~new_new_n17975__ & ~new_new_n17976__;
  assign new_new_n17978__ = po009 & new_new_n17977__;
  assign new_new_n17979__ = new_new_n17275__ & new_new_n17978__;
  assign new_new_n17980__ = ~new_new_n17275__ & ~new_new_n17978__;
  assign new_new_n17981__ = ~new_new_n17979__ & ~new_new_n17980__;
  assign new_new_n17982__ = ~new_new_n17974__ & ~new_new_n17981__;
  assign new_new_n17983__ = ~new_new_n17973__ & ~new_new_n17982__;
  assign new_new_n17984__ = ~new_new_n17896__ & ~new_new_n17983__;
  assign new_new_n17985__ = ~new_new_n17895__ & ~new_new_n17984__;
  assign new_new_n17986__ = ~new_new_n17887__ & ~new_new_n17985__;
  assign new_new_n17987__ = ~new_new_n17886__ & ~new_new_n17986__;
  assign new_new_n17988__ = ~new_new_n17880__ & ~new_new_n17987__;
  assign new_new_n17989__ = ~new_new_n17879__ & ~new_new_n17988__;
  assign new_new_n17990__ = ~new_new_n17871__ & new_new_n17989__;
  assign new_new_n17991__ = ~new_new_n17870__ & ~new_new_n17990__;
  assign new_new_n17992__ = ~new_new_n17862__ & ~new_new_n17991__;
  assign new_new_n17993__ = ~new_new_n17861__ & ~new_new_n17992__;
  assign new_new_n17994__ = ~new_new_n17853__ & new_new_n17993__;
  assign new_new_n17995__ = ~new_new_n17852__ & ~new_new_n17994__;
  assign new_new_n17996__ = ~new_new_n17844__ & ~new_new_n17995__;
  assign new_new_n17997__ = ~new_new_n17843__ & ~new_new_n17996__;
  assign new_new_n17998__ = ~new_new_n17835__ & ~new_new_n17997__;
  assign new_new_n17999__ = ~new_new_n17834__ & ~new_new_n17998__;
  assign new_new_n18000__ = ~new_new_n17826__ & ~new_new_n17999__;
  assign new_new_n18001__ = ~new_new_n17825__ & ~new_new_n18000__;
  assign new_new_n18002__ = ~new_new_n17817__ & ~new_new_n18001__;
  assign new_new_n18003__ = ~new_new_n17816__ & ~new_new_n18002__;
  assign new_new_n18004__ = ~new_new_n17808__ & ~new_new_n18003__;
  assign new_new_n18005__ = ~new_new_n17807__ & ~new_new_n18004__;
  assign new_new_n18006__ = ~new_new_n17799__ & new_new_n18005__;
  assign new_new_n18007__ = ~new_new_n17798__ & ~new_new_n18006__;
  assign new_new_n18008__ = ~new_new_n17790__ & ~new_new_n18007__;
  assign new_new_n18009__ = ~new_new_n17789__ & ~new_new_n18008__;
  assign new_new_n18010__ = ~new_new_n17781__ & new_new_n18009__;
  assign new_new_n18011__ = ~new_new_n17780__ & ~new_new_n18010__;
  assign new_new_n18012__ = ~new_new_n17772__ & ~new_new_n18011__;
  assign new_new_n18013__ = ~new_new_n17771__ & ~new_new_n18012__;
  assign new_new_n18014__ = ~new_new_n17763__ & new_new_n18013__;
  assign new_new_n18015__ = ~new_new_n17762__ & ~new_new_n18014__;
  assign new_new_n18016__ = ~new_new_n17754__ & new_new_n18015__;
  assign new_new_n18017__ = ~new_new_n17753__ & ~new_new_n18016__;
  assign new_new_n18018__ = ~new_new_n17745__ & ~new_new_n18017__;
  assign new_new_n18019__ = ~new_new_n17744__ & ~new_new_n18018__;
  assign new_new_n18020__ = ~new_new_n17736__ & new_new_n18019__;
  assign new_new_n18021__ = ~new_new_n17735__ & ~new_new_n18020__;
  assign new_new_n18022__ = ~new_new_n17727__ & ~new_new_n18021__;
  assign new_new_n18023__ = ~new_new_n17726__ & ~new_new_n18022__;
  assign new_new_n18024__ = ~new_new_n17718__ & ~new_new_n18023__;
  assign new_new_n18025__ = ~new_new_n17717__ & ~new_new_n18024__;
  assign new_new_n18026__ = ~new_new_n17709__ & new_new_n18025__;
  assign new_new_n18027__ = ~new_new_n17708__ & ~new_new_n18026__;
  assign new_new_n18028__ = ~new_new_n17700__ & ~new_new_n18027__;
  assign new_new_n18029__ = ~new_new_n17699__ & ~new_new_n18028__;
  assign new_new_n18030__ = ~new_new_n17691__ & new_new_n18029__;
  assign new_new_n18031__ = ~new_new_n17690__ & ~new_new_n18030__;
  assign new_new_n18032__ = ~new_new_n17682__ & ~new_new_n18031__;
  assign new_new_n18033__ = ~new_new_n17681__ & ~new_new_n18032__;
  assign new_new_n18034__ = ~new_new_n17673__ & ~new_new_n18033__;
  assign new_new_n18035__ = ~new_new_n17672__ & ~new_new_n18034__;
  assign new_new_n18036__ = ~new_new_n17664__ & new_new_n18035__;
  assign new_new_n18037__ = ~new_new_n17663__ & ~new_new_n18036__;
  assign new_new_n18038__ = ~new_new_n17655__ & ~new_new_n18037__;
  assign new_new_n18039__ = ~new_new_n17654__ & ~new_new_n18038__;
  assign new_new_n18040__ = ~new_new_n17646__ & new_new_n18039__;
  assign new_new_n18041__ = ~new_new_n17645__ & ~new_new_n18040__;
  assign new_new_n18042__ = ~new_new_n17637__ & new_new_n18041__;
  assign new_new_n18043__ = ~new_new_n17636__ & ~new_new_n18042__;
  assign new_new_n18044__ = ~new_new_n17628__ & ~new_new_n18043__;
  assign new_new_n18045__ = ~new_new_n17627__ & ~new_new_n18044__;
  assign new_new_n18046__ = ~new_new_n17619__ & new_new_n18045__;
  assign new_new_n18047__ = ~new_new_n17618__ & ~new_new_n18046__;
  assign new_new_n18048__ = ~new_new_n17610__ & ~new_new_n18047__;
  assign new_new_n18049__ = ~new_new_n17609__ & ~new_new_n18048__;
  assign new_new_n18050__ = ~new_new_n17601__ & new_new_n18049__;
  assign new_new_n18051__ = ~new_new_n17600__ & ~new_new_n18050__;
  assign new_new_n18052__ = ~new_new_n17592__ & ~new_new_n18051__;
  assign new_new_n18053__ = ~new_new_n17591__ & ~new_new_n18052__;
  assign new_new_n18054__ = ~new_new_n17583__ & ~new_new_n18053__;
  assign new_new_n18055__ = ~new_new_n17582__ & ~new_new_n18054__;
  assign new_new_n18056__ = ~new_new_n17574__ & ~new_new_n18055__;
  assign new_new_n18057__ = ~new_new_n17573__ & ~new_new_n18056__;
  assign new_new_n18058__ = ~new_new_n17565__ & ~new_new_n18057__;
  assign new_new_n18059__ = ~new_new_n17564__ & ~new_new_n18058__;
  assign new_new_n18060__ = ~new_new_n17556__ & ~new_new_n18059__;
  assign new_new_n18061__ = ~new_new_n17555__ & ~new_new_n18060__;
  assign new_new_n18062__ = ~new_new_n17547__ & ~new_new_n18061__;
  assign new_new_n18063__ = ~new_new_n17546__ & ~new_new_n18062__;
  assign new_new_n18064__ = ~new_new_n17538__ & new_new_n18063__;
  assign new_new_n18065__ = ~new_new_n17537__ & ~new_new_n18064__;
  assign new_new_n18066__ = ~new_new_n17529__ & ~new_new_n18065__;
  assign new_new_n18067__ = ~new_new_n17528__ & ~new_new_n18066__;
  assign new_new_n18068__ = ~new_new_n17522__ & ~new_new_n18067__;
  assign new_new_n18069__ = ~new_new_n17521__ & ~new_new_n18068__;
  assign new_new_n18070__ = ~new_new_n17513__ & ~new_new_n18069__;
  assign new_new_n18071__ = ~new_new_n17512__ & ~new_new_n18070__;
  assign new_new_n18072__ = ~new_new_n17504__ & new_new_n18071__;
  assign new_new_n18073__ = ~new_new_n17503__ & ~new_new_n18072__;
  assign new_new_n18074__ = ~new_new_n17495__ & new_new_n18073__;
  assign new_new_n18075__ = ~new_new_n17494__ & ~new_new_n18074__;
  assign new_new_n18076__ = ~new_new_n17486__ & ~new_new_n18075__;
  assign new_new_n18077__ = ~new_new_n17485__ & ~new_new_n18076__;
  assign new_new_n18078__ = ~new_new_n17477__ & new_new_n18077__;
  assign new_new_n18079__ = ~new_new_n17476__ & ~new_new_n18078__;
  assign new_new_n18080__ = ~new_new_n17468__ & ~new_new_n18079__;
  assign new_new_n18081__ = ~new_new_n17467__ & ~new_new_n18080__;
  assign new_new_n18082__ = ~pi119 & new_new_n17442__;
  assign new_new_n18083__ = ~new_new_n17455__ & ~new_new_n18081__;
  assign new_new_n18084__ = ~new_new_n17456__ & ~new_new_n18083__;
  assign new_new_n18085__ = ~new_new_n18082__ & new_new_n18084__;
  assign new_new_n18086__ = pi119 & ~new_new_n16229__;
  assign new_new_n18087__ = new_new_n16826__ & ~new_new_n18086__;
  assign po008 = ~new_new_n18085__ & new_new_n18087__;
  assign new_new_n18089__ = ~new_new_n18081__ & po008;
  assign new_new_n18090__ = ~pi118 & ~po008;
  assign new_new_n18091__ = ~new_new_n18089__ & ~new_new_n18090__;
  assign new_new_n18092__ = new_new_n17457__ & ~new_new_n18091__;
  assign new_new_n18093__ = ~new_new_n17457__ & new_new_n18091__;
  assign new_new_n18094__ = ~new_new_n18092__ & ~new_new_n18093__;
  assign new_new_n18095__ = pi119 & ~new_new_n18094__;
  assign new_new_n18096__ = ~pi119 & new_new_n18094__;
  assign new_new_n18097__ = ~new_new_n17467__ & ~new_new_n17468__;
  assign new_new_n18098__ = ~new_new_n18079__ & po008;
  assign new_new_n18099__ = ~pi117 & ~po008;
  assign new_new_n18100__ = ~new_new_n18098__ & ~new_new_n18099__;
  assign new_new_n18101__ = new_new_n18097__ & ~new_new_n18100__;
  assign new_new_n18102__ = ~new_new_n18097__ & new_new_n18100__;
  assign new_new_n18103__ = ~new_new_n18101__ & ~new_new_n18102__;
  assign new_new_n18104__ = ~pi118 & new_new_n18103__;
  assign new_new_n18105__ = pi118 & ~new_new_n18103__;
  assign new_new_n18106__ = ~new_new_n18077__ & po008;
  assign new_new_n18107__ = pi116 & ~po008;
  assign new_new_n18108__ = ~new_new_n18106__ & ~new_new_n18107__;
  assign new_new_n18109__ = ~new_new_n17476__ & ~new_new_n17477__;
  assign new_new_n18110__ = ~new_new_n18108__ & new_new_n18109__;
  assign new_new_n18111__ = new_new_n18108__ & ~new_new_n18109__;
  assign new_new_n18112__ = ~new_new_n18110__ & ~new_new_n18111__;
  assign new_new_n18113__ = ~pi117 & ~new_new_n18112__;
  assign new_new_n18114__ = pi117 & new_new_n18112__;
  assign new_new_n18115__ = pi115 & ~new_new_n18075__;
  assign new_new_n18116__ = ~pi115 & new_new_n18075__;
  assign new_new_n18117__ = ~new_new_n18115__ & ~new_new_n18116__;
  assign new_new_n18118__ = po008 & new_new_n18117__;
  assign new_new_n18119__ = new_new_n17484__ & new_new_n18118__;
  assign new_new_n18120__ = ~new_new_n17484__ & ~new_new_n18118__;
  assign new_new_n18121__ = ~new_new_n18119__ & ~new_new_n18120__;
  assign new_new_n18122__ = pi116 & ~new_new_n18121__;
  assign new_new_n18123__ = ~pi116 & new_new_n18121__;
  assign new_new_n18124__ = ~new_new_n17494__ & ~new_new_n17495__;
  assign new_new_n18125__ = ~new_new_n18073__ & po008;
  assign new_new_n18126__ = ~pi114 & ~po008;
  assign new_new_n18127__ = ~new_new_n18125__ & ~new_new_n18126__;
  assign new_new_n18128__ = new_new_n18124__ & ~new_new_n18127__;
  assign new_new_n18129__ = ~new_new_n18124__ & new_new_n18127__;
  assign new_new_n18130__ = ~new_new_n18128__ & ~new_new_n18129__;
  assign new_new_n18131__ = ~pi115 & new_new_n18130__;
  assign new_new_n18132__ = pi115 & ~new_new_n18130__;
  assign new_new_n18133__ = ~new_new_n17503__ & ~new_new_n17504__;
  assign new_new_n18134__ = new_new_n18071__ & po008;
  assign new_new_n18135__ = ~pi113 & ~po008;
  assign new_new_n18136__ = ~new_new_n18134__ & ~new_new_n18135__;
  assign new_new_n18137__ = ~new_new_n18133__ & ~new_new_n18136__;
  assign new_new_n18138__ = new_new_n18133__ & new_new_n18136__;
  assign new_new_n18139__ = ~new_new_n18137__ & ~new_new_n18138__;
  assign new_new_n18140__ = ~pi114 & ~new_new_n18139__;
  assign new_new_n18141__ = pi114 & new_new_n18139__;
  assign new_new_n18142__ = new_new_n18069__ & po008;
  assign new_new_n18143__ = ~pi112 & ~po008;
  assign new_new_n18144__ = ~new_new_n18142__ & ~new_new_n18143__;
  assign new_new_n18145__ = ~new_new_n17512__ & ~new_new_n17513__;
  assign new_new_n18146__ = ~new_new_n18144__ & ~new_new_n18145__;
  assign new_new_n18147__ = new_new_n18144__ & new_new_n18145__;
  assign new_new_n18148__ = ~new_new_n18146__ & ~new_new_n18147__;
  assign new_new_n18149__ = ~pi113 & ~new_new_n18148__;
  assign new_new_n18150__ = pi113 & new_new_n18148__;
  assign new_new_n18151__ = ~new_new_n18067__ & po008;
  assign new_new_n18152__ = pi111 & ~po008;
  assign new_new_n18153__ = ~new_new_n18151__ & ~new_new_n18152__;
  assign new_new_n18154__ = ~new_new_n17521__ & ~new_new_n17522__;
  assign new_new_n18155__ = ~new_new_n18153__ & new_new_n18154__;
  assign new_new_n18156__ = new_new_n18153__ & ~new_new_n18154__;
  assign new_new_n18157__ = ~new_new_n18155__ & ~new_new_n18156__;
  assign new_new_n18158__ = ~pi112 & ~new_new_n18157__;
  assign new_new_n18159__ = pi112 & new_new_n18157__;
  assign new_new_n18160__ = ~new_new_n17528__ & ~new_new_n17529__;
  assign new_new_n18161__ = pi110 & ~po008;
  assign new_new_n18162__ = ~new_new_n18065__ & po008;
  assign new_new_n18163__ = ~new_new_n18161__ & ~new_new_n18162__;
  assign new_new_n18164__ = new_new_n18160__ & ~new_new_n18163__;
  assign new_new_n18165__ = ~new_new_n18160__ & new_new_n18163__;
  assign new_new_n18166__ = ~new_new_n18164__ & ~new_new_n18165__;
  assign new_new_n18167__ = ~pi111 & ~new_new_n18166__;
  assign new_new_n18168__ = pi111 & new_new_n18166__;
  assign new_new_n18169__ = ~new_new_n17537__ & ~new_new_n17538__;
  assign new_new_n18170__ = ~new_new_n18063__ & po008;
  assign new_new_n18171__ = ~pi109 & ~po008;
  assign new_new_n18172__ = ~new_new_n18170__ & ~new_new_n18171__;
  assign new_new_n18173__ = new_new_n18169__ & ~new_new_n18172__;
  assign new_new_n18174__ = ~new_new_n18169__ & new_new_n18172__;
  assign new_new_n18175__ = ~new_new_n18173__ & ~new_new_n18174__;
  assign new_new_n18176__ = pi110 & ~new_new_n18175__;
  assign new_new_n18177__ = ~pi110 & new_new_n18175__;
  assign new_new_n18178__ = ~new_new_n17546__ & ~new_new_n17547__;
  assign new_new_n18179__ = ~new_new_n18061__ & po008;
  assign new_new_n18180__ = ~pi108 & ~po008;
  assign new_new_n18181__ = ~new_new_n18179__ & ~new_new_n18180__;
  assign new_new_n18182__ = new_new_n18178__ & ~new_new_n18181__;
  assign new_new_n18183__ = ~new_new_n18178__ & new_new_n18181__;
  assign new_new_n18184__ = ~new_new_n18182__ & ~new_new_n18183__;
  assign new_new_n18185__ = pi109 & ~new_new_n18184__;
  assign new_new_n18186__ = ~pi109 & new_new_n18184__;
  assign new_new_n18187__ = ~pi107 & ~new_new_n18059__;
  assign new_new_n18188__ = pi107 & new_new_n18059__;
  assign new_new_n18189__ = ~new_new_n18187__ & ~new_new_n18188__;
  assign new_new_n18190__ = po008 & new_new_n18189__;
  assign new_new_n18191__ = new_new_n17554__ & ~new_new_n18190__;
  assign new_new_n18192__ = ~new_new_n17554__ & new_new_n18190__;
  assign new_new_n18193__ = ~new_new_n18191__ & ~new_new_n18192__;
  assign new_new_n18194__ = ~pi108 & new_new_n18193__;
  assign new_new_n18195__ = pi108 & ~new_new_n18193__;
  assign new_new_n18196__ = ~new_new_n17564__ & ~new_new_n17565__;
  assign new_new_n18197__ = ~new_new_n18057__ & po008;
  assign new_new_n18198__ = ~pi106 & ~po008;
  assign new_new_n18199__ = ~new_new_n18197__ & ~new_new_n18198__;
  assign new_new_n18200__ = new_new_n18196__ & ~new_new_n18199__;
  assign new_new_n18201__ = ~new_new_n18196__ & new_new_n18199__;
  assign new_new_n18202__ = ~new_new_n18200__ & ~new_new_n18201__;
  assign new_new_n18203__ = ~pi107 & new_new_n18202__;
  assign new_new_n18204__ = pi107 & ~new_new_n18202__;
  assign new_new_n18205__ = ~pi105 & ~new_new_n18055__;
  assign new_new_n18206__ = pi105 & new_new_n18055__;
  assign new_new_n18207__ = ~new_new_n18205__ & ~new_new_n18206__;
  assign new_new_n18208__ = po008 & new_new_n18207__;
  assign new_new_n18209__ = new_new_n17572__ & new_new_n18208__;
  assign new_new_n18210__ = ~new_new_n17572__ & ~new_new_n18208__;
  assign new_new_n18211__ = ~new_new_n18209__ & ~new_new_n18210__;
  assign new_new_n18212__ = ~pi106 & ~new_new_n18211__;
  assign new_new_n18213__ = pi106 & new_new_n18211__;
  assign new_new_n18214__ = ~new_new_n17582__ & ~new_new_n17583__;
  assign new_new_n18215__ = ~new_new_n18053__ & po008;
  assign new_new_n18216__ = ~pi104 & ~po008;
  assign new_new_n18217__ = ~new_new_n18215__ & ~new_new_n18216__;
  assign new_new_n18218__ = new_new_n18214__ & ~new_new_n18217__;
  assign new_new_n18219__ = ~new_new_n18214__ & new_new_n18217__;
  assign new_new_n18220__ = ~new_new_n18218__ & ~new_new_n18219__;
  assign new_new_n18221__ = pi105 & ~new_new_n18220__;
  assign new_new_n18222__ = ~pi105 & new_new_n18220__;
  assign new_new_n18223__ = ~new_new_n17591__ & ~new_new_n17592__;
  assign new_new_n18224__ = ~new_new_n18051__ & po008;
  assign new_new_n18225__ = ~pi103 & ~po008;
  assign new_new_n18226__ = ~new_new_n18224__ & ~new_new_n18225__;
  assign new_new_n18227__ = new_new_n18223__ & ~new_new_n18226__;
  assign new_new_n18228__ = ~new_new_n18223__ & new_new_n18226__;
  assign new_new_n18229__ = ~new_new_n18227__ & ~new_new_n18228__;
  assign new_new_n18230__ = pi104 & ~new_new_n18229__;
  assign new_new_n18231__ = ~pi104 & new_new_n18229__;
  assign new_new_n18232__ = ~new_new_n17600__ & ~new_new_n17601__;
  assign new_new_n18233__ = pi102 & ~po008;
  assign new_new_n18234__ = ~new_new_n18049__ & po008;
  assign new_new_n18235__ = ~new_new_n18233__ & ~new_new_n18234__;
  assign new_new_n18236__ = new_new_n18232__ & ~new_new_n18235__;
  assign new_new_n18237__ = ~new_new_n18232__ & new_new_n18235__;
  assign new_new_n18238__ = ~new_new_n18236__ & ~new_new_n18237__;
  assign new_new_n18239__ = ~pi103 & ~new_new_n18238__;
  assign new_new_n18240__ = pi103 & new_new_n18238__;
  assign new_new_n18241__ = ~new_new_n17609__ & ~new_new_n17610__;
  assign new_new_n18242__ = pi101 & ~po008;
  assign new_new_n18243__ = ~new_new_n18047__ & po008;
  assign new_new_n18244__ = ~new_new_n18242__ & ~new_new_n18243__;
  assign new_new_n18245__ = new_new_n18241__ & ~new_new_n18244__;
  assign new_new_n18246__ = ~new_new_n18241__ & new_new_n18244__;
  assign new_new_n18247__ = ~new_new_n18245__ & ~new_new_n18246__;
  assign new_new_n18248__ = ~pi102 & ~new_new_n18247__;
  assign new_new_n18249__ = pi102 & new_new_n18247__;
  assign new_new_n18250__ = ~new_new_n17618__ & ~new_new_n17619__;
  assign new_new_n18251__ = ~new_new_n18045__ & po008;
  assign new_new_n18252__ = ~pi100 & ~po008;
  assign new_new_n18253__ = ~new_new_n18251__ & ~new_new_n18252__;
  assign new_new_n18254__ = new_new_n18250__ & new_new_n18253__;
  assign new_new_n18255__ = ~new_new_n18250__ & ~new_new_n18253__;
  assign new_new_n18256__ = ~new_new_n18254__ & ~new_new_n18255__;
  assign new_new_n18257__ = pi101 & new_new_n18256__;
  assign new_new_n18258__ = ~pi101 & ~new_new_n18256__;
  assign new_new_n18259__ = ~new_new_n17627__ & ~new_new_n17628__;
  assign new_new_n18260__ = ~new_new_n18043__ & po008;
  assign new_new_n18261__ = ~pi099 & ~po008;
  assign new_new_n18262__ = ~new_new_n18260__ & ~new_new_n18261__;
  assign new_new_n18263__ = new_new_n18259__ & ~new_new_n18262__;
  assign new_new_n18264__ = ~new_new_n18259__ & new_new_n18262__;
  assign new_new_n18265__ = ~new_new_n18263__ & ~new_new_n18264__;
  assign new_new_n18266__ = pi100 & ~new_new_n18265__;
  assign new_new_n18267__ = ~pi100 & new_new_n18265__;
  assign new_new_n18268__ = ~new_new_n18041__ & po008;
  assign new_new_n18269__ = pi098 & ~po008;
  assign new_new_n18270__ = ~new_new_n18268__ & ~new_new_n18269__;
  assign new_new_n18271__ = ~new_new_n17636__ & ~new_new_n17637__;
  assign new_new_n18272__ = ~new_new_n18270__ & new_new_n18271__;
  assign new_new_n18273__ = new_new_n18270__ & ~new_new_n18271__;
  assign new_new_n18274__ = ~new_new_n18272__ & ~new_new_n18273__;
  assign new_new_n18275__ = pi099 & new_new_n18274__;
  assign new_new_n18276__ = ~pi099 & ~new_new_n18274__;
  assign new_new_n18277__ = ~new_new_n17645__ & ~new_new_n17646__;
  assign new_new_n18278__ = ~new_new_n18039__ & po008;
  assign new_new_n18279__ = ~pi097 & ~po008;
  assign new_new_n18280__ = ~new_new_n18278__ & ~new_new_n18279__;
  assign new_new_n18281__ = new_new_n18277__ & ~new_new_n18280__;
  assign new_new_n18282__ = ~new_new_n18277__ & new_new_n18280__;
  assign new_new_n18283__ = ~new_new_n18281__ & ~new_new_n18282__;
  assign new_new_n18284__ = pi098 & ~new_new_n18283__;
  assign new_new_n18285__ = ~pi098 & new_new_n18283__;
  assign new_new_n18286__ = ~new_new_n17654__ & ~new_new_n17655__;
  assign new_new_n18287__ = ~new_new_n18037__ & po008;
  assign new_new_n18288__ = ~pi096 & ~po008;
  assign new_new_n18289__ = ~new_new_n18287__ & ~new_new_n18288__;
  assign new_new_n18290__ = ~new_new_n18286__ & ~new_new_n18289__;
  assign new_new_n18291__ = new_new_n18286__ & new_new_n18289__;
  assign new_new_n18292__ = ~new_new_n18290__ & ~new_new_n18291__;
  assign new_new_n18293__ = ~pi097 & ~new_new_n18292__;
  assign new_new_n18294__ = pi097 & new_new_n18292__;
  assign new_new_n18295__ = new_new_n18035__ & po008;
  assign new_new_n18296__ = ~pi095 & ~po008;
  assign new_new_n18297__ = ~new_new_n18295__ & ~new_new_n18296__;
  assign new_new_n18298__ = ~new_new_n17663__ & ~new_new_n17664__;
  assign new_new_n18299__ = ~new_new_n18297__ & ~new_new_n18298__;
  assign new_new_n18300__ = new_new_n18297__ & new_new_n18298__;
  assign new_new_n18301__ = ~new_new_n18299__ & ~new_new_n18300__;
  assign new_new_n18302__ = ~pi096 & ~new_new_n18301__;
  assign new_new_n18303__ = pi096 & new_new_n18301__;
  assign new_new_n18304__ = ~new_new_n17672__ & ~new_new_n17673__;
  assign new_new_n18305__ = ~new_new_n18033__ & po008;
  assign new_new_n18306__ = pi094 & ~po008;
  assign new_new_n18307__ = ~new_new_n18305__ & ~new_new_n18306__;
  assign new_new_n18308__ = new_new_n18304__ & ~new_new_n18307__;
  assign new_new_n18309__ = ~new_new_n18304__ & new_new_n18307__;
  assign new_new_n18310__ = ~new_new_n18308__ & ~new_new_n18309__;
  assign new_new_n18311__ = pi095 & new_new_n18310__;
  assign new_new_n18312__ = ~pi095 & ~new_new_n18310__;
  assign new_new_n18313__ = pi093 & ~new_new_n18031__;
  assign new_new_n18314__ = ~pi093 & new_new_n18031__;
  assign new_new_n18315__ = ~new_new_n18313__ & ~new_new_n18314__;
  assign new_new_n18316__ = po008 & new_new_n18315__;
  assign new_new_n18317__ = new_new_n17680__ & new_new_n18316__;
  assign new_new_n18318__ = ~new_new_n17680__ & ~new_new_n18316__;
  assign new_new_n18319__ = ~new_new_n18317__ & ~new_new_n18318__;
  assign new_new_n18320__ = pi094 & ~new_new_n18319__;
  assign new_new_n18321__ = ~pi094 & new_new_n18319__;
  assign new_new_n18322__ = ~new_new_n17690__ & ~new_new_n17691__;
  assign new_new_n18323__ = ~new_new_n18029__ & po008;
  assign new_new_n18324__ = ~pi092 & ~po008;
  assign new_new_n18325__ = ~new_new_n18323__ & ~new_new_n18324__;
  assign new_new_n18326__ = new_new_n18322__ & ~new_new_n18325__;
  assign new_new_n18327__ = ~new_new_n18322__ & new_new_n18325__;
  assign new_new_n18328__ = ~new_new_n18326__ & ~new_new_n18327__;
  assign new_new_n18329__ = pi093 & ~new_new_n18328__;
  assign new_new_n18330__ = ~pi093 & new_new_n18328__;
  assign new_new_n18331__ = ~new_new_n17699__ & ~new_new_n17700__;
  assign new_new_n18332__ = ~new_new_n18027__ & po008;
  assign new_new_n18333__ = ~pi091 & ~po008;
  assign new_new_n18334__ = ~new_new_n18332__ & ~new_new_n18333__;
  assign new_new_n18335__ = new_new_n18331__ & ~new_new_n18334__;
  assign new_new_n18336__ = ~new_new_n18331__ & new_new_n18334__;
  assign new_new_n18337__ = ~new_new_n18335__ & ~new_new_n18336__;
  assign new_new_n18338__ = ~pi092 & new_new_n18337__;
  assign new_new_n18339__ = pi092 & ~new_new_n18337__;
  assign new_new_n18340__ = ~new_new_n17708__ & ~new_new_n17709__;
  assign new_new_n18341__ = pi090 & ~po008;
  assign new_new_n18342__ = ~new_new_n18025__ & po008;
  assign new_new_n18343__ = ~new_new_n18341__ & ~new_new_n18342__;
  assign new_new_n18344__ = new_new_n18340__ & ~new_new_n18343__;
  assign new_new_n18345__ = ~new_new_n18340__ & new_new_n18343__;
  assign new_new_n18346__ = ~new_new_n18344__ & ~new_new_n18345__;
  assign new_new_n18347__ = ~pi091 & ~new_new_n18346__;
  assign new_new_n18348__ = pi091 & new_new_n18346__;
  assign new_new_n18349__ = ~new_new_n18023__ & po008;
  assign new_new_n18350__ = pi089 & ~po008;
  assign new_new_n18351__ = ~new_new_n18349__ & ~new_new_n18350__;
  assign new_new_n18352__ = ~new_new_n17717__ & ~new_new_n17718__;
  assign new_new_n18353__ = ~new_new_n18351__ & new_new_n18352__;
  assign new_new_n18354__ = new_new_n18351__ & ~new_new_n18352__;
  assign new_new_n18355__ = ~new_new_n18353__ & ~new_new_n18354__;
  assign new_new_n18356__ = ~pi090 & ~new_new_n18355__;
  assign new_new_n18357__ = pi090 & new_new_n18355__;
  assign new_new_n18358__ = pi088 & ~new_new_n18021__;
  assign new_new_n18359__ = ~pi088 & new_new_n18021__;
  assign new_new_n18360__ = ~new_new_n18358__ & ~new_new_n18359__;
  assign new_new_n18361__ = po008 & new_new_n18360__;
  assign new_new_n18362__ = ~new_new_n17725__ & ~new_new_n18361__;
  assign new_new_n18363__ = new_new_n17725__ & new_new_n18361__;
  assign new_new_n18364__ = ~new_new_n18362__ & ~new_new_n18363__;
  assign new_new_n18365__ = pi089 & ~new_new_n18364__;
  assign new_new_n18366__ = ~pi089 & new_new_n18364__;
  assign new_new_n18367__ = ~new_new_n17735__ & ~new_new_n17736__;
  assign new_new_n18368__ = ~new_new_n18019__ & po008;
  assign new_new_n18369__ = ~pi087 & ~po008;
  assign new_new_n18370__ = ~new_new_n18368__ & ~new_new_n18369__;
  assign new_new_n18371__ = new_new_n18367__ & ~new_new_n18370__;
  assign new_new_n18372__ = ~new_new_n18367__ & new_new_n18370__;
  assign new_new_n18373__ = ~new_new_n18371__ & ~new_new_n18372__;
  assign new_new_n18374__ = pi088 & ~new_new_n18373__;
  assign new_new_n18375__ = ~pi088 & new_new_n18373__;
  assign new_new_n18376__ = ~new_new_n17744__ & ~new_new_n17745__;
  assign new_new_n18377__ = ~new_new_n18017__ & po008;
  assign new_new_n18378__ = ~pi086 & ~po008;
  assign new_new_n18379__ = ~new_new_n18377__ & ~new_new_n18378__;
  assign new_new_n18380__ = new_new_n18376__ & ~new_new_n18379__;
  assign new_new_n18381__ = ~new_new_n18376__ & new_new_n18379__;
  assign new_new_n18382__ = ~new_new_n18380__ & ~new_new_n18381__;
  assign new_new_n18383__ = pi087 & ~new_new_n18382__;
  assign new_new_n18384__ = ~pi087 & new_new_n18382__;
  assign new_new_n18385__ = ~new_new_n17753__ & ~new_new_n17754__;
  assign new_new_n18386__ = pi085 & ~po008;
  assign new_new_n18387__ = ~new_new_n18015__ & po008;
  assign new_new_n18388__ = ~new_new_n18386__ & ~new_new_n18387__;
  assign new_new_n18389__ = new_new_n18385__ & ~new_new_n18388__;
  assign new_new_n18390__ = ~new_new_n18385__ & new_new_n18388__;
  assign new_new_n18391__ = ~new_new_n18389__ & ~new_new_n18390__;
  assign new_new_n18392__ = ~pi086 & ~new_new_n18391__;
  assign new_new_n18393__ = pi086 & new_new_n18391__;
  assign new_new_n18394__ = ~new_new_n17762__ & ~new_new_n17763__;
  assign new_new_n18395__ = ~new_new_n18013__ & po008;
  assign new_new_n18396__ = ~pi084 & ~po008;
  assign new_new_n18397__ = ~new_new_n18395__ & ~new_new_n18396__;
  assign new_new_n18398__ = new_new_n18394__ & ~new_new_n18397__;
  assign new_new_n18399__ = ~new_new_n18394__ & new_new_n18397__;
  assign new_new_n18400__ = ~new_new_n18398__ & ~new_new_n18399__;
  assign new_new_n18401__ = ~pi085 & new_new_n18400__;
  assign new_new_n18402__ = pi085 & ~new_new_n18400__;
  assign new_new_n18403__ = ~pi083 & ~new_new_n18011__;
  assign new_new_n18404__ = pi083 & new_new_n18011__;
  assign new_new_n18405__ = ~new_new_n18403__ & ~new_new_n18404__;
  assign new_new_n18406__ = po008 & new_new_n18405__;
  assign new_new_n18407__ = new_new_n17770__ & new_new_n18406__;
  assign new_new_n18408__ = ~new_new_n17770__ & ~new_new_n18406__;
  assign new_new_n18409__ = ~new_new_n18407__ & ~new_new_n18408__;
  assign new_new_n18410__ = ~pi084 & ~new_new_n18409__;
  assign new_new_n18411__ = pi084 & new_new_n18409__;
  assign new_new_n18412__ = ~new_new_n17780__ & ~new_new_n17781__;
  assign new_new_n18413__ = pi082 & ~po008;
  assign new_new_n18414__ = ~new_new_n18009__ & po008;
  assign new_new_n18415__ = ~new_new_n18413__ & ~new_new_n18414__;
  assign new_new_n18416__ = new_new_n18412__ & ~new_new_n18415__;
  assign new_new_n18417__ = ~new_new_n18412__ & new_new_n18415__;
  assign new_new_n18418__ = ~new_new_n18416__ & ~new_new_n18417__;
  assign new_new_n18419__ = ~pi083 & ~new_new_n18418__;
  assign new_new_n18420__ = pi083 & new_new_n18418__;
  assign new_new_n18421__ = ~new_new_n18007__ & po008;
  assign new_new_n18422__ = pi081 & ~po008;
  assign new_new_n18423__ = ~new_new_n18421__ & ~new_new_n18422__;
  assign new_new_n18424__ = ~new_new_n17789__ & ~new_new_n17790__;
  assign new_new_n18425__ = ~new_new_n18423__ & new_new_n18424__;
  assign new_new_n18426__ = new_new_n18423__ & ~new_new_n18424__;
  assign new_new_n18427__ = ~new_new_n18425__ & ~new_new_n18426__;
  assign new_new_n18428__ = pi082 & new_new_n18427__;
  assign new_new_n18429__ = ~pi082 & ~new_new_n18427__;
  assign new_new_n18430__ = ~new_new_n17798__ & ~new_new_n17799__;
  assign new_new_n18431__ = ~new_new_n18005__ & po008;
  assign new_new_n18432__ = ~pi080 & ~po008;
  assign new_new_n18433__ = ~new_new_n18431__ & ~new_new_n18432__;
  assign new_new_n18434__ = new_new_n18430__ & ~new_new_n18433__;
  assign new_new_n18435__ = ~new_new_n18430__ & new_new_n18433__;
  assign new_new_n18436__ = ~new_new_n18434__ & ~new_new_n18435__;
  assign new_new_n18437__ = pi081 & ~new_new_n18436__;
  assign new_new_n18438__ = ~pi081 & new_new_n18436__;
  assign new_new_n18439__ = ~pi079 & ~new_new_n18003__;
  assign new_new_n18440__ = pi079 & new_new_n18003__;
  assign new_new_n18441__ = ~new_new_n18439__ & ~new_new_n18440__;
  assign new_new_n18442__ = po008 & new_new_n18441__;
  assign new_new_n18443__ = ~new_new_n17806__ & new_new_n18442__;
  assign new_new_n18444__ = new_new_n17806__ & ~new_new_n18442__;
  assign new_new_n18445__ = ~new_new_n18443__ & ~new_new_n18444__;
  assign new_new_n18446__ = pi080 & ~new_new_n18445__;
  assign new_new_n18447__ = ~pi080 & new_new_n18445__;
  assign new_new_n18448__ = ~pi078 & ~new_new_n18001__;
  assign new_new_n18449__ = pi078 & new_new_n18001__;
  assign new_new_n18450__ = ~new_new_n18448__ & ~new_new_n18449__;
  assign new_new_n18451__ = po008 & new_new_n18450__;
  assign new_new_n18452__ = new_new_n17815__ & new_new_n18451__;
  assign new_new_n18453__ = ~new_new_n17815__ & ~new_new_n18451__;
  assign new_new_n18454__ = ~new_new_n18452__ & ~new_new_n18453__;
  assign new_new_n18455__ = ~pi079 & ~new_new_n18454__;
  assign new_new_n18456__ = pi079 & new_new_n18454__;
  assign new_new_n18457__ = ~pi077 & ~new_new_n17999__;
  assign new_new_n18458__ = pi077 & new_new_n17999__;
  assign new_new_n18459__ = ~new_new_n18457__ & ~new_new_n18458__;
  assign new_new_n18460__ = po008 & new_new_n18459__;
  assign new_new_n18461__ = new_new_n17824__ & new_new_n18460__;
  assign new_new_n18462__ = ~new_new_n17824__ & ~new_new_n18460__;
  assign new_new_n18463__ = ~new_new_n18461__ & ~new_new_n18462__;
  assign new_new_n18464__ = ~pi078 & ~new_new_n18463__;
  assign new_new_n18465__ = pi078 & new_new_n18463__;
  assign new_new_n18466__ = ~pi076 & ~new_new_n17997__;
  assign new_new_n18467__ = pi076 & new_new_n17997__;
  assign new_new_n18468__ = ~new_new_n18466__ & ~new_new_n18467__;
  assign new_new_n18469__ = po008 & new_new_n18468__;
  assign new_new_n18470__ = new_new_n17833__ & new_new_n18469__;
  assign new_new_n18471__ = ~new_new_n17833__ & ~new_new_n18469__;
  assign new_new_n18472__ = ~new_new_n18470__ & ~new_new_n18471__;
  assign new_new_n18473__ = ~pi077 & ~new_new_n18472__;
  assign new_new_n18474__ = pi077 & new_new_n18472__;
  assign new_new_n18475__ = ~new_new_n17843__ & ~new_new_n17844__;
  assign new_new_n18476__ = ~new_new_n17995__ & po008;
  assign new_new_n18477__ = ~pi075 & ~po008;
  assign new_new_n18478__ = ~new_new_n18476__ & ~new_new_n18477__;
  assign new_new_n18479__ = new_new_n18475__ & ~new_new_n18478__;
  assign new_new_n18480__ = ~new_new_n18475__ & new_new_n18478__;
  assign new_new_n18481__ = ~new_new_n18479__ & ~new_new_n18480__;
  assign new_new_n18482__ = ~pi076 & new_new_n18481__;
  assign new_new_n18483__ = pi076 & ~new_new_n18481__;
  assign new_new_n18484__ = ~new_new_n17993__ & po008;
  assign new_new_n18485__ = pi074 & ~po008;
  assign new_new_n18486__ = ~new_new_n18484__ & ~new_new_n18485__;
  assign new_new_n18487__ = ~new_new_n17852__ & ~new_new_n17853__;
  assign new_new_n18488__ = ~new_new_n18486__ & new_new_n18487__;
  assign new_new_n18489__ = new_new_n18486__ & ~new_new_n18487__;
  assign new_new_n18490__ = ~new_new_n18488__ & ~new_new_n18489__;
  assign new_new_n18491__ = ~pi075 & ~new_new_n18490__;
  assign new_new_n18492__ = pi075 & new_new_n18490__;
  assign new_new_n18493__ = ~new_new_n17861__ & ~new_new_n17862__;
  assign new_new_n18494__ = new_new_n17991__ & po008;
  assign new_new_n18495__ = ~pi073 & ~po008;
  assign new_new_n18496__ = ~new_new_n18494__ & ~new_new_n18495__;
  assign new_new_n18497__ = ~new_new_n18493__ & ~new_new_n18496__;
  assign new_new_n18498__ = new_new_n18493__ & new_new_n18496__;
  assign new_new_n18499__ = ~new_new_n18497__ & ~new_new_n18498__;
  assign new_new_n18500__ = pi074 & new_new_n18499__;
  assign new_new_n18501__ = ~pi074 & ~new_new_n18499__;
  assign new_new_n18502__ = new_new_n17989__ & po008;
  assign new_new_n18503__ = pi072 & ~po008;
  assign new_new_n18504__ = ~new_new_n18502__ & ~new_new_n18503__;
  assign new_new_n18505__ = ~new_new_n17870__ & ~new_new_n17871__;
  assign new_new_n18506__ = ~new_new_n18504__ & ~new_new_n18505__;
  assign new_new_n18507__ = new_new_n18504__ & new_new_n18505__;
  assign new_new_n18508__ = ~new_new_n18506__ & ~new_new_n18507__;
  assign new_new_n18509__ = pi073 & ~new_new_n18508__;
  assign new_new_n18510__ = ~pi073 & new_new_n18508__;
  assign new_new_n18511__ = ~new_new_n17879__ & ~new_new_n17880__;
  assign new_new_n18512__ = ~new_new_n17987__ & po008;
  assign new_new_n18513__ = ~pi071 & ~po008;
  assign new_new_n18514__ = ~new_new_n18512__ & ~new_new_n18513__;
  assign new_new_n18515__ = new_new_n18511__ & ~new_new_n18514__;
  assign new_new_n18516__ = ~new_new_n18511__ & new_new_n18514__;
  assign new_new_n18517__ = ~new_new_n18515__ & ~new_new_n18516__;
  assign new_new_n18518__ = pi072 & ~new_new_n18517__;
  assign new_new_n18519__ = ~pi072 & new_new_n18517__;
  assign new_new_n18520__ = ~pi070 & ~new_new_n17985__;
  assign new_new_n18521__ = pi070 & new_new_n17985__;
  assign new_new_n18522__ = ~new_new_n18520__ & ~new_new_n18521__;
  assign new_new_n18523__ = po008 & new_new_n18522__;
  assign new_new_n18524__ = new_new_n17885__ & ~new_new_n18523__;
  assign new_new_n18525__ = ~new_new_n17885__ & new_new_n18523__;
  assign new_new_n18526__ = ~new_new_n18524__ & ~new_new_n18525__;
  assign new_new_n18527__ = ~pi071 & new_new_n18526__;
  assign new_new_n18528__ = pi071 & ~new_new_n18526__;
  assign new_new_n18529__ = ~new_new_n17895__ & ~new_new_n17896__;
  assign new_new_n18530__ = ~new_new_n17983__ & po008;
  assign new_new_n18531__ = ~pi069 & ~po008;
  assign new_new_n18532__ = ~new_new_n18530__ & ~new_new_n18531__;
  assign new_new_n18533__ = new_new_n18529__ & ~new_new_n18532__;
  assign new_new_n18534__ = ~new_new_n18529__ & new_new_n18532__;
  assign new_new_n18535__ = ~new_new_n18533__ & ~new_new_n18534__;
  assign new_new_n18536__ = ~pi070 & new_new_n18535__;
  assign new_new_n18537__ = pi070 & ~new_new_n18535__;
  assign new_new_n18538__ = ~new_new_n17973__ & ~new_new_n17974__;
  assign new_new_n18539__ = po008 & new_new_n18538__;
  assign new_new_n18540__ = new_new_n17981__ & new_new_n18539__;
  assign new_new_n18541__ = ~new_new_n17981__ & ~new_new_n18539__;
  assign new_new_n18542__ = ~new_new_n18540__ & ~new_new_n18541__;
  assign new_new_n18543__ = ~pi069 & ~new_new_n18542__;
  assign new_new_n18544__ = pi069 & new_new_n18542__;
  assign new_new_n18545__ = ~new_new_n17930__ & ~new_new_n17970__;
  assign new_new_n18546__ = ~new_new_n17969__ & po008;
  assign new_new_n18547__ = pi067 & ~po008;
  assign new_new_n18548__ = ~new_new_n18546__ & ~new_new_n18547__;
  assign new_new_n18549__ = new_new_n18545__ & ~new_new_n18548__;
  assign new_new_n18550__ = ~new_new_n18545__ & new_new_n18548__;
  assign new_new_n18551__ = ~new_new_n18549__ & ~new_new_n18550__;
  assign new_new_n18552__ = ~pi068 & ~new_new_n18551__;
  assign new_new_n18553__ = pi068 & new_new_n18551__;
  assign new_new_n18554__ = ~new_new_n17942__ & ~new_new_n17967__;
  assign new_new_n18555__ = po008 & new_new_n18554__;
  assign new_new_n18556__ = new_new_n17966__ & ~new_new_n18555__;
  assign new_new_n18557__ = ~new_new_n17966__ & new_new_n18555__;
  assign new_new_n18558__ = ~new_new_n18556__ & ~new_new_n18557__;
  assign new_new_n18559__ = ~pi067 & ~new_new_n18558__;
  assign new_new_n18560__ = pi067 & new_new_n18558__;
  assign new_new_n18561__ = pi008 & po008;
  assign new_new_n18562__ = ~pi008 & ~po008;
  assign new_new_n18563__ = ~pi065 & ~new_new_n18561__;
  assign new_new_n18564__ = ~new_new_n18562__ & new_new_n18563__;
  assign new_new_n18565__ = ~pi007 & ~new_new_n18564__;
  assign new_new_n18566__ = pi065 & new_new_n18561__;
  assign new_new_n18567__ = ~new_new_n18565__ & ~new_new_n18566__;
  assign new_new_n18568__ = pi064 & ~new_new_n18567__;
  assign new_new_n18569__ = pi064 & po008;
  assign new_new_n18570__ = ~pi008 & pi065;
  assign new_new_n18571__ = ~new_new_n18569__ & new_new_n18570__;
  assign new_new_n18572__ = ~new_new_n18568__ & ~new_new_n18571__;
  assign new_new_n18573__ = ~pi066 & new_new_n18572__;
  assign new_new_n18574__ = pi066 & ~new_new_n18572__;
  assign new_new_n18575__ = new_new_n426__ & ~po009;
  assign new_new_n18576__ = ~pi065 & po008;
  assign new_new_n18577__ = po009 & new_new_n18576__;
  assign new_new_n18578__ = ~new_new_n18575__ & ~new_new_n18577__;
  assign new_new_n18579__ = ~pi008 & ~new_new_n18578__;
  assign new_new_n18580__ = ~new_new_n332__ & po008;
  assign new_new_n18581__ = ~new_new_n17939__ & ~new_new_n18580__;
  assign new_new_n18582__ = pi065 & po008;
  assign new_new_n18583__ = po009 & ~new_new_n18582__;
  assign new_new_n18584__ = pi065 & ~new_new_n17939__;
  assign new_new_n18585__ = pi008 & ~new_new_n18584__;
  assign new_new_n18586__ = ~new_new_n18583__ & new_new_n18585__;
  assign new_new_n18587__ = ~new_new_n18581__ & ~new_new_n18586__;
  assign new_new_n18588__ = ~new_new_n18579__ & new_new_n18587__;
  assign new_new_n18589__ = pi009 & ~new_new_n18588__;
  assign new_new_n18590__ = ~new_new_n17939__ & ~new_new_n18582__;
  assign new_new_n18591__ = pi008 & ~new_new_n17949__;
  assign new_new_n18592__ = pi064 & ~new_new_n18591__;
  assign new_new_n18593__ = ~new_new_n18590__ & ~new_new_n18592__;
  assign new_new_n18594__ = ~po009 & ~new_new_n18576__;
  assign new_new_n18595__ = pi064 & ~new_new_n18561__;
  assign new_new_n18596__ = ~new_new_n18577__ & new_new_n18595__;
  assign new_new_n18597__ = ~new_new_n18594__ & new_new_n18596__;
  assign new_new_n18598__ = ~new_new_n18593__ & ~new_new_n18597__;
  assign new_new_n18599__ = ~pi009 & ~new_new_n18598__;
  assign new_new_n18600__ = ~new_new_n18589__ & ~new_new_n18599__;
  assign new_new_n18601__ = ~new_new_n18574__ & ~new_new_n18600__;
  assign new_new_n18602__ = ~new_new_n18573__ & ~new_new_n18601__;
  assign new_new_n18603__ = ~new_new_n18560__ & ~new_new_n18602__;
  assign new_new_n18604__ = ~new_new_n18559__ & ~new_new_n18603__;
  assign new_new_n18605__ = ~new_new_n18553__ & ~new_new_n18604__;
  assign new_new_n18606__ = ~new_new_n18552__ & ~new_new_n18605__;
  assign new_new_n18607__ = ~new_new_n18544__ & ~new_new_n18606__;
  assign new_new_n18608__ = ~new_new_n18543__ & ~new_new_n18607__;
  assign new_new_n18609__ = ~new_new_n18537__ & ~new_new_n18608__;
  assign new_new_n18610__ = ~new_new_n18536__ & ~new_new_n18609__;
  assign new_new_n18611__ = ~new_new_n18528__ & ~new_new_n18610__;
  assign new_new_n18612__ = ~new_new_n18527__ & ~new_new_n18611__;
  assign new_new_n18613__ = ~new_new_n18519__ & new_new_n18612__;
  assign new_new_n18614__ = ~new_new_n18518__ & ~new_new_n18613__;
  assign new_new_n18615__ = ~new_new_n18510__ & ~new_new_n18614__;
  assign new_new_n18616__ = ~new_new_n18509__ & ~new_new_n18615__;
  assign new_new_n18617__ = ~new_new_n18501__ & ~new_new_n18616__;
  assign new_new_n18618__ = ~new_new_n18500__ & ~new_new_n18617__;
  assign new_new_n18619__ = ~new_new_n18492__ & new_new_n18618__;
  assign new_new_n18620__ = ~new_new_n18491__ & ~new_new_n18619__;
  assign new_new_n18621__ = ~new_new_n18483__ & ~new_new_n18620__;
  assign new_new_n18622__ = ~new_new_n18482__ & ~new_new_n18621__;
  assign new_new_n18623__ = ~new_new_n18474__ & ~new_new_n18622__;
  assign new_new_n18624__ = ~new_new_n18473__ & ~new_new_n18623__;
  assign new_new_n18625__ = ~new_new_n18465__ & ~new_new_n18624__;
  assign new_new_n18626__ = ~new_new_n18464__ & ~new_new_n18625__;
  assign new_new_n18627__ = ~new_new_n18456__ & ~new_new_n18626__;
  assign new_new_n18628__ = ~new_new_n18455__ & ~new_new_n18627__;
  assign new_new_n18629__ = ~new_new_n18447__ & new_new_n18628__;
  assign new_new_n18630__ = ~new_new_n18446__ & ~new_new_n18629__;
  assign new_new_n18631__ = ~new_new_n18438__ & ~new_new_n18630__;
  assign new_new_n18632__ = ~new_new_n18437__ & ~new_new_n18631__;
  assign new_new_n18633__ = ~new_new_n18429__ & ~new_new_n18632__;
  assign new_new_n18634__ = ~new_new_n18428__ & ~new_new_n18633__;
  assign new_new_n18635__ = ~new_new_n18420__ & new_new_n18634__;
  assign new_new_n18636__ = ~new_new_n18419__ & ~new_new_n18635__;
  assign new_new_n18637__ = ~new_new_n18411__ & ~new_new_n18636__;
  assign new_new_n18638__ = ~new_new_n18410__ & ~new_new_n18637__;
  assign new_new_n18639__ = ~new_new_n18402__ & ~new_new_n18638__;
  assign new_new_n18640__ = ~new_new_n18401__ & ~new_new_n18639__;
  assign new_new_n18641__ = ~new_new_n18393__ & ~new_new_n18640__;
  assign new_new_n18642__ = ~new_new_n18392__ & ~new_new_n18641__;
  assign new_new_n18643__ = ~new_new_n18384__ & new_new_n18642__;
  assign new_new_n18644__ = ~new_new_n18383__ & ~new_new_n18643__;
  assign new_new_n18645__ = ~new_new_n18375__ & ~new_new_n18644__;
  assign new_new_n18646__ = ~new_new_n18374__ & ~new_new_n18645__;
  assign new_new_n18647__ = ~new_new_n18366__ & ~new_new_n18646__;
  assign new_new_n18648__ = ~new_new_n18365__ & ~new_new_n18647__;
  assign new_new_n18649__ = ~new_new_n18357__ & new_new_n18648__;
  assign new_new_n18650__ = ~new_new_n18356__ & ~new_new_n18649__;
  assign new_new_n18651__ = ~new_new_n18348__ & ~new_new_n18650__;
  assign new_new_n18652__ = ~new_new_n18347__ & ~new_new_n18651__;
  assign new_new_n18653__ = ~new_new_n18339__ & ~new_new_n18652__;
  assign new_new_n18654__ = ~new_new_n18338__ & ~new_new_n18653__;
  assign new_new_n18655__ = ~new_new_n18330__ & new_new_n18654__;
  assign new_new_n18656__ = ~new_new_n18329__ & ~new_new_n18655__;
  assign new_new_n18657__ = ~new_new_n18321__ & ~new_new_n18656__;
  assign new_new_n18658__ = ~new_new_n18320__ & ~new_new_n18657__;
  assign new_new_n18659__ = ~new_new_n18312__ & ~new_new_n18658__;
  assign new_new_n18660__ = ~new_new_n18311__ & ~new_new_n18659__;
  assign new_new_n18661__ = ~new_new_n18303__ & new_new_n18660__;
  assign new_new_n18662__ = ~new_new_n18302__ & ~new_new_n18661__;
  assign new_new_n18663__ = ~new_new_n18294__ & ~new_new_n18662__;
  assign new_new_n18664__ = ~new_new_n18293__ & ~new_new_n18663__;
  assign new_new_n18665__ = ~new_new_n18285__ & new_new_n18664__;
  assign new_new_n18666__ = ~new_new_n18284__ & ~new_new_n18665__;
  assign new_new_n18667__ = ~new_new_n18276__ & ~new_new_n18666__;
  assign new_new_n18668__ = ~new_new_n18275__ & ~new_new_n18667__;
  assign new_new_n18669__ = ~new_new_n18267__ & ~new_new_n18668__;
  assign new_new_n18670__ = ~new_new_n18266__ & ~new_new_n18669__;
  assign new_new_n18671__ = ~new_new_n18258__ & ~new_new_n18670__;
  assign new_new_n18672__ = ~new_new_n18257__ & ~new_new_n18671__;
  assign new_new_n18673__ = ~new_new_n18249__ & new_new_n18672__;
  assign new_new_n18674__ = ~new_new_n18248__ & ~new_new_n18673__;
  assign new_new_n18675__ = ~new_new_n18240__ & ~new_new_n18674__;
  assign new_new_n18676__ = ~new_new_n18239__ & ~new_new_n18675__;
  assign new_new_n18677__ = ~new_new_n18231__ & new_new_n18676__;
  assign new_new_n18678__ = ~new_new_n18230__ & ~new_new_n18677__;
  assign new_new_n18679__ = ~new_new_n18222__ & ~new_new_n18678__;
  assign new_new_n18680__ = ~new_new_n18221__ & ~new_new_n18679__;
  assign new_new_n18681__ = ~new_new_n18213__ & new_new_n18680__;
  assign new_new_n18682__ = ~new_new_n18212__ & ~new_new_n18681__;
  assign new_new_n18683__ = ~new_new_n18204__ & ~new_new_n18682__;
  assign new_new_n18684__ = ~new_new_n18203__ & ~new_new_n18683__;
  assign new_new_n18685__ = ~new_new_n18195__ & ~new_new_n18684__;
  assign new_new_n18686__ = ~new_new_n18194__ & ~new_new_n18685__;
  assign new_new_n18687__ = ~new_new_n18186__ & new_new_n18686__;
  assign new_new_n18688__ = ~new_new_n18185__ & ~new_new_n18687__;
  assign new_new_n18689__ = ~new_new_n18177__ & ~new_new_n18688__;
  assign new_new_n18690__ = ~new_new_n18176__ & ~new_new_n18689__;
  assign new_new_n18691__ = ~new_new_n18168__ & new_new_n18690__;
  assign new_new_n18692__ = ~new_new_n18167__ & ~new_new_n18691__;
  assign new_new_n18693__ = ~new_new_n18159__ & ~new_new_n18692__;
  assign new_new_n18694__ = ~new_new_n18158__ & ~new_new_n18693__;
  assign new_new_n18695__ = ~new_new_n18150__ & ~new_new_n18694__;
  assign new_new_n18696__ = ~new_new_n18149__ & ~new_new_n18695__;
  assign new_new_n18697__ = ~new_new_n18141__ & ~new_new_n18696__;
  assign new_new_n18698__ = ~new_new_n18140__ & ~new_new_n18697__;
  assign new_new_n18699__ = ~new_new_n18132__ & ~new_new_n18698__;
  assign new_new_n18700__ = ~new_new_n18131__ & ~new_new_n18699__;
  assign new_new_n18701__ = ~new_new_n18123__ & new_new_n18700__;
  assign new_new_n18702__ = ~new_new_n18122__ & ~new_new_n18701__;
  assign new_new_n18703__ = ~new_new_n18114__ & new_new_n18702__;
  assign new_new_n18704__ = ~new_new_n18113__ & ~new_new_n18703__;
  assign new_new_n18705__ = ~new_new_n18105__ & ~new_new_n18704__;
  assign new_new_n18706__ = ~new_new_n18104__ & ~new_new_n18705__;
  assign new_new_n18707__ = ~new_new_n18096__ & new_new_n18706__;
  assign new_new_n18708__ = ~new_new_n18095__ & ~new_new_n18707__;
  assign new_new_n18709__ = pi120 & ~new_new_n18708__;
  assign new_new_n18710__ = ~pi119 & new_new_n18084__;
  assign new_new_n18711__ = pi119 & ~new_new_n18084__;
  assign new_new_n18712__ = ~new_new_n18710__ & ~new_new_n18711__;
  assign new_new_n18713__ = ~pi120 & new_new_n18712__;
  assign new_new_n18714__ = new_new_n18708__ & new_new_n18713__;
  assign new_new_n18715__ = new_new_n16825__ & ~new_new_n18709__;
  assign new_new_n18716__ = ~new_new_n18714__ & new_new_n18715__;
  assign new_new_n18717__ = new_new_n17442__ & ~new_new_n18716__;
  assign new_new_n18718__ = ~new_new_n18095__ & ~new_new_n18096__;
  assign new_new_n18719__ = new_new_n16826__ & ~new_new_n18712__;
  assign new_new_n18720__ = new_new_n17442__ & ~new_new_n18719__;
  assign new_new_n18721__ = ~pi120 & new_new_n18720__;
  assign new_new_n18722__ = pi120 & ~new_new_n16837__;
  assign new_new_n18723__ = new_new_n18708__ & ~new_new_n18722__;
  assign new_new_n18724__ = ~new_new_n18721__ & ~new_new_n18723__;
  assign po007 = new_new_n16825__ & ~new_new_n18724__;
  assign new_new_n18726__ = ~new_new_n18706__ & po007;
  assign new_new_n18727__ = ~pi119 & ~po007;
  assign new_new_n18728__ = ~new_new_n18726__ & ~new_new_n18727__;
  assign new_new_n18729__ = new_new_n18718__ & new_new_n18728__;
  assign new_new_n18730__ = ~new_new_n18718__ & ~new_new_n18728__;
  assign new_new_n18731__ = ~new_new_n18729__ & ~new_new_n18730__;
  assign new_new_n18732__ = pi120 & new_new_n18731__;
  assign new_new_n18733__ = ~pi120 & ~new_new_n18731__;
  assign new_new_n18734__ = new_new_n18704__ & po007;
  assign new_new_n18735__ = pi118 & ~po007;
  assign new_new_n18736__ = ~new_new_n18734__ & ~new_new_n18735__;
  assign new_new_n18737__ = ~new_new_n18104__ & ~new_new_n18105__;
  assign new_new_n18738__ = ~new_new_n18736__ & ~new_new_n18737__;
  assign new_new_n18739__ = new_new_n18736__ & new_new_n18737__;
  assign new_new_n18740__ = ~new_new_n18738__ & ~new_new_n18739__;
  assign new_new_n18741__ = pi119 & ~new_new_n18740__;
  assign new_new_n18742__ = ~pi119 & new_new_n18740__;
  assign new_new_n18743__ = new_new_n18702__ & po007;
  assign new_new_n18744__ = ~pi117 & ~po007;
  assign new_new_n18745__ = ~new_new_n18743__ & ~new_new_n18744__;
  assign new_new_n18746__ = ~new_new_n18113__ & ~new_new_n18114__;
  assign new_new_n18747__ = ~new_new_n18745__ & ~new_new_n18746__;
  assign new_new_n18748__ = new_new_n18745__ & new_new_n18746__;
  assign new_new_n18749__ = ~new_new_n18747__ & ~new_new_n18748__;
  assign new_new_n18750__ = ~pi118 & ~new_new_n18749__;
  assign new_new_n18751__ = pi118 & new_new_n18749__;
  assign new_new_n18752__ = new_new_n18700__ & po007;
  assign new_new_n18753__ = pi116 & ~po007;
  assign new_new_n18754__ = ~new_new_n18752__ & ~new_new_n18753__;
  assign new_new_n18755__ = ~new_new_n18122__ & ~new_new_n18123__;
  assign new_new_n18756__ = ~new_new_n18754__ & ~new_new_n18755__;
  assign new_new_n18757__ = new_new_n18754__ & new_new_n18755__;
  assign new_new_n18758__ = ~new_new_n18756__ & ~new_new_n18757__;
  assign new_new_n18759__ = pi117 & ~new_new_n18758__;
  assign new_new_n18760__ = ~pi117 & new_new_n18758__;
  assign new_new_n18761__ = ~new_new_n18131__ & ~new_new_n18132__;
  assign new_new_n18762__ = ~new_new_n18698__ & po007;
  assign new_new_n18763__ = ~pi115 & ~po007;
  assign new_new_n18764__ = ~new_new_n18762__ & ~new_new_n18763__;
  assign new_new_n18765__ = new_new_n18761__ & ~new_new_n18764__;
  assign new_new_n18766__ = ~new_new_n18761__ & new_new_n18764__;
  assign new_new_n18767__ = ~new_new_n18765__ & ~new_new_n18766__;
  assign new_new_n18768__ = pi116 & ~new_new_n18767__;
  assign new_new_n18769__ = ~pi116 & new_new_n18767__;
  assign new_new_n18770__ = ~new_new_n18140__ & ~new_new_n18141__;
  assign new_new_n18771__ = ~new_new_n18696__ & po007;
  assign new_new_n18772__ = ~pi114 & ~po007;
  assign new_new_n18773__ = ~new_new_n18771__ & ~new_new_n18772__;
  assign new_new_n18774__ = new_new_n18770__ & ~new_new_n18773__;
  assign new_new_n18775__ = ~new_new_n18770__ & new_new_n18773__;
  assign new_new_n18776__ = ~new_new_n18774__ & ~new_new_n18775__;
  assign new_new_n18777__ = pi115 & ~new_new_n18776__;
  assign new_new_n18778__ = ~pi115 & new_new_n18776__;
  assign new_new_n18779__ = ~pi113 & ~new_new_n18694__;
  assign new_new_n18780__ = pi113 & new_new_n18694__;
  assign new_new_n18781__ = ~new_new_n18779__ & ~new_new_n18780__;
  assign new_new_n18782__ = po007 & new_new_n18781__;
  assign new_new_n18783__ = ~new_new_n18148__ & new_new_n18782__;
  assign new_new_n18784__ = new_new_n18148__ & ~new_new_n18782__;
  assign new_new_n18785__ = ~new_new_n18783__ & ~new_new_n18784__;
  assign new_new_n18786__ = pi114 & ~new_new_n18785__;
  assign new_new_n18787__ = ~pi114 & new_new_n18785__;
  assign new_new_n18788__ = ~new_new_n18158__ & ~new_new_n18159__;
  assign new_new_n18789__ = ~new_new_n18692__ & po007;
  assign new_new_n18790__ = ~pi112 & ~po007;
  assign new_new_n18791__ = ~new_new_n18789__ & ~new_new_n18790__;
  assign new_new_n18792__ = new_new_n18788__ & ~new_new_n18791__;
  assign new_new_n18793__ = ~new_new_n18788__ & new_new_n18791__;
  assign new_new_n18794__ = ~new_new_n18792__ & ~new_new_n18793__;
  assign new_new_n18795__ = ~pi113 & new_new_n18794__;
  assign new_new_n18796__ = pi113 & ~new_new_n18794__;
  assign new_new_n18797__ = ~new_new_n18690__ & po007;
  assign new_new_n18798__ = pi111 & ~po007;
  assign new_new_n18799__ = ~new_new_n18797__ & ~new_new_n18798__;
  assign new_new_n18800__ = ~new_new_n18167__ & ~new_new_n18168__;
  assign new_new_n18801__ = ~new_new_n18799__ & new_new_n18800__;
  assign new_new_n18802__ = new_new_n18799__ & ~new_new_n18800__;
  assign new_new_n18803__ = ~new_new_n18801__ & ~new_new_n18802__;
  assign new_new_n18804__ = ~pi112 & ~new_new_n18803__;
  assign new_new_n18805__ = pi112 & new_new_n18803__;
  assign new_new_n18806__ = pi110 & ~new_new_n18688__;
  assign new_new_n18807__ = ~pi110 & new_new_n18688__;
  assign new_new_n18808__ = ~new_new_n18806__ & ~new_new_n18807__;
  assign new_new_n18809__ = po007 & new_new_n18808__;
  assign new_new_n18810__ = new_new_n18175__ & new_new_n18809__;
  assign new_new_n18811__ = ~new_new_n18175__ & ~new_new_n18809__;
  assign new_new_n18812__ = ~new_new_n18810__ & ~new_new_n18811__;
  assign new_new_n18813__ = pi111 & ~new_new_n18812__;
  assign new_new_n18814__ = ~pi111 & new_new_n18812__;
  assign new_new_n18815__ = ~new_new_n18194__ & ~new_new_n18195__;
  assign new_new_n18816__ = ~new_new_n18684__ & po007;
  assign new_new_n18817__ = ~pi108 & ~po007;
  assign new_new_n18818__ = ~new_new_n18816__ & ~new_new_n18817__;
  assign new_new_n18819__ = new_new_n18815__ & ~new_new_n18818__;
  assign new_new_n18820__ = ~new_new_n18815__ & new_new_n18818__;
  assign new_new_n18821__ = ~new_new_n18819__ & ~new_new_n18820__;
  assign new_new_n18822__ = ~pi109 & new_new_n18821__;
  assign new_new_n18823__ = pi109 & ~new_new_n18821__;
  assign new_new_n18824__ = ~new_new_n18203__ & ~new_new_n18204__;
  assign new_new_n18825__ = ~new_new_n18682__ & po007;
  assign new_new_n18826__ = ~pi107 & ~po007;
  assign new_new_n18827__ = ~new_new_n18825__ & ~new_new_n18826__;
  assign new_new_n18828__ = new_new_n18824__ & ~new_new_n18827__;
  assign new_new_n18829__ = ~new_new_n18824__ & new_new_n18827__;
  assign new_new_n18830__ = ~new_new_n18828__ & ~new_new_n18829__;
  assign new_new_n18831__ = ~pi108 & new_new_n18830__;
  assign new_new_n18832__ = pi108 & ~new_new_n18830__;
  assign new_new_n18833__ = ~new_new_n18680__ & po007;
  assign new_new_n18834__ = pi106 & ~po007;
  assign new_new_n18835__ = ~new_new_n18833__ & ~new_new_n18834__;
  assign new_new_n18836__ = ~new_new_n18212__ & ~new_new_n18213__;
  assign new_new_n18837__ = ~new_new_n18835__ & new_new_n18836__;
  assign new_new_n18838__ = new_new_n18835__ & ~new_new_n18836__;
  assign new_new_n18839__ = ~new_new_n18837__ & ~new_new_n18838__;
  assign new_new_n18840__ = ~pi107 & ~new_new_n18839__;
  assign new_new_n18841__ = pi107 & new_new_n18839__;
  assign new_new_n18842__ = ~new_new_n18221__ & ~new_new_n18222__;
  assign new_new_n18843__ = ~new_new_n18678__ & po007;
  assign new_new_n18844__ = pi105 & ~po007;
  assign new_new_n18845__ = ~new_new_n18843__ & ~new_new_n18844__;
  assign new_new_n18846__ = new_new_n18842__ & ~new_new_n18845__;
  assign new_new_n18847__ = ~new_new_n18842__ & new_new_n18845__;
  assign new_new_n18848__ = ~new_new_n18846__ & ~new_new_n18847__;
  assign new_new_n18849__ = ~pi106 & ~new_new_n18848__;
  assign new_new_n18850__ = pi106 & new_new_n18848__;
  assign new_new_n18851__ = ~new_new_n18230__ & ~new_new_n18231__;
  assign new_new_n18852__ = ~new_new_n18676__ & po007;
  assign new_new_n18853__ = ~pi104 & ~po007;
  assign new_new_n18854__ = ~new_new_n18852__ & ~new_new_n18853__;
  assign new_new_n18855__ = new_new_n18851__ & ~new_new_n18854__;
  assign new_new_n18856__ = ~new_new_n18851__ & new_new_n18854__;
  assign new_new_n18857__ = ~new_new_n18855__ & ~new_new_n18856__;
  assign new_new_n18858__ = ~pi105 & new_new_n18857__;
  assign new_new_n18859__ = pi105 & ~new_new_n18857__;
  assign new_new_n18860__ = ~pi103 & ~new_new_n18674__;
  assign new_new_n18861__ = pi103 & new_new_n18674__;
  assign new_new_n18862__ = ~new_new_n18860__ & ~new_new_n18861__;
  assign new_new_n18863__ = po007 & new_new_n18862__;
  assign new_new_n18864__ = new_new_n18238__ & new_new_n18863__;
  assign new_new_n18865__ = ~new_new_n18238__ & ~new_new_n18863__;
  assign new_new_n18866__ = ~new_new_n18864__ & ~new_new_n18865__;
  assign new_new_n18867__ = ~pi104 & ~new_new_n18866__;
  assign new_new_n18868__ = pi104 & new_new_n18866__;
  assign new_new_n18869__ = ~new_new_n18248__ & ~new_new_n18249__;
  assign new_new_n18870__ = ~new_new_n18672__ & po007;
  assign new_new_n18871__ = pi102 & ~po007;
  assign new_new_n18872__ = ~new_new_n18870__ & ~new_new_n18871__;
  assign new_new_n18873__ = new_new_n18869__ & ~new_new_n18872__;
  assign new_new_n18874__ = ~new_new_n18869__ & new_new_n18872__;
  assign new_new_n18875__ = ~new_new_n18873__ & ~new_new_n18874__;
  assign new_new_n18876__ = ~pi103 & ~new_new_n18875__;
  assign new_new_n18877__ = pi103 & new_new_n18875__;
  assign new_new_n18878__ = ~new_new_n18670__ & po007;
  assign new_new_n18879__ = pi101 & ~po007;
  assign new_new_n18880__ = ~new_new_n18878__ & ~new_new_n18879__;
  assign new_new_n18881__ = ~new_new_n18257__ & ~new_new_n18258__;
  assign new_new_n18882__ = ~new_new_n18880__ & new_new_n18881__;
  assign new_new_n18883__ = new_new_n18880__ & ~new_new_n18881__;
  assign new_new_n18884__ = ~new_new_n18882__ & ~new_new_n18883__;
  assign new_new_n18885__ = ~pi102 & ~new_new_n18884__;
  assign new_new_n18886__ = pi102 & new_new_n18884__;
  assign new_new_n18887__ = ~new_new_n18266__ & ~new_new_n18267__;
  assign new_new_n18888__ = ~new_new_n18668__ & po007;
  assign new_new_n18889__ = pi100 & ~po007;
  assign new_new_n18890__ = ~new_new_n18888__ & ~new_new_n18889__;
  assign new_new_n18891__ = new_new_n18887__ & new_new_n18890__;
  assign new_new_n18892__ = ~new_new_n18887__ & ~new_new_n18890__;
  assign new_new_n18893__ = ~new_new_n18891__ & ~new_new_n18892__;
  assign new_new_n18894__ = pi101 & ~new_new_n18893__;
  assign new_new_n18895__ = ~pi101 & new_new_n18893__;
  assign new_new_n18896__ = new_new_n18666__ & po007;
  assign new_new_n18897__ = ~pi099 & ~po007;
  assign new_new_n18898__ = ~new_new_n18896__ & ~new_new_n18897__;
  assign new_new_n18899__ = ~new_new_n18275__ & ~new_new_n18276__;
  assign new_new_n18900__ = ~new_new_n18898__ & ~new_new_n18899__;
  assign new_new_n18901__ = new_new_n18898__ & new_new_n18899__;
  assign new_new_n18902__ = ~new_new_n18900__ & ~new_new_n18901__;
  assign new_new_n18903__ = ~pi100 & ~new_new_n18902__;
  assign new_new_n18904__ = pi100 & new_new_n18902__;
  assign new_new_n18905__ = new_new_n18664__ & po007;
  assign new_new_n18906__ = pi098 & ~po007;
  assign new_new_n18907__ = ~new_new_n18905__ & ~new_new_n18906__;
  assign new_new_n18908__ = ~new_new_n18284__ & ~new_new_n18285__;
  assign new_new_n18909__ = ~new_new_n18907__ & ~new_new_n18908__;
  assign new_new_n18910__ = new_new_n18907__ & new_new_n18908__;
  assign new_new_n18911__ = ~new_new_n18909__ & ~new_new_n18910__;
  assign new_new_n18912__ = pi099 & ~new_new_n18911__;
  assign new_new_n18913__ = ~pi099 & new_new_n18911__;
  assign new_new_n18914__ = ~new_new_n18293__ & ~new_new_n18294__;
  assign new_new_n18915__ = ~new_new_n18662__ & po007;
  assign new_new_n18916__ = ~pi097 & ~po007;
  assign new_new_n18917__ = ~new_new_n18915__ & ~new_new_n18916__;
  assign new_new_n18918__ = ~new_new_n18914__ & ~new_new_n18917__;
  assign new_new_n18919__ = new_new_n18914__ & new_new_n18917__;
  assign new_new_n18920__ = ~new_new_n18918__ & ~new_new_n18919__;
  assign new_new_n18921__ = ~pi098 & ~new_new_n18920__;
  assign new_new_n18922__ = pi098 & new_new_n18920__;
  assign new_new_n18923__ = new_new_n18660__ & po007;
  assign new_new_n18924__ = ~pi096 & ~po007;
  assign new_new_n18925__ = ~new_new_n18923__ & ~new_new_n18924__;
  assign new_new_n18926__ = ~new_new_n18302__ & ~new_new_n18303__;
  assign new_new_n18927__ = ~new_new_n18925__ & ~new_new_n18926__;
  assign new_new_n18928__ = new_new_n18925__ & new_new_n18926__;
  assign new_new_n18929__ = ~new_new_n18927__ & ~new_new_n18928__;
  assign new_new_n18930__ = ~pi097 & ~new_new_n18929__;
  assign new_new_n18931__ = pi097 & new_new_n18929__;
  assign new_new_n18932__ = ~new_new_n18311__ & ~new_new_n18312__;
  assign new_new_n18933__ = ~new_new_n18658__ & po007;
  assign new_new_n18934__ = pi095 & ~po007;
  assign new_new_n18935__ = ~new_new_n18933__ & ~new_new_n18934__;
  assign new_new_n18936__ = new_new_n18932__ & ~new_new_n18935__;
  assign new_new_n18937__ = ~new_new_n18932__ & new_new_n18935__;
  assign new_new_n18938__ = ~new_new_n18936__ & ~new_new_n18937__;
  assign new_new_n18939__ = pi096 & new_new_n18938__;
  assign new_new_n18940__ = ~pi096 & ~new_new_n18938__;
  assign new_new_n18941__ = pi094 & ~new_new_n18656__;
  assign new_new_n18942__ = ~pi094 & new_new_n18656__;
  assign new_new_n18943__ = ~new_new_n18941__ & ~new_new_n18942__;
  assign new_new_n18944__ = po007 & new_new_n18943__;
  assign new_new_n18945__ = new_new_n18319__ & new_new_n18944__;
  assign new_new_n18946__ = ~new_new_n18319__ & ~new_new_n18944__;
  assign new_new_n18947__ = ~new_new_n18945__ & ~new_new_n18946__;
  assign new_new_n18948__ = pi095 & ~new_new_n18947__;
  assign new_new_n18949__ = ~pi095 & new_new_n18947__;
  assign new_new_n18950__ = ~new_new_n18329__ & ~new_new_n18330__;
  assign new_new_n18951__ = ~new_new_n18654__ & po007;
  assign new_new_n18952__ = ~pi093 & ~po007;
  assign new_new_n18953__ = ~new_new_n18951__ & ~new_new_n18952__;
  assign new_new_n18954__ = new_new_n18950__ & ~new_new_n18953__;
  assign new_new_n18955__ = ~new_new_n18950__ & new_new_n18953__;
  assign new_new_n18956__ = ~new_new_n18954__ & ~new_new_n18955__;
  assign new_new_n18957__ = pi094 & ~new_new_n18956__;
  assign new_new_n18958__ = ~pi094 & new_new_n18956__;
  assign new_new_n18959__ = ~new_new_n18338__ & ~new_new_n18339__;
  assign new_new_n18960__ = ~new_new_n18652__ & po007;
  assign new_new_n18961__ = ~pi092 & ~po007;
  assign new_new_n18962__ = ~new_new_n18960__ & ~new_new_n18961__;
  assign new_new_n18963__ = new_new_n18959__ & ~new_new_n18962__;
  assign new_new_n18964__ = ~new_new_n18959__ & new_new_n18962__;
  assign new_new_n18965__ = ~new_new_n18963__ & ~new_new_n18964__;
  assign new_new_n18966__ = pi093 & ~new_new_n18965__;
  assign new_new_n18967__ = ~pi093 & new_new_n18965__;
  assign new_new_n18968__ = ~pi091 & ~new_new_n18650__;
  assign new_new_n18969__ = pi091 & new_new_n18650__;
  assign new_new_n18970__ = ~new_new_n18968__ & ~new_new_n18969__;
  assign new_new_n18971__ = po007 & new_new_n18970__;
  assign new_new_n18972__ = new_new_n18346__ & new_new_n18971__;
  assign new_new_n18973__ = ~new_new_n18346__ & ~new_new_n18971__;
  assign new_new_n18974__ = ~new_new_n18972__ & ~new_new_n18973__;
  assign new_new_n18975__ = ~pi092 & ~new_new_n18974__;
  assign new_new_n18976__ = pi092 & new_new_n18974__;
  assign new_new_n18977__ = ~new_new_n18648__ & po007;
  assign new_new_n18978__ = pi090 & ~po007;
  assign new_new_n18979__ = ~new_new_n18977__ & ~new_new_n18978__;
  assign new_new_n18980__ = ~new_new_n18356__ & ~new_new_n18357__;
  assign new_new_n18981__ = ~new_new_n18979__ & new_new_n18980__;
  assign new_new_n18982__ = new_new_n18979__ & ~new_new_n18980__;
  assign new_new_n18983__ = ~new_new_n18981__ & ~new_new_n18982__;
  assign new_new_n18984__ = pi091 & new_new_n18983__;
  assign new_new_n18985__ = ~pi091 & ~new_new_n18983__;
  assign new_new_n18986__ = ~new_new_n18365__ & ~new_new_n18366__;
  assign new_new_n18987__ = ~new_new_n18646__ & po007;
  assign new_new_n18988__ = pi089 & ~po007;
  assign new_new_n18989__ = ~new_new_n18987__ & ~new_new_n18988__;
  assign new_new_n18990__ = new_new_n18986__ & new_new_n18989__;
  assign new_new_n18991__ = ~new_new_n18986__ & ~new_new_n18989__;
  assign new_new_n18992__ = ~new_new_n18990__ & ~new_new_n18991__;
  assign new_new_n18993__ = pi090 & ~new_new_n18992__;
  assign new_new_n18994__ = ~pi090 & new_new_n18992__;
  assign new_new_n18995__ = pi088 & ~new_new_n18644__;
  assign new_new_n18996__ = ~pi088 & new_new_n18644__;
  assign new_new_n18997__ = ~new_new_n18995__ & ~new_new_n18996__;
  assign new_new_n18998__ = po007 & new_new_n18997__;
  assign new_new_n18999__ = new_new_n18373__ & new_new_n18998__;
  assign new_new_n19000__ = ~new_new_n18373__ & ~new_new_n18998__;
  assign new_new_n19001__ = ~new_new_n18999__ & ~new_new_n19000__;
  assign new_new_n19002__ = pi089 & ~new_new_n19001__;
  assign new_new_n19003__ = ~pi089 & new_new_n19001__;
  assign new_new_n19004__ = ~new_new_n18383__ & ~new_new_n18384__;
  assign new_new_n19005__ = ~new_new_n18642__ & po007;
  assign new_new_n19006__ = ~pi087 & ~po007;
  assign new_new_n19007__ = ~new_new_n19005__ & ~new_new_n19006__;
  assign new_new_n19008__ = new_new_n19004__ & ~new_new_n19007__;
  assign new_new_n19009__ = ~new_new_n19004__ & new_new_n19007__;
  assign new_new_n19010__ = ~new_new_n19008__ & ~new_new_n19009__;
  assign new_new_n19011__ = pi088 & ~new_new_n19010__;
  assign new_new_n19012__ = ~pi088 & new_new_n19010__;
  assign new_new_n19013__ = ~pi086 & ~new_new_n18640__;
  assign new_new_n19014__ = pi086 & new_new_n18640__;
  assign new_new_n19015__ = ~new_new_n19013__ & ~new_new_n19014__;
  assign new_new_n19016__ = po007 & new_new_n19015__;
  assign new_new_n19017__ = new_new_n18391__ & new_new_n19016__;
  assign new_new_n19018__ = ~new_new_n18391__ & ~new_new_n19016__;
  assign new_new_n19019__ = ~new_new_n19017__ & ~new_new_n19018__;
  assign new_new_n19020__ = pi087 & new_new_n19019__;
  assign new_new_n19021__ = ~pi087 & ~new_new_n19019__;
  assign new_new_n19022__ = ~new_new_n18401__ & ~new_new_n18402__;
  assign new_new_n19023__ = ~new_new_n18638__ & po007;
  assign new_new_n19024__ = ~pi085 & ~po007;
  assign new_new_n19025__ = ~new_new_n19023__ & ~new_new_n19024__;
  assign new_new_n19026__ = new_new_n19022__ & ~new_new_n19025__;
  assign new_new_n19027__ = ~new_new_n19022__ & new_new_n19025__;
  assign new_new_n19028__ = ~new_new_n19026__ & ~new_new_n19027__;
  assign new_new_n19029__ = pi086 & ~new_new_n19028__;
  assign new_new_n19030__ = ~pi086 & new_new_n19028__;
  assign new_new_n19031__ = ~pi084 & ~new_new_n18636__;
  assign new_new_n19032__ = pi084 & new_new_n18636__;
  assign new_new_n19033__ = ~new_new_n19031__ & ~new_new_n19032__;
  assign new_new_n19034__ = po007 & new_new_n19033__;
  assign new_new_n19035__ = ~new_new_n18409__ & ~new_new_n19034__;
  assign new_new_n19036__ = new_new_n18409__ & new_new_n19034__;
  assign new_new_n19037__ = ~new_new_n19035__ & ~new_new_n19036__;
  assign new_new_n19038__ = ~pi085 & ~new_new_n19037__;
  assign new_new_n19039__ = pi085 & new_new_n19037__;
  assign new_new_n19040__ = ~new_new_n18419__ & ~new_new_n18420__;
  assign new_new_n19041__ = ~new_new_n18634__ & po007;
  assign new_new_n19042__ = pi083 & ~po007;
  assign new_new_n19043__ = ~new_new_n19041__ & ~new_new_n19042__;
  assign new_new_n19044__ = new_new_n19040__ & ~new_new_n19043__;
  assign new_new_n19045__ = ~new_new_n19040__ & new_new_n19043__;
  assign new_new_n19046__ = ~new_new_n19044__ & ~new_new_n19045__;
  assign new_new_n19047__ = pi084 & new_new_n19046__;
  assign new_new_n19048__ = ~pi084 & ~new_new_n19046__;
  assign new_new_n19049__ = ~new_new_n18632__ & po007;
  assign new_new_n19050__ = pi082 & ~po007;
  assign new_new_n19051__ = ~new_new_n19049__ & ~new_new_n19050__;
  assign new_new_n19052__ = ~new_new_n18428__ & ~new_new_n18429__;
  assign new_new_n19053__ = ~new_new_n19051__ & new_new_n19052__;
  assign new_new_n19054__ = new_new_n19051__ & ~new_new_n19052__;
  assign new_new_n19055__ = ~new_new_n19053__ & ~new_new_n19054__;
  assign new_new_n19056__ = pi083 & new_new_n19055__;
  assign new_new_n19057__ = ~pi083 & ~new_new_n19055__;
  assign new_new_n19058__ = ~new_new_n18437__ & ~new_new_n18438__;
  assign new_new_n19059__ = ~new_new_n18630__ & po007;
  assign new_new_n19060__ = pi081 & ~po007;
  assign new_new_n19061__ = ~new_new_n19059__ & ~new_new_n19060__;
  assign new_new_n19062__ = new_new_n19058__ & new_new_n19061__;
  assign new_new_n19063__ = ~new_new_n19058__ & ~new_new_n19061__;
  assign new_new_n19064__ = ~new_new_n19062__ & ~new_new_n19063__;
  assign new_new_n19065__ = pi082 & ~new_new_n19064__;
  assign new_new_n19066__ = ~pi082 & new_new_n19064__;
  assign new_new_n19067__ = new_new_n18628__ & po007;
  assign new_new_n19068__ = pi080 & ~po007;
  assign new_new_n19069__ = ~new_new_n19067__ & ~new_new_n19068__;
  assign new_new_n19070__ = ~new_new_n18446__ & ~new_new_n18447__;
  assign new_new_n19071__ = ~new_new_n19069__ & ~new_new_n19070__;
  assign new_new_n19072__ = new_new_n19069__ & new_new_n19070__;
  assign new_new_n19073__ = ~new_new_n19071__ & ~new_new_n19072__;
  assign new_new_n19074__ = pi081 & ~new_new_n19073__;
  assign new_new_n19075__ = ~pi081 & new_new_n19073__;
  assign new_new_n19076__ = ~pi079 & ~new_new_n18626__;
  assign new_new_n19077__ = pi079 & new_new_n18626__;
  assign new_new_n19078__ = ~new_new_n19076__ & ~new_new_n19077__;
  assign new_new_n19079__ = po007 & new_new_n19078__;
  assign new_new_n19080__ = ~new_new_n18454__ & ~new_new_n19079__;
  assign new_new_n19081__ = new_new_n18454__ & new_new_n19079__;
  assign new_new_n19082__ = ~new_new_n19080__ & ~new_new_n19081__;
  assign new_new_n19083__ = ~pi080 & ~new_new_n19082__;
  assign new_new_n19084__ = pi080 & new_new_n19082__;
  assign new_new_n19085__ = ~new_new_n18464__ & ~new_new_n18465__;
  assign new_new_n19086__ = ~new_new_n18624__ & po007;
  assign new_new_n19087__ = ~pi078 & ~po007;
  assign new_new_n19088__ = ~new_new_n19086__ & ~new_new_n19087__;
  assign new_new_n19089__ = new_new_n19085__ & ~new_new_n19088__;
  assign new_new_n19090__ = ~new_new_n19085__ & new_new_n19088__;
  assign new_new_n19091__ = ~new_new_n19089__ & ~new_new_n19090__;
  assign new_new_n19092__ = pi079 & ~new_new_n19091__;
  assign new_new_n19093__ = ~pi079 & new_new_n19091__;
  assign new_new_n19094__ = ~new_new_n18473__ & ~new_new_n18474__;
  assign new_new_n19095__ = ~new_new_n18622__ & po007;
  assign new_new_n19096__ = ~pi077 & ~po007;
  assign new_new_n19097__ = ~new_new_n19095__ & ~new_new_n19096__;
  assign new_new_n19098__ = ~new_new_n19094__ & ~new_new_n19097__;
  assign new_new_n19099__ = new_new_n19094__ & new_new_n19097__;
  assign new_new_n19100__ = ~new_new_n19098__ & ~new_new_n19099__;
  assign new_new_n19101__ = ~pi078 & ~new_new_n19100__;
  assign new_new_n19102__ = pi078 & new_new_n19100__;
  assign new_new_n19103__ = new_new_n18620__ & po007;
  assign new_new_n19104__ = pi076 & ~po007;
  assign new_new_n19105__ = ~new_new_n19103__ & ~new_new_n19104__;
  assign new_new_n19106__ = ~new_new_n18482__ & ~new_new_n18483__;
  assign new_new_n19107__ = ~new_new_n19105__ & ~new_new_n19106__;
  assign new_new_n19108__ = new_new_n19105__ & new_new_n19106__;
  assign new_new_n19109__ = ~new_new_n19107__ & ~new_new_n19108__;
  assign new_new_n19110__ = pi077 & ~new_new_n19109__;
  assign new_new_n19111__ = ~pi077 & new_new_n19109__;
  assign new_new_n19112__ = ~new_new_n18618__ & po007;
  assign new_new_n19113__ = pi075 & ~po007;
  assign new_new_n19114__ = ~new_new_n19112__ & ~new_new_n19113__;
  assign new_new_n19115__ = ~new_new_n18491__ & ~new_new_n18492__;
  assign new_new_n19116__ = ~new_new_n19114__ & new_new_n19115__;
  assign new_new_n19117__ = new_new_n19114__ & ~new_new_n19115__;
  assign new_new_n19118__ = ~new_new_n19116__ & ~new_new_n19117__;
  assign new_new_n19119__ = pi076 & new_new_n19118__;
  assign new_new_n19120__ = ~pi076 & ~new_new_n19118__;
  assign new_new_n19121__ = pi073 & ~new_new_n18614__;
  assign new_new_n19122__ = ~pi073 & new_new_n18614__;
  assign new_new_n19123__ = ~new_new_n19121__ & ~new_new_n19122__;
  assign new_new_n19124__ = po007 & new_new_n19123__;
  assign new_new_n19125__ = new_new_n18508__ & new_new_n19124__;
  assign new_new_n19126__ = ~new_new_n18508__ & ~new_new_n19124__;
  assign new_new_n19127__ = ~new_new_n19125__ & ~new_new_n19126__;
  assign new_new_n19128__ = pi074 & ~new_new_n19127__;
  assign new_new_n19129__ = ~pi074 & new_new_n19127__;
  assign new_new_n19130__ = new_new_n18612__ & po007;
  assign new_new_n19131__ = pi072 & ~po007;
  assign new_new_n19132__ = ~new_new_n19130__ & ~new_new_n19131__;
  assign new_new_n19133__ = ~new_new_n18518__ & ~new_new_n18519__;
  assign new_new_n19134__ = ~new_new_n19132__ & ~new_new_n19133__;
  assign new_new_n19135__ = new_new_n19132__ & new_new_n19133__;
  assign new_new_n19136__ = ~new_new_n19134__ & ~new_new_n19135__;
  assign new_new_n19137__ = pi073 & ~new_new_n19136__;
  assign new_new_n19138__ = ~pi073 & new_new_n19136__;
  assign new_new_n19139__ = ~new_new_n18527__ & ~new_new_n18528__;
  assign new_new_n19140__ = ~new_new_n18610__ & po007;
  assign new_new_n19141__ = ~pi071 & ~po007;
  assign new_new_n19142__ = ~new_new_n19140__ & ~new_new_n19141__;
  assign new_new_n19143__ = new_new_n19139__ & ~new_new_n19142__;
  assign new_new_n19144__ = ~new_new_n19139__ & new_new_n19142__;
  assign new_new_n19145__ = ~new_new_n19143__ & ~new_new_n19144__;
  assign new_new_n19146__ = pi072 & ~new_new_n19145__;
  assign new_new_n19147__ = ~pi072 & new_new_n19145__;
  assign new_new_n19148__ = new_new_n18608__ & po007;
  assign new_new_n19149__ = pi070 & ~po007;
  assign new_new_n19150__ = ~new_new_n19148__ & ~new_new_n19149__;
  assign new_new_n19151__ = ~new_new_n18536__ & ~new_new_n18537__;
  assign new_new_n19152__ = ~new_new_n19150__ & ~new_new_n19151__;
  assign new_new_n19153__ = new_new_n19150__ & new_new_n19151__;
  assign new_new_n19154__ = ~new_new_n19152__ & ~new_new_n19153__;
  assign new_new_n19155__ = ~pi071 & new_new_n19154__;
  assign new_new_n19156__ = pi071 & ~new_new_n19154__;
  assign new_new_n19157__ = ~pi069 & ~new_new_n18606__;
  assign new_new_n19158__ = pi069 & new_new_n18606__;
  assign new_new_n19159__ = ~new_new_n19157__ & ~new_new_n19158__;
  assign new_new_n19160__ = po007 & new_new_n19159__;
  assign new_new_n19161__ = ~new_new_n18542__ & new_new_n19160__;
  assign new_new_n19162__ = new_new_n18542__ & ~new_new_n19160__;
  assign new_new_n19163__ = ~new_new_n19161__ & ~new_new_n19162__;
  assign new_new_n19164__ = ~pi070 & new_new_n19163__;
  assign new_new_n19165__ = pi070 & ~new_new_n19163__;
  assign new_new_n19166__ = ~new_new_n18552__ & ~new_new_n18553__;
  assign new_new_n19167__ = ~new_new_n18604__ & po007;
  assign new_new_n19168__ = ~pi068 & ~po007;
  assign new_new_n19169__ = ~new_new_n19167__ & ~new_new_n19168__;
  assign new_new_n19170__ = ~new_new_n19166__ & ~new_new_n19169__;
  assign new_new_n19171__ = new_new_n19166__ & new_new_n19169__;
  assign new_new_n19172__ = ~new_new_n19170__ & ~new_new_n19171__;
  assign new_new_n19173__ = ~pi069 & ~new_new_n19172__;
  assign new_new_n19174__ = pi069 & new_new_n19172__;
  assign new_new_n19175__ = ~new_new_n18559__ & ~new_new_n18560__;
  assign new_new_n19176__ = ~new_new_n18602__ & po007;
  assign new_new_n19177__ = ~pi067 & ~po007;
  assign new_new_n19178__ = ~new_new_n19176__ & ~new_new_n19177__;
  assign new_new_n19179__ = new_new_n19175__ & ~new_new_n19178__;
  assign new_new_n19180__ = ~new_new_n19175__ & new_new_n19178__;
  assign new_new_n19181__ = ~new_new_n19179__ & ~new_new_n19180__;
  assign new_new_n19182__ = pi068 & ~new_new_n19181__;
  assign new_new_n19183__ = ~pi068 & new_new_n19181__;
  assign new_new_n19184__ = ~new_new_n18573__ & ~new_new_n18574__;
  assign new_new_n19185__ = po007 & new_new_n19184__;
  assign new_new_n19186__ = ~new_new_n18600__ & new_new_n19185__;
  assign new_new_n19187__ = new_new_n18600__ & ~new_new_n19185__;
  assign new_new_n19188__ = ~new_new_n19186__ & ~new_new_n19187__;
  assign new_new_n19189__ = pi067 & ~new_new_n19188__;
  assign new_new_n19190__ = ~pi067 & new_new_n19188__;
  assign new_new_n19191__ = pi007 & po007;
  assign new_new_n19192__ = ~pi007 & ~po007;
  assign new_new_n19193__ = ~pi065 & ~new_new_n19191__;
  assign new_new_n19194__ = ~new_new_n19192__ & new_new_n19193__;
  assign new_new_n19195__ = ~pi006 & ~new_new_n19194__;
  assign new_new_n19196__ = pi065 & new_new_n19191__;
  assign new_new_n19197__ = ~new_new_n19195__ & ~new_new_n19196__;
  assign new_new_n19198__ = pi064 & ~new_new_n19197__;
  assign new_new_n19199__ = pi064 & po007;
  assign new_new_n19200__ = ~pi007 & pi065;
  assign new_new_n19201__ = ~new_new_n19199__ & new_new_n19200__;
  assign new_new_n19202__ = ~new_new_n19198__ & ~new_new_n19201__;
  assign new_new_n19203__ = pi066 & ~new_new_n19202__;
  assign new_new_n19204__ = ~pi066 & new_new_n19202__;
  assign new_new_n19205__ = new_new_n426__ & ~po008;
  assign new_new_n19206__ = new_new_n18576__ & po007;
  assign new_new_n19207__ = ~new_new_n19205__ & ~new_new_n19206__;
  assign new_new_n19208__ = ~pi007 & ~new_new_n19207__;
  assign new_new_n19209__ = pi065 & po007;
  assign new_new_n19210__ = po008 & ~new_new_n19209__;
  assign new_new_n19211__ = pi065 & ~new_new_n18569__;
  assign new_new_n19212__ = pi007 & ~new_new_n19211__;
  assign new_new_n19213__ = ~new_new_n19210__ & new_new_n19212__;
  assign new_new_n19214__ = ~new_new_n332__ & po007;
  assign new_new_n19215__ = ~new_new_n18569__ & ~new_new_n19214__;
  assign new_new_n19216__ = ~new_new_n19208__ & ~new_new_n19215__;
  assign new_new_n19217__ = ~new_new_n19213__ & new_new_n19216__;
  assign new_new_n19218__ = pi008 & ~new_new_n19217__;
  assign new_new_n19219__ = ~new_new_n18569__ & ~new_new_n19209__;
  assign new_new_n19220__ = pi007 & ~new_new_n18582__;
  assign new_new_n19221__ = pi064 & ~new_new_n19220__;
  assign new_new_n19222__ = ~new_new_n19219__ & ~new_new_n19221__;
  assign new_new_n19223__ = ~pi065 & po007;
  assign new_new_n19224__ = ~po008 & ~new_new_n19223__;
  assign new_new_n19225__ = pi064 & ~new_new_n19191__;
  assign new_new_n19226__ = ~new_new_n19206__ & new_new_n19225__;
  assign new_new_n19227__ = ~new_new_n19224__ & new_new_n19226__;
  assign new_new_n19228__ = ~new_new_n19222__ & ~new_new_n19227__;
  assign new_new_n19229__ = ~pi008 & ~new_new_n19228__;
  assign new_new_n19230__ = ~new_new_n19218__ & ~new_new_n19229__;
  assign new_new_n19231__ = ~new_new_n19204__ & new_new_n19230__;
  assign new_new_n19232__ = ~new_new_n19203__ & ~new_new_n19231__;
  assign new_new_n19233__ = ~new_new_n19190__ & ~new_new_n19232__;
  assign new_new_n19234__ = ~new_new_n19189__ & ~new_new_n19233__;
  assign new_new_n19235__ = ~new_new_n19183__ & ~new_new_n19234__;
  assign new_new_n19236__ = ~new_new_n19182__ & ~new_new_n19235__;
  assign new_new_n19237__ = ~new_new_n19174__ & new_new_n19236__;
  assign new_new_n19238__ = ~new_new_n19173__ & ~new_new_n19237__;
  assign new_new_n19239__ = ~new_new_n19165__ & ~new_new_n19238__;
  assign new_new_n19240__ = ~new_new_n19164__ & ~new_new_n19239__;
  assign new_new_n19241__ = ~new_new_n19156__ & ~new_new_n19240__;
  assign new_new_n19242__ = ~new_new_n19155__ & ~new_new_n19241__;
  assign new_new_n19243__ = ~new_new_n19147__ & new_new_n19242__;
  assign new_new_n19244__ = ~new_new_n19146__ & ~new_new_n19243__;
  assign new_new_n19245__ = ~new_new_n19138__ & ~new_new_n19244__;
  assign new_new_n19246__ = ~new_new_n19137__ & ~new_new_n19245__;
  assign new_new_n19247__ = ~new_new_n19129__ & ~new_new_n19246__;
  assign new_new_n19248__ = ~new_new_n19128__ & ~new_new_n19247__;
  assign new_new_n19249__ = pi075 & ~new_new_n19248__;
  assign new_new_n19250__ = ~pi075 & new_new_n19248__;
  assign new_new_n19251__ = ~new_new_n18500__ & ~new_new_n18501__;
  assign new_new_n19252__ = new_new_n18616__ & po007;
  assign new_new_n19253__ = ~pi074 & ~po007;
  assign new_new_n19254__ = ~new_new_n19252__ & ~new_new_n19253__;
  assign new_new_n19255__ = ~new_new_n19251__ & ~new_new_n19254__;
  assign new_new_n19256__ = new_new_n19251__ & new_new_n19254__;
  assign new_new_n19257__ = ~new_new_n19255__ & ~new_new_n19256__;
  assign new_new_n19258__ = ~new_new_n19250__ & new_new_n19257__;
  assign new_new_n19259__ = ~new_new_n19249__ & ~new_new_n19258__;
  assign new_new_n19260__ = ~new_new_n19120__ & ~new_new_n19259__;
  assign new_new_n19261__ = ~new_new_n19119__ & ~new_new_n19260__;
  assign new_new_n19262__ = ~new_new_n19111__ & ~new_new_n19261__;
  assign new_new_n19263__ = ~new_new_n19110__ & ~new_new_n19262__;
  assign new_new_n19264__ = ~new_new_n19102__ & new_new_n19263__;
  assign new_new_n19265__ = ~new_new_n19101__ & ~new_new_n19264__;
  assign new_new_n19266__ = ~new_new_n19093__ & new_new_n19265__;
  assign new_new_n19267__ = ~new_new_n19092__ & ~new_new_n19266__;
  assign new_new_n19268__ = ~new_new_n19084__ & new_new_n19267__;
  assign new_new_n19269__ = ~new_new_n19083__ & ~new_new_n19268__;
  assign new_new_n19270__ = ~new_new_n19075__ & new_new_n19269__;
  assign new_new_n19271__ = ~new_new_n19074__ & ~new_new_n19270__;
  assign new_new_n19272__ = ~new_new_n19066__ & ~new_new_n19271__;
  assign new_new_n19273__ = ~new_new_n19065__ & ~new_new_n19272__;
  assign new_new_n19274__ = ~new_new_n19057__ & ~new_new_n19273__;
  assign new_new_n19275__ = ~new_new_n19056__ & ~new_new_n19274__;
  assign new_new_n19276__ = ~new_new_n19048__ & ~new_new_n19275__;
  assign new_new_n19277__ = ~new_new_n19047__ & ~new_new_n19276__;
  assign new_new_n19278__ = ~new_new_n19039__ & new_new_n19277__;
  assign new_new_n19279__ = ~new_new_n19038__ & ~new_new_n19278__;
  assign new_new_n19280__ = ~new_new_n19030__ & new_new_n19279__;
  assign new_new_n19281__ = ~new_new_n19029__ & ~new_new_n19280__;
  assign new_new_n19282__ = ~new_new_n19021__ & ~new_new_n19281__;
  assign new_new_n19283__ = ~new_new_n19020__ & ~new_new_n19282__;
  assign new_new_n19284__ = ~new_new_n19012__ & ~new_new_n19283__;
  assign new_new_n19285__ = ~new_new_n19011__ & ~new_new_n19284__;
  assign new_new_n19286__ = ~new_new_n19003__ & ~new_new_n19285__;
  assign new_new_n19287__ = ~new_new_n19002__ & ~new_new_n19286__;
  assign new_new_n19288__ = ~new_new_n18994__ & ~new_new_n19287__;
  assign new_new_n19289__ = ~new_new_n18993__ & ~new_new_n19288__;
  assign new_new_n19290__ = ~new_new_n18985__ & ~new_new_n19289__;
  assign new_new_n19291__ = ~new_new_n18984__ & ~new_new_n19290__;
  assign new_new_n19292__ = ~new_new_n18976__ & new_new_n19291__;
  assign new_new_n19293__ = ~new_new_n18975__ & ~new_new_n19292__;
  assign new_new_n19294__ = ~new_new_n18967__ & new_new_n19293__;
  assign new_new_n19295__ = ~new_new_n18966__ & ~new_new_n19294__;
  assign new_new_n19296__ = ~new_new_n18958__ & ~new_new_n19295__;
  assign new_new_n19297__ = ~new_new_n18957__ & ~new_new_n19296__;
  assign new_new_n19298__ = ~new_new_n18949__ & ~new_new_n19297__;
  assign new_new_n19299__ = ~new_new_n18948__ & ~new_new_n19298__;
  assign new_new_n19300__ = ~new_new_n18940__ & ~new_new_n19299__;
  assign new_new_n19301__ = ~new_new_n18939__ & ~new_new_n19300__;
  assign new_new_n19302__ = ~new_new_n18931__ & new_new_n19301__;
  assign new_new_n19303__ = ~new_new_n18930__ & ~new_new_n19302__;
  assign new_new_n19304__ = ~new_new_n18922__ & ~new_new_n19303__;
  assign new_new_n19305__ = ~new_new_n18921__ & ~new_new_n19304__;
  assign new_new_n19306__ = ~new_new_n18913__ & new_new_n19305__;
  assign new_new_n19307__ = ~new_new_n18912__ & ~new_new_n19306__;
  assign new_new_n19308__ = ~new_new_n18904__ & new_new_n19307__;
  assign new_new_n19309__ = ~new_new_n18903__ & ~new_new_n19308__;
  assign new_new_n19310__ = ~new_new_n18895__ & new_new_n19309__;
  assign new_new_n19311__ = ~new_new_n18894__ & ~new_new_n19310__;
  assign new_new_n19312__ = ~new_new_n18886__ & new_new_n19311__;
  assign new_new_n19313__ = ~new_new_n18885__ & ~new_new_n19312__;
  assign new_new_n19314__ = ~new_new_n18877__ & ~new_new_n19313__;
  assign new_new_n19315__ = ~new_new_n18876__ & ~new_new_n19314__;
  assign new_new_n19316__ = ~new_new_n18868__ & ~new_new_n19315__;
  assign new_new_n19317__ = ~new_new_n18867__ & ~new_new_n19316__;
  assign new_new_n19318__ = ~new_new_n18859__ & ~new_new_n19317__;
  assign new_new_n19319__ = ~new_new_n18858__ & ~new_new_n19318__;
  assign new_new_n19320__ = ~new_new_n18850__ & ~new_new_n19319__;
  assign new_new_n19321__ = ~new_new_n18849__ & ~new_new_n19320__;
  assign new_new_n19322__ = ~new_new_n18841__ & ~new_new_n19321__;
  assign new_new_n19323__ = ~new_new_n18840__ & ~new_new_n19322__;
  assign new_new_n19324__ = ~new_new_n18832__ & ~new_new_n19323__;
  assign new_new_n19325__ = ~new_new_n18831__ & ~new_new_n19324__;
  assign new_new_n19326__ = ~new_new_n18823__ & ~new_new_n19325__;
  assign new_new_n19327__ = ~new_new_n18822__ & ~new_new_n19326__;
  assign new_new_n19328__ = pi110 & new_new_n19327__;
  assign new_new_n19329__ = ~pi110 & ~new_new_n19327__;
  assign new_new_n19330__ = ~new_new_n18185__ & ~new_new_n18186__;
  assign new_new_n19331__ = ~new_new_n18686__ & po007;
  assign new_new_n19332__ = ~pi109 & ~po007;
  assign new_new_n19333__ = ~new_new_n19331__ & ~new_new_n19332__;
  assign new_new_n19334__ = new_new_n19330__ & ~new_new_n19333__;
  assign new_new_n19335__ = ~new_new_n19330__ & new_new_n19333__;
  assign new_new_n19336__ = ~new_new_n19334__ & ~new_new_n19335__;
  assign new_new_n19337__ = ~new_new_n19329__ & ~new_new_n19336__;
  assign new_new_n19338__ = ~new_new_n19328__ & ~new_new_n19337__;
  assign new_new_n19339__ = ~new_new_n18814__ & ~new_new_n19338__;
  assign new_new_n19340__ = ~new_new_n18813__ & ~new_new_n19339__;
  assign new_new_n19341__ = ~new_new_n18805__ & new_new_n19340__;
  assign new_new_n19342__ = ~new_new_n18804__ & ~new_new_n19341__;
  assign new_new_n19343__ = ~new_new_n18796__ & ~new_new_n19342__;
  assign new_new_n19344__ = ~new_new_n18795__ & ~new_new_n19343__;
  assign new_new_n19345__ = ~new_new_n18787__ & new_new_n19344__;
  assign new_new_n19346__ = ~new_new_n18786__ & ~new_new_n19345__;
  assign new_new_n19347__ = ~new_new_n18778__ & ~new_new_n19346__;
  assign new_new_n19348__ = ~new_new_n18777__ & ~new_new_n19347__;
  assign new_new_n19349__ = ~new_new_n18769__ & ~new_new_n19348__;
  assign new_new_n19350__ = ~new_new_n18768__ & ~new_new_n19349__;
  assign new_new_n19351__ = ~new_new_n18760__ & ~new_new_n19350__;
  assign new_new_n19352__ = ~new_new_n18759__ & ~new_new_n19351__;
  assign new_new_n19353__ = ~new_new_n18751__ & new_new_n19352__;
  assign new_new_n19354__ = ~new_new_n18750__ & ~new_new_n19353__;
  assign new_new_n19355__ = ~new_new_n18742__ & new_new_n19354__;
  assign new_new_n19356__ = ~new_new_n18741__ & ~new_new_n19355__;
  assign new_new_n19357__ = ~new_new_n18733__ & ~new_new_n19356__;
  assign new_new_n19358__ = ~new_new_n18732__ & ~new_new_n19357__;
  assign new_new_n19359__ = ~pi121 & new_new_n19358__;
  assign new_new_n19360__ = new_new_n264__ & ~new_new_n19359__;
  assign new_new_n19361__ = ~pi121 & new_new_n18717__;
  assign new_new_n19362__ = ~new_new_n19358__ & ~new_new_n19361__;
  assign new_new_n19363__ = pi121 & ~new_new_n17442__;
  assign new_new_n19364__ = new_new_n264__ & ~new_new_n19363__;
  assign po006 = ~new_new_n19362__ & new_new_n19364__;
  assign new_new_n19366__ = new_new_n19356__ & po006;
  assign new_new_n19367__ = ~pi120 & ~po006;
  assign new_new_n19368__ = ~new_new_n19366__ & ~new_new_n19367__;
  assign new_new_n19369__ = ~new_new_n18732__ & ~new_new_n18733__;
  assign new_new_n19370__ = ~new_new_n19368__ & ~new_new_n19369__;
  assign new_new_n19371__ = new_new_n19368__ & new_new_n19369__;
  assign new_new_n19372__ = ~new_new_n19370__ & ~new_new_n19371__;
  assign new_new_n19373__ = pi121 & new_new_n19372__;
  assign new_new_n19374__ = new_new_n19354__ & po006;
  assign new_new_n19375__ = pi119 & ~po006;
  assign new_new_n19376__ = ~new_new_n19374__ & ~new_new_n19375__;
  assign new_new_n19377__ = ~new_new_n18741__ & ~new_new_n18742__;
  assign new_new_n19378__ = ~new_new_n19376__ & ~new_new_n19377__;
  assign new_new_n19379__ = new_new_n19376__ & new_new_n19377__;
  assign new_new_n19380__ = ~new_new_n19378__ & ~new_new_n19379__;
  assign new_new_n19381__ = ~pi120 & new_new_n19380__;
  assign new_new_n19382__ = pi120 & ~new_new_n19380__;
  assign new_new_n19383__ = ~new_new_n18750__ & ~new_new_n18751__;
  assign new_new_n19384__ = new_new_n19352__ & po006;
  assign new_new_n19385__ = ~pi118 & ~po006;
  assign new_new_n19386__ = ~new_new_n19384__ & ~new_new_n19385__;
  assign new_new_n19387__ = ~new_new_n19383__ & ~new_new_n19386__;
  assign new_new_n19388__ = new_new_n19383__ & new_new_n19386__;
  assign new_new_n19389__ = ~new_new_n19387__ & ~new_new_n19388__;
  assign new_new_n19390__ = ~pi119 & ~new_new_n19389__;
  assign new_new_n19391__ = pi119 & new_new_n19389__;
  assign new_new_n19392__ = ~new_new_n19350__ & po006;
  assign new_new_n19393__ = pi117 & ~po006;
  assign new_new_n19394__ = ~new_new_n19392__ & ~new_new_n19393__;
  assign new_new_n19395__ = ~new_new_n18759__ & ~new_new_n18760__;
  assign new_new_n19396__ = ~new_new_n19394__ & new_new_n19395__;
  assign new_new_n19397__ = new_new_n19394__ & ~new_new_n19395__;
  assign new_new_n19398__ = ~new_new_n19396__ & ~new_new_n19397__;
  assign new_new_n19399__ = pi118 & new_new_n19398__;
  assign new_new_n19400__ = ~pi118 & ~new_new_n19398__;
  assign new_new_n19401__ = pi116 & ~new_new_n19348__;
  assign new_new_n19402__ = ~pi116 & new_new_n19348__;
  assign new_new_n19403__ = ~new_new_n19401__ & ~new_new_n19402__;
  assign new_new_n19404__ = po006 & new_new_n19403__;
  assign new_new_n19405__ = ~new_new_n18767__ & ~new_new_n19404__;
  assign new_new_n19406__ = new_new_n18767__ & new_new_n19404__;
  assign new_new_n19407__ = ~new_new_n19405__ & ~new_new_n19406__;
  assign new_new_n19408__ = pi117 & ~new_new_n19407__;
  assign new_new_n19409__ = ~pi117 & new_new_n19407__;
  assign new_new_n19410__ = ~new_new_n18777__ & ~new_new_n18778__;
  assign new_new_n19411__ = ~new_new_n19346__ & po006;
  assign new_new_n19412__ = pi115 & ~po006;
  assign new_new_n19413__ = ~new_new_n19411__ & ~new_new_n19412__;
  assign new_new_n19414__ = new_new_n19410__ & new_new_n19413__;
  assign new_new_n19415__ = ~new_new_n19410__ & ~new_new_n19413__;
  assign new_new_n19416__ = ~new_new_n19414__ & ~new_new_n19415__;
  assign new_new_n19417__ = pi116 & ~new_new_n19416__;
  assign new_new_n19418__ = ~pi116 & new_new_n19416__;
  assign new_new_n19419__ = new_new_n19344__ & po006;
  assign new_new_n19420__ = pi114 & ~po006;
  assign new_new_n19421__ = ~new_new_n19419__ & ~new_new_n19420__;
  assign new_new_n19422__ = ~new_new_n18786__ & ~new_new_n18787__;
  assign new_new_n19423__ = ~new_new_n19421__ & ~new_new_n19422__;
  assign new_new_n19424__ = new_new_n19421__ & new_new_n19422__;
  assign new_new_n19425__ = ~new_new_n19423__ & ~new_new_n19424__;
  assign new_new_n19426__ = pi115 & ~new_new_n19425__;
  assign new_new_n19427__ = ~pi115 & new_new_n19425__;
  assign new_new_n19428__ = ~new_new_n18795__ & ~new_new_n18796__;
  assign new_new_n19429__ = ~new_new_n19342__ & po006;
  assign new_new_n19430__ = ~pi113 & ~po006;
  assign new_new_n19431__ = ~new_new_n19429__ & ~new_new_n19430__;
  assign new_new_n19432__ = new_new_n19428__ & ~new_new_n19431__;
  assign new_new_n19433__ = ~new_new_n19428__ & new_new_n19431__;
  assign new_new_n19434__ = ~new_new_n19432__ & ~new_new_n19433__;
  assign new_new_n19435__ = pi114 & ~new_new_n19434__;
  assign new_new_n19436__ = ~pi114 & new_new_n19434__;
  assign new_new_n19437__ = ~new_new_n19340__ & po006;
  assign new_new_n19438__ = pi112 & ~po006;
  assign new_new_n19439__ = ~new_new_n19437__ & ~new_new_n19438__;
  assign new_new_n19440__ = ~new_new_n18804__ & ~new_new_n18805__;
  assign new_new_n19441__ = ~new_new_n19439__ & new_new_n19440__;
  assign new_new_n19442__ = new_new_n19439__ & ~new_new_n19440__;
  assign new_new_n19443__ = ~new_new_n19441__ & ~new_new_n19442__;
  assign new_new_n19444__ = ~pi113 & ~new_new_n19443__;
  assign new_new_n19445__ = pi113 & new_new_n19443__;
  assign new_new_n19446__ = ~new_new_n19338__ & po006;
  assign new_new_n19447__ = pi111 & ~po006;
  assign new_new_n19448__ = ~new_new_n19446__ & ~new_new_n19447__;
  assign new_new_n19449__ = ~new_new_n18813__ & ~new_new_n18814__;
  assign new_new_n19450__ = ~new_new_n19448__ & new_new_n19449__;
  assign new_new_n19451__ = new_new_n19448__ & ~new_new_n19449__;
  assign new_new_n19452__ = ~new_new_n19450__ & ~new_new_n19451__;
  assign new_new_n19453__ = ~pi112 & ~new_new_n19452__;
  assign new_new_n19454__ = pi112 & new_new_n19452__;
  assign new_new_n19455__ = ~new_new_n19328__ & ~new_new_n19329__;
  assign new_new_n19456__ = po006 & new_new_n19455__;
  assign new_new_n19457__ = ~new_new_n19336__ & ~new_new_n19456__;
  assign new_new_n19458__ = new_new_n19336__ & new_new_n19456__;
  assign new_new_n19459__ = ~new_new_n19457__ & ~new_new_n19458__;
  assign new_new_n19460__ = pi111 & ~new_new_n19459__;
  assign new_new_n19461__ = ~pi111 & new_new_n19459__;
  assign new_new_n19462__ = ~new_new_n18822__ & ~new_new_n18823__;
  assign new_new_n19463__ = ~new_new_n19325__ & po006;
  assign new_new_n19464__ = ~pi109 & ~po006;
  assign new_new_n19465__ = ~new_new_n19463__ & ~new_new_n19464__;
  assign new_new_n19466__ = new_new_n19462__ & ~new_new_n19465__;
  assign new_new_n19467__ = ~new_new_n19462__ & new_new_n19465__;
  assign new_new_n19468__ = ~new_new_n19466__ & ~new_new_n19467__;
  assign new_new_n19469__ = pi110 & ~new_new_n19468__;
  assign new_new_n19470__ = ~pi110 & new_new_n19468__;
  assign new_new_n19471__ = ~new_new_n18831__ & ~new_new_n18832__;
  assign new_new_n19472__ = ~new_new_n19323__ & po006;
  assign new_new_n19473__ = ~pi108 & ~po006;
  assign new_new_n19474__ = ~new_new_n19472__ & ~new_new_n19473__;
  assign new_new_n19475__ = new_new_n19471__ & ~new_new_n19474__;
  assign new_new_n19476__ = ~new_new_n19471__ & new_new_n19474__;
  assign new_new_n19477__ = ~new_new_n19475__ & ~new_new_n19476__;
  assign new_new_n19478__ = pi109 & ~new_new_n19477__;
  assign new_new_n19479__ = ~pi109 & new_new_n19477__;
  assign new_new_n19480__ = ~pi107 & ~new_new_n19321__;
  assign new_new_n19481__ = pi107 & new_new_n19321__;
  assign new_new_n19482__ = ~new_new_n19480__ & ~new_new_n19481__;
  assign new_new_n19483__ = po006 & new_new_n19482__;
  assign new_new_n19484__ = new_new_n18839__ & new_new_n19483__;
  assign new_new_n19485__ = ~new_new_n18839__ & ~new_new_n19483__;
  assign new_new_n19486__ = ~new_new_n19484__ & ~new_new_n19485__;
  assign new_new_n19487__ = ~pi108 & ~new_new_n19486__;
  assign new_new_n19488__ = pi108 & new_new_n19486__;
  assign new_new_n19489__ = ~pi106 & ~new_new_n19319__;
  assign new_new_n19490__ = pi106 & new_new_n19319__;
  assign new_new_n19491__ = ~new_new_n19489__ & ~new_new_n19490__;
  assign new_new_n19492__ = po006 & new_new_n19491__;
  assign new_new_n19493__ = new_new_n18848__ & new_new_n19492__;
  assign new_new_n19494__ = ~new_new_n18848__ & ~new_new_n19492__;
  assign new_new_n19495__ = ~new_new_n19493__ & ~new_new_n19494__;
  assign new_new_n19496__ = ~pi107 & ~new_new_n19495__;
  assign new_new_n19497__ = pi107 & new_new_n19495__;
  assign new_new_n19498__ = ~new_new_n18858__ & ~new_new_n18859__;
  assign new_new_n19499__ = ~new_new_n19317__ & po006;
  assign new_new_n19500__ = ~pi105 & ~po006;
  assign new_new_n19501__ = ~new_new_n19499__ & ~new_new_n19500__;
  assign new_new_n19502__ = new_new_n19498__ & ~new_new_n19501__;
  assign new_new_n19503__ = ~new_new_n19498__ & new_new_n19501__;
  assign new_new_n19504__ = ~new_new_n19502__ & ~new_new_n19503__;
  assign new_new_n19505__ = ~pi106 & new_new_n19504__;
  assign new_new_n19506__ = pi106 & ~new_new_n19504__;
  assign new_new_n19507__ = ~pi104 & ~new_new_n19315__;
  assign new_new_n19508__ = pi104 & new_new_n19315__;
  assign new_new_n19509__ = ~new_new_n19507__ & ~new_new_n19508__;
  assign new_new_n19510__ = po006 & new_new_n19509__;
  assign new_new_n19511__ = new_new_n18866__ & new_new_n19510__;
  assign new_new_n19512__ = ~new_new_n18866__ & ~new_new_n19510__;
  assign new_new_n19513__ = ~new_new_n19511__ & ~new_new_n19512__;
  assign new_new_n19514__ = ~pi105 & ~new_new_n19513__;
  assign new_new_n19515__ = pi105 & new_new_n19513__;
  assign new_new_n19516__ = ~pi103 & ~new_new_n19313__;
  assign new_new_n19517__ = pi103 & new_new_n19313__;
  assign new_new_n19518__ = ~new_new_n19516__ & ~new_new_n19517__;
  assign new_new_n19519__ = po006 & new_new_n19518__;
  assign new_new_n19520__ = new_new_n18875__ & new_new_n19519__;
  assign new_new_n19521__ = ~new_new_n18875__ & ~new_new_n19519__;
  assign new_new_n19522__ = ~new_new_n19520__ & ~new_new_n19521__;
  assign new_new_n19523__ = ~pi104 & ~new_new_n19522__;
  assign new_new_n19524__ = pi104 & new_new_n19522__;
  assign new_new_n19525__ = ~new_new_n18885__ & ~new_new_n18886__;
  assign new_new_n19526__ = ~new_new_n19311__ & po006;
  assign new_new_n19527__ = pi102 & ~po006;
  assign new_new_n19528__ = ~new_new_n19526__ & ~new_new_n19527__;
  assign new_new_n19529__ = new_new_n19525__ & ~new_new_n19528__;
  assign new_new_n19530__ = ~new_new_n19525__ & new_new_n19528__;
  assign new_new_n19531__ = ~new_new_n19529__ & ~new_new_n19530__;
  assign new_new_n19532__ = ~pi103 & ~new_new_n19531__;
  assign new_new_n19533__ = pi103 & new_new_n19531__;
  assign new_new_n19534__ = ~new_new_n18894__ & ~new_new_n18895__;
  assign new_new_n19535__ = ~new_new_n19309__ & po006;
  assign new_new_n19536__ = ~pi101 & ~po006;
  assign new_new_n19537__ = ~new_new_n19535__ & ~new_new_n19536__;
  assign new_new_n19538__ = new_new_n19534__ & ~new_new_n19537__;
  assign new_new_n19539__ = ~new_new_n19534__ & new_new_n19537__;
  assign new_new_n19540__ = ~new_new_n19538__ & ~new_new_n19539__;
  assign new_new_n19541__ = pi102 & ~new_new_n19540__;
  assign new_new_n19542__ = ~pi102 & new_new_n19540__;
  assign new_new_n19543__ = ~new_new_n18903__ & ~new_new_n18904__;
  assign new_new_n19544__ = new_new_n19307__ & po006;
  assign new_new_n19545__ = ~pi100 & ~po006;
  assign new_new_n19546__ = ~new_new_n19544__ & ~new_new_n19545__;
  assign new_new_n19547__ = ~new_new_n19543__ & ~new_new_n19546__;
  assign new_new_n19548__ = new_new_n19543__ & new_new_n19546__;
  assign new_new_n19549__ = ~new_new_n19547__ & ~new_new_n19548__;
  assign new_new_n19550__ = ~pi101 & ~new_new_n19549__;
  assign new_new_n19551__ = pi101 & new_new_n19549__;
  assign new_new_n19552__ = new_new_n19305__ & po006;
  assign new_new_n19553__ = pi099 & ~po006;
  assign new_new_n19554__ = ~new_new_n19552__ & ~new_new_n19553__;
  assign new_new_n19555__ = ~new_new_n18912__ & ~new_new_n18913__;
  assign new_new_n19556__ = ~new_new_n19554__ & ~new_new_n19555__;
  assign new_new_n19557__ = new_new_n19554__ & new_new_n19555__;
  assign new_new_n19558__ = ~new_new_n19556__ & ~new_new_n19557__;
  assign new_new_n19559__ = ~pi100 & new_new_n19558__;
  assign new_new_n19560__ = ~new_new_n18921__ & ~new_new_n18922__;
  assign new_new_n19561__ = ~new_new_n19303__ & po006;
  assign new_new_n19562__ = ~pi098 & ~po006;
  assign new_new_n19563__ = ~new_new_n19561__ & ~new_new_n19562__;
  assign new_new_n19564__ = ~new_new_n19560__ & ~new_new_n19563__;
  assign new_new_n19565__ = new_new_n19560__ & new_new_n19563__;
  assign new_new_n19566__ = ~new_new_n19564__ & ~new_new_n19565__;
  assign new_new_n19567__ = ~pi099 & ~new_new_n19566__;
  assign new_new_n19568__ = pi099 & new_new_n19566__;
  assign new_new_n19569__ = new_new_n19301__ & po006;
  assign new_new_n19570__ = ~pi097 & ~po006;
  assign new_new_n19571__ = ~new_new_n19569__ & ~new_new_n19570__;
  assign new_new_n19572__ = ~new_new_n18930__ & ~new_new_n18931__;
  assign new_new_n19573__ = ~new_new_n19571__ & ~new_new_n19572__;
  assign new_new_n19574__ = new_new_n19571__ & new_new_n19572__;
  assign new_new_n19575__ = ~new_new_n19573__ & ~new_new_n19574__;
  assign new_new_n19576__ = ~pi098 & ~new_new_n19575__;
  assign new_new_n19577__ = pi098 & new_new_n19575__;
  assign new_new_n19578__ = ~new_new_n18939__ & ~new_new_n18940__;
  assign new_new_n19579__ = ~new_new_n19299__ & po006;
  assign new_new_n19580__ = pi096 & ~po006;
  assign new_new_n19581__ = ~new_new_n19579__ & ~new_new_n19580__;
  assign new_new_n19582__ = new_new_n19578__ & ~new_new_n19581__;
  assign new_new_n19583__ = ~new_new_n19578__ & new_new_n19581__;
  assign new_new_n19584__ = ~new_new_n19582__ & ~new_new_n19583__;
  assign new_new_n19585__ = pi097 & new_new_n19584__;
  assign new_new_n19586__ = ~pi097 & ~new_new_n19584__;
  assign new_new_n19587__ = pi095 & ~new_new_n19297__;
  assign new_new_n19588__ = ~pi095 & new_new_n19297__;
  assign new_new_n19589__ = ~new_new_n19587__ & ~new_new_n19588__;
  assign new_new_n19590__ = po006 & new_new_n19589__;
  assign new_new_n19591__ = new_new_n18947__ & new_new_n19590__;
  assign new_new_n19592__ = ~new_new_n18947__ & ~new_new_n19590__;
  assign new_new_n19593__ = ~new_new_n19591__ & ~new_new_n19592__;
  assign new_new_n19594__ = pi096 & ~new_new_n19593__;
  assign new_new_n19595__ = ~pi096 & new_new_n19593__;
  assign new_new_n19596__ = pi094 & ~new_new_n19295__;
  assign new_new_n19597__ = ~pi094 & new_new_n19295__;
  assign new_new_n19598__ = ~new_new_n19596__ & ~new_new_n19597__;
  assign new_new_n19599__ = po006 & new_new_n19598__;
  assign new_new_n19600__ = new_new_n18956__ & new_new_n19599__;
  assign new_new_n19601__ = ~new_new_n18956__ & ~new_new_n19599__;
  assign new_new_n19602__ = ~new_new_n19600__ & ~new_new_n19601__;
  assign new_new_n19603__ = pi095 & ~new_new_n19602__;
  assign new_new_n19604__ = ~pi095 & new_new_n19602__;
  assign new_new_n19605__ = ~new_new_n18966__ & ~new_new_n18967__;
  assign new_new_n19606__ = ~new_new_n19293__ & po006;
  assign new_new_n19607__ = ~pi093 & ~po006;
  assign new_new_n19608__ = ~new_new_n19606__ & ~new_new_n19607__;
  assign new_new_n19609__ = new_new_n19605__ & ~new_new_n19608__;
  assign new_new_n19610__ = ~new_new_n19605__ & new_new_n19608__;
  assign new_new_n19611__ = ~new_new_n19609__ & ~new_new_n19610__;
  assign new_new_n19612__ = pi094 & ~new_new_n19611__;
  assign new_new_n19613__ = ~pi094 & new_new_n19611__;
  assign new_new_n19614__ = ~new_new_n18975__ & ~new_new_n18976__;
  assign new_new_n19615__ = ~new_new_n19291__ & po006;
  assign new_new_n19616__ = pi092 & ~po006;
  assign new_new_n19617__ = ~new_new_n19615__ & ~new_new_n19616__;
  assign new_new_n19618__ = new_new_n19614__ & ~new_new_n19617__;
  assign new_new_n19619__ = ~new_new_n19614__ & new_new_n19617__;
  assign new_new_n19620__ = ~new_new_n19618__ & ~new_new_n19619__;
  assign new_new_n19621__ = ~pi093 & ~new_new_n19620__;
  assign new_new_n19622__ = pi093 & new_new_n19620__;
  assign new_new_n19623__ = ~new_new_n19289__ & po006;
  assign new_new_n19624__ = pi091 & ~po006;
  assign new_new_n19625__ = ~new_new_n19623__ & ~new_new_n19624__;
  assign new_new_n19626__ = ~new_new_n18984__ & ~new_new_n18985__;
  assign new_new_n19627__ = ~new_new_n19625__ & new_new_n19626__;
  assign new_new_n19628__ = new_new_n19625__ & ~new_new_n19626__;
  assign new_new_n19629__ = ~new_new_n19627__ & ~new_new_n19628__;
  assign new_new_n19630__ = ~pi092 & ~new_new_n19629__;
  assign new_new_n19631__ = pi092 & new_new_n19629__;
  assign new_new_n19632__ = ~new_new_n18993__ & ~new_new_n18994__;
  assign new_new_n19633__ = pi090 & ~po006;
  assign new_new_n19634__ = ~new_new_n19287__ & po006;
  assign new_new_n19635__ = ~new_new_n19633__ & ~new_new_n19634__;
  assign new_new_n19636__ = new_new_n19632__ & new_new_n19635__;
  assign new_new_n19637__ = ~new_new_n19632__ & ~new_new_n19635__;
  assign new_new_n19638__ = ~new_new_n19636__ & ~new_new_n19637__;
  assign new_new_n19639__ = pi091 & ~new_new_n19638__;
  assign new_new_n19640__ = ~pi091 & new_new_n19638__;
  assign new_new_n19641__ = ~new_new_n19002__ & ~new_new_n19003__;
  assign new_new_n19642__ = pi089 & ~po006;
  assign new_new_n19643__ = ~new_new_n19285__ & po006;
  assign new_new_n19644__ = ~new_new_n19642__ & ~new_new_n19643__;
  assign new_new_n19645__ = new_new_n19641__ & new_new_n19644__;
  assign new_new_n19646__ = ~new_new_n19641__ & ~new_new_n19644__;
  assign new_new_n19647__ = ~new_new_n19645__ & ~new_new_n19646__;
  assign new_new_n19648__ = pi090 & ~new_new_n19647__;
  assign new_new_n19649__ = ~pi090 & new_new_n19647__;
  assign new_new_n19650__ = ~new_new_n19011__ & ~new_new_n19012__;
  assign new_new_n19651__ = ~new_new_n19283__ & po006;
  assign new_new_n19652__ = pi088 & ~po006;
  assign new_new_n19653__ = ~new_new_n19651__ & ~new_new_n19652__;
  assign new_new_n19654__ = new_new_n19650__ & new_new_n19653__;
  assign new_new_n19655__ = ~new_new_n19650__ & ~new_new_n19653__;
  assign new_new_n19656__ = ~new_new_n19654__ & ~new_new_n19655__;
  assign new_new_n19657__ = pi089 & ~new_new_n19656__;
  assign new_new_n19658__ = ~pi089 & new_new_n19656__;
  assign new_new_n19659__ = new_new_n19281__ & po006;
  assign new_new_n19660__ = ~pi087 & ~po006;
  assign new_new_n19661__ = ~new_new_n19659__ & ~new_new_n19660__;
  assign new_new_n19662__ = ~new_new_n19020__ & ~new_new_n19021__;
  assign new_new_n19663__ = ~new_new_n19661__ & ~new_new_n19662__;
  assign new_new_n19664__ = new_new_n19661__ & new_new_n19662__;
  assign new_new_n19665__ = ~new_new_n19663__ & ~new_new_n19664__;
  assign new_new_n19666__ = ~pi088 & ~new_new_n19665__;
  assign new_new_n19667__ = pi088 & new_new_n19665__;
  assign new_new_n19668__ = new_new_n19279__ & po006;
  assign new_new_n19669__ = pi086 & ~po006;
  assign new_new_n19670__ = ~new_new_n19668__ & ~new_new_n19669__;
  assign new_new_n19671__ = ~new_new_n19029__ & ~new_new_n19030__;
  assign new_new_n19672__ = ~new_new_n19670__ & ~new_new_n19671__;
  assign new_new_n19673__ = new_new_n19670__ & new_new_n19671__;
  assign new_new_n19674__ = ~new_new_n19672__ & ~new_new_n19673__;
  assign new_new_n19675__ = ~pi087 & new_new_n19674__;
  assign new_new_n19676__ = pi087 & ~new_new_n19674__;
  assign new_new_n19677__ = new_new_n19277__ & po006;
  assign new_new_n19678__ = ~pi085 & ~po006;
  assign new_new_n19679__ = ~new_new_n19677__ & ~new_new_n19678__;
  assign new_new_n19680__ = ~new_new_n19038__ & ~new_new_n19039__;
  assign new_new_n19681__ = ~new_new_n19679__ & ~new_new_n19680__;
  assign new_new_n19682__ = new_new_n19679__ & new_new_n19680__;
  assign new_new_n19683__ = ~new_new_n19681__ & ~new_new_n19682__;
  assign new_new_n19684__ = ~pi086 & ~new_new_n19683__;
  assign new_new_n19685__ = pi086 & new_new_n19683__;
  assign new_new_n19686__ = ~new_new_n19047__ & ~new_new_n19048__;
  assign new_new_n19687__ = ~new_new_n19275__ & po006;
  assign new_new_n19688__ = pi084 & ~po006;
  assign new_new_n19689__ = ~new_new_n19687__ & ~new_new_n19688__;
  assign new_new_n19690__ = new_new_n19686__ & ~new_new_n19689__;
  assign new_new_n19691__ = ~new_new_n19686__ & new_new_n19689__;
  assign new_new_n19692__ = ~new_new_n19690__ & ~new_new_n19691__;
  assign new_new_n19693__ = ~pi085 & ~new_new_n19692__;
  assign new_new_n19694__ = pi085 & new_new_n19692__;
  assign new_new_n19695__ = ~new_new_n19273__ & po006;
  assign new_new_n19696__ = pi083 & ~po006;
  assign new_new_n19697__ = ~new_new_n19695__ & ~new_new_n19696__;
  assign new_new_n19698__ = ~new_new_n19056__ & ~new_new_n19057__;
  assign new_new_n19699__ = ~new_new_n19697__ & new_new_n19698__;
  assign new_new_n19700__ = new_new_n19697__ & ~new_new_n19698__;
  assign new_new_n19701__ = ~new_new_n19699__ & ~new_new_n19700__;
  assign new_new_n19702__ = ~pi084 & ~new_new_n19701__;
  assign new_new_n19703__ = pi084 & new_new_n19701__;
  assign new_new_n19704__ = ~new_new_n19065__ & ~new_new_n19066__;
  assign new_new_n19705__ = ~new_new_n19271__ & po006;
  assign new_new_n19706__ = pi082 & ~po006;
  assign new_new_n19707__ = ~new_new_n19705__ & ~new_new_n19706__;
  assign new_new_n19708__ = new_new_n19704__ & new_new_n19707__;
  assign new_new_n19709__ = ~new_new_n19704__ & ~new_new_n19707__;
  assign new_new_n19710__ = ~new_new_n19708__ & ~new_new_n19709__;
  assign new_new_n19711__ = ~pi083 & new_new_n19710__;
  assign new_new_n19712__ = pi083 & ~new_new_n19710__;
  assign new_new_n19713__ = new_new_n19269__ & po006;
  assign new_new_n19714__ = pi081 & ~po006;
  assign new_new_n19715__ = ~new_new_n19713__ & ~new_new_n19714__;
  assign new_new_n19716__ = ~new_new_n19074__ & ~new_new_n19075__;
  assign new_new_n19717__ = ~new_new_n19715__ & ~new_new_n19716__;
  assign new_new_n19718__ = new_new_n19715__ & new_new_n19716__;
  assign new_new_n19719__ = ~new_new_n19717__ & ~new_new_n19718__;
  assign new_new_n19720__ = ~pi082 & new_new_n19719__;
  assign new_new_n19721__ = pi082 & ~new_new_n19719__;
  assign new_new_n19722__ = ~new_new_n19083__ & ~new_new_n19084__;
  assign new_new_n19723__ = new_new_n19267__ & po006;
  assign new_new_n19724__ = ~pi080 & ~po006;
  assign new_new_n19725__ = ~new_new_n19723__ & ~new_new_n19724__;
  assign new_new_n19726__ = ~new_new_n19722__ & ~new_new_n19725__;
  assign new_new_n19727__ = new_new_n19722__ & new_new_n19725__;
  assign new_new_n19728__ = ~new_new_n19726__ & ~new_new_n19727__;
  assign new_new_n19729__ = ~pi081 & ~new_new_n19728__;
  assign new_new_n19730__ = pi081 & new_new_n19728__;
  assign new_new_n19731__ = new_new_n19265__ & po006;
  assign new_new_n19732__ = pi079 & ~po006;
  assign new_new_n19733__ = ~new_new_n19731__ & ~new_new_n19732__;
  assign new_new_n19734__ = ~new_new_n19092__ & ~new_new_n19093__;
  assign new_new_n19735__ = ~new_new_n19733__ & ~new_new_n19734__;
  assign new_new_n19736__ = new_new_n19733__ & new_new_n19734__;
  assign new_new_n19737__ = ~new_new_n19735__ & ~new_new_n19736__;
  assign new_new_n19738__ = pi080 & ~new_new_n19737__;
  assign new_new_n19739__ = ~pi080 & new_new_n19737__;
  assign new_new_n19740__ = ~new_new_n19263__ & po006;
  assign new_new_n19741__ = pi078 & ~po006;
  assign new_new_n19742__ = ~new_new_n19740__ & ~new_new_n19741__;
  assign new_new_n19743__ = ~new_new_n19101__ & ~new_new_n19102__;
  assign new_new_n19744__ = ~new_new_n19742__ & new_new_n19743__;
  assign new_new_n19745__ = new_new_n19742__ & ~new_new_n19743__;
  assign new_new_n19746__ = ~new_new_n19744__ & ~new_new_n19745__;
  assign new_new_n19747__ = ~pi079 & ~new_new_n19746__;
  assign new_new_n19748__ = pi079 & new_new_n19746__;
  assign new_new_n19749__ = pi077 & ~new_new_n19261__;
  assign new_new_n19750__ = ~pi077 & new_new_n19261__;
  assign new_new_n19751__ = ~new_new_n19749__ & ~new_new_n19750__;
  assign new_new_n19752__ = po006 & new_new_n19751__;
  assign new_new_n19753__ = new_new_n19109__ & new_new_n19752__;
  assign new_new_n19754__ = ~new_new_n19109__ & ~new_new_n19752__;
  assign new_new_n19755__ = ~new_new_n19753__ & ~new_new_n19754__;
  assign new_new_n19756__ = pi078 & ~new_new_n19755__;
  assign new_new_n19757__ = ~pi078 & new_new_n19755__;
  assign new_new_n19758__ = ~new_new_n19259__ & po006;
  assign new_new_n19759__ = pi076 & ~po006;
  assign new_new_n19760__ = ~new_new_n19758__ & ~new_new_n19759__;
  assign new_new_n19761__ = ~new_new_n19119__ & ~new_new_n19120__;
  assign new_new_n19762__ = ~new_new_n19760__ & new_new_n19761__;
  assign new_new_n19763__ = new_new_n19760__ & ~new_new_n19761__;
  assign new_new_n19764__ = ~new_new_n19762__ & ~new_new_n19763__;
  assign new_new_n19765__ = ~pi077 & ~new_new_n19764__;
  assign new_new_n19766__ = pi077 & new_new_n19764__;
  assign new_new_n19767__ = ~new_new_n19249__ & ~new_new_n19250__;
  assign new_new_n19768__ = po006 & new_new_n19767__;
  assign new_new_n19769__ = new_new_n19257__ & ~new_new_n19768__;
  assign new_new_n19770__ = ~new_new_n19257__ & new_new_n19768__;
  assign new_new_n19771__ = ~new_new_n19769__ & ~new_new_n19770__;
  assign new_new_n19772__ = ~pi076 & new_new_n19771__;
  assign new_new_n19773__ = pi076 & ~new_new_n19771__;
  assign new_new_n19774__ = pi074 & ~new_new_n19246__;
  assign new_new_n19775__ = ~pi074 & new_new_n19246__;
  assign new_new_n19776__ = ~new_new_n19774__ & ~new_new_n19775__;
  assign new_new_n19777__ = po006 & new_new_n19776__;
  assign new_new_n19778__ = ~new_new_n19127__ & new_new_n19777__;
  assign new_new_n19779__ = new_new_n19127__ & ~new_new_n19777__;
  assign new_new_n19780__ = ~new_new_n19778__ & ~new_new_n19779__;
  assign new_new_n19781__ = ~pi075 & ~new_new_n19780__;
  assign new_new_n19782__ = pi075 & new_new_n19780__;
  assign new_new_n19783__ = ~new_new_n19137__ & ~new_new_n19138__;
  assign new_new_n19784__ = ~new_new_n19244__ & po006;
  assign new_new_n19785__ = pi073 & ~po006;
  assign new_new_n19786__ = ~new_new_n19784__ & ~new_new_n19785__;
  assign new_new_n19787__ = new_new_n19783__ & ~new_new_n19786__;
  assign new_new_n19788__ = ~new_new_n19783__ & new_new_n19786__;
  assign new_new_n19789__ = ~new_new_n19787__ & ~new_new_n19788__;
  assign new_new_n19790__ = ~pi074 & ~new_new_n19789__;
  assign new_new_n19791__ = pi074 & new_new_n19789__;
  assign new_new_n19792__ = ~new_new_n19146__ & ~new_new_n19147__;
  assign new_new_n19793__ = ~new_new_n19242__ & po006;
  assign new_new_n19794__ = ~pi072 & ~po006;
  assign new_new_n19795__ = ~new_new_n19793__ & ~new_new_n19794__;
  assign new_new_n19796__ = new_new_n19792__ & ~new_new_n19795__;
  assign new_new_n19797__ = ~new_new_n19792__ & new_new_n19795__;
  assign new_new_n19798__ = ~new_new_n19796__ & ~new_new_n19797__;
  assign new_new_n19799__ = pi073 & ~new_new_n19798__;
  assign new_new_n19800__ = ~pi073 & new_new_n19798__;
  assign new_new_n19801__ = ~new_new_n19164__ & ~new_new_n19165__;
  assign new_new_n19802__ = ~new_new_n19238__ & po006;
  assign new_new_n19803__ = ~pi070 & ~po006;
  assign new_new_n19804__ = ~new_new_n19802__ & ~new_new_n19803__;
  assign new_new_n19805__ = new_new_n19801__ & ~new_new_n19804__;
  assign new_new_n19806__ = ~new_new_n19801__ & new_new_n19804__;
  assign new_new_n19807__ = ~new_new_n19805__ & ~new_new_n19806__;
  assign new_new_n19808__ = pi071 & ~new_new_n19807__;
  assign new_new_n19809__ = ~pi071 & new_new_n19807__;
  assign new_new_n19810__ = ~new_new_n19173__ & ~new_new_n19174__;
  assign new_new_n19811__ = ~new_new_n19236__ & po006;
  assign new_new_n19812__ = pi069 & ~po006;
  assign new_new_n19813__ = ~new_new_n19811__ & ~new_new_n19812__;
  assign new_new_n19814__ = new_new_n19810__ & ~new_new_n19813__;
  assign new_new_n19815__ = ~new_new_n19810__ & new_new_n19813__;
  assign new_new_n19816__ = ~new_new_n19814__ & ~new_new_n19815__;
  assign new_new_n19817__ = pi070 & new_new_n19816__;
  assign new_new_n19818__ = ~pi070 & ~new_new_n19816__;
  assign new_new_n19819__ = ~new_new_n19182__ & ~new_new_n19183__;
  assign new_new_n19820__ = ~new_new_n19234__ & po006;
  assign new_new_n19821__ = pi068 & ~po006;
  assign new_new_n19822__ = ~new_new_n19820__ & ~new_new_n19821__;
  assign new_new_n19823__ = new_new_n19819__ & ~new_new_n19822__;
  assign new_new_n19824__ = ~new_new_n19819__ & new_new_n19822__;
  assign new_new_n19825__ = ~new_new_n19823__ & ~new_new_n19824__;
  assign new_new_n19826__ = pi069 & new_new_n19825__;
  assign new_new_n19827__ = ~pi069 & ~new_new_n19825__;
  assign new_new_n19828__ = ~new_new_n19189__ & ~new_new_n19190__;
  assign new_new_n19829__ = ~new_new_n19232__ & po006;
  assign new_new_n19830__ = pi067 & ~po006;
  assign new_new_n19831__ = ~new_new_n19829__ & ~new_new_n19830__;
  assign new_new_n19832__ = new_new_n19828__ & ~new_new_n19831__;
  assign new_new_n19833__ = ~new_new_n19828__ & new_new_n19831__;
  assign new_new_n19834__ = ~new_new_n19832__ & ~new_new_n19833__;
  assign new_new_n19835__ = pi068 & new_new_n19834__;
  assign new_new_n19836__ = ~pi068 & ~new_new_n19834__;
  assign new_new_n19837__ = ~new_new_n19203__ & ~new_new_n19204__;
  assign new_new_n19838__ = po006 & new_new_n19837__;
  assign new_new_n19839__ = new_new_n19230__ & ~new_new_n19838__;
  assign new_new_n19840__ = ~new_new_n19230__ & new_new_n19838__;
  assign new_new_n19841__ = ~new_new_n19839__ & ~new_new_n19840__;
  assign new_new_n19842__ = pi067 & ~new_new_n19841__;
  assign new_new_n19843__ = ~pi067 & new_new_n19841__;
  assign new_new_n19844__ = pi006 & po006;
  assign new_new_n19845__ = ~pi006 & ~po006;
  assign new_new_n19846__ = ~pi065 & ~new_new_n19844__;
  assign new_new_n19847__ = ~new_new_n19845__ & new_new_n19846__;
  assign new_new_n19848__ = ~pi005 & ~new_new_n19847__;
  assign new_new_n19849__ = pi065 & new_new_n19844__;
  assign new_new_n19850__ = ~new_new_n19848__ & ~new_new_n19849__;
  assign new_new_n19851__ = pi064 & ~new_new_n19850__;
  assign new_new_n19852__ = pi064 & po006;
  assign new_new_n19853__ = ~pi006 & pi065;
  assign new_new_n19854__ = ~new_new_n19852__ & new_new_n19853__;
  assign new_new_n19855__ = ~new_new_n19851__ & ~new_new_n19854__;
  assign new_new_n19856__ = pi066 & ~new_new_n19855__;
  assign new_new_n19857__ = new_new_n426__ & ~po007;
  assign new_new_n19858__ = new_new_n19223__ & po006;
  assign new_new_n19859__ = ~new_new_n19857__ & ~new_new_n19858__;
  assign new_new_n19860__ = ~pi006 & ~new_new_n19859__;
  assign new_new_n19861__ = pi065 & po006;
  assign new_new_n19862__ = po007 & ~new_new_n19861__;
  assign new_new_n19863__ = pi065 & ~new_new_n19199__;
  assign new_new_n19864__ = pi006 & ~new_new_n19863__;
  assign new_new_n19865__ = ~new_new_n19862__ & new_new_n19864__;
  assign new_new_n19866__ = ~new_new_n332__ & po006;
  assign new_new_n19867__ = ~new_new_n19199__ & ~new_new_n19866__;
  assign new_new_n19868__ = ~new_new_n19860__ & ~new_new_n19867__;
  assign new_new_n19869__ = ~new_new_n19865__ & new_new_n19868__;
  assign new_new_n19870__ = ~pi007 & ~new_new_n19869__;
  assign new_new_n19871__ = ~new_new_n19199__ & ~new_new_n19861__;
  assign new_new_n19872__ = pi006 & ~new_new_n19209__;
  assign new_new_n19873__ = pi064 & ~new_new_n19872__;
  assign new_new_n19874__ = ~new_new_n19871__ & ~new_new_n19873__;
  assign new_new_n19875__ = ~pi065 & po006;
  assign new_new_n19876__ = ~po007 & ~new_new_n19875__;
  assign new_new_n19877__ = pi064 & ~new_new_n19844__;
  assign new_new_n19878__ = ~new_new_n19858__ & new_new_n19877__;
  assign new_new_n19879__ = ~new_new_n19876__ & new_new_n19878__;
  assign new_new_n19880__ = ~new_new_n19874__ & ~new_new_n19879__;
  assign new_new_n19881__ = pi007 & ~new_new_n19880__;
  assign new_new_n19882__ = ~new_new_n19870__ & ~new_new_n19881__;
  assign new_new_n19883__ = ~pi066 & new_new_n19855__;
  assign new_new_n19884__ = ~new_new_n19882__ & ~new_new_n19883__;
  assign new_new_n19885__ = ~new_new_n19856__ & ~new_new_n19884__;
  assign new_new_n19886__ = ~new_new_n19843__ & ~new_new_n19885__;
  assign new_new_n19887__ = ~new_new_n19842__ & ~new_new_n19886__;
  assign new_new_n19888__ = ~new_new_n19836__ & ~new_new_n19887__;
  assign new_new_n19889__ = ~new_new_n19835__ & ~new_new_n19888__;
  assign new_new_n19890__ = ~new_new_n19827__ & ~new_new_n19889__;
  assign new_new_n19891__ = ~new_new_n19826__ & ~new_new_n19890__;
  assign new_new_n19892__ = ~new_new_n19818__ & ~new_new_n19891__;
  assign new_new_n19893__ = ~new_new_n19817__ & ~new_new_n19892__;
  assign new_new_n19894__ = ~new_new_n19809__ & ~new_new_n19893__;
  assign new_new_n19895__ = ~new_new_n19808__ & ~new_new_n19894__;
  assign new_new_n19896__ = ~pi072 & new_new_n19895__;
  assign new_new_n19897__ = pi072 & ~new_new_n19895__;
  assign new_new_n19898__ = ~new_new_n19155__ & ~new_new_n19156__;
  assign new_new_n19899__ = ~new_new_n19240__ & po006;
  assign new_new_n19900__ = ~pi071 & ~po006;
  assign new_new_n19901__ = ~new_new_n19899__ & ~new_new_n19900__;
  assign new_new_n19902__ = new_new_n19898__ & ~new_new_n19901__;
  assign new_new_n19903__ = ~new_new_n19898__ & new_new_n19901__;
  assign new_new_n19904__ = ~new_new_n19902__ & ~new_new_n19903__;
  assign new_new_n19905__ = ~new_new_n19897__ & new_new_n19904__;
  assign new_new_n19906__ = ~new_new_n19896__ & ~new_new_n19905__;
  assign new_new_n19907__ = ~new_new_n19800__ & new_new_n19906__;
  assign new_new_n19908__ = ~new_new_n19799__ & ~new_new_n19907__;
  assign new_new_n19909__ = ~new_new_n19791__ & new_new_n19908__;
  assign new_new_n19910__ = ~new_new_n19790__ & ~new_new_n19909__;
  assign new_new_n19911__ = ~new_new_n19782__ & ~new_new_n19910__;
  assign new_new_n19912__ = ~new_new_n19781__ & ~new_new_n19911__;
  assign new_new_n19913__ = ~new_new_n19773__ & ~new_new_n19912__;
  assign new_new_n19914__ = ~new_new_n19772__ & ~new_new_n19913__;
  assign new_new_n19915__ = ~new_new_n19766__ & ~new_new_n19914__;
  assign new_new_n19916__ = ~new_new_n19765__ & ~new_new_n19915__;
  assign new_new_n19917__ = ~new_new_n19757__ & new_new_n19916__;
  assign new_new_n19918__ = ~new_new_n19756__ & ~new_new_n19917__;
  assign new_new_n19919__ = ~new_new_n19748__ & new_new_n19918__;
  assign new_new_n19920__ = ~new_new_n19747__ & ~new_new_n19919__;
  assign new_new_n19921__ = ~new_new_n19739__ & new_new_n19920__;
  assign new_new_n19922__ = ~new_new_n19738__ & ~new_new_n19921__;
  assign new_new_n19923__ = ~new_new_n19730__ & new_new_n19922__;
  assign new_new_n19924__ = ~new_new_n19729__ & ~new_new_n19923__;
  assign new_new_n19925__ = ~new_new_n19721__ & ~new_new_n19924__;
  assign new_new_n19926__ = ~new_new_n19720__ & ~new_new_n19925__;
  assign new_new_n19927__ = ~new_new_n19712__ & ~new_new_n19926__;
  assign new_new_n19928__ = ~new_new_n19711__ & ~new_new_n19927__;
  assign new_new_n19929__ = ~new_new_n19703__ & ~new_new_n19928__;
  assign new_new_n19930__ = ~new_new_n19702__ & ~new_new_n19929__;
  assign new_new_n19931__ = ~new_new_n19694__ & ~new_new_n19930__;
  assign new_new_n19932__ = ~new_new_n19693__ & ~new_new_n19931__;
  assign new_new_n19933__ = ~new_new_n19685__ & ~new_new_n19932__;
  assign new_new_n19934__ = ~new_new_n19684__ & ~new_new_n19933__;
  assign new_new_n19935__ = ~new_new_n19676__ & ~new_new_n19934__;
  assign new_new_n19936__ = ~new_new_n19675__ & ~new_new_n19935__;
  assign new_new_n19937__ = ~new_new_n19667__ & ~new_new_n19936__;
  assign new_new_n19938__ = ~new_new_n19666__ & ~new_new_n19937__;
  assign new_new_n19939__ = ~new_new_n19658__ & new_new_n19938__;
  assign new_new_n19940__ = ~new_new_n19657__ & ~new_new_n19939__;
  assign new_new_n19941__ = ~new_new_n19649__ & ~new_new_n19940__;
  assign new_new_n19942__ = ~new_new_n19648__ & ~new_new_n19941__;
  assign new_new_n19943__ = ~new_new_n19640__ & ~new_new_n19942__;
  assign new_new_n19944__ = ~new_new_n19639__ & ~new_new_n19943__;
  assign new_new_n19945__ = ~new_new_n19631__ & new_new_n19944__;
  assign new_new_n19946__ = ~new_new_n19630__ & ~new_new_n19945__;
  assign new_new_n19947__ = ~new_new_n19622__ & ~new_new_n19946__;
  assign new_new_n19948__ = ~new_new_n19621__ & ~new_new_n19947__;
  assign new_new_n19949__ = ~new_new_n19613__ & new_new_n19948__;
  assign new_new_n19950__ = ~new_new_n19612__ & ~new_new_n19949__;
  assign new_new_n19951__ = ~new_new_n19604__ & ~new_new_n19950__;
  assign new_new_n19952__ = ~new_new_n19603__ & ~new_new_n19951__;
  assign new_new_n19953__ = ~new_new_n19595__ & ~new_new_n19952__;
  assign new_new_n19954__ = ~new_new_n19594__ & ~new_new_n19953__;
  assign new_new_n19955__ = ~new_new_n19586__ & ~new_new_n19954__;
  assign new_new_n19956__ = ~new_new_n19585__ & ~new_new_n19955__;
  assign new_new_n19957__ = ~new_new_n19577__ & new_new_n19956__;
  assign new_new_n19958__ = ~new_new_n19576__ & ~new_new_n19957__;
  assign new_new_n19959__ = ~new_new_n19568__ & ~new_new_n19958__;
  assign new_new_n19960__ = ~new_new_n19567__ & ~new_new_n19959__;
  assign new_new_n19961__ = pi100 & ~new_new_n19558__;
  assign new_new_n19962__ = ~new_new_n19960__ & ~new_new_n19961__;
  assign new_new_n19963__ = ~new_new_n19559__ & ~new_new_n19962__;
  assign new_new_n19964__ = ~new_new_n19551__ & ~new_new_n19963__;
  assign new_new_n19965__ = ~new_new_n19550__ & ~new_new_n19964__;
  assign new_new_n19966__ = ~new_new_n19542__ & new_new_n19965__;
  assign new_new_n19967__ = ~new_new_n19541__ & ~new_new_n19966__;
  assign new_new_n19968__ = ~new_new_n19533__ & new_new_n19967__;
  assign new_new_n19969__ = ~new_new_n19532__ & ~new_new_n19968__;
  assign new_new_n19970__ = ~new_new_n19524__ & ~new_new_n19969__;
  assign new_new_n19971__ = ~new_new_n19523__ & ~new_new_n19970__;
  assign new_new_n19972__ = ~new_new_n19515__ & ~new_new_n19971__;
  assign new_new_n19973__ = ~new_new_n19514__ & ~new_new_n19972__;
  assign new_new_n19974__ = ~new_new_n19506__ & ~new_new_n19973__;
  assign new_new_n19975__ = ~new_new_n19505__ & ~new_new_n19974__;
  assign new_new_n19976__ = ~new_new_n19497__ & ~new_new_n19975__;
  assign new_new_n19977__ = ~new_new_n19496__ & ~new_new_n19976__;
  assign new_new_n19978__ = ~new_new_n19488__ & ~new_new_n19977__;
  assign new_new_n19979__ = ~new_new_n19487__ & ~new_new_n19978__;
  assign new_new_n19980__ = ~new_new_n19479__ & new_new_n19979__;
  assign new_new_n19981__ = ~new_new_n19478__ & ~new_new_n19980__;
  assign new_new_n19982__ = ~new_new_n19470__ & ~new_new_n19981__;
  assign new_new_n19983__ = ~new_new_n19469__ & ~new_new_n19982__;
  assign new_new_n19984__ = ~new_new_n19461__ & ~new_new_n19983__;
  assign new_new_n19985__ = ~new_new_n19460__ & ~new_new_n19984__;
  assign new_new_n19986__ = ~new_new_n19454__ & new_new_n19985__;
  assign new_new_n19987__ = ~new_new_n19453__ & ~new_new_n19986__;
  assign new_new_n19988__ = ~new_new_n19445__ & ~new_new_n19987__;
  assign new_new_n19989__ = ~new_new_n19444__ & ~new_new_n19988__;
  assign new_new_n19990__ = ~new_new_n19436__ & new_new_n19989__;
  assign new_new_n19991__ = ~new_new_n19435__ & ~new_new_n19990__;
  assign new_new_n19992__ = ~new_new_n19427__ & ~new_new_n19991__;
  assign new_new_n19993__ = ~new_new_n19426__ & ~new_new_n19992__;
  assign new_new_n19994__ = ~new_new_n19418__ & ~new_new_n19993__;
  assign new_new_n19995__ = ~new_new_n19417__ & ~new_new_n19994__;
  assign new_new_n19996__ = ~new_new_n19409__ & ~new_new_n19995__;
  assign new_new_n19997__ = ~new_new_n19408__ & ~new_new_n19996__;
  assign new_new_n19998__ = ~new_new_n19400__ & ~new_new_n19997__;
  assign new_new_n19999__ = ~new_new_n19399__ & ~new_new_n19998__;
  assign new_new_n20000__ = ~new_new_n19391__ & new_new_n19999__;
  assign new_new_n20001__ = ~new_new_n19390__ & ~new_new_n20000__;
  assign new_new_n20002__ = ~new_new_n19382__ & ~new_new_n20001__;
  assign new_new_n20003__ = ~new_new_n19381__ & ~new_new_n20002__;
  assign new_new_n20004__ = ~new_new_n19373__ & ~new_new_n20003__;
  assign new_new_n20005__ = ~pi121 & ~new_new_n19372__;
  assign new_new_n20006__ = pi121 & ~new_new_n19358__;
  assign new_new_n20007__ = ~new_new_n19359__ & ~new_new_n20006__;
  assign new_new_n20008__ = ~pi122 & new_new_n18717__;
  assign new_new_n20009__ = ~new_new_n20007__ & new_new_n20008__;
  assign new_new_n20010__ = ~new_new_n20005__ & ~new_new_n20009__;
  assign new_new_n20011__ = ~new_new_n20004__ & new_new_n20010__;
  assign new_new_n20012__ = pi122 & ~new_new_n18720__;
  assign new_new_n20013__ = ~pi123 & new_new_n262__;
  assign new_new_n20014__ = ~new_new_n20012__ & new_new_n20013__;
  assign po005 = ~new_new_n20011__ & new_new_n20014__;
  assign new_new_n20016__ = ~new_new_n264__ & po005;
  assign new_new_n20017__ = new_new_n18717__ & ~new_new_n19360__;
  assign new_new_n20018__ = ~new_new_n20016__ & new_new_n20017__;
  assign new_new_n20019__ = pi127 & ~new_new_n20018__;
  assign new_new_n20020__ = ~new_new_n19381__ & ~new_new_n19382__;
  assign new_new_n20021__ = ~new_new_n20001__ & po005;
  assign new_new_n20022__ = ~pi120 & ~po005;
  assign new_new_n20023__ = ~new_new_n20021__ & ~new_new_n20022__;
  assign new_new_n20024__ = new_new_n20020__ & new_new_n20023__;
  assign new_new_n20025__ = ~new_new_n20020__ & ~new_new_n20023__;
  assign new_new_n20026__ = ~new_new_n20024__ & ~new_new_n20025__;
  assign new_new_n20027__ = ~pi121 & ~new_new_n20026__;
  assign new_new_n20028__ = pi121 & new_new_n20026__;
  assign new_new_n20029__ = new_new_n19999__ & po005;
  assign new_new_n20030__ = ~pi119 & ~po005;
  assign new_new_n20031__ = ~new_new_n20029__ & ~new_new_n20030__;
  assign new_new_n20032__ = ~new_new_n19390__ & ~new_new_n19391__;
  assign new_new_n20033__ = ~new_new_n20031__ & ~new_new_n20032__;
  assign new_new_n20034__ = new_new_n20031__ & new_new_n20032__;
  assign new_new_n20035__ = ~new_new_n20033__ & ~new_new_n20034__;
  assign new_new_n20036__ = ~pi120 & ~new_new_n20035__;
  assign new_new_n20037__ = pi120 & new_new_n20035__;
  assign new_new_n20038__ = ~new_new_n19997__ & po005;
  assign new_new_n20039__ = pi118 & ~po005;
  assign new_new_n20040__ = ~new_new_n20038__ & ~new_new_n20039__;
  assign new_new_n20041__ = ~new_new_n19399__ & ~new_new_n19400__;
  assign new_new_n20042__ = ~new_new_n20040__ & new_new_n20041__;
  assign new_new_n20043__ = new_new_n20040__ & ~new_new_n20041__;
  assign new_new_n20044__ = ~new_new_n20042__ & ~new_new_n20043__;
  assign new_new_n20045__ = ~pi119 & ~new_new_n20044__;
  assign new_new_n20046__ = pi119 & new_new_n20044__;
  assign new_new_n20047__ = ~new_new_n19995__ & po005;
  assign new_new_n20048__ = pi117 & ~po005;
  assign new_new_n20049__ = ~new_new_n20047__ & ~new_new_n20048__;
  assign new_new_n20050__ = ~new_new_n19408__ & ~new_new_n19409__;
  assign new_new_n20051__ = ~new_new_n20049__ & new_new_n20050__;
  assign new_new_n20052__ = new_new_n20049__ & ~new_new_n20050__;
  assign new_new_n20053__ = ~new_new_n20051__ & ~new_new_n20052__;
  assign new_new_n20054__ = ~pi118 & ~new_new_n20053__;
  assign new_new_n20055__ = pi118 & new_new_n20053__;
  assign new_new_n20056__ = ~new_new_n19417__ & ~new_new_n19418__;
  assign new_new_n20057__ = pi116 & ~po005;
  assign new_new_n20058__ = ~new_new_n19993__ & po005;
  assign new_new_n20059__ = ~new_new_n20057__ & ~new_new_n20058__;
  assign new_new_n20060__ = new_new_n20056__ & new_new_n20059__;
  assign new_new_n20061__ = ~new_new_n20056__ & ~new_new_n20059__;
  assign new_new_n20062__ = ~new_new_n20060__ & ~new_new_n20061__;
  assign new_new_n20063__ = pi117 & ~new_new_n20062__;
  assign new_new_n20064__ = ~pi117 & new_new_n20062__;
  assign new_new_n20065__ = ~new_new_n19991__ & po005;
  assign new_new_n20066__ = pi115 & ~po005;
  assign new_new_n20067__ = ~new_new_n20065__ & ~new_new_n20066__;
  assign new_new_n20068__ = ~new_new_n19426__ & ~new_new_n19427__;
  assign new_new_n20069__ = ~new_new_n20067__ & new_new_n20068__;
  assign new_new_n20070__ = new_new_n20067__ & ~new_new_n20068__;
  assign new_new_n20071__ = ~new_new_n20069__ & ~new_new_n20070__;
  assign new_new_n20072__ = pi116 & new_new_n20071__;
  assign new_new_n20073__ = ~pi116 & ~new_new_n20071__;
  assign new_new_n20074__ = ~new_new_n19435__ & ~new_new_n19436__;
  assign new_new_n20075__ = ~new_new_n19989__ & po005;
  assign new_new_n20076__ = ~pi114 & ~po005;
  assign new_new_n20077__ = ~new_new_n20075__ & ~new_new_n20076__;
  assign new_new_n20078__ = new_new_n20074__ & ~new_new_n20077__;
  assign new_new_n20079__ = ~new_new_n20074__ & new_new_n20077__;
  assign new_new_n20080__ = ~new_new_n20078__ & ~new_new_n20079__;
  assign new_new_n20081__ = pi115 & ~new_new_n20080__;
  assign new_new_n20082__ = ~pi115 & new_new_n20080__;
  assign new_new_n20083__ = ~new_new_n19444__ & ~new_new_n19445__;
  assign new_new_n20084__ = ~new_new_n19987__ & po005;
  assign new_new_n20085__ = ~pi113 & ~po005;
  assign new_new_n20086__ = ~new_new_n20084__ & ~new_new_n20085__;
  assign new_new_n20087__ = ~new_new_n20083__ & ~new_new_n20086__;
  assign new_new_n20088__ = new_new_n20083__ & new_new_n20086__;
  assign new_new_n20089__ = ~new_new_n20087__ & ~new_new_n20088__;
  assign new_new_n20090__ = pi114 & new_new_n20089__;
  assign new_new_n20091__ = ~pi114 & ~new_new_n20089__;
  assign new_new_n20092__ = ~new_new_n19453__ & ~new_new_n19454__;
  assign new_new_n20093__ = pi112 & ~po005;
  assign new_new_n20094__ = ~new_new_n19985__ & po005;
  assign new_new_n20095__ = ~new_new_n20093__ & ~new_new_n20094__;
  assign new_new_n20096__ = new_new_n20092__ & ~new_new_n20095__;
  assign new_new_n20097__ = ~new_new_n20092__ & new_new_n20095__;
  assign new_new_n20098__ = ~new_new_n20096__ & ~new_new_n20097__;
  assign new_new_n20099__ = pi113 & new_new_n20098__;
  assign new_new_n20100__ = ~pi113 & ~new_new_n20098__;
  assign new_new_n20101__ = pi111 & ~new_new_n19983__;
  assign new_new_n20102__ = ~pi111 & new_new_n19983__;
  assign new_new_n20103__ = ~new_new_n20101__ & ~new_new_n20102__;
  assign new_new_n20104__ = po005 & new_new_n20103__;
  assign new_new_n20105__ = new_new_n19459__ & new_new_n20104__;
  assign new_new_n20106__ = ~new_new_n19459__ & ~new_new_n20104__;
  assign new_new_n20107__ = ~new_new_n20105__ & ~new_new_n20106__;
  assign new_new_n20108__ = pi112 & ~new_new_n20107__;
  assign new_new_n20109__ = ~pi112 & new_new_n20107__;
  assign new_new_n20110__ = pi110 & ~new_new_n19981__;
  assign new_new_n20111__ = ~pi110 & new_new_n19981__;
  assign new_new_n20112__ = ~new_new_n20110__ & ~new_new_n20111__;
  assign new_new_n20113__ = po005 & new_new_n20112__;
  assign new_new_n20114__ = new_new_n19468__ & new_new_n20113__;
  assign new_new_n20115__ = ~new_new_n19468__ & ~new_new_n20113__;
  assign new_new_n20116__ = ~new_new_n20114__ & ~new_new_n20115__;
  assign new_new_n20117__ = pi111 & ~new_new_n20116__;
  assign new_new_n20118__ = ~pi111 & new_new_n20116__;
  assign new_new_n20119__ = ~new_new_n19478__ & ~new_new_n19479__;
  assign new_new_n20120__ = ~new_new_n19979__ & po005;
  assign new_new_n20121__ = ~pi109 & ~po005;
  assign new_new_n20122__ = ~new_new_n20120__ & ~new_new_n20121__;
  assign new_new_n20123__ = new_new_n20119__ & ~new_new_n20122__;
  assign new_new_n20124__ = ~new_new_n20119__ & new_new_n20122__;
  assign new_new_n20125__ = ~new_new_n20123__ & ~new_new_n20124__;
  assign new_new_n20126__ = pi110 & ~new_new_n20125__;
  assign new_new_n20127__ = ~pi108 & ~new_new_n19977__;
  assign new_new_n20128__ = pi108 & new_new_n19977__;
  assign new_new_n20129__ = ~new_new_n20127__ & ~new_new_n20128__;
  assign new_new_n20130__ = po005 & new_new_n20129__;
  assign new_new_n20131__ = new_new_n19486__ & new_new_n20130__;
  assign new_new_n20132__ = ~new_new_n19486__ & ~new_new_n20130__;
  assign new_new_n20133__ = ~new_new_n20131__ & ~new_new_n20132__;
  assign new_new_n20134__ = ~pi109 & ~new_new_n20133__;
  assign new_new_n20135__ = pi109 & new_new_n20133__;
  assign new_new_n20136__ = ~new_new_n19496__ & ~new_new_n19497__;
  assign new_new_n20137__ = ~new_new_n19975__ & po005;
  assign new_new_n20138__ = ~pi107 & ~po005;
  assign new_new_n20139__ = ~new_new_n20137__ & ~new_new_n20138__;
  assign new_new_n20140__ = ~new_new_n20136__ & ~new_new_n20139__;
  assign new_new_n20141__ = new_new_n20136__ & new_new_n20139__;
  assign new_new_n20142__ = ~new_new_n20140__ & ~new_new_n20141__;
  assign new_new_n20143__ = ~pi108 & ~new_new_n20142__;
  assign new_new_n20144__ = pi108 & new_new_n20142__;
  assign new_new_n20145__ = new_new_n19973__ & po005;
  assign new_new_n20146__ = pi106 & ~po005;
  assign new_new_n20147__ = ~new_new_n20145__ & ~new_new_n20146__;
  assign new_new_n20148__ = ~new_new_n19505__ & ~new_new_n19506__;
  assign new_new_n20149__ = ~new_new_n20147__ & ~new_new_n20148__;
  assign new_new_n20150__ = new_new_n20147__ & new_new_n20148__;
  assign new_new_n20151__ = ~new_new_n20149__ & ~new_new_n20150__;
  assign new_new_n20152__ = ~pi107 & new_new_n20151__;
  assign new_new_n20153__ = pi107 & ~new_new_n20151__;
  assign new_new_n20154__ = ~new_new_n19514__ & ~new_new_n19515__;
  assign new_new_n20155__ = ~new_new_n19971__ & po005;
  assign new_new_n20156__ = ~pi105 & ~po005;
  assign new_new_n20157__ = ~new_new_n20155__ & ~new_new_n20156__;
  assign new_new_n20158__ = new_new_n20154__ & ~new_new_n20157__;
  assign new_new_n20159__ = ~new_new_n20154__ & new_new_n20157__;
  assign new_new_n20160__ = ~new_new_n20158__ & ~new_new_n20159__;
  assign new_new_n20161__ = ~pi106 & new_new_n20160__;
  assign new_new_n20162__ = pi106 & ~new_new_n20160__;
  assign new_new_n20163__ = ~pi104 & ~new_new_n19969__;
  assign new_new_n20164__ = pi104 & new_new_n19969__;
  assign new_new_n20165__ = ~new_new_n20163__ & ~new_new_n20164__;
  assign new_new_n20166__ = po005 & new_new_n20165__;
  assign new_new_n20167__ = new_new_n19522__ & new_new_n20166__;
  assign new_new_n20168__ = ~new_new_n19522__ & ~new_new_n20166__;
  assign new_new_n20169__ = ~new_new_n20167__ & ~new_new_n20168__;
  assign new_new_n20170__ = ~pi105 & ~new_new_n20169__;
  assign new_new_n20171__ = pi105 & new_new_n20169__;
  assign new_new_n20172__ = ~new_new_n19532__ & ~new_new_n19533__;
  assign new_new_n20173__ = pi103 & ~po005;
  assign new_new_n20174__ = ~new_new_n19967__ & po005;
  assign new_new_n20175__ = ~new_new_n20173__ & ~new_new_n20174__;
  assign new_new_n20176__ = new_new_n20172__ & ~new_new_n20175__;
  assign new_new_n20177__ = ~new_new_n20172__ & new_new_n20175__;
  assign new_new_n20178__ = ~new_new_n20176__ & ~new_new_n20177__;
  assign new_new_n20179__ = pi104 & new_new_n20178__;
  assign new_new_n20180__ = ~pi104 & ~new_new_n20178__;
  assign new_new_n20181__ = ~new_new_n19541__ & ~new_new_n19542__;
  assign new_new_n20182__ = ~new_new_n19965__ & po005;
  assign new_new_n20183__ = ~pi102 & ~po005;
  assign new_new_n20184__ = ~new_new_n20182__ & ~new_new_n20183__;
  assign new_new_n20185__ = new_new_n20181__ & ~new_new_n20184__;
  assign new_new_n20186__ = ~new_new_n20181__ & new_new_n20184__;
  assign new_new_n20187__ = ~new_new_n20185__ & ~new_new_n20186__;
  assign new_new_n20188__ = pi103 & ~new_new_n20187__;
  assign new_new_n20189__ = ~pi103 & new_new_n20187__;
  assign new_new_n20190__ = ~new_new_n19550__ & ~new_new_n19551__;
  assign new_new_n20191__ = ~new_new_n19963__ & po005;
  assign new_new_n20192__ = ~pi101 & ~po005;
  assign new_new_n20193__ = ~new_new_n20191__ & ~new_new_n20192__;
  assign new_new_n20194__ = new_new_n20190__ & ~new_new_n20193__;
  assign new_new_n20195__ = ~new_new_n20190__ & new_new_n20193__;
  assign new_new_n20196__ = ~new_new_n20194__ & ~new_new_n20195__;
  assign new_new_n20197__ = pi102 & ~new_new_n20196__;
  assign new_new_n20198__ = ~pi102 & new_new_n20196__;
  assign new_new_n20199__ = ~new_new_n19559__ & ~new_new_n19961__;
  assign new_new_n20200__ = ~new_new_n19960__ & po005;
  assign new_new_n20201__ = ~pi100 & ~po005;
  assign new_new_n20202__ = ~new_new_n20200__ & ~new_new_n20201__;
  assign new_new_n20203__ = new_new_n20199__ & ~new_new_n20202__;
  assign new_new_n20204__ = ~new_new_n20199__ & new_new_n20202__;
  assign new_new_n20205__ = ~new_new_n20203__ & ~new_new_n20204__;
  assign new_new_n20206__ = pi101 & ~new_new_n20205__;
  assign new_new_n20207__ = ~pi101 & new_new_n20205__;
  assign new_new_n20208__ = ~pi099 & ~new_new_n19958__;
  assign new_new_n20209__ = pi099 & new_new_n19958__;
  assign new_new_n20210__ = ~new_new_n20208__ & ~new_new_n20209__;
  assign new_new_n20211__ = po005 & new_new_n20210__;
  assign new_new_n20212__ = new_new_n19566__ & ~new_new_n20211__;
  assign new_new_n20213__ = ~new_new_n19566__ & new_new_n20211__;
  assign new_new_n20214__ = ~new_new_n20212__ & ~new_new_n20213__;
  assign new_new_n20215__ = pi100 & ~new_new_n20214__;
  assign new_new_n20216__ = ~pi100 & new_new_n20214__;
  assign new_new_n20217__ = ~new_new_n19576__ & ~new_new_n19577__;
  assign new_new_n20218__ = new_new_n19956__ & po005;
  assign new_new_n20219__ = ~pi098 & ~po005;
  assign new_new_n20220__ = ~new_new_n20218__ & ~new_new_n20219__;
  assign new_new_n20221__ = ~new_new_n20217__ & ~new_new_n20220__;
  assign new_new_n20222__ = new_new_n20217__ & new_new_n20220__;
  assign new_new_n20223__ = ~new_new_n20221__ & ~new_new_n20222__;
  assign new_new_n20224__ = pi099 & new_new_n20223__;
  assign new_new_n20225__ = ~pi099 & ~new_new_n20223__;
  assign new_new_n20226__ = new_new_n19954__ & po005;
  assign new_new_n20227__ = ~pi097 & ~po005;
  assign new_new_n20228__ = ~new_new_n20226__ & ~new_new_n20227__;
  assign new_new_n20229__ = ~new_new_n19585__ & ~new_new_n19586__;
  assign new_new_n20230__ = ~new_new_n20228__ & ~new_new_n20229__;
  assign new_new_n20231__ = new_new_n20228__ & new_new_n20229__;
  assign new_new_n20232__ = ~new_new_n20230__ & ~new_new_n20231__;
  assign new_new_n20233__ = pi098 & new_new_n20232__;
  assign new_new_n20234__ = ~pi098 & ~new_new_n20232__;
  assign new_new_n20235__ = ~new_new_n19952__ & po005;
  assign new_new_n20236__ = pi096 & ~po005;
  assign new_new_n20237__ = ~new_new_n20235__ & ~new_new_n20236__;
  assign new_new_n20238__ = ~new_new_n19594__ & ~new_new_n19595__;
  assign new_new_n20239__ = ~new_new_n20237__ & new_new_n20238__;
  assign new_new_n20240__ = new_new_n20237__ & ~new_new_n20238__;
  assign new_new_n20241__ = ~new_new_n20239__ & ~new_new_n20240__;
  assign new_new_n20242__ = pi097 & new_new_n20241__;
  assign new_new_n20243__ = ~pi097 & ~new_new_n20241__;
  assign new_new_n20244__ = pi095 & ~new_new_n19950__;
  assign new_new_n20245__ = ~pi095 & new_new_n19950__;
  assign new_new_n20246__ = ~new_new_n20244__ & ~new_new_n20245__;
  assign new_new_n20247__ = po005 & new_new_n20246__;
  assign new_new_n20248__ = new_new_n19602__ & new_new_n20247__;
  assign new_new_n20249__ = ~new_new_n19602__ & ~new_new_n20247__;
  assign new_new_n20250__ = ~new_new_n20248__ & ~new_new_n20249__;
  assign new_new_n20251__ = pi096 & ~new_new_n20250__;
  assign new_new_n20252__ = ~pi096 & new_new_n20250__;
  assign new_new_n20253__ = ~new_new_n19612__ & ~new_new_n19613__;
  assign new_new_n20254__ = ~new_new_n19948__ & po005;
  assign new_new_n20255__ = ~pi094 & ~po005;
  assign new_new_n20256__ = ~new_new_n20254__ & ~new_new_n20255__;
  assign new_new_n20257__ = new_new_n20253__ & ~new_new_n20256__;
  assign new_new_n20258__ = ~new_new_n20253__ & new_new_n20256__;
  assign new_new_n20259__ = ~new_new_n20257__ & ~new_new_n20258__;
  assign new_new_n20260__ = pi095 & ~new_new_n20259__;
  assign new_new_n20261__ = ~pi095 & new_new_n20259__;
  assign new_new_n20262__ = ~pi093 & ~new_new_n19946__;
  assign new_new_n20263__ = pi093 & new_new_n19946__;
  assign new_new_n20264__ = ~new_new_n20262__ & ~new_new_n20263__;
  assign new_new_n20265__ = po005 & new_new_n20264__;
  assign new_new_n20266__ = new_new_n19620__ & new_new_n20265__;
  assign new_new_n20267__ = ~new_new_n19620__ & ~new_new_n20265__;
  assign new_new_n20268__ = ~new_new_n20266__ & ~new_new_n20267__;
  assign new_new_n20269__ = ~pi094 & ~new_new_n20268__;
  assign new_new_n20270__ = pi094 & new_new_n20268__;
  assign new_new_n20271__ = ~new_new_n19944__ & po005;
  assign new_new_n20272__ = pi092 & ~po005;
  assign new_new_n20273__ = ~new_new_n20271__ & ~new_new_n20272__;
  assign new_new_n20274__ = ~new_new_n19630__ & ~new_new_n19631__;
  assign new_new_n20275__ = ~new_new_n20273__ & new_new_n20274__;
  assign new_new_n20276__ = new_new_n20273__ & ~new_new_n20274__;
  assign new_new_n20277__ = ~new_new_n20275__ & ~new_new_n20276__;
  assign new_new_n20278__ = ~pi093 & ~new_new_n20277__;
  assign new_new_n20279__ = pi093 & new_new_n20277__;
  assign new_new_n20280__ = pi091 & ~new_new_n19942__;
  assign new_new_n20281__ = ~pi091 & new_new_n19942__;
  assign new_new_n20282__ = ~new_new_n20280__ & ~new_new_n20281__;
  assign new_new_n20283__ = po005 & new_new_n20282__;
  assign new_new_n20284__ = new_new_n19638__ & new_new_n20283__;
  assign new_new_n20285__ = ~new_new_n19638__ & ~new_new_n20283__;
  assign new_new_n20286__ = ~new_new_n20284__ & ~new_new_n20285__;
  assign new_new_n20287__ = pi092 & ~new_new_n20286__;
  assign new_new_n20288__ = ~pi092 & new_new_n20286__;
  assign new_new_n20289__ = ~new_new_n19648__ & ~new_new_n19649__;
  assign new_new_n20290__ = pi090 & ~po005;
  assign new_new_n20291__ = ~new_new_n19940__ & po005;
  assign new_new_n20292__ = ~new_new_n20290__ & ~new_new_n20291__;
  assign new_new_n20293__ = new_new_n20289__ & ~new_new_n20292__;
  assign new_new_n20294__ = ~new_new_n20289__ & new_new_n20292__;
  assign new_new_n20295__ = ~new_new_n20293__ & ~new_new_n20294__;
  assign new_new_n20296__ = ~pi091 & ~new_new_n20295__;
  assign new_new_n20297__ = pi091 & new_new_n20295__;
  assign new_new_n20298__ = ~new_new_n19657__ & ~new_new_n19658__;
  assign new_new_n20299__ = ~new_new_n19938__ & po005;
  assign new_new_n20300__ = ~pi089 & ~po005;
  assign new_new_n20301__ = ~new_new_n20299__ & ~new_new_n20300__;
  assign new_new_n20302__ = new_new_n20298__ & ~new_new_n20301__;
  assign new_new_n20303__ = ~new_new_n20298__ & new_new_n20301__;
  assign new_new_n20304__ = ~new_new_n20302__ & ~new_new_n20303__;
  assign new_new_n20305__ = ~pi090 & new_new_n20304__;
  assign new_new_n20306__ = pi090 & ~new_new_n20304__;
  assign new_new_n20307__ = ~pi088 & ~new_new_n19936__;
  assign new_new_n20308__ = pi088 & new_new_n19936__;
  assign new_new_n20309__ = ~new_new_n20307__ & ~new_new_n20308__;
  assign new_new_n20310__ = po005 & new_new_n20309__;
  assign new_new_n20311__ = new_new_n19665__ & new_new_n20310__;
  assign new_new_n20312__ = ~new_new_n19665__ & ~new_new_n20310__;
  assign new_new_n20313__ = ~new_new_n20311__ & ~new_new_n20312__;
  assign new_new_n20314__ = ~pi089 & ~new_new_n20313__;
  assign new_new_n20315__ = pi089 & new_new_n20313__;
  assign new_new_n20316__ = ~new_new_n19675__ & ~new_new_n19676__;
  assign new_new_n20317__ = ~new_new_n19934__ & po005;
  assign new_new_n20318__ = ~pi087 & ~po005;
  assign new_new_n20319__ = ~new_new_n20317__ & ~new_new_n20318__;
  assign new_new_n20320__ = new_new_n20316__ & ~new_new_n20319__;
  assign new_new_n20321__ = ~new_new_n20316__ & new_new_n20319__;
  assign new_new_n20322__ = ~new_new_n20320__ & ~new_new_n20321__;
  assign new_new_n20323__ = pi088 & ~new_new_n20322__;
  assign new_new_n20324__ = ~pi088 & new_new_n20322__;
  assign new_new_n20325__ = ~new_new_n19684__ & ~new_new_n19685__;
  assign new_new_n20326__ = ~new_new_n19932__ & po005;
  assign new_new_n20327__ = ~pi086 & ~po005;
  assign new_new_n20328__ = ~new_new_n20326__ & ~new_new_n20327__;
  assign new_new_n20329__ = new_new_n20325__ & ~new_new_n20328__;
  assign new_new_n20330__ = ~new_new_n20325__ & new_new_n20328__;
  assign new_new_n20331__ = ~new_new_n20329__ & ~new_new_n20330__;
  assign new_new_n20332__ = pi087 & ~new_new_n20331__;
  assign new_new_n20333__ = ~pi087 & new_new_n20331__;
  assign new_new_n20334__ = ~pi085 & ~new_new_n19930__;
  assign new_new_n20335__ = pi085 & new_new_n19930__;
  assign new_new_n20336__ = ~new_new_n20334__ & ~new_new_n20335__;
  assign new_new_n20337__ = po005 & new_new_n20336__;
  assign new_new_n20338__ = new_new_n19692__ & new_new_n20337__;
  assign new_new_n20339__ = ~new_new_n19692__ & ~new_new_n20337__;
  assign new_new_n20340__ = ~new_new_n20338__ & ~new_new_n20339__;
  assign new_new_n20341__ = pi086 & new_new_n20340__;
  assign new_new_n20342__ = ~pi086 & ~new_new_n20340__;
  assign new_new_n20343__ = ~pi084 & ~new_new_n19928__;
  assign new_new_n20344__ = pi084 & new_new_n19928__;
  assign new_new_n20345__ = ~new_new_n20343__ & ~new_new_n20344__;
  assign new_new_n20346__ = po005 & new_new_n20345__;
  assign new_new_n20347__ = new_new_n19701__ & new_new_n20346__;
  assign new_new_n20348__ = ~new_new_n19701__ & ~new_new_n20346__;
  assign new_new_n20349__ = ~new_new_n20347__ & ~new_new_n20348__;
  assign new_new_n20350__ = pi085 & new_new_n20349__;
  assign new_new_n20351__ = ~pi085 & ~new_new_n20349__;
  assign new_new_n20352__ = ~new_new_n19711__ & ~new_new_n19712__;
  assign new_new_n20353__ = ~new_new_n19926__ & po005;
  assign new_new_n20354__ = ~pi083 & ~po005;
  assign new_new_n20355__ = ~new_new_n20353__ & ~new_new_n20354__;
  assign new_new_n20356__ = new_new_n20352__ & ~new_new_n20355__;
  assign new_new_n20357__ = ~new_new_n20352__ & new_new_n20355__;
  assign new_new_n20358__ = ~new_new_n20356__ & ~new_new_n20357__;
  assign new_new_n20359__ = pi084 & ~new_new_n20358__;
  assign new_new_n20360__ = ~pi084 & new_new_n20358__;
  assign new_new_n20361__ = ~new_new_n19720__ & ~new_new_n19721__;
  assign new_new_n20362__ = ~new_new_n19924__ & po005;
  assign new_new_n20363__ = ~pi082 & ~po005;
  assign new_new_n20364__ = ~new_new_n20362__ & ~new_new_n20363__;
  assign new_new_n20365__ = new_new_n20361__ & ~new_new_n20364__;
  assign new_new_n20366__ = ~new_new_n20361__ & new_new_n20364__;
  assign new_new_n20367__ = ~new_new_n20365__ & ~new_new_n20366__;
  assign new_new_n20368__ = pi083 & ~new_new_n20367__;
  assign new_new_n20369__ = ~pi083 & new_new_n20367__;
  assign new_new_n20370__ = ~new_new_n19729__ & ~new_new_n19730__;
  assign new_new_n20371__ = new_new_n19922__ & po005;
  assign new_new_n20372__ = ~pi081 & ~po005;
  assign new_new_n20373__ = ~new_new_n20371__ & ~new_new_n20372__;
  assign new_new_n20374__ = ~new_new_n20370__ & ~new_new_n20373__;
  assign new_new_n20375__ = new_new_n20370__ & new_new_n20373__;
  assign new_new_n20376__ = ~new_new_n20374__ & ~new_new_n20375__;
  assign new_new_n20377__ = pi082 & new_new_n20376__;
  assign new_new_n20378__ = ~pi082 & ~new_new_n20376__;
  assign new_new_n20379__ = new_new_n19920__ & po005;
  assign new_new_n20380__ = pi080 & ~po005;
  assign new_new_n20381__ = ~new_new_n20379__ & ~new_new_n20380__;
  assign new_new_n20382__ = ~new_new_n19738__ & ~new_new_n19739__;
  assign new_new_n20383__ = ~new_new_n20381__ & ~new_new_n20382__;
  assign new_new_n20384__ = new_new_n20381__ & new_new_n20382__;
  assign new_new_n20385__ = ~new_new_n20383__ & ~new_new_n20384__;
  assign new_new_n20386__ = pi081 & ~new_new_n20385__;
  assign new_new_n20387__ = ~pi081 & new_new_n20385__;
  assign new_new_n20388__ = ~new_new_n19747__ & ~new_new_n19748__;
  assign new_new_n20389__ = pi079 & ~po005;
  assign new_new_n20390__ = ~new_new_n19918__ & po005;
  assign new_new_n20391__ = ~new_new_n20389__ & ~new_new_n20390__;
  assign new_new_n20392__ = new_new_n20388__ & ~new_new_n20391__;
  assign new_new_n20393__ = ~new_new_n20388__ & new_new_n20391__;
  assign new_new_n20394__ = ~new_new_n20392__ & ~new_new_n20393__;
  assign new_new_n20395__ = pi080 & new_new_n20394__;
  assign new_new_n20396__ = ~pi080 & ~new_new_n20394__;
  assign new_new_n20397__ = new_new_n19916__ & po005;
  assign new_new_n20398__ = pi078 & ~po005;
  assign new_new_n20399__ = ~new_new_n20397__ & ~new_new_n20398__;
  assign new_new_n20400__ = ~new_new_n19756__ & ~new_new_n19757__;
  assign new_new_n20401__ = ~new_new_n20399__ & ~new_new_n20400__;
  assign new_new_n20402__ = new_new_n20399__ & new_new_n20400__;
  assign new_new_n20403__ = ~new_new_n20401__ & ~new_new_n20402__;
  assign new_new_n20404__ = pi079 & ~new_new_n20403__;
  assign new_new_n20405__ = ~pi079 & new_new_n20403__;
  assign new_new_n20406__ = ~pi077 & ~new_new_n19914__;
  assign new_new_n20407__ = pi077 & new_new_n19914__;
  assign new_new_n20408__ = ~new_new_n20406__ & ~new_new_n20407__;
  assign new_new_n20409__ = po005 & new_new_n20408__;
  assign new_new_n20410__ = new_new_n19764__ & new_new_n20409__;
  assign new_new_n20411__ = ~new_new_n19764__ & ~new_new_n20409__;
  assign new_new_n20412__ = ~new_new_n20410__ & ~new_new_n20411__;
  assign new_new_n20413__ = pi078 & new_new_n20412__;
  assign new_new_n20414__ = ~pi078 & ~new_new_n20412__;
  assign new_new_n20415__ = ~new_new_n19772__ & ~new_new_n19773__;
  assign new_new_n20416__ = ~new_new_n19912__ & po005;
  assign new_new_n20417__ = ~pi076 & ~po005;
  assign new_new_n20418__ = ~new_new_n20416__ & ~new_new_n20417__;
  assign new_new_n20419__ = new_new_n20415__ & ~new_new_n20418__;
  assign new_new_n20420__ = ~new_new_n20415__ & new_new_n20418__;
  assign new_new_n20421__ = ~new_new_n20419__ & ~new_new_n20420__;
  assign new_new_n20422__ = pi077 & ~new_new_n20421__;
  assign new_new_n20423__ = ~pi077 & new_new_n20421__;
  assign new_new_n20424__ = ~new_new_n19781__ & ~new_new_n19782__;
  assign new_new_n20425__ = ~new_new_n19910__ & po005;
  assign new_new_n20426__ = ~pi075 & ~po005;
  assign new_new_n20427__ = ~new_new_n20425__ & ~new_new_n20426__;
  assign new_new_n20428__ = new_new_n20424__ & ~new_new_n20427__;
  assign new_new_n20429__ = ~new_new_n20424__ & new_new_n20427__;
  assign new_new_n20430__ = ~new_new_n20428__ & ~new_new_n20429__;
  assign new_new_n20431__ = pi076 & ~new_new_n20430__;
  assign new_new_n20432__ = ~pi076 & new_new_n20430__;
  assign new_new_n20433__ = ~new_new_n19908__ & po005;
  assign new_new_n20434__ = pi074 & ~po005;
  assign new_new_n20435__ = ~new_new_n20433__ & ~new_new_n20434__;
  assign new_new_n20436__ = ~new_new_n19790__ & ~new_new_n19791__;
  assign new_new_n20437__ = ~new_new_n20435__ & new_new_n20436__;
  assign new_new_n20438__ = new_new_n20435__ & ~new_new_n20436__;
  assign new_new_n20439__ = ~new_new_n20437__ & ~new_new_n20438__;
  assign new_new_n20440__ = pi075 & new_new_n20439__;
  assign new_new_n20441__ = ~pi075 & ~new_new_n20439__;
  assign new_new_n20442__ = ~new_new_n19799__ & ~new_new_n19800__;
  assign new_new_n20443__ = ~new_new_n19906__ & po005;
  assign new_new_n20444__ = ~pi073 & ~po005;
  assign new_new_n20445__ = ~new_new_n20443__ & ~new_new_n20444__;
  assign new_new_n20446__ = new_new_n20442__ & ~new_new_n20445__;
  assign new_new_n20447__ = ~new_new_n20442__ & new_new_n20445__;
  assign new_new_n20448__ = ~new_new_n20446__ & ~new_new_n20447__;
  assign new_new_n20449__ = pi074 & ~new_new_n20448__;
  assign new_new_n20450__ = ~pi074 & new_new_n20448__;
  assign new_new_n20451__ = ~new_new_n19896__ & ~new_new_n19897__;
  assign new_new_n20452__ = po005 & new_new_n20451__;
  assign new_new_n20453__ = new_new_n19904__ & new_new_n20452__;
  assign new_new_n20454__ = ~new_new_n19904__ & ~new_new_n20452__;
  assign new_new_n20455__ = ~new_new_n20453__ & ~new_new_n20454__;
  assign new_new_n20456__ = pi073 & ~new_new_n20455__;
  assign new_new_n20457__ = ~pi073 & new_new_n20455__;
  assign new_new_n20458__ = ~new_new_n19808__ & ~new_new_n19809__;
  assign new_new_n20459__ = pi071 & ~po005;
  assign new_new_n20460__ = ~new_new_n19893__ & po005;
  assign new_new_n20461__ = ~new_new_n20459__ & ~new_new_n20460__;
  assign new_new_n20462__ = new_new_n20458__ & new_new_n20461__;
  assign new_new_n20463__ = ~new_new_n20458__ & ~new_new_n20461__;
  assign new_new_n20464__ = ~new_new_n20462__ & ~new_new_n20463__;
  assign new_new_n20465__ = pi072 & ~new_new_n20464__;
  assign new_new_n20466__ = ~pi072 & new_new_n20464__;
  assign new_new_n20467__ = new_new_n19891__ & po005;
  assign new_new_n20468__ = ~pi070 & ~po005;
  assign new_new_n20469__ = ~new_new_n20467__ & ~new_new_n20468__;
  assign new_new_n20470__ = ~new_new_n19817__ & ~new_new_n19818__;
  assign new_new_n20471__ = ~new_new_n20469__ & ~new_new_n20470__;
  assign new_new_n20472__ = new_new_n20469__ & new_new_n20470__;
  assign new_new_n20473__ = ~new_new_n20471__ & ~new_new_n20472__;
  assign new_new_n20474__ = ~pi071 & ~new_new_n20473__;
  assign new_new_n20475__ = pi071 & new_new_n20473__;
  assign new_new_n20476__ = new_new_n19889__ & po005;
  assign new_new_n20477__ = ~pi069 & ~po005;
  assign new_new_n20478__ = ~new_new_n20476__ & ~new_new_n20477__;
  assign new_new_n20479__ = ~new_new_n19826__ & ~new_new_n19827__;
  assign new_new_n20480__ = ~new_new_n20478__ & ~new_new_n20479__;
  assign new_new_n20481__ = new_new_n20478__ & new_new_n20479__;
  assign new_new_n20482__ = ~new_new_n20480__ & ~new_new_n20481__;
  assign new_new_n20483__ = ~pi070 & ~new_new_n20482__;
  assign new_new_n20484__ = pi070 & new_new_n20482__;
  assign new_new_n20485__ = new_new_n19887__ & po005;
  assign new_new_n20486__ = ~pi068 & ~po005;
  assign new_new_n20487__ = ~new_new_n20485__ & ~new_new_n20486__;
  assign new_new_n20488__ = ~new_new_n19835__ & ~new_new_n19836__;
  assign new_new_n20489__ = ~new_new_n20487__ & ~new_new_n20488__;
  assign new_new_n20490__ = new_new_n20487__ & new_new_n20488__;
  assign new_new_n20491__ = ~new_new_n20489__ & ~new_new_n20490__;
  assign new_new_n20492__ = ~pi069 & ~new_new_n20491__;
  assign new_new_n20493__ = pi069 & new_new_n20491__;
  assign new_new_n20494__ = ~pi067 & ~new_new_n19885__;
  assign new_new_n20495__ = pi067 & new_new_n19885__;
  assign new_new_n20496__ = ~new_new_n20494__ & ~new_new_n20495__;
  assign new_new_n20497__ = po005 & ~new_new_n20496__;
  assign new_new_n20498__ = new_new_n19841__ & new_new_n20497__;
  assign new_new_n20499__ = ~new_new_n19841__ & ~new_new_n20497__;
  assign new_new_n20500__ = ~new_new_n20498__ & ~new_new_n20499__;
  assign new_new_n20501__ = pi068 & ~new_new_n20500__;
  assign new_new_n20502__ = ~pi068 & new_new_n20500__;
  assign new_new_n20503__ = ~new_new_n19856__ & ~new_new_n19883__;
  assign new_new_n20504__ = po005 & new_new_n20503__;
  assign new_new_n20505__ = new_new_n19882__ & ~new_new_n20504__;
  assign new_new_n20506__ = ~new_new_n19882__ & new_new_n20504__;
  assign new_new_n20507__ = ~new_new_n20505__ & ~new_new_n20506__;
  assign new_new_n20508__ = pi067 & new_new_n20507__;
  assign new_new_n20509__ = ~pi067 & ~new_new_n20507__;
  assign new_new_n20510__ = ~pi005 & ~po005;
  assign new_new_n20511__ = ~pi065 & ~new_new_n20510__;
  assign new_new_n20512__ = ~pi004 & ~new_new_n20511__;
  assign new_new_n20513__ = pi004 & ~pi065;
  assign new_new_n20514__ = pi005 & ~new_new_n20513__;
  assign new_new_n20515__ = po005 & new_new_n20514__;
  assign new_new_n20516__ = ~new_new_n20512__ & ~new_new_n20515__;
  assign new_new_n20517__ = pi064 & ~new_new_n20516__;
  assign new_new_n20518__ = pi064 & po005;
  assign new_new_n20519__ = pi065 & ~new_new_n20518__;
  assign new_new_n20520__ = ~pi005 & new_new_n20519__;
  assign new_new_n20521__ = ~new_new_n20517__ & ~new_new_n20520__;
  assign new_new_n20522__ = ~new_new_n332__ & po005;
  assign new_new_n20523__ = ~new_new_n19852__ & ~new_new_n20522__;
  assign new_new_n20524__ = po006 & ~po005;
  assign new_new_n20525__ = ~pi065 & ~po006;
  assign new_new_n20526__ = ~new_new_n19861__ & ~new_new_n20525__;
  assign new_new_n20527__ = ~pi005 & ~new_new_n403__;
  assign new_new_n20528__ = new_new_n20526__ & new_new_n20527__;
  assign new_new_n20529__ = ~new_new_n20524__ & new_new_n20528__;
  assign new_new_n20530__ = pi005 & ~new_new_n20526__;
  assign new_new_n20531__ = ~new_new_n20519__ & new_new_n20530__;
  assign new_new_n20532__ = ~new_new_n20523__ & ~new_new_n20529__;
  assign new_new_n20533__ = ~new_new_n20531__ & new_new_n20532__;
  assign new_new_n20534__ = ~pi006 & ~new_new_n20533__;
  assign new_new_n20535__ = ~pi065 & ~po005;
  assign new_new_n20536__ = ~pi005 & ~new_new_n20526__;
  assign new_new_n20537__ = ~new_new_n20535__ & new_new_n20536__;
  assign new_new_n20538__ = ~new_new_n20524__ & ~new_new_n20537__;
  assign new_new_n20539__ = pi064 & ~new_new_n20538__;
  assign new_new_n20540__ = pi065 & po005;
  assign new_new_n20541__ = ~new_new_n19852__ & ~new_new_n20540__;
  assign new_new_n20542__ = pi005 & ~new_new_n19861__;
  assign new_new_n20543__ = pi064 & ~new_new_n20542__;
  assign new_new_n20544__ = ~new_new_n20541__ & ~new_new_n20543__;
  assign new_new_n20545__ = ~new_new_n20539__ & ~new_new_n20544__;
  assign new_new_n20546__ = pi006 & ~new_new_n20545__;
  assign new_new_n20547__ = ~new_new_n20534__ & ~new_new_n20546__;
  assign new_new_n20548__ = ~pi066 & new_new_n20547__;
  assign new_new_n20549__ = ~new_new_n20521__ & ~new_new_n20548__;
  assign new_new_n20550__ = pi066 & ~new_new_n20547__;
  assign new_new_n20551__ = ~new_new_n20549__ & ~new_new_n20550__;
  assign new_new_n20552__ = ~new_new_n20509__ & ~new_new_n20551__;
  assign new_new_n20553__ = ~new_new_n20508__ & ~new_new_n20552__;
  assign new_new_n20554__ = ~new_new_n20502__ & ~new_new_n20553__;
  assign new_new_n20555__ = ~new_new_n20501__ & ~new_new_n20554__;
  assign new_new_n20556__ = ~new_new_n20493__ & new_new_n20555__;
  assign new_new_n20557__ = ~new_new_n20492__ & ~new_new_n20556__;
  assign new_new_n20558__ = ~new_new_n20484__ & ~new_new_n20557__;
  assign new_new_n20559__ = ~new_new_n20483__ & ~new_new_n20558__;
  assign new_new_n20560__ = ~new_new_n20475__ & ~new_new_n20559__;
  assign new_new_n20561__ = ~new_new_n20474__ & ~new_new_n20560__;
  assign new_new_n20562__ = ~new_new_n20466__ & new_new_n20561__;
  assign new_new_n20563__ = ~new_new_n20465__ & ~new_new_n20562__;
  assign new_new_n20564__ = ~new_new_n20457__ & ~new_new_n20563__;
  assign new_new_n20565__ = ~new_new_n20456__ & ~new_new_n20564__;
  assign new_new_n20566__ = ~new_new_n20450__ & ~new_new_n20565__;
  assign new_new_n20567__ = ~new_new_n20449__ & ~new_new_n20566__;
  assign new_new_n20568__ = ~new_new_n20441__ & ~new_new_n20567__;
  assign new_new_n20569__ = ~new_new_n20440__ & ~new_new_n20568__;
  assign new_new_n20570__ = ~new_new_n20432__ & ~new_new_n20569__;
  assign new_new_n20571__ = ~new_new_n20431__ & ~new_new_n20570__;
  assign new_new_n20572__ = ~new_new_n20423__ & ~new_new_n20571__;
  assign new_new_n20573__ = ~new_new_n20422__ & ~new_new_n20572__;
  assign new_new_n20574__ = ~new_new_n20414__ & ~new_new_n20573__;
  assign new_new_n20575__ = ~new_new_n20413__ & ~new_new_n20574__;
  assign new_new_n20576__ = ~new_new_n20405__ & ~new_new_n20575__;
  assign new_new_n20577__ = ~new_new_n20404__ & ~new_new_n20576__;
  assign new_new_n20578__ = ~new_new_n20396__ & ~new_new_n20577__;
  assign new_new_n20579__ = ~new_new_n20395__ & ~new_new_n20578__;
  assign new_new_n20580__ = ~new_new_n20387__ & ~new_new_n20579__;
  assign new_new_n20581__ = ~new_new_n20386__ & ~new_new_n20580__;
  assign new_new_n20582__ = ~new_new_n20378__ & ~new_new_n20581__;
  assign new_new_n20583__ = ~new_new_n20377__ & ~new_new_n20582__;
  assign new_new_n20584__ = ~new_new_n20369__ & ~new_new_n20583__;
  assign new_new_n20585__ = ~new_new_n20368__ & ~new_new_n20584__;
  assign new_new_n20586__ = ~new_new_n20360__ & ~new_new_n20585__;
  assign new_new_n20587__ = ~new_new_n20359__ & ~new_new_n20586__;
  assign new_new_n20588__ = ~new_new_n20351__ & ~new_new_n20587__;
  assign new_new_n20589__ = ~new_new_n20350__ & ~new_new_n20588__;
  assign new_new_n20590__ = ~new_new_n20342__ & ~new_new_n20589__;
  assign new_new_n20591__ = ~new_new_n20341__ & ~new_new_n20590__;
  assign new_new_n20592__ = ~new_new_n20333__ & ~new_new_n20591__;
  assign new_new_n20593__ = ~new_new_n20332__ & ~new_new_n20592__;
  assign new_new_n20594__ = ~new_new_n20324__ & ~new_new_n20593__;
  assign new_new_n20595__ = ~new_new_n20323__ & ~new_new_n20594__;
  assign new_new_n20596__ = ~new_new_n20315__ & new_new_n20595__;
  assign new_new_n20597__ = ~new_new_n20314__ & ~new_new_n20596__;
  assign new_new_n20598__ = ~new_new_n20306__ & ~new_new_n20597__;
  assign new_new_n20599__ = ~new_new_n20305__ & ~new_new_n20598__;
  assign new_new_n20600__ = ~new_new_n20297__ & ~new_new_n20599__;
  assign new_new_n20601__ = ~new_new_n20296__ & ~new_new_n20600__;
  assign new_new_n20602__ = ~new_new_n20288__ & new_new_n20601__;
  assign new_new_n20603__ = ~new_new_n20287__ & ~new_new_n20602__;
  assign new_new_n20604__ = ~new_new_n20279__ & new_new_n20603__;
  assign new_new_n20605__ = ~new_new_n20278__ & ~new_new_n20604__;
  assign new_new_n20606__ = ~new_new_n20270__ & ~new_new_n20605__;
  assign new_new_n20607__ = ~new_new_n20269__ & ~new_new_n20606__;
  assign new_new_n20608__ = ~new_new_n20261__ & new_new_n20607__;
  assign new_new_n20609__ = ~new_new_n20260__ & ~new_new_n20608__;
  assign new_new_n20610__ = ~new_new_n20252__ & ~new_new_n20609__;
  assign new_new_n20611__ = ~new_new_n20251__ & ~new_new_n20610__;
  assign new_new_n20612__ = ~new_new_n20243__ & ~new_new_n20611__;
  assign new_new_n20613__ = ~new_new_n20242__ & ~new_new_n20612__;
  assign new_new_n20614__ = ~new_new_n20234__ & ~new_new_n20613__;
  assign new_new_n20615__ = ~new_new_n20233__ & ~new_new_n20614__;
  assign new_new_n20616__ = ~new_new_n20225__ & ~new_new_n20615__;
  assign new_new_n20617__ = ~new_new_n20224__ & ~new_new_n20616__;
  assign new_new_n20618__ = ~new_new_n20216__ & ~new_new_n20617__;
  assign new_new_n20619__ = ~new_new_n20215__ & ~new_new_n20618__;
  assign new_new_n20620__ = ~new_new_n20207__ & ~new_new_n20619__;
  assign new_new_n20621__ = ~new_new_n20206__ & ~new_new_n20620__;
  assign new_new_n20622__ = ~new_new_n20198__ & ~new_new_n20621__;
  assign new_new_n20623__ = ~new_new_n20197__ & ~new_new_n20622__;
  assign new_new_n20624__ = ~new_new_n20189__ & ~new_new_n20623__;
  assign new_new_n20625__ = ~new_new_n20188__ & ~new_new_n20624__;
  assign new_new_n20626__ = ~new_new_n20180__ & ~new_new_n20625__;
  assign new_new_n20627__ = ~new_new_n20179__ & ~new_new_n20626__;
  assign new_new_n20628__ = ~new_new_n20171__ & new_new_n20627__;
  assign new_new_n20629__ = ~new_new_n20170__ & ~new_new_n20628__;
  assign new_new_n20630__ = ~new_new_n20162__ & ~new_new_n20629__;
  assign new_new_n20631__ = ~new_new_n20161__ & ~new_new_n20630__;
  assign new_new_n20632__ = ~new_new_n20153__ & ~new_new_n20631__;
  assign new_new_n20633__ = ~new_new_n20152__ & ~new_new_n20632__;
  assign new_new_n20634__ = ~new_new_n20144__ & ~new_new_n20633__;
  assign new_new_n20635__ = ~new_new_n20143__ & ~new_new_n20634__;
  assign new_new_n20636__ = ~new_new_n20135__ & ~new_new_n20635__;
  assign new_new_n20637__ = ~new_new_n20134__ & ~new_new_n20636__;
  assign new_new_n20638__ = ~pi110 & new_new_n20125__;
  assign new_new_n20639__ = new_new_n20637__ & ~new_new_n20638__;
  assign new_new_n20640__ = ~new_new_n20126__ & ~new_new_n20639__;
  assign new_new_n20641__ = ~new_new_n20118__ & ~new_new_n20640__;
  assign new_new_n20642__ = ~new_new_n20117__ & ~new_new_n20641__;
  assign new_new_n20643__ = ~new_new_n20109__ & ~new_new_n20642__;
  assign new_new_n20644__ = ~new_new_n20108__ & ~new_new_n20643__;
  assign new_new_n20645__ = ~new_new_n20100__ & ~new_new_n20644__;
  assign new_new_n20646__ = ~new_new_n20099__ & ~new_new_n20645__;
  assign new_new_n20647__ = ~new_new_n20091__ & ~new_new_n20646__;
  assign new_new_n20648__ = ~new_new_n20090__ & ~new_new_n20647__;
  assign new_new_n20649__ = ~new_new_n20082__ & ~new_new_n20648__;
  assign new_new_n20650__ = ~new_new_n20081__ & ~new_new_n20649__;
  assign new_new_n20651__ = ~new_new_n20073__ & ~new_new_n20650__;
  assign new_new_n20652__ = ~new_new_n20072__ & ~new_new_n20651__;
  assign new_new_n20653__ = ~new_new_n20064__ & ~new_new_n20652__;
  assign new_new_n20654__ = ~new_new_n20063__ & ~new_new_n20653__;
  assign new_new_n20655__ = ~new_new_n20055__ & new_new_n20654__;
  assign new_new_n20656__ = ~new_new_n20054__ & ~new_new_n20655__;
  assign new_new_n20657__ = ~new_new_n20046__ & ~new_new_n20656__;
  assign new_new_n20658__ = ~new_new_n20045__ & ~new_new_n20657__;
  assign new_new_n20659__ = ~new_new_n20037__ & ~new_new_n20658__;
  assign new_new_n20660__ = ~new_new_n20036__ & ~new_new_n20659__;
  assign new_new_n20661__ = ~new_new_n20028__ & ~new_new_n20660__;
  assign new_new_n20662__ = ~new_new_n20027__ & ~new_new_n20661__;
  assign new_new_n20663__ = ~pi123 & new_new_n20018__;
  assign new_new_n20664__ = pi123 & ~new_new_n18720__;
  assign new_new_n20665__ = ~pi121 & ~new_new_n20003__;
  assign new_new_n20666__ = pi121 & new_new_n20003__;
  assign new_new_n20667__ = ~new_new_n20665__ & ~new_new_n20666__;
  assign new_new_n20668__ = po005 & new_new_n20667__;
  assign new_new_n20669__ = ~new_new_n19372__ & new_new_n20668__;
  assign new_new_n20670__ = new_new_n19372__ & ~new_new_n20668__;
  assign new_new_n20671__ = ~new_new_n20669__ & ~new_new_n20670__;
  assign new_new_n20672__ = pi122 & ~new_new_n20671__;
  assign new_new_n20673__ = ~pi122 & new_new_n20671__;
  assign new_new_n20674__ = new_new_n20662__ & ~new_new_n20673__;
  assign new_new_n20675__ = ~new_new_n20672__ & ~new_new_n20674__;
  assign new_new_n20676__ = ~new_new_n20664__ & new_new_n20675__;
  assign new_new_n20677__ = ~new_new_n20663__ & ~new_new_n20676__;
  assign po004 = new_new_n262__ & ~new_new_n20677__;
  assign new_new_n20679__ = new_new_n20662__ & po004;
  assign new_new_n20680__ = pi122 & ~po004;
  assign new_new_n20681__ = ~new_new_n20679__ & ~new_new_n20680__;
  assign new_new_n20682__ = ~new_new_n20672__ & ~new_new_n20673__;
  assign new_new_n20683__ = ~new_new_n20681__ & ~new_new_n20682__;
  assign new_new_n20684__ = new_new_n20681__ & new_new_n20682__;
  assign new_new_n20685__ = ~new_new_n20683__ & ~new_new_n20684__;
  assign new_new_n20686__ = pi123 & ~new_new_n20685__;
  assign new_new_n20687__ = ~pi123 & new_new_n20685__;
  assign new_new_n20688__ = ~new_new_n20027__ & ~new_new_n20028__;
  assign new_new_n20689__ = ~new_new_n20660__ & po004;
  assign new_new_n20690__ = ~pi121 & ~po004;
  assign new_new_n20691__ = ~new_new_n20689__ & ~new_new_n20690__;
  assign new_new_n20692__ = new_new_n20688__ & ~new_new_n20691__;
  assign new_new_n20693__ = ~new_new_n20688__ & new_new_n20691__;
  assign new_new_n20694__ = ~new_new_n20692__ & ~new_new_n20693__;
  assign new_new_n20695__ = pi122 & ~new_new_n20694__;
  assign new_new_n20696__ = ~pi122 & new_new_n20694__;
  assign new_new_n20697__ = ~new_new_n20036__ & ~new_new_n20037__;
  assign new_new_n20698__ = ~new_new_n20658__ & po004;
  assign new_new_n20699__ = ~pi120 & ~po004;
  assign new_new_n20700__ = ~new_new_n20698__ & ~new_new_n20699__;
  assign new_new_n20701__ = new_new_n20697__ & ~new_new_n20700__;
  assign new_new_n20702__ = ~new_new_n20697__ & new_new_n20700__;
  assign new_new_n20703__ = ~new_new_n20701__ & ~new_new_n20702__;
  assign new_new_n20704__ = pi121 & ~new_new_n20703__;
  assign new_new_n20705__ = ~pi121 & new_new_n20703__;
  assign new_new_n20706__ = ~new_new_n20045__ & ~new_new_n20046__;
  assign new_new_n20707__ = ~new_new_n20656__ & po004;
  assign new_new_n20708__ = ~pi119 & ~po004;
  assign new_new_n20709__ = ~new_new_n20707__ & ~new_new_n20708__;
  assign new_new_n20710__ = new_new_n20706__ & ~new_new_n20709__;
  assign new_new_n20711__ = ~new_new_n20706__ & new_new_n20709__;
  assign new_new_n20712__ = ~new_new_n20710__ & ~new_new_n20711__;
  assign new_new_n20713__ = pi120 & ~new_new_n20712__;
  assign new_new_n20714__ = ~pi120 & new_new_n20712__;
  assign new_new_n20715__ = ~new_new_n20654__ & po004;
  assign new_new_n20716__ = pi118 & ~po004;
  assign new_new_n20717__ = ~new_new_n20715__ & ~new_new_n20716__;
  assign new_new_n20718__ = ~new_new_n20054__ & ~new_new_n20055__;
  assign new_new_n20719__ = ~new_new_n20717__ & new_new_n20718__;
  assign new_new_n20720__ = new_new_n20717__ & ~new_new_n20718__;
  assign new_new_n20721__ = ~new_new_n20719__ & ~new_new_n20720__;
  assign new_new_n20722__ = ~pi119 & ~new_new_n20721__;
  assign new_new_n20723__ = pi119 & new_new_n20721__;
  assign new_new_n20724__ = pi117 & ~new_new_n20652__;
  assign new_new_n20725__ = ~pi117 & new_new_n20652__;
  assign new_new_n20726__ = ~new_new_n20724__ & ~new_new_n20725__;
  assign new_new_n20727__ = po004 & new_new_n20726__;
  assign new_new_n20728__ = new_new_n20062__ & new_new_n20727__;
  assign new_new_n20729__ = ~new_new_n20062__ & ~new_new_n20727__;
  assign new_new_n20730__ = ~new_new_n20728__ & ~new_new_n20729__;
  assign new_new_n20731__ = ~pi118 & new_new_n20730__;
  assign new_new_n20732__ = pi118 & ~new_new_n20730__;
  assign new_new_n20733__ = ~new_new_n20650__ & po004;
  assign new_new_n20734__ = pi116 & ~po004;
  assign new_new_n20735__ = ~new_new_n20733__ & ~new_new_n20734__;
  assign new_new_n20736__ = ~new_new_n20072__ & ~new_new_n20073__;
  assign new_new_n20737__ = ~new_new_n20735__ & new_new_n20736__;
  assign new_new_n20738__ = new_new_n20735__ & ~new_new_n20736__;
  assign new_new_n20739__ = ~new_new_n20737__ & ~new_new_n20738__;
  assign new_new_n20740__ = ~pi117 & ~new_new_n20739__;
  assign new_new_n20741__ = pi117 & new_new_n20739__;
  assign new_new_n20742__ = ~new_new_n20081__ & ~new_new_n20082__;
  assign new_new_n20743__ = ~new_new_n20648__ & po004;
  assign new_new_n20744__ = pi115 & ~po004;
  assign new_new_n20745__ = ~new_new_n20743__ & ~new_new_n20744__;
  assign new_new_n20746__ = new_new_n20742__ & new_new_n20745__;
  assign new_new_n20747__ = ~new_new_n20742__ & ~new_new_n20745__;
  assign new_new_n20748__ = ~new_new_n20746__ & ~new_new_n20747__;
  assign new_new_n20749__ = ~pi116 & new_new_n20748__;
  assign new_new_n20750__ = pi116 & ~new_new_n20748__;
  assign new_new_n20751__ = new_new_n20646__ & po004;
  assign new_new_n20752__ = ~pi114 & ~po004;
  assign new_new_n20753__ = ~new_new_n20751__ & ~new_new_n20752__;
  assign new_new_n20754__ = ~new_new_n20090__ & ~new_new_n20091__;
  assign new_new_n20755__ = ~new_new_n20753__ & ~new_new_n20754__;
  assign new_new_n20756__ = new_new_n20753__ & new_new_n20754__;
  assign new_new_n20757__ = ~new_new_n20755__ & ~new_new_n20756__;
  assign new_new_n20758__ = ~pi115 & ~new_new_n20757__;
  assign new_new_n20759__ = pi115 & new_new_n20757__;
  assign new_new_n20760__ = new_new_n20644__ & po004;
  assign new_new_n20761__ = ~pi113 & ~po004;
  assign new_new_n20762__ = ~new_new_n20760__ & ~new_new_n20761__;
  assign new_new_n20763__ = ~new_new_n20099__ & ~new_new_n20100__;
  assign new_new_n20764__ = ~new_new_n20762__ & ~new_new_n20763__;
  assign new_new_n20765__ = new_new_n20762__ & new_new_n20763__;
  assign new_new_n20766__ = ~new_new_n20764__ & ~new_new_n20765__;
  assign new_new_n20767__ = ~pi114 & ~new_new_n20766__;
  assign new_new_n20768__ = pi114 & new_new_n20766__;
  assign new_new_n20769__ = ~new_new_n20642__ & po004;
  assign new_new_n20770__ = pi112 & ~po004;
  assign new_new_n20771__ = ~new_new_n20769__ & ~new_new_n20770__;
  assign new_new_n20772__ = ~new_new_n20108__ & ~new_new_n20109__;
  assign new_new_n20773__ = ~new_new_n20771__ & new_new_n20772__;
  assign new_new_n20774__ = new_new_n20771__ & ~new_new_n20772__;
  assign new_new_n20775__ = ~new_new_n20773__ & ~new_new_n20774__;
  assign new_new_n20776__ = ~pi113 & ~new_new_n20775__;
  assign new_new_n20777__ = pi113 & new_new_n20775__;
  assign new_new_n20778__ = pi111 & ~new_new_n20640__;
  assign new_new_n20779__ = ~pi111 & new_new_n20640__;
  assign new_new_n20780__ = ~new_new_n20778__ & ~new_new_n20779__;
  assign new_new_n20781__ = po004 & new_new_n20780__;
  assign new_new_n20782__ = new_new_n20116__ & new_new_n20781__;
  assign new_new_n20783__ = ~new_new_n20116__ & ~new_new_n20781__;
  assign new_new_n20784__ = ~new_new_n20782__ & ~new_new_n20783__;
  assign new_new_n20785__ = pi112 & ~new_new_n20784__;
  assign new_new_n20786__ = ~pi112 & new_new_n20784__;
  assign new_new_n20787__ = ~new_new_n20126__ & ~new_new_n20638__;
  assign new_new_n20788__ = ~new_new_n20637__ & po004;
  assign new_new_n20789__ = ~pi110 & ~po004;
  assign new_new_n20790__ = ~new_new_n20788__ & ~new_new_n20789__;
  assign new_new_n20791__ = new_new_n20787__ & ~new_new_n20790__;
  assign new_new_n20792__ = ~new_new_n20787__ & new_new_n20790__;
  assign new_new_n20793__ = ~new_new_n20791__ & ~new_new_n20792__;
  assign new_new_n20794__ = pi111 & ~new_new_n20793__;
  assign new_new_n20795__ = ~pi111 & new_new_n20793__;
  assign new_new_n20796__ = ~new_new_n20134__ & ~new_new_n20135__;
  assign new_new_n20797__ = ~new_new_n20635__ & po004;
  assign new_new_n20798__ = ~pi109 & ~po004;
  assign new_new_n20799__ = ~new_new_n20797__ & ~new_new_n20798__;
  assign new_new_n20800__ = new_new_n20796__ & ~new_new_n20799__;
  assign new_new_n20801__ = ~new_new_n20796__ & new_new_n20799__;
  assign new_new_n20802__ = ~new_new_n20800__ & ~new_new_n20801__;
  assign new_new_n20803__ = pi110 & ~new_new_n20802__;
  assign new_new_n20804__ = ~pi110 & new_new_n20802__;
  assign new_new_n20805__ = ~new_new_n20143__ & ~new_new_n20144__;
  assign new_new_n20806__ = ~new_new_n20633__ & po004;
  assign new_new_n20807__ = ~pi108 & ~po004;
  assign new_new_n20808__ = ~new_new_n20806__ & ~new_new_n20807__;
  assign new_new_n20809__ = new_new_n20805__ & ~new_new_n20808__;
  assign new_new_n20810__ = ~new_new_n20805__ & new_new_n20808__;
  assign new_new_n20811__ = ~new_new_n20809__ & ~new_new_n20810__;
  assign new_new_n20812__ = pi109 & ~new_new_n20811__;
  assign new_new_n20813__ = ~pi109 & new_new_n20811__;
  assign new_new_n20814__ = ~new_new_n20152__ & ~new_new_n20153__;
  assign new_new_n20815__ = ~new_new_n20631__ & po004;
  assign new_new_n20816__ = ~pi107 & ~po004;
  assign new_new_n20817__ = ~new_new_n20815__ & ~new_new_n20816__;
  assign new_new_n20818__ = new_new_n20814__ & ~new_new_n20817__;
  assign new_new_n20819__ = ~new_new_n20814__ & new_new_n20817__;
  assign new_new_n20820__ = ~new_new_n20818__ & ~new_new_n20819__;
  assign new_new_n20821__ = pi108 & ~new_new_n20820__;
  assign new_new_n20822__ = ~pi108 & new_new_n20820__;
  assign new_new_n20823__ = new_new_n20629__ & po004;
  assign new_new_n20824__ = pi106 & ~po004;
  assign new_new_n20825__ = ~new_new_n20823__ & ~new_new_n20824__;
  assign new_new_n20826__ = ~new_new_n20161__ & ~new_new_n20162__;
  assign new_new_n20827__ = ~new_new_n20825__ & ~new_new_n20826__;
  assign new_new_n20828__ = new_new_n20825__ & new_new_n20826__;
  assign new_new_n20829__ = ~new_new_n20827__ & ~new_new_n20828__;
  assign new_new_n20830__ = pi107 & ~new_new_n20829__;
  assign new_new_n20831__ = ~pi107 & new_new_n20829__;
  assign new_new_n20832__ = new_new_n20627__ & po004;
  assign new_new_n20833__ = ~pi105 & ~po004;
  assign new_new_n20834__ = ~new_new_n20832__ & ~new_new_n20833__;
  assign new_new_n20835__ = ~new_new_n20170__ & ~new_new_n20171__;
  assign new_new_n20836__ = ~new_new_n20834__ & ~new_new_n20835__;
  assign new_new_n20837__ = new_new_n20834__ & new_new_n20835__;
  assign new_new_n20838__ = ~new_new_n20836__ & ~new_new_n20837__;
  assign new_new_n20839__ = pi106 & new_new_n20838__;
  assign new_new_n20840__ = ~pi106 & ~new_new_n20838__;
  assign new_new_n20841__ = new_new_n20625__ & po004;
  assign new_new_n20842__ = ~pi104 & ~po004;
  assign new_new_n20843__ = ~new_new_n20841__ & ~new_new_n20842__;
  assign new_new_n20844__ = ~new_new_n20179__ & ~new_new_n20180__;
  assign new_new_n20845__ = ~new_new_n20843__ & ~new_new_n20844__;
  assign new_new_n20846__ = new_new_n20843__ & new_new_n20844__;
  assign new_new_n20847__ = ~new_new_n20845__ & ~new_new_n20846__;
  assign new_new_n20848__ = pi105 & new_new_n20847__;
  assign new_new_n20849__ = ~pi105 & ~new_new_n20847__;
  assign new_new_n20850__ = ~new_new_n20188__ & ~new_new_n20189__;
  assign new_new_n20851__ = ~new_new_n20623__ & po004;
  assign new_new_n20852__ = pi103 & ~po004;
  assign new_new_n20853__ = ~new_new_n20851__ & ~new_new_n20852__;
  assign new_new_n20854__ = new_new_n20850__ & ~new_new_n20853__;
  assign new_new_n20855__ = ~new_new_n20850__ & new_new_n20853__;
  assign new_new_n20856__ = ~new_new_n20854__ & ~new_new_n20855__;
  assign new_new_n20857__ = pi104 & new_new_n20856__;
  assign new_new_n20858__ = ~pi104 & ~new_new_n20856__;
  assign new_new_n20859__ = ~pi102 & new_new_n20621__;
  assign new_new_n20860__ = pi102 & ~new_new_n20621__;
  assign new_new_n20861__ = ~new_new_n20859__ & ~new_new_n20860__;
  assign new_new_n20862__ = po004 & new_new_n20861__;
  assign new_new_n20863__ = new_new_n20196__ & new_new_n20862__;
  assign new_new_n20864__ = ~new_new_n20196__ & ~new_new_n20862__;
  assign new_new_n20865__ = ~new_new_n20863__ & ~new_new_n20864__;
  assign new_new_n20866__ = pi103 & ~new_new_n20865__;
  assign new_new_n20867__ = ~pi103 & new_new_n20865__;
  assign new_new_n20868__ = ~new_new_n20619__ & po004;
  assign new_new_n20869__ = pi101 & ~po004;
  assign new_new_n20870__ = ~new_new_n20868__ & ~new_new_n20869__;
  assign new_new_n20871__ = ~new_new_n20206__ & ~new_new_n20207__;
  assign new_new_n20872__ = new_new_n20870__ & new_new_n20871__;
  assign new_new_n20873__ = ~new_new_n20870__ & ~new_new_n20871__;
  assign new_new_n20874__ = ~new_new_n20872__ & ~new_new_n20873__;
  assign new_new_n20875__ = pi102 & ~new_new_n20874__;
  assign new_new_n20876__ = ~pi102 & new_new_n20874__;
  assign new_new_n20877__ = ~new_new_n20215__ & ~new_new_n20216__;
  assign new_new_n20878__ = ~new_new_n20617__ & po004;
  assign new_new_n20879__ = pi100 & ~po004;
  assign new_new_n20880__ = ~new_new_n20878__ & ~new_new_n20879__;
  assign new_new_n20881__ = new_new_n20877__ & new_new_n20880__;
  assign new_new_n20882__ = ~new_new_n20877__ & ~new_new_n20880__;
  assign new_new_n20883__ = ~new_new_n20881__ & ~new_new_n20882__;
  assign new_new_n20884__ = pi101 & ~new_new_n20883__;
  assign new_new_n20885__ = ~pi101 & new_new_n20883__;
  assign new_new_n20886__ = ~new_new_n20224__ & ~new_new_n20225__;
  assign new_new_n20887__ = ~new_new_n20615__ & po004;
  assign new_new_n20888__ = pi099 & ~po004;
  assign new_new_n20889__ = ~new_new_n20887__ & ~new_new_n20888__;
  assign new_new_n20890__ = new_new_n20886__ & ~new_new_n20889__;
  assign new_new_n20891__ = ~new_new_n20886__ & new_new_n20889__;
  assign new_new_n20892__ = ~new_new_n20890__ & ~new_new_n20891__;
  assign new_new_n20893__ = ~pi100 & ~new_new_n20892__;
  assign new_new_n20894__ = pi100 & new_new_n20892__;
  assign new_new_n20895__ = ~new_new_n20613__ & po004;
  assign new_new_n20896__ = pi098 & ~po004;
  assign new_new_n20897__ = ~new_new_n20895__ & ~new_new_n20896__;
  assign new_new_n20898__ = ~new_new_n20233__ & ~new_new_n20234__;
  assign new_new_n20899__ = ~new_new_n20897__ & new_new_n20898__;
  assign new_new_n20900__ = new_new_n20897__ & ~new_new_n20898__;
  assign new_new_n20901__ = ~new_new_n20899__ & ~new_new_n20900__;
  assign new_new_n20902__ = ~pi099 & ~new_new_n20901__;
  assign new_new_n20903__ = pi099 & new_new_n20901__;
  assign new_new_n20904__ = ~new_new_n20611__ & po004;
  assign new_new_n20905__ = pi097 & ~po004;
  assign new_new_n20906__ = ~new_new_n20904__ & ~new_new_n20905__;
  assign new_new_n20907__ = ~new_new_n20242__ & ~new_new_n20243__;
  assign new_new_n20908__ = ~new_new_n20906__ & new_new_n20907__;
  assign new_new_n20909__ = new_new_n20906__ & ~new_new_n20907__;
  assign new_new_n20910__ = ~new_new_n20908__ & ~new_new_n20909__;
  assign new_new_n20911__ = ~pi098 & ~new_new_n20910__;
  assign new_new_n20912__ = pi098 & new_new_n20910__;
  assign new_new_n20913__ = pi096 & ~new_new_n20609__;
  assign new_new_n20914__ = ~pi096 & new_new_n20609__;
  assign new_new_n20915__ = ~new_new_n20913__ & ~new_new_n20914__;
  assign new_new_n20916__ = po004 & new_new_n20915__;
  assign new_new_n20917__ = new_new_n20250__ & new_new_n20916__;
  assign new_new_n20918__ = ~new_new_n20250__ & ~new_new_n20916__;
  assign new_new_n20919__ = ~new_new_n20917__ & ~new_new_n20918__;
  assign new_new_n20920__ = pi097 & ~new_new_n20919__;
  assign new_new_n20921__ = ~pi097 & new_new_n20919__;
  assign new_new_n20922__ = ~new_new_n20260__ & ~new_new_n20261__;
  assign new_new_n20923__ = ~new_new_n20607__ & po004;
  assign new_new_n20924__ = ~pi095 & ~po004;
  assign new_new_n20925__ = ~new_new_n20923__ & ~new_new_n20924__;
  assign new_new_n20926__ = new_new_n20922__ & ~new_new_n20925__;
  assign new_new_n20927__ = ~new_new_n20922__ & new_new_n20925__;
  assign new_new_n20928__ = ~new_new_n20926__ & ~new_new_n20927__;
  assign new_new_n20929__ = ~pi096 & new_new_n20928__;
  assign new_new_n20930__ = pi096 & ~new_new_n20928__;
  assign new_new_n20931__ = ~pi094 & ~new_new_n20605__;
  assign new_new_n20932__ = pi094 & new_new_n20605__;
  assign new_new_n20933__ = ~new_new_n20931__ & ~new_new_n20932__;
  assign new_new_n20934__ = po004 & new_new_n20933__;
  assign new_new_n20935__ = new_new_n20268__ & new_new_n20934__;
  assign new_new_n20936__ = ~new_new_n20268__ & ~new_new_n20934__;
  assign new_new_n20937__ = ~new_new_n20935__ & ~new_new_n20936__;
  assign new_new_n20938__ = ~pi095 & ~new_new_n20937__;
  assign new_new_n20939__ = pi095 & new_new_n20937__;
  assign new_new_n20940__ = ~new_new_n20278__ & ~new_new_n20279__;
  assign new_new_n20941__ = ~new_new_n20603__ & po004;
  assign new_new_n20942__ = pi093 & ~po004;
  assign new_new_n20943__ = ~new_new_n20941__ & ~new_new_n20942__;
  assign new_new_n20944__ = new_new_n20940__ & ~new_new_n20943__;
  assign new_new_n20945__ = ~new_new_n20940__ & new_new_n20943__;
  assign new_new_n20946__ = ~new_new_n20944__ & ~new_new_n20945__;
  assign new_new_n20947__ = ~pi094 & ~new_new_n20946__;
  assign new_new_n20948__ = pi094 & new_new_n20946__;
  assign new_new_n20949__ = ~new_new_n20287__ & ~new_new_n20288__;
  assign new_new_n20950__ = ~new_new_n20601__ & po004;
  assign new_new_n20951__ = ~pi092 & ~po004;
  assign new_new_n20952__ = ~new_new_n20950__ & ~new_new_n20951__;
  assign new_new_n20953__ = new_new_n20949__ & ~new_new_n20952__;
  assign new_new_n20954__ = ~new_new_n20949__ & new_new_n20952__;
  assign new_new_n20955__ = ~new_new_n20953__ & ~new_new_n20954__;
  assign new_new_n20956__ = pi093 & ~new_new_n20955__;
  assign new_new_n20957__ = ~pi093 & new_new_n20955__;
  assign new_new_n20958__ = ~new_new_n20296__ & ~new_new_n20297__;
  assign new_new_n20959__ = ~new_new_n20599__ & po004;
  assign new_new_n20960__ = ~pi091 & ~po004;
  assign new_new_n20961__ = ~new_new_n20959__ & ~new_new_n20960__;
  assign new_new_n20962__ = ~new_new_n20958__ & ~new_new_n20961__;
  assign new_new_n20963__ = new_new_n20958__ & new_new_n20961__;
  assign new_new_n20964__ = ~new_new_n20962__ & ~new_new_n20963__;
  assign new_new_n20965__ = pi092 & new_new_n20964__;
  assign new_new_n20966__ = ~pi092 & ~new_new_n20964__;
  assign new_new_n20967__ = new_new_n20597__ & po004;
  assign new_new_n20968__ = pi090 & ~po004;
  assign new_new_n20969__ = ~new_new_n20967__ & ~new_new_n20968__;
  assign new_new_n20970__ = ~new_new_n20305__ & ~new_new_n20306__;
  assign new_new_n20971__ = ~new_new_n20969__ & ~new_new_n20970__;
  assign new_new_n20972__ = new_new_n20969__ & new_new_n20970__;
  assign new_new_n20973__ = ~new_new_n20971__ & ~new_new_n20972__;
  assign new_new_n20974__ = pi091 & ~new_new_n20973__;
  assign new_new_n20975__ = ~pi091 & new_new_n20973__;
  assign new_new_n20976__ = new_new_n20595__ & po004;
  assign new_new_n20977__ = ~pi089 & ~po004;
  assign new_new_n20978__ = ~new_new_n20976__ & ~new_new_n20977__;
  assign new_new_n20979__ = ~new_new_n20314__ & ~new_new_n20315__;
  assign new_new_n20980__ = ~new_new_n20978__ & ~new_new_n20979__;
  assign new_new_n20981__ = new_new_n20978__ & new_new_n20979__;
  assign new_new_n20982__ = ~new_new_n20980__ & ~new_new_n20981__;
  assign new_new_n20983__ = pi090 & new_new_n20982__;
  assign new_new_n20984__ = ~pi090 & ~new_new_n20982__;
  assign new_new_n20985__ = pi088 & ~new_new_n20593__;
  assign new_new_n20986__ = ~pi088 & new_new_n20593__;
  assign new_new_n20987__ = ~new_new_n20985__ & ~new_new_n20986__;
  assign new_new_n20988__ = po004 & new_new_n20987__;
  assign new_new_n20989__ = ~new_new_n20322__ & ~new_new_n20988__;
  assign new_new_n20990__ = new_new_n20322__ & new_new_n20988__;
  assign new_new_n20991__ = ~new_new_n20989__ & ~new_new_n20990__;
  assign new_new_n20992__ = pi089 & ~new_new_n20991__;
  assign new_new_n20993__ = ~pi089 & new_new_n20991__;
  assign new_new_n20994__ = pi087 & ~new_new_n20591__;
  assign new_new_n20995__ = ~pi087 & new_new_n20591__;
  assign new_new_n20996__ = ~new_new_n20994__ & ~new_new_n20995__;
  assign new_new_n20997__ = po004 & new_new_n20996__;
  assign new_new_n20998__ = new_new_n20331__ & new_new_n20997__;
  assign new_new_n20999__ = ~new_new_n20331__ & ~new_new_n20997__;
  assign new_new_n21000__ = ~new_new_n20998__ & ~new_new_n20999__;
  assign new_new_n21001__ = pi088 & ~new_new_n21000__;
  assign new_new_n21002__ = ~pi088 & new_new_n21000__;
  assign new_new_n21003__ = ~new_new_n20589__ & po004;
  assign new_new_n21004__ = pi086 & ~po004;
  assign new_new_n21005__ = ~new_new_n21003__ & ~new_new_n21004__;
  assign new_new_n21006__ = ~new_new_n20341__ & ~new_new_n20342__;
  assign new_new_n21007__ = ~new_new_n21005__ & new_new_n21006__;
  assign new_new_n21008__ = new_new_n21005__ & ~new_new_n21006__;
  assign new_new_n21009__ = ~new_new_n21007__ & ~new_new_n21008__;
  assign new_new_n21010__ = ~pi087 & ~new_new_n21009__;
  assign new_new_n21011__ = pi087 & new_new_n21009__;
  assign new_new_n21012__ = ~new_new_n20587__ & po004;
  assign new_new_n21013__ = pi085 & ~po004;
  assign new_new_n21014__ = ~new_new_n21012__ & ~new_new_n21013__;
  assign new_new_n21015__ = ~new_new_n20350__ & ~new_new_n20351__;
  assign new_new_n21016__ = ~new_new_n21014__ & new_new_n21015__;
  assign new_new_n21017__ = new_new_n21014__ & ~new_new_n21015__;
  assign new_new_n21018__ = ~new_new_n21016__ & ~new_new_n21017__;
  assign new_new_n21019__ = ~pi086 & ~new_new_n21018__;
  assign new_new_n21020__ = pi086 & new_new_n21018__;
  assign new_new_n21021__ = pi084 & ~new_new_n20585__;
  assign new_new_n21022__ = ~pi084 & new_new_n20585__;
  assign new_new_n21023__ = ~new_new_n21021__ & ~new_new_n21022__;
  assign new_new_n21024__ = po004 & new_new_n21023__;
  assign new_new_n21025__ = ~new_new_n20358__ & ~new_new_n21024__;
  assign new_new_n21026__ = new_new_n20358__ & new_new_n21024__;
  assign new_new_n21027__ = ~new_new_n21025__ & ~new_new_n21026__;
  assign new_new_n21028__ = pi085 & ~new_new_n21027__;
  assign new_new_n21029__ = ~pi085 & new_new_n21027__;
  assign new_new_n21030__ = pi083 & ~new_new_n20583__;
  assign new_new_n21031__ = ~pi083 & new_new_n20583__;
  assign new_new_n21032__ = ~new_new_n21030__ & ~new_new_n21031__;
  assign new_new_n21033__ = po004 & new_new_n21032__;
  assign new_new_n21034__ = new_new_n20367__ & new_new_n21033__;
  assign new_new_n21035__ = ~new_new_n20367__ & ~new_new_n21033__;
  assign new_new_n21036__ = ~new_new_n21034__ & ~new_new_n21035__;
  assign new_new_n21037__ = ~pi084 & new_new_n21036__;
  assign new_new_n21038__ = pi084 & ~new_new_n21036__;
  assign new_new_n21039__ = ~new_new_n20377__ & ~new_new_n20378__;
  assign new_new_n21040__ = new_new_n20581__ & po004;
  assign new_new_n21041__ = ~pi082 & ~po004;
  assign new_new_n21042__ = ~new_new_n21040__ & ~new_new_n21041__;
  assign new_new_n21043__ = ~new_new_n21039__ & ~new_new_n21042__;
  assign new_new_n21044__ = new_new_n21039__ & new_new_n21042__;
  assign new_new_n21045__ = ~new_new_n21043__ & ~new_new_n21044__;
  assign new_new_n21046__ = ~pi083 & ~new_new_n21045__;
  assign new_new_n21047__ = pi083 & new_new_n21045__;
  assign new_new_n21048__ = ~new_new_n20386__ & ~new_new_n20387__;
  assign new_new_n21049__ = ~new_new_n20579__ & po004;
  assign new_new_n21050__ = pi081 & ~po004;
  assign new_new_n21051__ = ~new_new_n21049__ & ~new_new_n21050__;
  assign new_new_n21052__ = new_new_n21048__ & new_new_n21051__;
  assign new_new_n21053__ = ~new_new_n21048__ & ~new_new_n21051__;
  assign new_new_n21054__ = ~new_new_n21052__ & ~new_new_n21053__;
  assign new_new_n21055__ = ~pi082 & new_new_n21054__;
  assign new_new_n21056__ = pi082 & ~new_new_n21054__;
  assign new_new_n21057__ = new_new_n20577__ & po004;
  assign new_new_n21058__ = ~pi080 & ~po004;
  assign new_new_n21059__ = ~new_new_n21057__ & ~new_new_n21058__;
  assign new_new_n21060__ = ~new_new_n20395__ & ~new_new_n20396__;
  assign new_new_n21061__ = ~new_new_n21059__ & ~new_new_n21060__;
  assign new_new_n21062__ = new_new_n21059__ & new_new_n21060__;
  assign new_new_n21063__ = ~new_new_n21061__ & ~new_new_n21062__;
  assign new_new_n21064__ = ~pi081 & ~new_new_n21063__;
  assign new_new_n21065__ = pi081 & new_new_n21063__;
  assign new_new_n21066__ = pi079 & ~new_new_n20575__;
  assign new_new_n21067__ = ~pi079 & new_new_n20575__;
  assign new_new_n21068__ = ~new_new_n21066__ & ~new_new_n21067__;
  assign new_new_n21069__ = po004 & new_new_n21068__;
  assign new_new_n21070__ = new_new_n20403__ & new_new_n21069__;
  assign new_new_n21071__ = ~new_new_n20403__ & ~new_new_n21069__;
  assign new_new_n21072__ = ~new_new_n21070__ & ~new_new_n21071__;
  assign new_new_n21073__ = ~pi080 & new_new_n21072__;
  assign new_new_n21074__ = pi080 & ~new_new_n21072__;
  assign new_new_n21075__ = new_new_n20573__ & po004;
  assign new_new_n21076__ = ~pi078 & ~po004;
  assign new_new_n21077__ = ~new_new_n21075__ & ~new_new_n21076__;
  assign new_new_n21078__ = ~new_new_n20413__ & ~new_new_n20414__;
  assign new_new_n21079__ = ~new_new_n21077__ & ~new_new_n21078__;
  assign new_new_n21080__ = new_new_n21077__ & new_new_n21078__;
  assign new_new_n21081__ = ~new_new_n21079__ & ~new_new_n21080__;
  assign new_new_n21082__ = ~pi079 & ~new_new_n21081__;
  assign new_new_n21083__ = pi079 & new_new_n21081__;
  assign new_new_n21084__ = ~new_new_n20422__ & ~new_new_n20423__;
  assign new_new_n21085__ = ~new_new_n20571__ & po004;
  assign new_new_n21086__ = pi077 & ~po004;
  assign new_new_n21087__ = ~new_new_n21085__ & ~new_new_n21086__;
  assign new_new_n21088__ = new_new_n21084__ & new_new_n21087__;
  assign new_new_n21089__ = ~new_new_n21084__ & ~new_new_n21087__;
  assign new_new_n21090__ = ~new_new_n21088__ & ~new_new_n21089__;
  assign new_new_n21091__ = pi078 & ~new_new_n21090__;
  assign new_new_n21092__ = ~pi078 & new_new_n21090__;
  assign new_new_n21093__ = pi076 & ~new_new_n20569__;
  assign new_new_n21094__ = ~pi076 & new_new_n20569__;
  assign new_new_n21095__ = ~new_new_n21093__ & ~new_new_n21094__;
  assign new_new_n21096__ = po004 & new_new_n21095__;
  assign new_new_n21097__ = new_new_n20430__ & new_new_n21096__;
  assign new_new_n21098__ = ~new_new_n20430__ & ~new_new_n21096__;
  assign new_new_n21099__ = ~new_new_n21097__ & ~new_new_n21098__;
  assign new_new_n21100__ = pi077 & ~new_new_n21099__;
  assign new_new_n21101__ = ~pi077 & new_new_n21099__;
  assign new_new_n21102__ = ~new_new_n20567__ & po004;
  assign new_new_n21103__ = pi075 & ~po004;
  assign new_new_n21104__ = ~new_new_n21102__ & ~new_new_n21103__;
  assign new_new_n21105__ = ~new_new_n20440__ & ~new_new_n20441__;
  assign new_new_n21106__ = ~new_new_n21104__ & new_new_n21105__;
  assign new_new_n21107__ = new_new_n21104__ & ~new_new_n21105__;
  assign new_new_n21108__ = ~new_new_n21106__ & ~new_new_n21107__;
  assign new_new_n21109__ = pi076 & new_new_n21108__;
  assign new_new_n21110__ = ~pi076 & ~new_new_n21108__;
  assign new_new_n21111__ = pi074 & ~new_new_n20565__;
  assign new_new_n21112__ = ~pi074 & new_new_n20565__;
  assign new_new_n21113__ = ~new_new_n21111__ & ~new_new_n21112__;
  assign new_new_n21114__ = po004 & new_new_n21113__;
  assign new_new_n21115__ = new_new_n20448__ & new_new_n21114__;
  assign new_new_n21116__ = ~new_new_n20448__ & ~new_new_n21114__;
  assign new_new_n21117__ = ~new_new_n21115__ & ~new_new_n21116__;
  assign new_new_n21118__ = pi075 & ~new_new_n21117__;
  assign new_new_n21119__ = ~pi075 & new_new_n21117__;
  assign new_new_n21120__ = ~new_new_n20456__ & ~new_new_n20457__;
  assign new_new_n21121__ = ~new_new_n20563__ & po004;
  assign new_new_n21122__ = pi073 & ~po004;
  assign new_new_n21123__ = ~new_new_n21121__ & ~new_new_n21122__;
  assign new_new_n21124__ = new_new_n21120__ & ~new_new_n21123__;
  assign new_new_n21125__ = ~new_new_n21120__ & new_new_n21123__;
  assign new_new_n21126__ = ~new_new_n21124__ & ~new_new_n21125__;
  assign new_new_n21127__ = pi074 & new_new_n21126__;
  assign new_new_n21128__ = ~pi074 & ~new_new_n21126__;
  assign new_new_n21129__ = ~new_new_n20465__ & ~new_new_n20466__;
  assign new_new_n21130__ = ~new_new_n20561__ & po004;
  assign new_new_n21131__ = ~pi072 & ~po004;
  assign new_new_n21132__ = ~new_new_n21130__ & ~new_new_n21131__;
  assign new_new_n21133__ = new_new_n21129__ & ~new_new_n21132__;
  assign new_new_n21134__ = ~new_new_n21129__ & new_new_n21132__;
  assign new_new_n21135__ = ~new_new_n21133__ & ~new_new_n21134__;
  assign new_new_n21136__ = pi073 & ~new_new_n21135__;
  assign new_new_n21137__ = ~pi073 & new_new_n21135__;
  assign new_new_n21138__ = ~new_new_n20474__ & ~new_new_n20475__;
  assign new_new_n21139__ = ~new_new_n20559__ & po004;
  assign new_new_n21140__ = ~pi071 & ~po004;
  assign new_new_n21141__ = ~new_new_n21139__ & ~new_new_n21140__;
  assign new_new_n21142__ = new_new_n21138__ & ~new_new_n21141__;
  assign new_new_n21143__ = ~new_new_n21138__ & new_new_n21141__;
  assign new_new_n21144__ = ~new_new_n21142__ & ~new_new_n21143__;
  assign new_new_n21145__ = pi072 & ~new_new_n21144__;
  assign new_new_n21146__ = ~pi072 & new_new_n21144__;
  assign new_new_n21147__ = ~pi070 & ~new_new_n20557__;
  assign new_new_n21148__ = pi070 & new_new_n20557__;
  assign new_new_n21149__ = ~new_new_n21147__ & ~new_new_n21148__;
  assign new_new_n21150__ = po004 & new_new_n21149__;
  assign new_new_n21151__ = ~new_new_n20482__ & new_new_n21150__;
  assign new_new_n21152__ = new_new_n20482__ & ~new_new_n21150__;
  assign new_new_n21153__ = ~new_new_n21151__ & ~new_new_n21152__;
  assign new_new_n21154__ = pi071 & ~new_new_n21153__;
  assign new_new_n21155__ = ~pi071 & new_new_n21153__;
  assign new_new_n21156__ = ~new_new_n20555__ & po004;
  assign new_new_n21157__ = pi069 & ~po004;
  assign new_new_n21158__ = ~new_new_n21156__ & ~new_new_n21157__;
  assign new_new_n21159__ = ~new_new_n20492__ & ~new_new_n20493__;
  assign new_new_n21160__ = ~new_new_n21158__ & new_new_n21159__;
  assign new_new_n21161__ = new_new_n21158__ & ~new_new_n21159__;
  assign new_new_n21162__ = ~new_new_n21160__ & ~new_new_n21161__;
  assign new_new_n21163__ = ~pi070 & ~new_new_n21162__;
  assign new_new_n21164__ = pi070 & new_new_n21162__;
  assign new_new_n21165__ = ~new_new_n20553__ & po004;
  assign new_new_n21166__ = pi068 & ~po004;
  assign new_new_n21167__ = ~new_new_n21165__ & ~new_new_n21166__;
  assign new_new_n21168__ = ~new_new_n20501__ & ~new_new_n20502__;
  assign new_new_n21169__ = ~new_new_n21167__ & new_new_n21168__;
  assign new_new_n21170__ = new_new_n21167__ & ~new_new_n21168__;
  assign new_new_n21171__ = ~new_new_n21169__ & ~new_new_n21170__;
  assign new_new_n21172__ = ~pi069 & ~new_new_n21171__;
  assign new_new_n21173__ = pi069 & new_new_n21171__;
  assign new_new_n21174__ = ~new_new_n20508__ & ~new_new_n20509__;
  assign new_new_n21175__ = new_new_n20551__ & po004;
  assign new_new_n21176__ = ~pi067 & ~po004;
  assign new_new_n21177__ = ~new_new_n21175__ & ~new_new_n21176__;
  assign new_new_n21178__ = ~new_new_n21174__ & ~new_new_n21177__;
  assign new_new_n21179__ = new_new_n21174__ & new_new_n21177__;
  assign new_new_n21180__ = ~new_new_n21178__ & ~new_new_n21179__;
  assign new_new_n21181__ = ~pi068 & ~new_new_n21180__;
  assign new_new_n21182__ = pi068 & new_new_n21180__;
  assign new_new_n21183__ = pi066 & ~new_new_n20521__;
  assign new_new_n21184__ = ~pi066 & new_new_n20521__;
  assign new_new_n21185__ = ~new_new_n21183__ & ~new_new_n21184__;
  assign new_new_n21186__ = po004 & new_new_n21185__;
  assign new_new_n21187__ = new_new_n20547__ & ~new_new_n21186__;
  assign new_new_n21188__ = ~new_new_n20547__ & new_new_n21186__;
  assign new_new_n21189__ = ~new_new_n21187__ & ~new_new_n21188__;
  assign new_new_n21190__ = ~pi067 & ~new_new_n21189__;
  assign new_new_n21191__ = pi067 & new_new_n21189__;
  assign new_new_n21192__ = ~pi004 & ~po004;
  assign new_new_n21193__ = ~pi065 & ~new_new_n21192__;
  assign new_new_n21194__ = ~pi003 & ~new_new_n21193__;
  assign new_new_n21195__ = pi003 & ~pi065;
  assign new_new_n21196__ = pi004 & ~new_new_n21195__;
  assign new_new_n21197__ = po004 & new_new_n21196__;
  assign new_new_n21198__ = ~new_new_n21194__ & ~new_new_n21197__;
  assign new_new_n21199__ = pi064 & ~new_new_n21198__;
  assign new_new_n21200__ = ~pi004 & pi065;
  assign new_new_n21201__ = pi064 & po004;
  assign new_new_n21202__ = new_new_n21200__ & ~new_new_n21201__;
  assign new_new_n21203__ = ~new_new_n21199__ & ~new_new_n21202__;
  assign new_new_n21204__ = ~pi066 & new_new_n21203__;
  assign new_new_n21205__ = pi066 & ~new_new_n21203__;
  assign new_new_n21206__ = ~new_new_n20677__ & ~new_new_n21200__;
  assign new_new_n21207__ = new_new_n20518__ & ~new_new_n21206__;
  assign new_new_n21208__ = ~pi004 & new_new_n20535__;
  assign new_new_n21209__ = pi064 & ~new_new_n21208__;
  assign new_new_n21210__ = ~new_new_n332__ & ~new_new_n21209__;
  assign new_new_n21211__ = po004 & new_new_n21210__;
  assign new_new_n21212__ = pi065 & po004;
  assign new_new_n21213__ = ~new_new_n20518__ & ~new_new_n21212__;
  assign new_new_n21214__ = pi004 & ~new_new_n20540__;
  assign new_new_n21215__ = ~new_new_n21213__ & new_new_n21214__;
  assign new_new_n21216__ = ~new_new_n21207__ & ~new_new_n21211__;
  assign new_new_n21217__ = ~new_new_n21215__ & new_new_n21216__;
  assign new_new_n21218__ = pi005 & ~new_new_n21217__;
  assign new_new_n21219__ = ~pi005 & new_new_n21217__;
  assign new_new_n21220__ = ~new_new_n21218__ & ~new_new_n21219__;
  assign new_new_n21221__ = ~new_new_n21205__ & new_new_n21220__;
  assign new_new_n21222__ = ~new_new_n21204__ & ~new_new_n21221__;
  assign new_new_n21223__ = ~new_new_n21191__ & ~new_new_n21222__;
  assign new_new_n21224__ = ~new_new_n21190__ & ~new_new_n21223__;
  assign new_new_n21225__ = ~new_new_n21182__ & ~new_new_n21224__;
  assign new_new_n21226__ = ~new_new_n21181__ & ~new_new_n21225__;
  assign new_new_n21227__ = ~new_new_n21173__ & ~new_new_n21226__;
  assign new_new_n21228__ = ~new_new_n21172__ & ~new_new_n21227__;
  assign new_new_n21229__ = ~new_new_n21164__ & ~new_new_n21228__;
  assign new_new_n21230__ = ~new_new_n21163__ & ~new_new_n21229__;
  assign new_new_n21231__ = ~new_new_n21155__ & new_new_n21230__;
  assign new_new_n21232__ = ~new_new_n21154__ & ~new_new_n21231__;
  assign new_new_n21233__ = ~new_new_n21146__ & ~new_new_n21232__;
  assign new_new_n21234__ = ~new_new_n21145__ & ~new_new_n21233__;
  assign new_new_n21235__ = ~new_new_n21137__ & ~new_new_n21234__;
  assign new_new_n21236__ = ~new_new_n21136__ & ~new_new_n21235__;
  assign new_new_n21237__ = ~new_new_n21128__ & ~new_new_n21236__;
  assign new_new_n21238__ = ~new_new_n21127__ & ~new_new_n21237__;
  assign new_new_n21239__ = ~new_new_n21119__ & ~new_new_n21238__;
  assign new_new_n21240__ = ~new_new_n21118__ & ~new_new_n21239__;
  assign new_new_n21241__ = ~new_new_n21110__ & ~new_new_n21240__;
  assign new_new_n21242__ = ~new_new_n21109__ & ~new_new_n21241__;
  assign new_new_n21243__ = ~new_new_n21101__ & ~new_new_n21242__;
  assign new_new_n21244__ = ~new_new_n21100__ & ~new_new_n21243__;
  assign new_new_n21245__ = ~new_new_n21092__ & ~new_new_n21244__;
  assign new_new_n21246__ = ~new_new_n21091__ & ~new_new_n21245__;
  assign new_new_n21247__ = ~new_new_n21083__ & new_new_n21246__;
  assign new_new_n21248__ = ~new_new_n21082__ & ~new_new_n21247__;
  assign new_new_n21249__ = ~new_new_n21074__ & ~new_new_n21248__;
  assign new_new_n21250__ = ~new_new_n21073__ & ~new_new_n21249__;
  assign new_new_n21251__ = ~new_new_n21065__ & ~new_new_n21250__;
  assign new_new_n21252__ = ~new_new_n21064__ & ~new_new_n21251__;
  assign new_new_n21253__ = ~new_new_n21056__ & ~new_new_n21252__;
  assign new_new_n21254__ = ~new_new_n21055__ & ~new_new_n21253__;
  assign new_new_n21255__ = ~new_new_n21047__ & ~new_new_n21254__;
  assign new_new_n21256__ = ~new_new_n21046__ & ~new_new_n21255__;
  assign new_new_n21257__ = ~new_new_n21038__ & ~new_new_n21256__;
  assign new_new_n21258__ = ~new_new_n21037__ & ~new_new_n21257__;
  assign new_new_n21259__ = ~new_new_n21029__ & new_new_n21258__;
  assign new_new_n21260__ = ~new_new_n21028__ & ~new_new_n21259__;
  assign new_new_n21261__ = ~new_new_n21020__ & new_new_n21260__;
  assign new_new_n21262__ = ~new_new_n21019__ & ~new_new_n21261__;
  assign new_new_n21263__ = ~new_new_n21011__ & ~new_new_n21262__;
  assign new_new_n21264__ = ~new_new_n21010__ & ~new_new_n21263__;
  assign new_new_n21265__ = ~new_new_n21002__ & new_new_n21264__;
  assign new_new_n21266__ = ~new_new_n21001__ & ~new_new_n21265__;
  assign new_new_n21267__ = ~new_new_n20993__ & ~new_new_n21266__;
  assign new_new_n21268__ = ~new_new_n20992__ & ~new_new_n21267__;
  assign new_new_n21269__ = ~new_new_n20984__ & ~new_new_n21268__;
  assign new_new_n21270__ = ~new_new_n20983__ & ~new_new_n21269__;
  assign new_new_n21271__ = ~new_new_n20975__ & ~new_new_n21270__;
  assign new_new_n21272__ = ~new_new_n20974__ & ~new_new_n21271__;
  assign new_new_n21273__ = ~new_new_n20966__ & ~new_new_n21272__;
  assign new_new_n21274__ = ~new_new_n20965__ & ~new_new_n21273__;
  assign new_new_n21275__ = ~new_new_n20957__ & ~new_new_n21274__;
  assign new_new_n21276__ = ~new_new_n20956__ & ~new_new_n21275__;
  assign new_new_n21277__ = ~new_new_n20948__ & new_new_n21276__;
  assign new_new_n21278__ = ~new_new_n20947__ & ~new_new_n21277__;
  assign new_new_n21279__ = ~new_new_n20939__ & ~new_new_n21278__;
  assign new_new_n21280__ = ~new_new_n20938__ & ~new_new_n21279__;
  assign new_new_n21281__ = ~new_new_n20930__ & ~new_new_n21280__;
  assign new_new_n21282__ = ~new_new_n20929__ & ~new_new_n21281__;
  assign new_new_n21283__ = ~new_new_n20921__ & new_new_n21282__;
  assign new_new_n21284__ = ~new_new_n20920__ & ~new_new_n21283__;
  assign new_new_n21285__ = ~new_new_n20912__ & new_new_n21284__;
  assign new_new_n21286__ = ~new_new_n20911__ & ~new_new_n21285__;
  assign new_new_n21287__ = ~new_new_n20903__ & ~new_new_n21286__;
  assign new_new_n21288__ = ~new_new_n20902__ & ~new_new_n21287__;
  assign new_new_n21289__ = ~new_new_n20894__ & ~new_new_n21288__;
  assign new_new_n21290__ = ~new_new_n20893__ & ~new_new_n21289__;
  assign new_new_n21291__ = ~new_new_n20885__ & new_new_n21290__;
  assign new_new_n21292__ = ~new_new_n20884__ & ~new_new_n21291__;
  assign new_new_n21293__ = ~new_new_n20876__ & ~new_new_n21292__;
  assign new_new_n21294__ = ~new_new_n20875__ & ~new_new_n21293__;
  assign new_new_n21295__ = ~new_new_n20867__ & ~new_new_n21294__;
  assign new_new_n21296__ = ~new_new_n20866__ & ~new_new_n21295__;
  assign new_new_n21297__ = ~new_new_n20858__ & ~new_new_n21296__;
  assign new_new_n21298__ = ~new_new_n20857__ & ~new_new_n21297__;
  assign new_new_n21299__ = ~new_new_n20849__ & ~new_new_n21298__;
  assign new_new_n21300__ = ~new_new_n20848__ & ~new_new_n21299__;
  assign new_new_n21301__ = ~new_new_n20840__ & ~new_new_n21300__;
  assign new_new_n21302__ = ~new_new_n20839__ & ~new_new_n21301__;
  assign new_new_n21303__ = ~new_new_n20831__ & ~new_new_n21302__;
  assign new_new_n21304__ = ~new_new_n20830__ & ~new_new_n21303__;
  assign new_new_n21305__ = ~new_new_n20822__ & ~new_new_n21304__;
  assign new_new_n21306__ = ~new_new_n20821__ & ~new_new_n21305__;
  assign new_new_n21307__ = ~new_new_n20813__ & ~new_new_n21306__;
  assign new_new_n21308__ = ~new_new_n20812__ & ~new_new_n21307__;
  assign new_new_n21309__ = ~new_new_n20804__ & ~new_new_n21308__;
  assign new_new_n21310__ = ~new_new_n20803__ & ~new_new_n21309__;
  assign new_new_n21311__ = ~new_new_n20795__ & ~new_new_n21310__;
  assign new_new_n21312__ = ~new_new_n20794__ & ~new_new_n21311__;
  assign new_new_n21313__ = ~new_new_n20786__ & ~new_new_n21312__;
  assign new_new_n21314__ = ~new_new_n20785__ & ~new_new_n21313__;
  assign new_new_n21315__ = ~new_new_n20777__ & new_new_n21314__;
  assign new_new_n21316__ = ~new_new_n20776__ & ~new_new_n21315__;
  assign new_new_n21317__ = ~new_new_n20768__ & ~new_new_n21316__;
  assign new_new_n21318__ = ~new_new_n20767__ & ~new_new_n21317__;
  assign new_new_n21319__ = ~new_new_n20759__ & ~new_new_n21318__;
  assign new_new_n21320__ = ~new_new_n20758__ & ~new_new_n21319__;
  assign new_new_n21321__ = ~new_new_n20750__ & ~new_new_n21320__;
  assign new_new_n21322__ = ~new_new_n20749__ & ~new_new_n21321__;
  assign new_new_n21323__ = ~new_new_n20741__ & ~new_new_n21322__;
  assign new_new_n21324__ = ~new_new_n20740__ & ~new_new_n21323__;
  assign new_new_n21325__ = ~new_new_n20732__ & ~new_new_n21324__;
  assign new_new_n21326__ = ~new_new_n20731__ & ~new_new_n21325__;
  assign new_new_n21327__ = ~new_new_n20723__ & ~new_new_n21326__;
  assign new_new_n21328__ = ~new_new_n20722__ & ~new_new_n21327__;
  assign new_new_n21329__ = ~new_new_n20714__ & new_new_n21328__;
  assign new_new_n21330__ = ~new_new_n20713__ & ~new_new_n21329__;
  assign new_new_n21331__ = ~new_new_n20705__ & ~new_new_n21330__;
  assign new_new_n21332__ = ~new_new_n20704__ & ~new_new_n21331__;
  assign new_new_n21333__ = ~new_new_n20696__ & ~new_new_n21332__;
  assign new_new_n21334__ = ~new_new_n20695__ & ~new_new_n21333__;
  assign new_new_n21335__ = ~new_new_n20687__ & ~new_new_n21334__;
  assign new_new_n21336__ = ~new_new_n20686__ & ~new_new_n21335__;
  assign new_new_n21337__ = ~pi124 & new_new_n21336__;
  assign new_new_n21338__ = ~new_new_n20018__ & ~new_new_n21337__;
  assign new_new_n21339__ = ~pi125 & new_new_n260__;
  assign new_new_n21340__ = ~pi124 & new_new_n20677__;
  assign new_new_n21341__ = ~new_new_n21336__ & ~new_new_n21340__;
  assign new_new_n21342__ = new_new_n21339__ & ~new_new_n21341__;
  assign po003 = ~new_new_n21338__ & new_new_n21342__;
  assign new_new_n21344__ = pi123 & ~new_new_n21334__;
  assign new_new_n21345__ = ~pi123 & new_new_n21334__;
  assign new_new_n21346__ = ~new_new_n21344__ & ~new_new_n21345__;
  assign new_new_n21347__ = po003 & new_new_n21346__;
  assign new_new_n21348__ = new_new_n20685__ & new_new_n21347__;
  assign new_new_n21349__ = ~new_new_n20685__ & ~new_new_n21347__;
  assign new_new_n21350__ = ~new_new_n21348__ & ~new_new_n21349__;
  assign new_new_n21351__ = ~pi124 & new_new_n21350__;
  assign new_new_n21352__ = pi124 & ~new_new_n21350__;
  assign new_new_n21353__ = ~new_new_n21351__ & ~new_new_n21352__;
  assign new_new_n21354__ = ~new_new_n20695__ & ~new_new_n20696__;
  assign new_new_n21355__ = ~new_new_n21332__ & po003;
  assign new_new_n21356__ = pi122 & ~po003;
  assign new_new_n21357__ = ~new_new_n21355__ & ~new_new_n21356__;
  assign new_new_n21358__ = new_new_n21354__ & ~new_new_n21357__;
  assign new_new_n21359__ = ~new_new_n21354__ & new_new_n21357__;
  assign new_new_n21360__ = ~new_new_n21358__ & ~new_new_n21359__;
  assign new_new_n21361__ = ~pi123 & ~new_new_n21360__;
  assign new_new_n21362__ = pi123 & new_new_n21360__;
  assign new_new_n21363__ = ~new_new_n20704__ & ~new_new_n20705__;
  assign new_new_n21364__ = ~new_new_n21330__ & po003;
  assign new_new_n21365__ = pi121 & ~po003;
  assign new_new_n21366__ = ~new_new_n21364__ & ~new_new_n21365__;
  assign new_new_n21367__ = new_new_n21363__ & ~new_new_n21366__;
  assign new_new_n21368__ = ~new_new_n21363__ & new_new_n21366__;
  assign new_new_n21369__ = ~new_new_n21367__ & ~new_new_n21368__;
  assign new_new_n21370__ = ~pi122 & ~new_new_n21369__;
  assign new_new_n21371__ = pi122 & new_new_n21369__;
  assign new_new_n21372__ = ~new_new_n20713__ & ~new_new_n20714__;
  assign new_new_n21373__ = ~new_new_n21328__ & po003;
  assign new_new_n21374__ = ~pi120 & ~po003;
  assign new_new_n21375__ = ~new_new_n21373__ & ~new_new_n21374__;
  assign new_new_n21376__ = new_new_n21372__ & ~new_new_n21375__;
  assign new_new_n21377__ = ~new_new_n21372__ & new_new_n21375__;
  assign new_new_n21378__ = ~new_new_n21376__ & ~new_new_n21377__;
  assign new_new_n21379__ = pi121 & ~new_new_n21378__;
  assign new_new_n21380__ = ~pi121 & new_new_n21378__;
  assign new_new_n21381__ = ~new_new_n20722__ & ~new_new_n20723__;
  assign new_new_n21382__ = ~new_new_n21326__ & po003;
  assign new_new_n21383__ = ~pi119 & ~po003;
  assign new_new_n21384__ = ~new_new_n21382__ & ~new_new_n21383__;
  assign new_new_n21385__ = new_new_n21381__ & ~new_new_n21384__;
  assign new_new_n21386__ = ~new_new_n21381__ & new_new_n21384__;
  assign new_new_n21387__ = ~new_new_n21385__ & ~new_new_n21386__;
  assign new_new_n21388__ = pi120 & ~new_new_n21387__;
  assign new_new_n21389__ = ~pi120 & new_new_n21387__;
  assign new_new_n21390__ = ~new_new_n20731__ & ~new_new_n20732__;
  assign new_new_n21391__ = ~new_new_n21324__ & po003;
  assign new_new_n21392__ = ~pi118 & ~po003;
  assign new_new_n21393__ = ~new_new_n21391__ & ~new_new_n21392__;
  assign new_new_n21394__ = new_new_n21390__ & ~new_new_n21393__;
  assign new_new_n21395__ = ~new_new_n21390__ & new_new_n21393__;
  assign new_new_n21396__ = ~new_new_n21394__ & ~new_new_n21395__;
  assign new_new_n21397__ = pi119 & ~new_new_n21396__;
  assign new_new_n21398__ = ~pi119 & new_new_n21396__;
  assign new_new_n21399__ = ~new_new_n20740__ & ~new_new_n20741__;
  assign new_new_n21400__ = ~new_new_n21322__ & po003;
  assign new_new_n21401__ = ~pi117 & ~po003;
  assign new_new_n21402__ = ~new_new_n21400__ & ~new_new_n21401__;
  assign new_new_n21403__ = new_new_n21399__ & ~new_new_n21402__;
  assign new_new_n21404__ = ~new_new_n21399__ & new_new_n21402__;
  assign new_new_n21405__ = ~new_new_n21403__ & ~new_new_n21404__;
  assign new_new_n21406__ = pi118 & ~new_new_n21405__;
  assign new_new_n21407__ = ~pi118 & new_new_n21405__;
  assign new_new_n21408__ = ~new_new_n20749__ & ~new_new_n20750__;
  assign new_new_n21409__ = ~new_new_n21320__ & po003;
  assign new_new_n21410__ = ~pi116 & ~po003;
  assign new_new_n21411__ = ~new_new_n21409__ & ~new_new_n21410__;
  assign new_new_n21412__ = new_new_n21408__ & ~new_new_n21411__;
  assign new_new_n21413__ = ~new_new_n21408__ & new_new_n21411__;
  assign new_new_n21414__ = ~new_new_n21412__ & ~new_new_n21413__;
  assign new_new_n21415__ = pi117 & ~new_new_n21414__;
  assign new_new_n21416__ = ~pi117 & new_new_n21414__;
  assign new_new_n21417__ = ~pi115 & ~new_new_n21318__;
  assign new_new_n21418__ = pi115 & new_new_n21318__;
  assign new_new_n21419__ = ~new_new_n21417__ & ~new_new_n21418__;
  assign new_new_n21420__ = po003 & new_new_n21419__;
  assign new_new_n21421__ = new_new_n20757__ & new_new_n21420__;
  assign new_new_n21422__ = ~new_new_n20757__ & ~new_new_n21420__;
  assign new_new_n21423__ = ~new_new_n21421__ & ~new_new_n21422__;
  assign new_new_n21424__ = ~pi116 & ~new_new_n21423__;
  assign new_new_n21425__ = pi116 & new_new_n21423__;
  assign new_new_n21426__ = ~pi114 & ~new_new_n21316__;
  assign new_new_n21427__ = pi114 & new_new_n21316__;
  assign new_new_n21428__ = ~new_new_n21426__ & ~new_new_n21427__;
  assign new_new_n21429__ = po003 & new_new_n21428__;
  assign new_new_n21430__ = ~new_new_n20766__ & ~new_new_n21429__;
  assign new_new_n21431__ = new_new_n20766__ & new_new_n21429__;
  assign new_new_n21432__ = ~new_new_n21430__ & ~new_new_n21431__;
  assign new_new_n21433__ = ~pi115 & ~new_new_n21432__;
  assign new_new_n21434__ = pi115 & new_new_n21432__;
  assign new_new_n21435__ = ~new_new_n20776__ & ~new_new_n20777__;
  assign new_new_n21436__ = ~new_new_n21314__ & po003;
  assign new_new_n21437__ = pi113 & ~po003;
  assign new_new_n21438__ = ~new_new_n21436__ & ~new_new_n21437__;
  assign new_new_n21439__ = new_new_n21435__ & ~new_new_n21438__;
  assign new_new_n21440__ = ~new_new_n21435__ & new_new_n21438__;
  assign new_new_n21441__ = ~new_new_n21439__ & ~new_new_n21440__;
  assign new_new_n21442__ = ~pi114 & ~new_new_n21441__;
  assign new_new_n21443__ = pi114 & new_new_n21441__;
  assign new_new_n21444__ = pi112 & ~new_new_n21312__;
  assign new_new_n21445__ = ~pi112 & new_new_n21312__;
  assign new_new_n21446__ = ~new_new_n21444__ & ~new_new_n21445__;
  assign new_new_n21447__ = po003 & new_new_n21446__;
  assign new_new_n21448__ = ~new_new_n20784__ & new_new_n21447__;
  assign new_new_n21449__ = new_new_n20784__ & ~new_new_n21447__;
  assign new_new_n21450__ = ~new_new_n21448__ & ~new_new_n21449__;
  assign new_new_n21451__ = ~pi113 & ~new_new_n21450__;
  assign new_new_n21452__ = pi113 & new_new_n21450__;
  assign new_new_n21453__ = ~new_new_n21310__ & po003;
  assign new_new_n21454__ = pi111 & ~po003;
  assign new_new_n21455__ = ~new_new_n21453__ & ~new_new_n21454__;
  assign new_new_n21456__ = ~new_new_n20794__ & ~new_new_n20795__;
  assign new_new_n21457__ = ~new_new_n21455__ & new_new_n21456__;
  assign new_new_n21458__ = new_new_n21455__ & ~new_new_n21456__;
  assign new_new_n21459__ = ~new_new_n21457__ & ~new_new_n21458__;
  assign new_new_n21460__ = ~pi112 & ~new_new_n21459__;
  assign new_new_n21461__ = pi112 & new_new_n21459__;
  assign new_new_n21462__ = ~new_new_n20803__ & ~new_new_n20804__;
  assign new_new_n21463__ = ~new_new_n21308__ & po003;
  assign new_new_n21464__ = pi110 & ~po003;
  assign new_new_n21465__ = ~new_new_n21463__ & ~new_new_n21464__;
  assign new_new_n21466__ = new_new_n21462__ & ~new_new_n21465__;
  assign new_new_n21467__ = ~new_new_n21462__ & new_new_n21465__;
  assign new_new_n21468__ = ~new_new_n21466__ & ~new_new_n21467__;
  assign new_new_n21469__ = pi111 & new_new_n21468__;
  assign new_new_n21470__ = ~pi111 & ~new_new_n21468__;
  assign new_new_n21471__ = ~pi109 & ~new_new_n21306__;
  assign new_new_n21472__ = pi109 & new_new_n21306__;
  assign new_new_n21473__ = ~new_new_n21471__ & ~new_new_n21472__;
  assign new_new_n21474__ = po003 & ~new_new_n21473__;
  assign new_new_n21475__ = new_new_n20811__ & new_new_n21474__;
  assign new_new_n21476__ = ~new_new_n20811__ & ~new_new_n21474__;
  assign new_new_n21477__ = ~new_new_n21475__ & ~new_new_n21476__;
  assign new_new_n21478__ = pi110 & ~new_new_n21477__;
  assign new_new_n21479__ = ~pi110 & new_new_n21477__;
  assign new_new_n21480__ = ~new_new_n20821__ & ~new_new_n20822__;
  assign new_new_n21481__ = ~new_new_n21304__ & po003;
  assign new_new_n21482__ = pi108 & ~po003;
  assign new_new_n21483__ = ~new_new_n21481__ & ~new_new_n21482__;
  assign new_new_n21484__ = new_new_n21480__ & new_new_n21483__;
  assign new_new_n21485__ = ~new_new_n21480__ & ~new_new_n21483__;
  assign new_new_n21486__ = ~new_new_n21484__ & ~new_new_n21485__;
  assign new_new_n21487__ = pi109 & ~new_new_n21486__;
  assign new_new_n21488__ = ~pi109 & new_new_n21486__;
  assign new_new_n21489__ = ~new_new_n20830__ & ~new_new_n20831__;
  assign new_new_n21490__ = ~new_new_n21302__ & po003;
  assign new_new_n21491__ = pi107 & ~po003;
  assign new_new_n21492__ = ~new_new_n21490__ & ~new_new_n21491__;
  assign new_new_n21493__ = new_new_n21489__ & ~new_new_n21492__;
  assign new_new_n21494__ = ~new_new_n21489__ & new_new_n21492__;
  assign new_new_n21495__ = ~new_new_n21493__ & ~new_new_n21494__;
  assign new_new_n21496__ = ~pi108 & ~new_new_n21495__;
  assign new_new_n21497__ = pi108 & new_new_n21495__;
  assign new_new_n21498__ = ~new_new_n21300__ & po003;
  assign new_new_n21499__ = pi106 & ~po003;
  assign new_new_n21500__ = ~new_new_n21498__ & ~new_new_n21499__;
  assign new_new_n21501__ = ~new_new_n20839__ & ~new_new_n20840__;
  assign new_new_n21502__ = ~new_new_n21500__ & new_new_n21501__;
  assign new_new_n21503__ = new_new_n21500__ & ~new_new_n21501__;
  assign new_new_n21504__ = ~new_new_n21502__ & ~new_new_n21503__;
  assign new_new_n21505__ = ~pi107 & ~new_new_n21504__;
  assign new_new_n21506__ = pi107 & new_new_n21504__;
  assign new_new_n21507__ = ~new_new_n21298__ & po003;
  assign new_new_n21508__ = pi105 & ~po003;
  assign new_new_n21509__ = ~new_new_n21507__ & ~new_new_n21508__;
  assign new_new_n21510__ = ~new_new_n20848__ & ~new_new_n20849__;
  assign new_new_n21511__ = ~new_new_n21509__ & new_new_n21510__;
  assign new_new_n21512__ = new_new_n21509__ & ~new_new_n21510__;
  assign new_new_n21513__ = ~new_new_n21511__ & ~new_new_n21512__;
  assign new_new_n21514__ = ~pi106 & ~new_new_n21513__;
  assign new_new_n21515__ = pi106 & new_new_n21513__;
  assign new_new_n21516__ = ~new_new_n21296__ & po003;
  assign new_new_n21517__ = pi104 & ~po003;
  assign new_new_n21518__ = ~new_new_n21516__ & ~new_new_n21517__;
  assign new_new_n21519__ = ~new_new_n20857__ & ~new_new_n20858__;
  assign new_new_n21520__ = ~new_new_n21518__ & new_new_n21519__;
  assign new_new_n21521__ = new_new_n21518__ & ~new_new_n21519__;
  assign new_new_n21522__ = ~new_new_n21520__ & ~new_new_n21521__;
  assign new_new_n21523__ = ~pi105 & ~new_new_n21522__;
  assign new_new_n21524__ = pi105 & new_new_n21522__;
  assign new_new_n21525__ = pi103 & ~new_new_n21294__;
  assign new_new_n21526__ = ~pi103 & new_new_n21294__;
  assign new_new_n21527__ = ~new_new_n21525__ & ~new_new_n21526__;
  assign new_new_n21528__ = po003 & new_new_n21527__;
  assign new_new_n21529__ = new_new_n20865__ & new_new_n21528__;
  assign new_new_n21530__ = ~new_new_n20865__ & ~new_new_n21528__;
  assign new_new_n21531__ = ~new_new_n21529__ & ~new_new_n21530__;
  assign new_new_n21532__ = ~pi104 & new_new_n21531__;
  assign new_new_n21533__ = pi104 & ~new_new_n21531__;
  assign new_new_n21534__ = pi102 & ~new_new_n21292__;
  assign new_new_n21535__ = ~pi102 & new_new_n21292__;
  assign new_new_n21536__ = ~new_new_n21534__ & ~new_new_n21535__;
  assign new_new_n21537__ = po003 & new_new_n21536__;
  assign new_new_n21538__ = new_new_n20874__ & new_new_n21537__;
  assign new_new_n21539__ = ~new_new_n20874__ & ~new_new_n21537__;
  assign new_new_n21540__ = ~new_new_n21538__ & ~new_new_n21539__;
  assign new_new_n21541__ = ~pi103 & new_new_n21540__;
  assign new_new_n21542__ = pi103 & ~new_new_n21540__;
  assign new_new_n21543__ = ~new_new_n20884__ & ~new_new_n20885__;
  assign new_new_n21544__ = ~new_new_n21290__ & po003;
  assign new_new_n21545__ = ~pi101 & ~po003;
  assign new_new_n21546__ = ~new_new_n21544__ & ~new_new_n21545__;
  assign new_new_n21547__ = new_new_n21543__ & ~new_new_n21546__;
  assign new_new_n21548__ = ~new_new_n21543__ & new_new_n21546__;
  assign new_new_n21549__ = ~new_new_n21547__ & ~new_new_n21548__;
  assign new_new_n21550__ = ~pi102 & new_new_n21549__;
  assign new_new_n21551__ = pi102 & ~new_new_n21549__;
  assign new_new_n21552__ = ~new_new_n20893__ & ~new_new_n20894__;
  assign new_new_n21553__ = ~new_new_n21288__ & po003;
  assign new_new_n21554__ = ~pi100 & ~po003;
  assign new_new_n21555__ = ~new_new_n21553__ & ~new_new_n21554__;
  assign new_new_n21556__ = new_new_n21552__ & ~new_new_n21555__;
  assign new_new_n21557__ = ~new_new_n21552__ & new_new_n21555__;
  assign new_new_n21558__ = ~new_new_n21556__ & ~new_new_n21557__;
  assign new_new_n21559__ = ~pi101 & new_new_n21558__;
  assign new_new_n21560__ = pi101 & ~new_new_n21558__;
  assign new_new_n21561__ = ~pi099 & ~new_new_n21286__;
  assign new_new_n21562__ = pi099 & new_new_n21286__;
  assign new_new_n21563__ = ~new_new_n21561__ & ~new_new_n21562__;
  assign new_new_n21564__ = po003 & new_new_n21563__;
  assign new_new_n21565__ = new_new_n20901__ & new_new_n21564__;
  assign new_new_n21566__ = ~new_new_n20901__ & ~new_new_n21564__;
  assign new_new_n21567__ = ~new_new_n21565__ & ~new_new_n21566__;
  assign new_new_n21568__ = ~pi100 & ~new_new_n21567__;
  assign new_new_n21569__ = pi100 & new_new_n21567__;
  assign new_new_n21570__ = ~new_new_n20911__ & ~new_new_n20912__;
  assign new_new_n21571__ = new_new_n21284__ & po003;
  assign new_new_n21572__ = ~pi098 & ~po003;
  assign new_new_n21573__ = ~new_new_n21571__ & ~new_new_n21572__;
  assign new_new_n21574__ = ~new_new_n21570__ & ~new_new_n21573__;
  assign new_new_n21575__ = new_new_n21570__ & new_new_n21573__;
  assign new_new_n21576__ = ~new_new_n21574__ & ~new_new_n21575__;
  assign new_new_n21577__ = ~pi099 & ~new_new_n21576__;
  assign new_new_n21578__ = pi099 & new_new_n21576__;
  assign new_new_n21579__ = new_new_n21282__ & po003;
  assign new_new_n21580__ = pi097 & ~po003;
  assign new_new_n21581__ = ~new_new_n21579__ & ~new_new_n21580__;
  assign new_new_n21582__ = ~new_new_n20920__ & ~new_new_n20921__;
  assign new_new_n21583__ = ~new_new_n21581__ & ~new_new_n21582__;
  assign new_new_n21584__ = new_new_n21581__ & new_new_n21582__;
  assign new_new_n21585__ = ~new_new_n21583__ & ~new_new_n21584__;
  assign new_new_n21586__ = pi098 & ~new_new_n21585__;
  assign new_new_n21587__ = ~pi098 & new_new_n21585__;
  assign new_new_n21588__ = ~new_new_n20929__ & ~new_new_n20930__;
  assign new_new_n21589__ = ~new_new_n21280__ & po003;
  assign new_new_n21590__ = ~pi096 & ~po003;
  assign new_new_n21591__ = ~new_new_n21589__ & ~new_new_n21590__;
  assign new_new_n21592__ = new_new_n21588__ & ~new_new_n21591__;
  assign new_new_n21593__ = ~new_new_n21588__ & new_new_n21591__;
  assign new_new_n21594__ = ~new_new_n21592__ & ~new_new_n21593__;
  assign new_new_n21595__ = pi097 & ~new_new_n21594__;
  assign new_new_n21596__ = ~pi097 & new_new_n21594__;
  assign new_new_n21597__ = ~pi095 & ~new_new_n21278__;
  assign new_new_n21598__ = pi095 & new_new_n21278__;
  assign new_new_n21599__ = ~new_new_n21597__ & ~new_new_n21598__;
  assign new_new_n21600__ = po003 & new_new_n21599__;
  assign new_new_n21601__ = new_new_n20937__ & ~new_new_n21600__;
  assign new_new_n21602__ = ~new_new_n20937__ & new_new_n21600__;
  assign new_new_n21603__ = ~new_new_n21601__ & ~new_new_n21602__;
  assign new_new_n21604__ = pi096 & ~new_new_n21603__;
  assign new_new_n21605__ = ~pi096 & new_new_n21603__;
  assign new_new_n21606__ = ~new_new_n21276__ & po003;
  assign new_new_n21607__ = pi094 & ~po003;
  assign new_new_n21608__ = ~new_new_n21606__ & ~new_new_n21607__;
  assign new_new_n21609__ = ~new_new_n20947__ & ~new_new_n20948__;
  assign new_new_n21610__ = ~new_new_n21608__ & new_new_n21609__;
  assign new_new_n21611__ = new_new_n21608__ & ~new_new_n21609__;
  assign new_new_n21612__ = ~new_new_n21610__ & ~new_new_n21611__;
  assign new_new_n21613__ = pi095 & new_new_n21612__;
  assign new_new_n21614__ = ~pi095 & ~new_new_n21612__;
  assign new_new_n21615__ = pi093 & ~new_new_n21274__;
  assign new_new_n21616__ = ~pi093 & new_new_n21274__;
  assign new_new_n21617__ = ~new_new_n21615__ & ~new_new_n21616__;
  assign new_new_n21618__ = po003 & new_new_n21617__;
  assign new_new_n21619__ = new_new_n20955__ & new_new_n21618__;
  assign new_new_n21620__ = ~new_new_n20955__ & ~new_new_n21618__;
  assign new_new_n21621__ = ~new_new_n21619__ & ~new_new_n21620__;
  assign new_new_n21622__ = pi094 & ~new_new_n21621__;
  assign new_new_n21623__ = ~pi094 & new_new_n21621__;
  assign new_new_n21624__ = ~new_new_n21272__ & po003;
  assign new_new_n21625__ = pi092 & ~po003;
  assign new_new_n21626__ = ~new_new_n21624__ & ~new_new_n21625__;
  assign new_new_n21627__ = ~new_new_n20965__ & ~new_new_n20966__;
  assign new_new_n21628__ = ~new_new_n21626__ & new_new_n21627__;
  assign new_new_n21629__ = new_new_n21626__ & ~new_new_n21627__;
  assign new_new_n21630__ = ~new_new_n21628__ & ~new_new_n21629__;
  assign new_new_n21631__ = ~pi093 & ~new_new_n21630__;
  assign new_new_n21632__ = pi093 & new_new_n21630__;
  assign new_new_n21633__ = ~new_new_n20974__ & ~new_new_n20975__;
  assign new_new_n21634__ = ~new_new_n21270__ & po003;
  assign new_new_n21635__ = pi091 & ~po003;
  assign new_new_n21636__ = ~new_new_n21634__ & ~new_new_n21635__;
  assign new_new_n21637__ = new_new_n21633__ & ~new_new_n21636__;
  assign new_new_n21638__ = ~new_new_n21633__ & new_new_n21636__;
  assign new_new_n21639__ = ~new_new_n21637__ & ~new_new_n21638__;
  assign new_new_n21640__ = ~pi092 & ~new_new_n21639__;
  assign new_new_n21641__ = pi092 & new_new_n21639__;
  assign new_new_n21642__ = ~new_new_n20983__ & ~new_new_n20984__;
  assign new_new_n21643__ = new_new_n21268__ & po003;
  assign new_new_n21644__ = ~pi090 & ~po003;
  assign new_new_n21645__ = ~new_new_n21643__ & ~new_new_n21644__;
  assign new_new_n21646__ = ~new_new_n21642__ & ~new_new_n21645__;
  assign new_new_n21647__ = new_new_n21642__ & new_new_n21645__;
  assign new_new_n21648__ = ~new_new_n21646__ & ~new_new_n21647__;
  assign new_new_n21649__ = pi091 & new_new_n21648__;
  assign new_new_n21650__ = ~pi091 & ~new_new_n21648__;
  assign new_new_n21651__ = ~new_new_n20992__ & ~new_new_n20993__;
  assign new_new_n21652__ = ~new_new_n21266__ & po003;
  assign new_new_n21653__ = pi089 & ~po003;
  assign new_new_n21654__ = ~new_new_n21652__ & ~new_new_n21653__;
  assign new_new_n21655__ = new_new_n21651__ & new_new_n21654__;
  assign new_new_n21656__ = ~new_new_n21651__ & ~new_new_n21654__;
  assign new_new_n21657__ = ~new_new_n21655__ & ~new_new_n21656__;
  assign new_new_n21658__ = pi090 & ~new_new_n21657__;
  assign new_new_n21659__ = ~pi090 & new_new_n21657__;
  assign new_new_n21660__ = new_new_n21264__ & po003;
  assign new_new_n21661__ = pi088 & ~po003;
  assign new_new_n21662__ = ~new_new_n21660__ & ~new_new_n21661__;
  assign new_new_n21663__ = ~new_new_n21001__ & ~new_new_n21002__;
  assign new_new_n21664__ = ~new_new_n21662__ & ~new_new_n21663__;
  assign new_new_n21665__ = new_new_n21662__ & new_new_n21663__;
  assign new_new_n21666__ = ~new_new_n21664__ & ~new_new_n21665__;
  assign new_new_n21667__ = pi089 & ~new_new_n21666__;
  assign new_new_n21668__ = ~pi089 & new_new_n21666__;
  assign new_new_n21669__ = ~pi087 & ~new_new_n21262__;
  assign new_new_n21670__ = pi087 & new_new_n21262__;
  assign new_new_n21671__ = ~new_new_n21669__ & ~new_new_n21670__;
  assign new_new_n21672__ = po003 & new_new_n21671__;
  assign new_new_n21673__ = new_new_n21009__ & new_new_n21672__;
  assign new_new_n21674__ = ~new_new_n21009__ & ~new_new_n21672__;
  assign new_new_n21675__ = ~new_new_n21673__ & ~new_new_n21674__;
  assign new_new_n21676__ = ~pi088 & ~new_new_n21675__;
  assign new_new_n21677__ = pi088 & new_new_n21675__;
  assign new_new_n21678__ = ~new_new_n21019__ & ~new_new_n21020__;
  assign new_new_n21679__ = ~new_new_n21260__ & po003;
  assign new_new_n21680__ = pi086 & ~po003;
  assign new_new_n21681__ = ~new_new_n21679__ & ~new_new_n21680__;
  assign new_new_n21682__ = new_new_n21678__ & ~new_new_n21681__;
  assign new_new_n21683__ = ~new_new_n21678__ & new_new_n21681__;
  assign new_new_n21684__ = ~new_new_n21682__ & ~new_new_n21683__;
  assign new_new_n21685__ = ~pi087 & ~new_new_n21684__;
  assign new_new_n21686__ = pi087 & new_new_n21684__;
  assign new_new_n21687__ = ~new_new_n21028__ & ~new_new_n21029__;
  assign new_new_n21688__ = ~new_new_n21258__ & po003;
  assign new_new_n21689__ = ~pi085 & ~po003;
  assign new_new_n21690__ = ~new_new_n21688__ & ~new_new_n21689__;
  assign new_new_n21691__ = new_new_n21687__ & new_new_n21690__;
  assign new_new_n21692__ = ~new_new_n21687__ & ~new_new_n21690__;
  assign new_new_n21693__ = ~new_new_n21691__ & ~new_new_n21692__;
  assign new_new_n21694__ = ~pi086 & ~new_new_n21693__;
  assign new_new_n21695__ = pi086 & new_new_n21693__;
  assign new_new_n21696__ = new_new_n21256__ & po003;
  assign new_new_n21697__ = pi084 & ~po003;
  assign new_new_n21698__ = ~new_new_n21696__ & ~new_new_n21697__;
  assign new_new_n21699__ = ~new_new_n21037__ & ~new_new_n21038__;
  assign new_new_n21700__ = ~new_new_n21698__ & ~new_new_n21699__;
  assign new_new_n21701__ = new_new_n21698__ & new_new_n21699__;
  assign new_new_n21702__ = ~new_new_n21700__ & ~new_new_n21701__;
  assign new_new_n21703__ = pi085 & ~new_new_n21702__;
  assign new_new_n21704__ = ~pi085 & new_new_n21702__;
  assign new_new_n21705__ = ~new_new_n21046__ & ~new_new_n21047__;
  assign new_new_n21706__ = ~new_new_n21254__ & po003;
  assign new_new_n21707__ = ~pi083 & ~po003;
  assign new_new_n21708__ = ~new_new_n21706__ & ~new_new_n21707__;
  assign new_new_n21709__ = new_new_n21705__ & ~new_new_n21708__;
  assign new_new_n21710__ = ~new_new_n21705__ & new_new_n21708__;
  assign new_new_n21711__ = ~new_new_n21709__ & ~new_new_n21710__;
  assign new_new_n21712__ = pi084 & ~new_new_n21711__;
  assign new_new_n21713__ = ~pi084 & new_new_n21711__;
  assign new_new_n21714__ = ~new_new_n21055__ & ~new_new_n21056__;
  assign new_new_n21715__ = ~new_new_n21252__ & po003;
  assign new_new_n21716__ = ~pi082 & ~po003;
  assign new_new_n21717__ = ~new_new_n21715__ & ~new_new_n21716__;
  assign new_new_n21718__ = new_new_n21714__ & ~new_new_n21717__;
  assign new_new_n21719__ = ~new_new_n21714__ & new_new_n21717__;
  assign new_new_n21720__ = ~new_new_n21718__ & ~new_new_n21719__;
  assign new_new_n21721__ = pi083 & ~new_new_n21720__;
  assign new_new_n21722__ = ~pi083 & new_new_n21720__;
  assign new_new_n21723__ = ~new_new_n21064__ & ~new_new_n21065__;
  assign new_new_n21724__ = ~new_new_n21250__ & po003;
  assign new_new_n21725__ = ~pi081 & ~po003;
  assign new_new_n21726__ = ~new_new_n21724__ & ~new_new_n21725__;
  assign new_new_n21727__ = new_new_n21723__ & ~new_new_n21726__;
  assign new_new_n21728__ = ~new_new_n21723__ & new_new_n21726__;
  assign new_new_n21729__ = ~new_new_n21727__ & ~new_new_n21728__;
  assign new_new_n21730__ = pi082 & ~new_new_n21729__;
  assign new_new_n21731__ = ~pi082 & new_new_n21729__;
  assign new_new_n21732__ = ~new_new_n21073__ & ~new_new_n21074__;
  assign new_new_n21733__ = ~new_new_n21248__ & po003;
  assign new_new_n21734__ = ~pi080 & ~po003;
  assign new_new_n21735__ = ~new_new_n21733__ & ~new_new_n21734__;
  assign new_new_n21736__ = new_new_n21732__ & ~new_new_n21735__;
  assign new_new_n21737__ = ~new_new_n21732__ & new_new_n21735__;
  assign new_new_n21738__ = ~new_new_n21736__ & ~new_new_n21737__;
  assign new_new_n21739__ = pi081 & ~new_new_n21738__;
  assign new_new_n21740__ = ~pi081 & new_new_n21738__;
  assign new_new_n21741__ = ~new_new_n21246__ & po003;
  assign new_new_n21742__ = pi079 & ~po003;
  assign new_new_n21743__ = ~new_new_n21741__ & ~new_new_n21742__;
  assign new_new_n21744__ = ~new_new_n21082__ & ~new_new_n21083__;
  assign new_new_n21745__ = ~new_new_n21743__ & new_new_n21744__;
  assign new_new_n21746__ = new_new_n21743__ & ~new_new_n21744__;
  assign new_new_n21747__ = ~new_new_n21745__ & ~new_new_n21746__;
  assign new_new_n21748__ = ~pi080 & ~new_new_n21747__;
  assign new_new_n21749__ = pi080 & new_new_n21747__;
  assign new_new_n21750__ = pi078 & ~new_new_n21244__;
  assign new_new_n21751__ = ~pi078 & new_new_n21244__;
  assign new_new_n21752__ = ~new_new_n21750__ & ~new_new_n21751__;
  assign new_new_n21753__ = po003 & new_new_n21752__;
  assign new_new_n21754__ = new_new_n21090__ & new_new_n21753__;
  assign new_new_n21755__ = ~new_new_n21090__ & ~new_new_n21753__;
  assign new_new_n21756__ = ~new_new_n21754__ & ~new_new_n21755__;
  assign new_new_n21757__ = pi079 & ~new_new_n21756__;
  assign new_new_n21758__ = ~pi079 & new_new_n21756__;
  assign new_new_n21759__ = ~new_new_n21100__ & ~new_new_n21101__;
  assign new_new_n21760__ = ~new_new_n21242__ & po003;
  assign new_new_n21761__ = pi077 & ~po003;
  assign new_new_n21762__ = ~new_new_n21760__ & ~new_new_n21761__;
  assign new_new_n21763__ = new_new_n21759__ & new_new_n21762__;
  assign new_new_n21764__ = ~new_new_n21759__ & ~new_new_n21762__;
  assign new_new_n21765__ = ~new_new_n21763__ & ~new_new_n21764__;
  assign new_new_n21766__ = pi078 & ~new_new_n21765__;
  assign new_new_n21767__ = ~pi078 & new_new_n21765__;
  assign new_new_n21768__ = new_new_n21240__ & po003;
  assign new_new_n21769__ = ~pi076 & ~po003;
  assign new_new_n21770__ = ~new_new_n21768__ & ~new_new_n21769__;
  assign new_new_n21771__ = ~new_new_n21109__ & ~new_new_n21110__;
  assign new_new_n21772__ = ~new_new_n21770__ & ~new_new_n21771__;
  assign new_new_n21773__ = new_new_n21770__ & new_new_n21771__;
  assign new_new_n21774__ = ~new_new_n21772__ & ~new_new_n21773__;
  assign new_new_n21775__ = pi077 & new_new_n21774__;
  assign new_new_n21776__ = ~pi077 & ~new_new_n21774__;
  assign new_new_n21777__ = ~new_new_n21118__ & ~new_new_n21119__;
  assign new_new_n21778__ = ~new_new_n21238__ & po003;
  assign new_new_n21779__ = pi075 & ~po003;
  assign new_new_n21780__ = ~new_new_n21778__ & ~new_new_n21779__;
  assign new_new_n21781__ = new_new_n21777__ & new_new_n21780__;
  assign new_new_n21782__ = ~new_new_n21777__ & ~new_new_n21780__;
  assign new_new_n21783__ = ~new_new_n21781__ & ~new_new_n21782__;
  assign new_new_n21784__ = pi076 & ~new_new_n21783__;
  assign new_new_n21785__ = ~pi076 & new_new_n21783__;
  assign new_new_n21786__ = new_new_n21236__ & po003;
  assign new_new_n21787__ = ~pi074 & ~po003;
  assign new_new_n21788__ = ~new_new_n21786__ & ~new_new_n21787__;
  assign new_new_n21789__ = ~new_new_n21127__ & ~new_new_n21128__;
  assign new_new_n21790__ = ~new_new_n21788__ & ~new_new_n21789__;
  assign new_new_n21791__ = new_new_n21788__ & new_new_n21789__;
  assign new_new_n21792__ = ~new_new_n21790__ & ~new_new_n21791__;
  assign new_new_n21793__ = pi075 & new_new_n21792__;
  assign new_new_n21794__ = ~pi075 & ~new_new_n21792__;
  assign new_new_n21795__ = ~new_new_n21136__ & ~new_new_n21137__;
  assign new_new_n21796__ = ~new_new_n21234__ & po003;
  assign new_new_n21797__ = pi073 & ~po003;
  assign new_new_n21798__ = ~new_new_n21796__ & ~new_new_n21797__;
  assign new_new_n21799__ = new_new_n21795__ & new_new_n21798__;
  assign new_new_n21800__ = ~new_new_n21795__ & ~new_new_n21798__;
  assign new_new_n21801__ = ~new_new_n21799__ & ~new_new_n21800__;
  assign new_new_n21802__ = pi074 & ~new_new_n21801__;
  assign new_new_n21803__ = ~pi074 & new_new_n21801__;
  assign new_new_n21804__ = pi072 & ~new_new_n21232__;
  assign new_new_n21805__ = ~pi072 & new_new_n21232__;
  assign new_new_n21806__ = ~new_new_n21804__ & ~new_new_n21805__;
  assign new_new_n21807__ = po003 & new_new_n21806__;
  assign new_new_n21808__ = new_new_n21144__ & new_new_n21807__;
  assign new_new_n21809__ = ~new_new_n21144__ & ~new_new_n21807__;
  assign new_new_n21810__ = ~new_new_n21808__ & ~new_new_n21809__;
  assign new_new_n21811__ = pi073 & ~new_new_n21810__;
  assign new_new_n21812__ = ~pi073 & new_new_n21810__;
  assign new_new_n21813__ = ~new_new_n21163__ & ~new_new_n21164__;
  assign new_new_n21814__ = ~new_new_n21228__ & po003;
  assign new_new_n21815__ = ~pi070 & ~po003;
  assign new_new_n21816__ = ~new_new_n21814__ & ~new_new_n21815__;
  assign new_new_n21817__ = ~new_new_n21813__ & ~new_new_n21816__;
  assign new_new_n21818__ = new_new_n21813__ & new_new_n21816__;
  assign new_new_n21819__ = ~new_new_n21817__ & ~new_new_n21818__;
  assign new_new_n21820__ = ~pi071 & ~new_new_n21819__;
  assign new_new_n21821__ = pi071 & new_new_n21819__;
  assign new_new_n21822__ = ~pi069 & ~new_new_n21226__;
  assign new_new_n21823__ = pi069 & new_new_n21226__;
  assign new_new_n21824__ = ~new_new_n21822__ & ~new_new_n21823__;
  assign new_new_n21825__ = po003 & new_new_n21824__;
  assign new_new_n21826__ = new_new_n21171__ & new_new_n21825__;
  assign new_new_n21827__ = ~new_new_n21171__ & ~new_new_n21825__;
  assign new_new_n21828__ = ~new_new_n21826__ & ~new_new_n21827__;
  assign new_new_n21829__ = pi070 & new_new_n21828__;
  assign new_new_n21830__ = ~pi070 & ~new_new_n21828__;
  assign new_new_n21831__ = ~new_new_n21181__ & ~new_new_n21182__;
  assign new_new_n21832__ = ~new_new_n21224__ & po003;
  assign new_new_n21833__ = ~pi068 & ~po003;
  assign new_new_n21834__ = ~new_new_n21832__ & ~new_new_n21833__;
  assign new_new_n21835__ = new_new_n21831__ & ~new_new_n21834__;
  assign new_new_n21836__ = ~new_new_n21831__ & new_new_n21834__;
  assign new_new_n21837__ = ~new_new_n21835__ & ~new_new_n21836__;
  assign new_new_n21838__ = pi069 & ~new_new_n21837__;
  assign new_new_n21839__ = ~pi069 & new_new_n21837__;
  assign new_new_n21840__ = ~new_new_n21204__ & ~new_new_n21205__;
  assign new_new_n21841__ = po003 & new_new_n21840__;
  assign new_new_n21842__ = new_new_n21220__ & new_new_n21841__;
  assign new_new_n21843__ = ~new_new_n21220__ & ~new_new_n21841__;
  assign new_new_n21844__ = ~new_new_n21842__ & ~new_new_n21843__;
  assign new_new_n21845__ = pi067 & ~new_new_n21844__;
  assign new_new_n21846__ = ~pi067 & new_new_n21844__;
  assign new_new_n21847__ = pi002 & ~pi065;
  assign new_new_n21848__ = pi003 & po003;
  assign new_new_n21849__ = ~pi004 & ~new_new_n21201__;
  assign new_new_n21850__ = pi004 & new_new_n21201__;
  assign new_new_n21851__ = ~new_new_n21849__ & ~new_new_n21850__;
  assign new_new_n21852__ = pi065 & new_new_n21851__;
  assign new_new_n21853__ = ~pi065 & ~new_new_n21851__;
  assign new_new_n21854__ = ~new_new_n21852__ & ~new_new_n21853__;
  assign new_new_n21855__ = ~new_new_n21847__ & ~new_new_n21854__;
  assign new_new_n21856__ = new_new_n21848__ & new_new_n21855__;
  assign new_new_n21857__ = ~pi003 & pi065;
  assign new_new_n21858__ = po003 & ~new_new_n21857__;
  assign new_new_n21859__ = ~pi002 & ~new_new_n21195__;
  assign new_new_n21860__ = ~new_new_n21851__ & new_new_n21859__;
  assign new_new_n21861__ = ~new_new_n21858__ & new_new_n21860__;
  assign new_new_n21862__ = ~new_new_n21856__ & ~new_new_n21861__;
  assign new_new_n21863__ = pi064 & ~new_new_n21862__;
  assign new_new_n21864__ = po003 & ~new_new_n21851__;
  assign new_new_n21865__ = pi064 & po003;
  assign new_new_n21866__ = new_new_n21857__ & ~new_new_n21865__;
  assign new_new_n21867__ = ~po003 & new_new_n21851__;
  assign new_new_n21868__ = ~new_new_n21864__ & ~new_new_n21867__;
  assign new_new_n21869__ = new_new_n21866__ & new_new_n21868__;
  assign new_new_n21870__ = ~pi066 & ~new_new_n21869__;
  assign new_new_n21871__ = ~new_new_n21863__ & new_new_n21870__;
  assign new_new_n21872__ = ~pi002 & pi065;
  assign new_new_n21873__ = ~pi003 & pi064;
  assign new_new_n21874__ = ~new_new_n21872__ & new_new_n21873__;
  assign new_new_n21875__ = ~new_new_n21854__ & new_new_n21874__;
  assign new_new_n21876__ = pi003 & new_new_n403__;
  assign new_new_n21877__ = ~new_new_n21851__ & new_new_n21876__;
  assign new_new_n21878__ = ~new_new_n21875__ & ~new_new_n21877__;
  assign new_new_n21879__ = po003 & ~new_new_n21878__;
  assign new_new_n21880__ = ~new_new_n21195__ & po003;
  assign new_new_n21881__ = pi002 & ~new_new_n21880__;
  assign new_new_n21882__ = ~new_new_n332__ & po003;
  assign new_new_n21883__ = pi064 & ~new_new_n21195__;
  assign new_new_n21884__ = ~new_new_n21882__ & ~new_new_n21883__;
  assign new_new_n21885__ = ~new_new_n21881__ & ~new_new_n21884__;
  assign new_new_n21886__ = new_new_n21851__ & ~new_new_n21857__;
  assign new_new_n21887__ = ~new_new_n21885__ & new_new_n21886__;
  assign new_new_n21888__ = ~new_new_n21879__ & ~new_new_n21887__;
  assign new_new_n21889__ = ~new_new_n21871__ & new_new_n21888__;
  assign new_new_n21890__ = ~new_new_n21846__ & new_new_n21889__;
  assign new_new_n21891__ = ~new_new_n21845__ & ~new_new_n21890__;
  assign new_new_n21892__ = pi068 & ~new_new_n21891__;
  assign new_new_n21893__ = ~pi068 & new_new_n21891__;
  assign new_new_n21894__ = ~new_new_n21190__ & ~new_new_n21191__;
  assign new_new_n21895__ = ~new_new_n21222__ & po003;
  assign new_new_n21896__ = ~pi067 & ~po003;
  assign new_new_n21897__ = ~new_new_n21895__ & ~new_new_n21896__;
  assign new_new_n21898__ = new_new_n21894__ & ~new_new_n21897__;
  assign new_new_n21899__ = ~new_new_n21894__ & new_new_n21897__;
  assign new_new_n21900__ = ~new_new_n21898__ & ~new_new_n21899__;
  assign new_new_n21901__ = ~new_new_n21893__ & ~new_new_n21900__;
  assign new_new_n21902__ = ~new_new_n21892__ & ~new_new_n21901__;
  assign new_new_n21903__ = ~new_new_n21839__ & ~new_new_n21902__;
  assign new_new_n21904__ = ~new_new_n21838__ & ~new_new_n21903__;
  assign new_new_n21905__ = ~new_new_n21830__ & ~new_new_n21904__;
  assign new_new_n21906__ = ~new_new_n21829__ & ~new_new_n21905__;
  assign new_new_n21907__ = ~new_new_n21821__ & new_new_n21906__;
  assign new_new_n21908__ = ~new_new_n21820__ & ~new_new_n21907__;
  assign new_new_n21909__ = pi072 & new_new_n21908__;
  assign new_new_n21910__ = ~pi072 & ~new_new_n21908__;
  assign new_new_n21911__ = ~new_new_n21154__ & ~new_new_n21155__;
  assign new_new_n21912__ = ~new_new_n21230__ & po003;
  assign new_new_n21913__ = ~pi071 & ~po003;
  assign new_new_n21914__ = ~new_new_n21912__ & ~new_new_n21913__;
  assign new_new_n21915__ = new_new_n21911__ & new_new_n21914__;
  assign new_new_n21916__ = ~new_new_n21911__ & ~new_new_n21914__;
  assign new_new_n21917__ = ~new_new_n21915__ & ~new_new_n21916__;
  assign new_new_n21918__ = ~new_new_n21910__ & new_new_n21917__;
  assign new_new_n21919__ = ~new_new_n21909__ & ~new_new_n21918__;
  assign new_new_n21920__ = ~new_new_n21812__ & ~new_new_n21919__;
  assign new_new_n21921__ = ~new_new_n21811__ & ~new_new_n21920__;
  assign new_new_n21922__ = ~new_new_n21803__ & ~new_new_n21921__;
  assign new_new_n21923__ = ~new_new_n21802__ & ~new_new_n21922__;
  assign new_new_n21924__ = ~new_new_n21794__ & ~new_new_n21923__;
  assign new_new_n21925__ = ~new_new_n21793__ & ~new_new_n21924__;
  assign new_new_n21926__ = ~new_new_n21785__ & ~new_new_n21925__;
  assign new_new_n21927__ = ~new_new_n21784__ & ~new_new_n21926__;
  assign new_new_n21928__ = ~new_new_n21776__ & ~new_new_n21927__;
  assign new_new_n21929__ = ~new_new_n21775__ & ~new_new_n21928__;
  assign new_new_n21930__ = ~new_new_n21767__ & ~new_new_n21929__;
  assign new_new_n21931__ = ~new_new_n21766__ & ~new_new_n21930__;
  assign new_new_n21932__ = ~new_new_n21758__ & ~new_new_n21931__;
  assign new_new_n21933__ = ~new_new_n21757__ & ~new_new_n21932__;
  assign new_new_n21934__ = ~new_new_n21749__ & new_new_n21933__;
  assign new_new_n21935__ = ~new_new_n21748__ & ~new_new_n21934__;
  assign new_new_n21936__ = ~new_new_n21740__ & new_new_n21935__;
  assign new_new_n21937__ = ~new_new_n21739__ & ~new_new_n21936__;
  assign new_new_n21938__ = ~new_new_n21731__ & ~new_new_n21937__;
  assign new_new_n21939__ = ~new_new_n21730__ & ~new_new_n21938__;
  assign new_new_n21940__ = ~new_new_n21722__ & ~new_new_n21939__;
  assign new_new_n21941__ = ~new_new_n21721__ & ~new_new_n21940__;
  assign new_new_n21942__ = ~new_new_n21713__ & ~new_new_n21941__;
  assign new_new_n21943__ = ~new_new_n21712__ & ~new_new_n21942__;
  assign new_new_n21944__ = ~new_new_n21704__ & ~new_new_n21943__;
  assign new_new_n21945__ = ~new_new_n21703__ & ~new_new_n21944__;
  assign new_new_n21946__ = ~new_new_n21695__ & new_new_n21945__;
  assign new_new_n21947__ = ~new_new_n21694__ & ~new_new_n21946__;
  assign new_new_n21948__ = ~new_new_n21686__ & ~new_new_n21947__;
  assign new_new_n21949__ = ~new_new_n21685__ & ~new_new_n21948__;
  assign new_new_n21950__ = ~new_new_n21677__ & ~new_new_n21949__;
  assign new_new_n21951__ = ~new_new_n21676__ & ~new_new_n21950__;
  assign new_new_n21952__ = ~new_new_n21668__ & new_new_n21951__;
  assign new_new_n21953__ = ~new_new_n21667__ & ~new_new_n21952__;
  assign new_new_n21954__ = ~new_new_n21659__ & ~new_new_n21953__;
  assign new_new_n21955__ = ~new_new_n21658__ & ~new_new_n21954__;
  assign new_new_n21956__ = ~new_new_n21650__ & ~new_new_n21955__;
  assign new_new_n21957__ = ~new_new_n21649__ & ~new_new_n21956__;
  assign new_new_n21958__ = ~new_new_n21641__ & new_new_n21957__;
  assign new_new_n21959__ = ~new_new_n21640__ & ~new_new_n21958__;
  assign new_new_n21960__ = ~new_new_n21632__ & ~new_new_n21959__;
  assign new_new_n21961__ = ~new_new_n21631__ & ~new_new_n21960__;
  assign new_new_n21962__ = ~new_new_n21623__ & new_new_n21961__;
  assign new_new_n21963__ = ~new_new_n21622__ & ~new_new_n21962__;
  assign new_new_n21964__ = ~new_new_n21614__ & ~new_new_n21963__;
  assign new_new_n21965__ = ~new_new_n21613__ & ~new_new_n21964__;
  assign new_new_n21966__ = ~new_new_n21605__ & ~new_new_n21965__;
  assign new_new_n21967__ = ~new_new_n21604__ & ~new_new_n21966__;
  assign new_new_n21968__ = ~new_new_n21596__ & ~new_new_n21967__;
  assign new_new_n21969__ = ~new_new_n21595__ & ~new_new_n21968__;
  assign new_new_n21970__ = ~new_new_n21587__ & ~new_new_n21969__;
  assign new_new_n21971__ = ~new_new_n21586__ & ~new_new_n21970__;
  assign new_new_n21972__ = ~new_new_n21578__ & new_new_n21971__;
  assign new_new_n21973__ = ~new_new_n21577__ & ~new_new_n21972__;
  assign new_new_n21974__ = ~new_new_n21569__ & ~new_new_n21973__;
  assign new_new_n21975__ = ~new_new_n21568__ & ~new_new_n21974__;
  assign new_new_n21976__ = ~new_new_n21560__ & ~new_new_n21975__;
  assign new_new_n21977__ = ~new_new_n21559__ & ~new_new_n21976__;
  assign new_new_n21978__ = ~new_new_n21551__ & ~new_new_n21977__;
  assign new_new_n21979__ = ~new_new_n21550__ & ~new_new_n21978__;
  assign new_new_n21980__ = ~new_new_n21542__ & ~new_new_n21979__;
  assign new_new_n21981__ = ~new_new_n21541__ & ~new_new_n21980__;
  assign new_new_n21982__ = ~new_new_n21533__ & ~new_new_n21981__;
  assign new_new_n21983__ = ~new_new_n21532__ & ~new_new_n21982__;
  assign new_new_n21984__ = ~new_new_n21524__ & ~new_new_n21983__;
  assign new_new_n21985__ = ~new_new_n21523__ & ~new_new_n21984__;
  assign new_new_n21986__ = ~new_new_n21515__ & ~new_new_n21985__;
  assign new_new_n21987__ = ~new_new_n21514__ & ~new_new_n21986__;
  assign new_new_n21988__ = ~new_new_n21506__ & ~new_new_n21987__;
  assign new_new_n21989__ = ~new_new_n21505__ & ~new_new_n21988__;
  assign new_new_n21990__ = ~new_new_n21497__ & ~new_new_n21989__;
  assign new_new_n21991__ = ~new_new_n21496__ & ~new_new_n21990__;
  assign new_new_n21992__ = ~new_new_n21488__ & new_new_n21991__;
  assign new_new_n21993__ = ~new_new_n21487__ & ~new_new_n21992__;
  assign new_new_n21994__ = ~new_new_n21479__ & ~new_new_n21993__;
  assign new_new_n21995__ = ~new_new_n21478__ & ~new_new_n21994__;
  assign new_new_n21996__ = ~new_new_n21470__ & ~new_new_n21995__;
  assign new_new_n21997__ = ~new_new_n21469__ & ~new_new_n21996__;
  assign new_new_n21998__ = ~new_new_n21461__ & new_new_n21997__;
  assign new_new_n21999__ = ~new_new_n21460__ & ~new_new_n21998__;
  assign new_new_n22000__ = ~new_new_n21452__ & ~new_new_n21999__;
  assign new_new_n22001__ = ~new_new_n21451__ & ~new_new_n22000__;
  assign new_new_n22002__ = ~new_new_n21443__ & ~new_new_n22001__;
  assign new_new_n22003__ = ~new_new_n21442__ & ~new_new_n22002__;
  assign new_new_n22004__ = ~new_new_n21434__ & ~new_new_n22003__;
  assign new_new_n22005__ = ~new_new_n21433__ & ~new_new_n22004__;
  assign new_new_n22006__ = ~new_new_n21425__ & ~new_new_n22005__;
  assign new_new_n22007__ = ~new_new_n21424__ & ~new_new_n22006__;
  assign new_new_n22008__ = ~new_new_n21416__ & new_new_n22007__;
  assign new_new_n22009__ = ~new_new_n21415__ & ~new_new_n22008__;
  assign new_new_n22010__ = ~new_new_n21407__ & ~new_new_n22009__;
  assign new_new_n22011__ = ~new_new_n21406__ & ~new_new_n22010__;
  assign new_new_n22012__ = ~new_new_n21398__ & ~new_new_n22011__;
  assign new_new_n22013__ = ~new_new_n21397__ & ~new_new_n22012__;
  assign new_new_n22014__ = ~new_new_n21389__ & ~new_new_n22013__;
  assign new_new_n22015__ = ~new_new_n21388__ & ~new_new_n22014__;
  assign new_new_n22016__ = ~new_new_n21380__ & ~new_new_n22015__;
  assign new_new_n22017__ = ~new_new_n21379__ & ~new_new_n22016__;
  assign new_new_n22018__ = ~new_new_n21371__ & new_new_n22017__;
  assign new_new_n22019__ = ~new_new_n21370__ & ~new_new_n22018__;
  assign new_new_n22020__ = ~new_new_n21362__ & ~new_new_n22019__;
  assign new_new_n22021__ = ~new_new_n21361__ & ~new_new_n22020__;
  assign new_new_n22022__ = pi125 & ~new_new_n18717__;
  assign new_new_n22023__ = pi124 & ~new_new_n21336__;
  assign new_new_n22024__ = ~pi123 & ~new_new_n20675__;
  assign new_new_n22025__ = pi123 & new_new_n20675__;
  assign new_new_n22026__ = ~new_new_n22024__ & ~new_new_n22025__;
  assign new_new_n22027__ = new_new_n21337__ & new_new_n22026__;
  assign new_new_n22028__ = new_new_n21339__ & ~new_new_n22023__;
  assign new_new_n22029__ = ~new_new_n22027__ & new_new_n22028__;
  assign new_new_n22030__ = new_new_n20018__ & ~new_new_n22029__;
  assign new_new_n22031__ = ~pi125 & new_new_n22030__;
  assign new_new_n22032__ = ~new_new_n21352__ & ~new_new_n22021__;
  assign new_new_n22033__ = ~new_new_n21351__ & ~new_new_n22032__;
  assign new_new_n22034__ = ~new_new_n22031__ & new_new_n22033__;
  assign new_new_n22035__ = ~new_new_n22022__ & ~new_new_n22034__;
  assign po002 = new_new_n260__ & new_new_n22035__;
  assign new_new_n22037__ = ~new_new_n22021__ & po002;
  assign new_new_n22038__ = ~pi124 & ~po002;
  assign new_new_n22039__ = ~new_new_n22037__ & ~new_new_n22038__;
  assign new_new_n22040__ = new_new_n21353__ & ~new_new_n22039__;
  assign new_new_n22041__ = ~new_new_n21353__ & new_new_n22039__;
  assign new_new_n22042__ = ~new_new_n22040__ & ~new_new_n22041__;
  assign new_new_n22043__ = ~pi123 & ~new_new_n22019__;
  assign new_new_n22044__ = pi123 & new_new_n22019__;
  assign new_new_n22045__ = ~new_new_n22043__ & ~new_new_n22044__;
  assign new_new_n22046__ = po002 & new_new_n22045__;
  assign new_new_n22047__ = new_new_n21360__ & new_new_n22046__;
  assign new_new_n22048__ = ~new_new_n21360__ & ~new_new_n22046__;
  assign new_new_n22049__ = ~new_new_n22047__ & ~new_new_n22048__;
  assign new_new_n22050__ = ~pi124 & ~new_new_n22049__;
  assign new_new_n22051__ = pi124 & new_new_n22049__;
  assign new_new_n22052__ = ~new_new_n22017__ & po002;
  assign new_new_n22053__ = pi122 & ~po002;
  assign new_new_n22054__ = ~new_new_n22052__ & ~new_new_n22053__;
  assign new_new_n22055__ = ~new_new_n21370__ & ~new_new_n21371__;
  assign new_new_n22056__ = ~new_new_n22054__ & new_new_n22055__;
  assign new_new_n22057__ = new_new_n22054__ & ~new_new_n22055__;
  assign new_new_n22058__ = ~new_new_n22056__ & ~new_new_n22057__;
  assign new_new_n22059__ = ~pi123 & ~new_new_n22058__;
  assign new_new_n22060__ = pi123 & new_new_n22058__;
  assign new_new_n22061__ = ~new_new_n21379__ & ~new_new_n21380__;
  assign new_new_n22062__ = ~new_new_n22015__ & po002;
  assign new_new_n22063__ = pi121 & ~po002;
  assign new_new_n22064__ = ~new_new_n22062__ & ~new_new_n22063__;
  assign new_new_n22065__ = new_new_n22061__ & ~new_new_n22064__;
  assign new_new_n22066__ = ~new_new_n22061__ & new_new_n22064__;
  assign new_new_n22067__ = ~new_new_n22065__ & ~new_new_n22066__;
  assign new_new_n22068__ = pi122 & new_new_n22067__;
  assign new_new_n22069__ = ~pi122 & ~new_new_n22067__;
  assign new_new_n22070__ = ~new_new_n21388__ & ~new_new_n21389__;
  assign new_new_n22071__ = ~new_new_n22013__ & po002;
  assign new_new_n22072__ = pi120 & ~po002;
  assign new_new_n22073__ = ~new_new_n22071__ & ~new_new_n22072__;
  assign new_new_n22074__ = new_new_n22070__ & new_new_n22073__;
  assign new_new_n22075__ = ~new_new_n22070__ & ~new_new_n22073__;
  assign new_new_n22076__ = ~new_new_n22074__ & ~new_new_n22075__;
  assign new_new_n22077__ = pi121 & ~new_new_n22076__;
  assign new_new_n22078__ = ~pi121 & new_new_n22076__;
  assign new_new_n22079__ = pi119 & ~new_new_n22011__;
  assign new_new_n22080__ = ~pi119 & new_new_n22011__;
  assign new_new_n22081__ = ~new_new_n22079__ & ~new_new_n22080__;
  assign new_new_n22082__ = po002 & new_new_n22081__;
  assign new_new_n22083__ = ~new_new_n21396__ & ~new_new_n22082__;
  assign new_new_n22084__ = new_new_n21396__ & new_new_n22082__;
  assign new_new_n22085__ = ~new_new_n22083__ & ~new_new_n22084__;
  assign new_new_n22086__ = pi120 & ~new_new_n22085__;
  assign new_new_n22087__ = ~pi120 & new_new_n22085__;
  assign new_new_n22088__ = pi118 & ~new_new_n22009__;
  assign new_new_n22089__ = ~pi118 & new_new_n22009__;
  assign new_new_n22090__ = ~new_new_n22088__ & ~new_new_n22089__;
  assign new_new_n22091__ = po002 & new_new_n22090__;
  assign new_new_n22092__ = new_new_n21405__ & new_new_n22091__;
  assign new_new_n22093__ = ~new_new_n21405__ & ~new_new_n22091__;
  assign new_new_n22094__ = ~new_new_n22092__ & ~new_new_n22093__;
  assign new_new_n22095__ = pi119 & ~new_new_n22094__;
  assign new_new_n22096__ = ~pi119 & new_new_n22094__;
  assign new_new_n22097__ = ~new_new_n21415__ & ~new_new_n21416__;
  assign new_new_n22098__ = ~new_new_n22007__ & po002;
  assign new_new_n22099__ = ~pi117 & ~po002;
  assign new_new_n22100__ = ~new_new_n22098__ & ~new_new_n22099__;
  assign new_new_n22101__ = new_new_n22097__ & new_new_n22100__;
  assign new_new_n22102__ = ~new_new_n22097__ & ~new_new_n22100__;
  assign new_new_n22103__ = ~new_new_n22101__ & ~new_new_n22102__;
  assign new_new_n22104__ = ~pi118 & ~new_new_n22103__;
  assign new_new_n22105__ = pi118 & new_new_n22103__;
  assign new_new_n22106__ = ~pi116 & ~new_new_n22005__;
  assign new_new_n22107__ = pi116 & new_new_n22005__;
  assign new_new_n22108__ = ~new_new_n22106__ & ~new_new_n22107__;
  assign new_new_n22109__ = po002 & new_new_n22108__;
  assign new_new_n22110__ = new_new_n21423__ & new_new_n22109__;
  assign new_new_n22111__ = ~new_new_n21423__ & ~new_new_n22109__;
  assign new_new_n22112__ = ~new_new_n22110__ & ~new_new_n22111__;
  assign new_new_n22113__ = pi117 & new_new_n22112__;
  assign new_new_n22114__ = ~pi117 & ~new_new_n22112__;
  assign new_new_n22115__ = ~new_new_n21433__ & ~new_new_n21434__;
  assign new_new_n22116__ = ~new_new_n22003__ & po002;
  assign new_new_n22117__ = ~pi115 & ~po002;
  assign new_new_n22118__ = ~new_new_n22116__ & ~new_new_n22117__;
  assign new_new_n22119__ = new_new_n22115__ & ~new_new_n22118__;
  assign new_new_n22120__ = ~new_new_n22115__ & new_new_n22118__;
  assign new_new_n22121__ = ~new_new_n22119__ & ~new_new_n22120__;
  assign new_new_n22122__ = pi116 & ~new_new_n22121__;
  assign new_new_n22123__ = ~pi116 & new_new_n22121__;
  assign new_new_n22124__ = ~new_new_n21442__ & ~new_new_n21443__;
  assign new_new_n22125__ = ~new_new_n22001__ & po002;
  assign new_new_n22126__ = ~pi114 & ~po002;
  assign new_new_n22127__ = ~new_new_n22125__ & ~new_new_n22126__;
  assign new_new_n22128__ = new_new_n22124__ & ~new_new_n22127__;
  assign new_new_n22129__ = ~new_new_n22124__ & new_new_n22127__;
  assign new_new_n22130__ = ~new_new_n22128__ & ~new_new_n22129__;
  assign new_new_n22131__ = pi115 & ~new_new_n22130__;
  assign new_new_n22132__ = ~pi115 & new_new_n22130__;
  assign new_new_n22133__ = ~new_new_n21451__ & ~new_new_n21452__;
  assign new_new_n22134__ = ~new_new_n21999__ & po002;
  assign new_new_n22135__ = ~pi113 & ~po002;
  assign new_new_n22136__ = ~new_new_n22134__ & ~new_new_n22135__;
  assign new_new_n22137__ = new_new_n22133__ & ~new_new_n22136__;
  assign new_new_n22138__ = ~new_new_n22133__ & new_new_n22136__;
  assign new_new_n22139__ = ~new_new_n22137__ & ~new_new_n22138__;
  assign new_new_n22140__ = pi114 & ~new_new_n22139__;
  assign new_new_n22141__ = ~pi114 & new_new_n22139__;
  assign new_new_n22142__ = ~new_new_n21460__ & ~new_new_n21461__;
  assign new_new_n22143__ = ~new_new_n21997__ & po002;
  assign new_new_n22144__ = pi112 & ~po002;
  assign new_new_n22145__ = ~new_new_n22143__ & ~new_new_n22144__;
  assign new_new_n22146__ = new_new_n22142__ & ~new_new_n22145__;
  assign new_new_n22147__ = ~new_new_n22142__ & new_new_n22145__;
  assign new_new_n22148__ = ~new_new_n22146__ & ~new_new_n22147__;
  assign new_new_n22149__ = ~pi113 & ~new_new_n22148__;
  assign new_new_n22150__ = pi113 & new_new_n22148__;
  assign new_new_n22151__ = ~new_new_n21469__ & ~new_new_n21470__;
  assign new_new_n22152__ = ~new_new_n21995__ & po002;
  assign new_new_n22153__ = pi111 & ~po002;
  assign new_new_n22154__ = ~new_new_n22152__ & ~new_new_n22153__;
  assign new_new_n22155__ = new_new_n22151__ & ~new_new_n22154__;
  assign new_new_n22156__ = ~new_new_n22151__ & new_new_n22154__;
  assign new_new_n22157__ = ~new_new_n22155__ & ~new_new_n22156__;
  assign new_new_n22158__ = ~pi112 & ~new_new_n22157__;
  assign new_new_n22159__ = pi112 & new_new_n22157__;
  assign new_new_n22160__ = pi110 & ~new_new_n21993__;
  assign new_new_n22161__ = ~pi110 & new_new_n21993__;
  assign new_new_n22162__ = ~new_new_n22160__ & ~new_new_n22161__;
  assign new_new_n22163__ = po002 & new_new_n22162__;
  assign new_new_n22164__ = new_new_n21477__ & new_new_n22163__;
  assign new_new_n22165__ = ~new_new_n21477__ & ~new_new_n22163__;
  assign new_new_n22166__ = ~new_new_n22164__ & ~new_new_n22165__;
  assign new_new_n22167__ = pi111 & ~new_new_n22166__;
  assign new_new_n22168__ = ~pi111 & new_new_n22166__;
  assign new_new_n22169__ = ~new_new_n21487__ & ~new_new_n21488__;
  assign new_new_n22170__ = ~new_new_n21991__ & po002;
  assign new_new_n22171__ = ~pi109 & ~po002;
  assign new_new_n22172__ = ~new_new_n22170__ & ~new_new_n22171__;
  assign new_new_n22173__ = new_new_n22169__ & ~new_new_n22172__;
  assign new_new_n22174__ = ~new_new_n22169__ & new_new_n22172__;
  assign new_new_n22175__ = ~new_new_n22173__ & ~new_new_n22174__;
  assign new_new_n22176__ = pi110 & ~new_new_n22175__;
  assign new_new_n22177__ = ~pi110 & new_new_n22175__;
  assign new_new_n22178__ = ~pi108 & ~new_new_n21989__;
  assign new_new_n22179__ = pi108 & new_new_n21989__;
  assign new_new_n22180__ = ~new_new_n22178__ & ~new_new_n22179__;
  assign new_new_n22181__ = po002 & new_new_n22180__;
  assign new_new_n22182__ = new_new_n21495__ & new_new_n22181__;
  assign new_new_n22183__ = ~new_new_n21495__ & ~new_new_n22181__;
  assign new_new_n22184__ = ~new_new_n22182__ & ~new_new_n22183__;
  assign new_new_n22185__ = ~pi109 & ~new_new_n22184__;
  assign new_new_n22186__ = pi109 & new_new_n22184__;
  assign new_new_n22187__ = ~new_new_n21505__ & ~new_new_n21506__;
  assign new_new_n22188__ = ~new_new_n21987__ & po002;
  assign new_new_n22189__ = ~pi107 & ~po002;
  assign new_new_n22190__ = ~new_new_n22188__ & ~new_new_n22189__;
  assign new_new_n22191__ = ~new_new_n22187__ & ~new_new_n22190__;
  assign new_new_n22192__ = new_new_n22187__ & new_new_n22190__;
  assign new_new_n22193__ = ~new_new_n22191__ & ~new_new_n22192__;
  assign new_new_n22194__ = pi108 & new_new_n22193__;
  assign new_new_n22195__ = ~pi108 & ~new_new_n22193__;
  assign new_new_n22196__ = ~new_new_n21514__ & ~new_new_n21515__;
  assign new_new_n22197__ = ~new_new_n21985__ & po002;
  assign new_new_n22198__ = ~pi106 & ~po002;
  assign new_new_n22199__ = ~new_new_n22197__ & ~new_new_n22198__;
  assign new_new_n22200__ = new_new_n22196__ & ~new_new_n22199__;
  assign new_new_n22201__ = ~new_new_n22196__ & new_new_n22199__;
  assign new_new_n22202__ = ~new_new_n22200__ & ~new_new_n22201__;
  assign new_new_n22203__ = pi107 & ~new_new_n22202__;
  assign new_new_n22204__ = ~pi107 & new_new_n22202__;
  assign new_new_n22205__ = ~pi105 & ~new_new_n21983__;
  assign new_new_n22206__ = pi105 & new_new_n21983__;
  assign new_new_n22207__ = ~new_new_n22205__ & ~new_new_n22206__;
  assign new_new_n22208__ = po002 & new_new_n22207__;
  assign new_new_n22209__ = new_new_n21522__ & new_new_n22208__;
  assign new_new_n22210__ = ~new_new_n21522__ & ~new_new_n22208__;
  assign new_new_n22211__ = ~new_new_n22209__ & ~new_new_n22210__;
  assign new_new_n22212__ = ~pi106 & ~new_new_n22211__;
  assign new_new_n22213__ = pi106 & new_new_n22211__;
  assign new_new_n22214__ = ~new_new_n21532__ & ~new_new_n21533__;
  assign new_new_n22215__ = ~new_new_n21981__ & po002;
  assign new_new_n22216__ = ~pi104 & ~po002;
  assign new_new_n22217__ = ~new_new_n22215__ & ~new_new_n22216__;
  assign new_new_n22218__ = new_new_n22214__ & ~new_new_n22217__;
  assign new_new_n22219__ = ~new_new_n22214__ & new_new_n22217__;
  assign new_new_n22220__ = ~new_new_n22218__ & ~new_new_n22219__;
  assign new_new_n22221__ = pi105 & ~new_new_n22220__;
  assign new_new_n22222__ = ~pi105 & new_new_n22220__;
  assign new_new_n22223__ = ~new_new_n21541__ & ~new_new_n21542__;
  assign new_new_n22224__ = ~new_new_n21979__ & po002;
  assign new_new_n22225__ = ~pi103 & ~po002;
  assign new_new_n22226__ = ~new_new_n22224__ & ~new_new_n22225__;
  assign new_new_n22227__ = new_new_n22223__ & ~new_new_n22226__;
  assign new_new_n22228__ = ~new_new_n22223__ & new_new_n22226__;
  assign new_new_n22229__ = ~new_new_n22227__ & ~new_new_n22228__;
  assign new_new_n22230__ = ~pi104 & new_new_n22229__;
  assign new_new_n22231__ = pi104 & ~new_new_n22229__;
  assign new_new_n22232__ = ~new_new_n21550__ & ~new_new_n21551__;
  assign new_new_n22233__ = ~new_new_n21977__ & po002;
  assign new_new_n22234__ = ~pi102 & ~po002;
  assign new_new_n22235__ = ~new_new_n22233__ & ~new_new_n22234__;
  assign new_new_n22236__ = new_new_n22232__ & ~new_new_n22235__;
  assign new_new_n22237__ = ~new_new_n22232__ & new_new_n22235__;
  assign new_new_n22238__ = ~new_new_n22236__ & ~new_new_n22237__;
  assign new_new_n22239__ = ~pi103 & new_new_n22238__;
  assign new_new_n22240__ = pi103 & ~new_new_n22238__;
  assign new_new_n22241__ = ~new_new_n21559__ & ~new_new_n21560__;
  assign new_new_n22242__ = ~new_new_n21975__ & po002;
  assign new_new_n22243__ = ~pi101 & ~po002;
  assign new_new_n22244__ = ~new_new_n22242__ & ~new_new_n22243__;
  assign new_new_n22245__ = new_new_n22241__ & ~new_new_n22244__;
  assign new_new_n22246__ = ~new_new_n22241__ & new_new_n22244__;
  assign new_new_n22247__ = ~new_new_n22245__ & ~new_new_n22246__;
  assign new_new_n22248__ = ~pi102 & new_new_n22247__;
  assign new_new_n22249__ = pi102 & ~new_new_n22247__;
  assign new_new_n22250__ = ~pi100 & ~new_new_n21973__;
  assign new_new_n22251__ = pi100 & new_new_n21973__;
  assign new_new_n22252__ = ~new_new_n22250__ & ~new_new_n22251__;
  assign new_new_n22253__ = po002 & new_new_n22252__;
  assign new_new_n22254__ = new_new_n21567__ & new_new_n22253__;
  assign new_new_n22255__ = ~new_new_n21567__ & ~new_new_n22253__;
  assign new_new_n22256__ = ~new_new_n22254__ & ~new_new_n22255__;
  assign new_new_n22257__ = ~pi101 & ~new_new_n22256__;
  assign new_new_n22258__ = pi101 & new_new_n22256__;
  assign new_new_n22259__ = ~new_new_n21577__ & ~new_new_n21578__;
  assign new_new_n22260__ = new_new_n21971__ & po002;
  assign new_new_n22261__ = ~pi099 & ~po002;
  assign new_new_n22262__ = ~new_new_n22260__ & ~new_new_n22261__;
  assign new_new_n22263__ = ~new_new_n22259__ & ~new_new_n22262__;
  assign new_new_n22264__ = new_new_n22259__ & new_new_n22262__;
  assign new_new_n22265__ = ~new_new_n22263__ & ~new_new_n22264__;
  assign new_new_n22266__ = ~pi100 & ~new_new_n22265__;
  assign new_new_n22267__ = pi100 & new_new_n22265__;
  assign new_new_n22268__ = ~new_new_n21969__ & po002;
  assign new_new_n22269__ = pi098 & ~po002;
  assign new_new_n22270__ = ~new_new_n22268__ & ~new_new_n22269__;
  assign new_new_n22271__ = ~new_new_n21586__ & ~new_new_n21587__;
  assign new_new_n22272__ = new_new_n22270__ & new_new_n22271__;
  assign new_new_n22273__ = ~new_new_n22270__ & ~new_new_n22271__;
  assign new_new_n22274__ = ~new_new_n22272__ & ~new_new_n22273__;
  assign new_new_n22275__ = pi099 & ~new_new_n22274__;
  assign new_new_n22276__ = ~pi099 & new_new_n22274__;
  assign new_new_n22277__ = ~new_new_n21595__ & ~new_new_n21596__;
  assign new_new_n22278__ = ~new_new_n21967__ & po002;
  assign new_new_n22279__ = pi097 & ~po002;
  assign new_new_n22280__ = ~new_new_n22278__ & ~new_new_n22279__;
  assign new_new_n22281__ = new_new_n22277__ & new_new_n22280__;
  assign new_new_n22282__ = ~new_new_n22277__ & ~new_new_n22280__;
  assign new_new_n22283__ = ~new_new_n22281__ & ~new_new_n22282__;
  assign new_new_n22284__ = pi098 & ~new_new_n22283__;
  assign new_new_n22285__ = ~pi098 & new_new_n22283__;
  assign new_new_n22286__ = ~new_new_n21965__ & po002;
  assign new_new_n22287__ = pi096 & ~po002;
  assign new_new_n22288__ = ~new_new_n22286__ & ~new_new_n22287__;
  assign new_new_n22289__ = ~new_new_n21604__ & ~new_new_n21605__;
  assign new_new_n22290__ = ~new_new_n22288__ & new_new_n22289__;
  assign new_new_n22291__ = new_new_n22288__ & ~new_new_n22289__;
  assign new_new_n22292__ = ~new_new_n22290__ & ~new_new_n22291__;
  assign new_new_n22293__ = ~pi097 & ~new_new_n22292__;
  assign new_new_n22294__ = pi097 & new_new_n22292__;
  assign new_new_n22295__ = ~new_new_n21613__ & ~new_new_n21614__;
  assign new_new_n22296__ = ~new_new_n21963__ & po002;
  assign new_new_n22297__ = pi095 & ~po002;
  assign new_new_n22298__ = ~new_new_n22296__ & ~new_new_n22297__;
  assign new_new_n22299__ = new_new_n22295__ & ~new_new_n22298__;
  assign new_new_n22300__ = ~new_new_n22295__ & new_new_n22298__;
  assign new_new_n22301__ = ~new_new_n22299__ & ~new_new_n22300__;
  assign new_new_n22302__ = ~pi096 & ~new_new_n22301__;
  assign new_new_n22303__ = pi096 & new_new_n22301__;
  assign new_new_n22304__ = ~new_new_n21622__ & ~new_new_n21623__;
  assign new_new_n22305__ = ~new_new_n21961__ & po002;
  assign new_new_n22306__ = ~pi094 & ~po002;
  assign new_new_n22307__ = ~new_new_n22305__ & ~new_new_n22306__;
  assign new_new_n22308__ = new_new_n22304__ & ~new_new_n22307__;
  assign new_new_n22309__ = ~new_new_n22304__ & new_new_n22307__;
  assign new_new_n22310__ = ~new_new_n22308__ & ~new_new_n22309__;
  assign new_new_n22311__ = ~pi095 & new_new_n22310__;
  assign new_new_n22312__ = pi095 & ~new_new_n22310__;
  assign new_new_n22313__ = ~pi093 & ~new_new_n21959__;
  assign new_new_n22314__ = pi093 & new_new_n21959__;
  assign new_new_n22315__ = ~new_new_n22313__ & ~new_new_n22314__;
  assign new_new_n22316__ = po002 & new_new_n22315__;
  assign new_new_n22317__ = new_new_n21630__ & new_new_n22316__;
  assign new_new_n22318__ = ~new_new_n21630__ & ~new_new_n22316__;
  assign new_new_n22319__ = ~new_new_n22317__ & ~new_new_n22318__;
  assign new_new_n22320__ = ~pi094 & ~new_new_n22319__;
  assign new_new_n22321__ = pi094 & new_new_n22319__;
  assign new_new_n22322__ = ~new_new_n21640__ & ~new_new_n21641__;
  assign new_new_n22323__ = ~new_new_n21957__ & po002;
  assign new_new_n22324__ = pi092 & ~po002;
  assign new_new_n22325__ = ~new_new_n22323__ & ~new_new_n22324__;
  assign new_new_n22326__ = new_new_n22322__ & ~new_new_n22325__;
  assign new_new_n22327__ = ~new_new_n22322__ & new_new_n22325__;
  assign new_new_n22328__ = ~new_new_n22326__ & ~new_new_n22327__;
  assign new_new_n22329__ = ~pi093 & ~new_new_n22328__;
  assign new_new_n22330__ = pi093 & new_new_n22328__;
  assign new_new_n22331__ = ~new_new_n21649__ & ~new_new_n21650__;
  assign new_new_n22332__ = ~new_new_n21955__ & po002;
  assign new_new_n22333__ = pi091 & ~po002;
  assign new_new_n22334__ = ~new_new_n22332__ & ~new_new_n22333__;
  assign new_new_n22335__ = new_new_n22331__ & ~new_new_n22334__;
  assign new_new_n22336__ = ~new_new_n22331__ & new_new_n22334__;
  assign new_new_n22337__ = ~new_new_n22335__ & ~new_new_n22336__;
  assign new_new_n22338__ = ~pi092 & ~new_new_n22337__;
  assign new_new_n22339__ = pi092 & new_new_n22337__;
  assign new_new_n22340__ = ~new_new_n21658__ & ~new_new_n21659__;
  assign new_new_n22341__ = ~new_new_n21953__ & po002;
  assign new_new_n22342__ = pi090 & ~po002;
  assign new_new_n22343__ = ~new_new_n22341__ & ~new_new_n22342__;
  assign new_new_n22344__ = new_new_n22340__ & new_new_n22343__;
  assign new_new_n22345__ = ~new_new_n22340__ & ~new_new_n22343__;
  assign new_new_n22346__ = ~new_new_n22344__ & ~new_new_n22345__;
  assign new_new_n22347__ = pi091 & ~new_new_n22346__;
  assign new_new_n22348__ = ~pi091 & new_new_n22346__;
  assign new_new_n22349__ = new_new_n21951__ & po002;
  assign new_new_n22350__ = pi089 & ~po002;
  assign new_new_n22351__ = ~new_new_n22349__ & ~new_new_n22350__;
  assign new_new_n22352__ = ~new_new_n21667__ & ~new_new_n21668__;
  assign new_new_n22353__ = ~new_new_n22351__ & ~new_new_n22352__;
  assign new_new_n22354__ = new_new_n22351__ & new_new_n22352__;
  assign new_new_n22355__ = ~new_new_n22353__ & ~new_new_n22354__;
  assign new_new_n22356__ = pi090 & ~new_new_n22355__;
  assign new_new_n22357__ = ~pi090 & new_new_n22355__;
  assign new_new_n22358__ = ~new_new_n21676__ & ~new_new_n21677__;
  assign new_new_n22359__ = ~new_new_n21949__ & po002;
  assign new_new_n22360__ = ~pi088 & ~po002;
  assign new_new_n22361__ = ~new_new_n22359__ & ~new_new_n22360__;
  assign new_new_n22362__ = new_new_n22358__ & ~new_new_n22361__;
  assign new_new_n22363__ = ~new_new_n22358__ & new_new_n22361__;
  assign new_new_n22364__ = ~new_new_n22362__ & ~new_new_n22363__;
  assign new_new_n22365__ = pi089 & ~new_new_n22364__;
  assign new_new_n22366__ = ~pi089 & new_new_n22364__;
  assign new_new_n22367__ = ~pi087 & ~new_new_n21947__;
  assign new_new_n22368__ = pi087 & new_new_n21947__;
  assign new_new_n22369__ = ~new_new_n22367__ & ~new_new_n22368__;
  assign new_new_n22370__ = po002 & new_new_n22369__;
  assign new_new_n22371__ = new_new_n21684__ & new_new_n22370__;
  assign new_new_n22372__ = ~new_new_n21684__ & ~new_new_n22370__;
  assign new_new_n22373__ = ~new_new_n22371__ & ~new_new_n22372__;
  assign new_new_n22374__ = pi088 & new_new_n22373__;
  assign new_new_n22375__ = ~pi088 & ~new_new_n22373__;
  assign new_new_n22376__ = ~new_new_n21945__ & po002;
  assign new_new_n22377__ = pi086 & ~po002;
  assign new_new_n22378__ = ~new_new_n22376__ & ~new_new_n22377__;
  assign new_new_n22379__ = ~new_new_n21694__ & ~new_new_n21695__;
  assign new_new_n22380__ = ~new_new_n22378__ & new_new_n22379__;
  assign new_new_n22381__ = new_new_n22378__ & ~new_new_n22379__;
  assign new_new_n22382__ = ~new_new_n22380__ & ~new_new_n22381__;
  assign new_new_n22383__ = pi087 & new_new_n22382__;
  assign new_new_n22384__ = ~pi087 & ~new_new_n22382__;
  assign new_new_n22385__ = pi085 & ~new_new_n21943__;
  assign new_new_n22386__ = ~pi085 & new_new_n21943__;
  assign new_new_n22387__ = ~new_new_n22385__ & ~new_new_n22386__;
  assign new_new_n22388__ = po002 & new_new_n22387__;
  assign new_new_n22389__ = new_new_n21702__ & new_new_n22388__;
  assign new_new_n22390__ = ~new_new_n21702__ & ~new_new_n22388__;
  assign new_new_n22391__ = ~new_new_n22389__ & ~new_new_n22390__;
  assign new_new_n22392__ = pi086 & ~new_new_n22391__;
  assign new_new_n22393__ = ~pi086 & new_new_n22391__;
  assign new_new_n22394__ = ~new_new_n21712__ & ~new_new_n21713__;
  assign new_new_n22395__ = ~new_new_n21941__ & po002;
  assign new_new_n22396__ = pi084 & ~po002;
  assign new_new_n22397__ = ~new_new_n22395__ & ~new_new_n22396__;
  assign new_new_n22398__ = new_new_n22394__ & new_new_n22397__;
  assign new_new_n22399__ = ~new_new_n22394__ & ~new_new_n22397__;
  assign new_new_n22400__ = ~new_new_n22398__ & ~new_new_n22399__;
  assign new_new_n22401__ = pi085 & ~new_new_n22400__;
  assign new_new_n22402__ = ~pi085 & new_new_n22400__;
  assign new_new_n22403__ = ~new_new_n21721__ & ~new_new_n21722__;
  assign new_new_n22404__ = ~new_new_n21939__ & po002;
  assign new_new_n22405__ = pi083 & ~po002;
  assign new_new_n22406__ = ~new_new_n22404__ & ~new_new_n22405__;
  assign new_new_n22407__ = new_new_n22403__ & ~new_new_n22406__;
  assign new_new_n22408__ = ~new_new_n22403__ & new_new_n22406__;
  assign new_new_n22409__ = ~new_new_n22407__ & ~new_new_n22408__;
  assign new_new_n22410__ = ~pi084 & ~new_new_n22409__;
  assign new_new_n22411__ = pi084 & new_new_n22409__;
  assign new_new_n22412__ = pi082 & ~new_new_n21937__;
  assign new_new_n22413__ = ~pi082 & new_new_n21937__;
  assign new_new_n22414__ = ~new_new_n22412__ & ~new_new_n22413__;
  assign new_new_n22415__ = po002 & new_new_n22414__;
  assign new_new_n22416__ = new_new_n21729__ & new_new_n22415__;
  assign new_new_n22417__ = ~new_new_n21729__ & ~new_new_n22415__;
  assign new_new_n22418__ = ~new_new_n22416__ & ~new_new_n22417__;
  assign new_new_n22419__ = pi083 & ~new_new_n22418__;
  assign new_new_n22420__ = ~pi083 & new_new_n22418__;
  assign new_new_n22421__ = ~new_new_n21739__ & ~new_new_n21740__;
  assign new_new_n22422__ = ~new_new_n21935__ & po002;
  assign new_new_n22423__ = ~pi081 & ~po002;
  assign new_new_n22424__ = ~new_new_n22422__ & ~new_new_n22423__;
  assign new_new_n22425__ = new_new_n22421__ & ~new_new_n22424__;
  assign new_new_n22426__ = ~new_new_n22421__ & new_new_n22424__;
  assign new_new_n22427__ = ~new_new_n22425__ & ~new_new_n22426__;
  assign new_new_n22428__ = pi082 & ~new_new_n22427__;
  assign new_new_n22429__ = ~pi082 & new_new_n22427__;
  assign new_new_n22430__ = ~new_new_n21933__ & po002;
  assign new_new_n22431__ = pi080 & ~po002;
  assign new_new_n22432__ = ~new_new_n22430__ & ~new_new_n22431__;
  assign new_new_n22433__ = ~new_new_n21748__ & ~new_new_n21749__;
  assign new_new_n22434__ = ~new_new_n22432__ & new_new_n22433__;
  assign new_new_n22435__ = new_new_n22432__ & ~new_new_n22433__;
  assign new_new_n22436__ = ~new_new_n22434__ & ~new_new_n22435__;
  assign new_new_n22437__ = ~pi081 & ~new_new_n22436__;
  assign new_new_n22438__ = pi081 & new_new_n22436__;
  assign new_new_n22439__ = ~new_new_n21757__ & ~new_new_n21758__;
  assign new_new_n22440__ = ~new_new_n21931__ & po002;
  assign new_new_n22441__ = pi079 & ~po002;
  assign new_new_n22442__ = ~new_new_n22440__ & ~new_new_n22441__;
  assign new_new_n22443__ = new_new_n22439__ & ~new_new_n22442__;
  assign new_new_n22444__ = ~new_new_n22439__ & new_new_n22442__;
  assign new_new_n22445__ = ~new_new_n22443__ & ~new_new_n22444__;
  assign new_new_n22446__ = ~pi080 & ~new_new_n22445__;
  assign new_new_n22447__ = pi080 & new_new_n22445__;
  assign new_new_n22448__ = ~new_new_n21766__ & ~new_new_n21767__;
  assign new_new_n22449__ = ~new_new_n21929__ & po002;
  assign new_new_n22450__ = pi078 & ~po002;
  assign new_new_n22451__ = ~new_new_n22449__ & ~new_new_n22450__;
  assign new_new_n22452__ = new_new_n22448__ & ~new_new_n22451__;
  assign new_new_n22453__ = ~new_new_n22448__ & new_new_n22451__;
  assign new_new_n22454__ = ~new_new_n22452__ & ~new_new_n22453__;
  assign new_new_n22455__ = ~pi079 & ~new_new_n22454__;
  assign new_new_n22456__ = pi079 & new_new_n22454__;
  assign new_new_n22457__ = ~new_new_n21927__ & po002;
  assign new_new_n22458__ = pi077 & ~po002;
  assign new_new_n22459__ = ~new_new_n22457__ & ~new_new_n22458__;
  assign new_new_n22460__ = ~new_new_n21775__ & ~new_new_n21776__;
  assign new_new_n22461__ = ~new_new_n22459__ & new_new_n22460__;
  assign new_new_n22462__ = new_new_n22459__ & ~new_new_n22460__;
  assign new_new_n22463__ = ~new_new_n22461__ & ~new_new_n22462__;
  assign new_new_n22464__ = ~pi078 & ~new_new_n22463__;
  assign new_new_n22465__ = pi078 & new_new_n22463__;
  assign new_new_n22466__ = ~new_new_n21784__ & ~new_new_n21785__;
  assign new_new_n22467__ = ~new_new_n21925__ & po002;
  assign new_new_n22468__ = pi076 & ~po002;
  assign new_new_n22469__ = ~new_new_n22467__ & ~new_new_n22468__;
  assign new_new_n22470__ = new_new_n22466__ & ~new_new_n22469__;
  assign new_new_n22471__ = ~new_new_n22466__ & new_new_n22469__;
  assign new_new_n22472__ = ~new_new_n22470__ & ~new_new_n22471__;
  assign new_new_n22473__ = ~pi077 & ~new_new_n22472__;
  assign new_new_n22474__ = pi077 & new_new_n22472__;
  assign new_new_n22475__ = ~new_new_n21923__ & po002;
  assign new_new_n22476__ = pi075 & ~po002;
  assign new_new_n22477__ = ~new_new_n22475__ & ~new_new_n22476__;
  assign new_new_n22478__ = ~new_new_n21793__ & ~new_new_n21794__;
  assign new_new_n22479__ = ~new_new_n22477__ & new_new_n22478__;
  assign new_new_n22480__ = new_new_n22477__ & ~new_new_n22478__;
  assign new_new_n22481__ = ~new_new_n22479__ & ~new_new_n22480__;
  assign new_new_n22482__ = ~pi076 & ~new_new_n22481__;
  assign new_new_n22483__ = pi076 & new_new_n22481__;
  assign new_new_n22484__ = pi074 & ~new_new_n21921__;
  assign new_new_n22485__ = ~pi074 & new_new_n21921__;
  assign new_new_n22486__ = ~new_new_n22484__ & ~new_new_n22485__;
  assign new_new_n22487__ = po002 & new_new_n22486__;
  assign new_new_n22488__ = new_new_n21801__ & new_new_n22487__;
  assign new_new_n22489__ = ~new_new_n21801__ & ~new_new_n22487__;
  assign new_new_n22490__ = ~new_new_n22488__ & ~new_new_n22489__;
  assign new_new_n22491__ = pi075 & ~new_new_n22490__;
  assign new_new_n22492__ = ~pi075 & new_new_n22490__;
  assign new_new_n22493__ = pi073 & ~new_new_n21919__;
  assign new_new_n22494__ = ~pi073 & new_new_n21919__;
  assign new_new_n22495__ = ~new_new_n22493__ & ~new_new_n22494__;
  assign new_new_n22496__ = po002 & new_new_n22495__;
  assign new_new_n22497__ = new_new_n21810__ & new_new_n22496__;
  assign new_new_n22498__ = ~new_new_n21810__ & ~new_new_n22496__;
  assign new_new_n22499__ = ~new_new_n22497__ & ~new_new_n22498__;
  assign new_new_n22500__ = ~pi074 & new_new_n22499__;
  assign new_new_n22501__ = pi074 & ~new_new_n22499__;
  assign new_new_n22502__ = ~new_new_n21909__ & ~new_new_n21910__;
  assign new_new_n22503__ = po002 & new_new_n22502__;
  assign new_new_n22504__ = new_new_n21917__ & new_new_n22503__;
  assign new_new_n22505__ = ~new_new_n21917__ & ~new_new_n22503__;
  assign new_new_n22506__ = ~new_new_n22504__ & ~new_new_n22505__;
  assign new_new_n22507__ = ~pi073 & ~new_new_n22506__;
  assign new_new_n22508__ = pi073 & new_new_n22506__;
  assign new_new_n22509__ = ~new_new_n21906__ & po002;
  assign new_new_n22510__ = pi071 & ~po002;
  assign new_new_n22511__ = ~new_new_n22509__ & ~new_new_n22510__;
  assign new_new_n22512__ = ~new_new_n21820__ & ~new_new_n21821__;
  assign new_new_n22513__ = ~new_new_n22511__ & new_new_n22512__;
  assign new_new_n22514__ = new_new_n22511__ & ~new_new_n22512__;
  assign new_new_n22515__ = ~new_new_n22513__ & ~new_new_n22514__;
  assign new_new_n22516__ = ~pi072 & ~new_new_n22515__;
  assign new_new_n22517__ = pi072 & new_new_n22515__;
  assign new_new_n22518__ = ~new_new_n21829__ & ~new_new_n21830__;
  assign new_new_n22519__ = new_new_n21904__ & po002;
  assign new_new_n22520__ = ~pi070 & ~po002;
  assign new_new_n22521__ = ~new_new_n22519__ & ~new_new_n22520__;
  assign new_new_n22522__ = ~new_new_n22518__ & ~new_new_n22521__;
  assign new_new_n22523__ = new_new_n22518__ & new_new_n22521__;
  assign new_new_n22524__ = ~new_new_n22522__ & ~new_new_n22523__;
  assign new_new_n22525__ = ~pi071 & ~new_new_n22524__;
  assign new_new_n22526__ = pi071 & new_new_n22524__;
  assign new_new_n22527__ = ~new_new_n21838__ & ~new_new_n21839__;
  assign new_new_n22528__ = ~new_new_n21902__ & po002;
  assign new_new_n22529__ = pi069 & ~po002;
  assign new_new_n22530__ = ~new_new_n22528__ & ~new_new_n22529__;
  assign new_new_n22531__ = new_new_n22527__ & new_new_n22530__;
  assign new_new_n22532__ = ~new_new_n22527__ & ~new_new_n22530__;
  assign new_new_n22533__ = ~new_new_n22531__ & ~new_new_n22532__;
  assign new_new_n22534__ = pi070 & ~new_new_n22533__;
  assign new_new_n22535__ = ~pi070 & new_new_n22533__;
  assign new_new_n22536__ = ~new_new_n21892__ & ~new_new_n21893__;
  assign new_new_n22537__ = po002 & new_new_n22536__;
  assign new_new_n22538__ = new_new_n21900__ & new_new_n22537__;
  assign new_new_n22539__ = ~new_new_n21900__ & ~new_new_n22537__;
  assign new_new_n22540__ = ~new_new_n22538__ & ~new_new_n22539__;
  assign new_new_n22541__ = pi069 & ~new_new_n22540__;
  assign new_new_n22542__ = ~pi069 & new_new_n22540__;
  assign new_new_n22543__ = ~new_new_n21845__ & ~new_new_n21846__;
  assign new_new_n22544__ = ~new_new_n21889__ & po002;
  assign new_new_n22545__ = ~pi067 & ~po002;
  assign new_new_n22546__ = ~new_new_n22544__ & ~new_new_n22545__;
  assign new_new_n22547__ = new_new_n22543__ & new_new_n22546__;
  assign new_new_n22548__ = ~new_new_n22543__ & ~new_new_n22546__;
  assign new_new_n22549__ = ~new_new_n22547__ & ~new_new_n22548__;
  assign new_new_n22550__ = pi068 & new_new_n22549__;
  assign new_new_n22551__ = ~pi068 & ~new_new_n22549__;
  assign new_new_n22552__ = pi002 & po002;
  assign new_new_n22553__ = ~pi002 & ~po002;
  assign new_new_n22554__ = ~pi065 & ~new_new_n22552__;
  assign new_new_n22555__ = ~new_new_n22553__ & new_new_n22554__;
  assign new_new_n22556__ = ~pi001 & ~new_new_n22555__;
  assign new_new_n22557__ = pi065 & new_new_n22552__;
  assign new_new_n22558__ = ~new_new_n22556__ & ~new_new_n22557__;
  assign new_new_n22559__ = pi064 & ~new_new_n22558__;
  assign new_new_n22560__ = pi064 & po002;
  assign new_new_n22561__ = new_new_n21872__ & ~new_new_n22560__;
  assign new_new_n22562__ = ~new_new_n22559__ & ~new_new_n22561__;
  assign new_new_n22563__ = pi066 & ~new_new_n22562__;
  assign new_new_n22564__ = ~pi066 & new_new_n22562__;
  assign new_new_n22565__ = po003 & ~new_new_n22035__;
  assign new_new_n22566__ = ~pi065 & ~po002;
  assign new_new_n22567__ = pi065 & po003;
  assign new_new_n22568__ = ~pi065 & ~po003;
  assign new_new_n22569__ = ~new_new_n22567__ & ~new_new_n22568__;
  assign new_new_n22570__ = ~pi002 & ~new_new_n22569__;
  assign new_new_n22571__ = ~new_new_n22566__ & new_new_n22570__;
  assign new_new_n22572__ = ~new_new_n22565__ & ~new_new_n22571__;
  assign new_new_n22573__ = pi064 & ~new_new_n22572__;
  assign new_new_n22574__ = pi065 & po002;
  assign new_new_n22575__ = ~new_new_n21865__ & ~new_new_n22574__;
  assign new_new_n22576__ = pi002 & ~new_new_n22567__;
  assign new_new_n22577__ = pi064 & ~new_new_n22576__;
  assign new_new_n22578__ = ~new_new_n22575__ & ~new_new_n22577__;
  assign new_new_n22579__ = ~new_new_n22573__ & ~new_new_n22578__;
  assign new_new_n22580__ = pi003 & ~new_new_n22579__;
  assign new_new_n22581__ = ~pi003 & new_new_n22579__;
  assign new_new_n22582__ = ~new_new_n22580__ & ~new_new_n22581__;
  assign new_new_n22583__ = ~new_new_n22564__ & ~new_new_n22582__;
  assign new_new_n22584__ = ~new_new_n22563__ & ~new_new_n22583__;
  assign new_new_n22585__ = pi067 & ~new_new_n22584__;
  assign new_new_n22586__ = ~pi067 & new_new_n22584__;
  assign new_new_n22587__ = ~new_new_n21201__ & ~new_new_n21882__;
  assign new_new_n22588__ = ~pi065 & ~po004;
  assign new_new_n22589__ = new_new_n21201__ & new_new_n22567__;
  assign new_new_n22590__ = ~new_new_n22588__ & ~new_new_n22589__;
  assign new_new_n22591__ = pi003 & ~new_new_n22590__;
  assign new_new_n22592__ = po004 & ~po003;
  assign new_new_n22593__ = ~new_new_n426__ & ~po004;
  assign new_new_n22594__ = ~pi003 & ~new_new_n21212__;
  assign new_new_n22595__ = ~new_new_n22593__ & new_new_n22594__;
  assign new_new_n22596__ = ~new_new_n22592__ & new_new_n22595__;
  assign new_new_n22597__ = ~new_new_n22587__ & ~new_new_n22596__;
  assign new_new_n22598__ = ~new_new_n22591__ & new_new_n22597__;
  assign new_new_n22599__ = pi004 & ~new_new_n22598__;
  assign new_new_n22600__ = ~new_new_n21212__ & ~new_new_n22588__;
  assign new_new_n22601__ = ~pi003 & ~new_new_n22600__;
  assign new_new_n22602__ = ~new_new_n22568__ & new_new_n22601__;
  assign new_new_n22603__ = ~new_new_n22592__ & ~new_new_n22602__;
  assign new_new_n22604__ = pi064 & ~new_new_n22603__;
  assign new_new_n22605__ = ~new_new_n21201__ & ~new_new_n22567__;
  assign new_new_n22606__ = pi003 & ~new_new_n21212__;
  assign new_new_n22607__ = pi064 & ~new_new_n22606__;
  assign new_new_n22608__ = ~new_new_n22605__ & ~new_new_n22607__;
  assign new_new_n22609__ = ~new_new_n22604__ & ~new_new_n22608__;
  assign new_new_n22610__ = ~pi004 & ~new_new_n22609__;
  assign new_new_n22611__ = ~new_new_n22599__ & ~new_new_n22610__;
  assign new_new_n22612__ = ~new_new_n21847__ & new_new_n21848__;
  assign new_new_n22613__ = ~pi003 & ~po003;
  assign new_new_n22614__ = ~pi065 & ~new_new_n22613__;
  assign new_new_n22615__ = ~pi002 & ~new_new_n22614__;
  assign new_new_n22616__ = ~new_new_n22612__ & ~new_new_n22615__;
  assign new_new_n22617__ = pi064 & ~new_new_n22616__;
  assign new_new_n22618__ = ~new_new_n21866__ & ~new_new_n22617__;
  assign new_new_n22619__ = ~pi066 & new_new_n22618__;
  assign new_new_n22620__ = pi066 & ~new_new_n22618__;
  assign new_new_n22621__ = ~new_new_n22619__ & ~new_new_n22620__;
  assign new_new_n22622__ = po002 & new_new_n22621__;
  assign new_new_n22623__ = ~new_new_n22611__ & new_new_n22622__;
  assign new_new_n22624__ = new_new_n22611__ & ~new_new_n22622__;
  assign new_new_n22625__ = ~new_new_n22623__ & ~new_new_n22624__;
  assign new_new_n22626__ = ~new_new_n22586__ & ~new_new_n22625__;
  assign new_new_n22627__ = ~new_new_n22585__ & ~new_new_n22626__;
  assign new_new_n22628__ = ~new_new_n22551__ & ~new_new_n22627__;
  assign new_new_n22629__ = ~new_new_n22550__ & ~new_new_n22628__;
  assign new_new_n22630__ = ~new_new_n22542__ & ~new_new_n22629__;
  assign new_new_n22631__ = ~new_new_n22541__ & ~new_new_n22630__;
  assign new_new_n22632__ = ~new_new_n22535__ & ~new_new_n22631__;
  assign new_new_n22633__ = ~new_new_n22534__ & ~new_new_n22632__;
  assign new_new_n22634__ = ~new_new_n22526__ & new_new_n22633__;
  assign new_new_n22635__ = ~new_new_n22525__ & ~new_new_n22634__;
  assign new_new_n22636__ = ~new_new_n22517__ & ~new_new_n22635__;
  assign new_new_n22637__ = ~new_new_n22516__ & ~new_new_n22636__;
  assign new_new_n22638__ = ~new_new_n22508__ & ~new_new_n22637__;
  assign new_new_n22639__ = ~new_new_n22507__ & ~new_new_n22638__;
  assign new_new_n22640__ = ~new_new_n22501__ & ~new_new_n22639__;
  assign new_new_n22641__ = ~new_new_n22500__ & ~new_new_n22640__;
  assign new_new_n22642__ = ~new_new_n22492__ & new_new_n22641__;
  assign new_new_n22643__ = ~new_new_n22491__ & ~new_new_n22642__;
  assign new_new_n22644__ = ~new_new_n22483__ & new_new_n22643__;
  assign new_new_n22645__ = ~new_new_n22482__ & ~new_new_n22644__;
  assign new_new_n22646__ = ~new_new_n22474__ & ~new_new_n22645__;
  assign new_new_n22647__ = ~new_new_n22473__ & ~new_new_n22646__;
  assign new_new_n22648__ = ~new_new_n22465__ & ~new_new_n22647__;
  assign new_new_n22649__ = ~new_new_n22464__ & ~new_new_n22648__;
  assign new_new_n22650__ = ~new_new_n22456__ & ~new_new_n22649__;
  assign new_new_n22651__ = ~new_new_n22455__ & ~new_new_n22650__;
  assign new_new_n22652__ = ~new_new_n22447__ & ~new_new_n22651__;
  assign new_new_n22653__ = ~new_new_n22446__ & ~new_new_n22652__;
  assign new_new_n22654__ = ~new_new_n22438__ & ~new_new_n22653__;
  assign new_new_n22655__ = ~new_new_n22437__ & ~new_new_n22654__;
  assign new_new_n22656__ = ~new_new_n22429__ & new_new_n22655__;
  assign new_new_n22657__ = ~new_new_n22428__ & ~new_new_n22656__;
  assign new_new_n22658__ = ~new_new_n22420__ & ~new_new_n22657__;
  assign new_new_n22659__ = ~new_new_n22419__ & ~new_new_n22658__;
  assign new_new_n22660__ = ~new_new_n22411__ & new_new_n22659__;
  assign new_new_n22661__ = ~new_new_n22410__ & ~new_new_n22660__;
  assign new_new_n22662__ = ~new_new_n22402__ & new_new_n22661__;
  assign new_new_n22663__ = ~new_new_n22401__ & ~new_new_n22662__;
  assign new_new_n22664__ = ~new_new_n22393__ & ~new_new_n22663__;
  assign new_new_n22665__ = ~new_new_n22392__ & ~new_new_n22664__;
  assign new_new_n22666__ = ~new_new_n22384__ & ~new_new_n22665__;
  assign new_new_n22667__ = ~new_new_n22383__ & ~new_new_n22666__;
  assign new_new_n22668__ = ~new_new_n22375__ & ~new_new_n22667__;
  assign new_new_n22669__ = ~new_new_n22374__ & ~new_new_n22668__;
  assign new_new_n22670__ = ~new_new_n22366__ & ~new_new_n22669__;
  assign new_new_n22671__ = ~new_new_n22365__ & ~new_new_n22670__;
  assign new_new_n22672__ = ~new_new_n22357__ & ~new_new_n22671__;
  assign new_new_n22673__ = ~new_new_n22356__ & ~new_new_n22672__;
  assign new_new_n22674__ = ~new_new_n22348__ & ~new_new_n22673__;
  assign new_new_n22675__ = ~new_new_n22347__ & ~new_new_n22674__;
  assign new_new_n22676__ = ~new_new_n22339__ & new_new_n22675__;
  assign new_new_n22677__ = ~new_new_n22338__ & ~new_new_n22676__;
  assign new_new_n22678__ = ~new_new_n22330__ & ~new_new_n22677__;
  assign new_new_n22679__ = ~new_new_n22329__ & ~new_new_n22678__;
  assign new_new_n22680__ = ~new_new_n22321__ & ~new_new_n22679__;
  assign new_new_n22681__ = ~new_new_n22320__ & ~new_new_n22680__;
  assign new_new_n22682__ = ~new_new_n22312__ & ~new_new_n22681__;
  assign new_new_n22683__ = ~new_new_n22311__ & ~new_new_n22682__;
  assign new_new_n22684__ = ~new_new_n22303__ & ~new_new_n22683__;
  assign new_new_n22685__ = ~new_new_n22302__ & ~new_new_n22684__;
  assign new_new_n22686__ = ~new_new_n22294__ & ~new_new_n22685__;
  assign new_new_n22687__ = ~new_new_n22293__ & ~new_new_n22686__;
  assign new_new_n22688__ = ~new_new_n22285__ & new_new_n22687__;
  assign new_new_n22689__ = ~new_new_n22284__ & ~new_new_n22688__;
  assign new_new_n22690__ = ~new_new_n22276__ & ~new_new_n22689__;
  assign new_new_n22691__ = ~new_new_n22275__ & ~new_new_n22690__;
  assign new_new_n22692__ = ~new_new_n22267__ & new_new_n22691__;
  assign new_new_n22693__ = ~new_new_n22266__ & ~new_new_n22692__;
  assign new_new_n22694__ = ~new_new_n22258__ & ~new_new_n22693__;
  assign new_new_n22695__ = ~new_new_n22257__ & ~new_new_n22694__;
  assign new_new_n22696__ = ~new_new_n22249__ & ~new_new_n22695__;
  assign new_new_n22697__ = ~new_new_n22248__ & ~new_new_n22696__;
  assign new_new_n22698__ = ~new_new_n22240__ & ~new_new_n22697__;
  assign new_new_n22699__ = ~new_new_n22239__ & ~new_new_n22698__;
  assign new_new_n22700__ = ~new_new_n22231__ & ~new_new_n22699__;
  assign new_new_n22701__ = ~new_new_n22230__ & ~new_new_n22700__;
  assign new_new_n22702__ = ~new_new_n22222__ & new_new_n22701__;
  assign new_new_n22703__ = ~new_new_n22221__ & ~new_new_n22702__;
  assign new_new_n22704__ = ~new_new_n22213__ & new_new_n22703__;
  assign new_new_n22705__ = ~new_new_n22212__ & ~new_new_n22704__;
  assign new_new_n22706__ = ~new_new_n22204__ & new_new_n22705__;
  assign new_new_n22707__ = ~new_new_n22203__ & ~new_new_n22706__;
  assign new_new_n22708__ = ~new_new_n22195__ & ~new_new_n22707__;
  assign new_new_n22709__ = ~new_new_n22194__ & ~new_new_n22708__;
  assign new_new_n22710__ = ~new_new_n22186__ & new_new_n22709__;
  assign new_new_n22711__ = ~new_new_n22185__ & ~new_new_n22710__;
  assign new_new_n22712__ = ~new_new_n22177__ & new_new_n22711__;
  assign new_new_n22713__ = ~new_new_n22176__ & ~new_new_n22712__;
  assign new_new_n22714__ = ~new_new_n22168__ & ~new_new_n22713__;
  assign new_new_n22715__ = ~new_new_n22167__ & ~new_new_n22714__;
  assign new_new_n22716__ = ~new_new_n22159__ & new_new_n22715__;
  assign new_new_n22717__ = ~new_new_n22158__ & ~new_new_n22716__;
  assign new_new_n22718__ = ~new_new_n22150__ & ~new_new_n22717__;
  assign new_new_n22719__ = ~new_new_n22149__ & ~new_new_n22718__;
  assign new_new_n22720__ = ~new_new_n22141__ & new_new_n22719__;
  assign new_new_n22721__ = ~new_new_n22140__ & ~new_new_n22720__;
  assign new_new_n22722__ = ~new_new_n22132__ & ~new_new_n22721__;
  assign new_new_n22723__ = ~new_new_n22131__ & ~new_new_n22722__;
  assign new_new_n22724__ = ~new_new_n22123__ & ~new_new_n22723__;
  assign new_new_n22725__ = ~new_new_n22122__ & ~new_new_n22724__;
  assign new_new_n22726__ = ~new_new_n22114__ & ~new_new_n22725__;
  assign new_new_n22727__ = ~new_new_n22113__ & ~new_new_n22726__;
  assign new_new_n22728__ = ~new_new_n22105__ & new_new_n22727__;
  assign new_new_n22729__ = ~new_new_n22104__ & ~new_new_n22728__;
  assign new_new_n22730__ = ~new_new_n22096__ & new_new_n22729__;
  assign new_new_n22731__ = ~new_new_n22095__ & ~new_new_n22730__;
  assign new_new_n22732__ = ~new_new_n22087__ & ~new_new_n22731__;
  assign new_new_n22733__ = ~new_new_n22086__ & ~new_new_n22732__;
  assign new_new_n22734__ = ~new_new_n22078__ & ~new_new_n22733__;
  assign new_new_n22735__ = ~new_new_n22077__ & ~new_new_n22734__;
  assign new_new_n22736__ = ~new_new_n22069__ & ~new_new_n22735__;
  assign new_new_n22737__ = ~new_new_n22068__ & ~new_new_n22736__;
  assign new_new_n22738__ = ~new_new_n22060__ & new_new_n22737__;
  assign new_new_n22739__ = ~new_new_n22059__ & ~new_new_n22738__;
  assign new_new_n22740__ = ~new_new_n22051__ & ~new_new_n22739__;
  assign new_new_n22741__ = ~new_new_n22050__ & ~new_new_n22740__;
  assign new_new_n22742__ = ~pi125 & new_new_n22741__;
  assign new_new_n22743__ = pi125 & ~new_new_n22741__;
  assign new_new_n22744__ = ~new_new_n22742__ & ~new_new_n22743__;
  assign new_new_n22745__ = pi126 & ~new_new_n22030__;
  assign new_new_n22746__ = ~pi127 & ~new_new_n22745__;
  assign new_new_n22747__ = ~new_new_n22744__ & new_new_n22746__;
  assign new_new_n22748__ = new_new_n22042__ & ~new_new_n22747__;
  assign new_new_n22749__ = pi125 & new_new_n22033__;
  assign new_new_n22750__ = ~pi125 & ~new_new_n22033__;
  assign new_new_n22751__ = new_new_n260__ & ~new_new_n22749__;
  assign new_new_n22752__ = ~new_new_n22750__ & new_new_n22751__;
  assign new_new_n22753__ = new_new_n22030__ & ~new_new_n22752__;
  assign new_new_n22754__ = new_new_n260__ & new_new_n22753__;
  assign new_new_n22755__ = ~new_new_n22042__ & new_new_n22754__;
  assign new_new_n22756__ = ~new_new_n22744__ & new_new_n22755__;
  assign new_new_n22757__ = ~new_new_n22748__ & ~new_new_n22756__;
  assign new_new_n22758__ = pi126 & new_new_n22757__;
  assign new_new_n22759__ = ~pi126 & ~new_new_n22757__;
  assign new_new_n22760__ = ~new_new_n22050__ & ~new_new_n22051__;
  assign new_new_n22761__ = pi125 & ~new_new_n22042__;
  assign new_new_n22762__ = ~pi125 & new_new_n22042__;
  assign new_new_n22763__ = new_new_n22741__ & ~new_new_n22762__;
  assign new_new_n22764__ = ~new_new_n22761__ & ~new_new_n22763__;
  assign new_new_n22765__ = ~pi126 & new_new_n22764__;
  assign new_new_n22766__ = ~new_new_n22753__ & ~new_new_n22765__;
  assign new_new_n22767__ = pi126 & ~new_new_n22764__;
  assign new_new_n22768__ = ~pi127 & ~new_new_n22767__;
  assign po001 = ~new_new_n22766__ & new_new_n22768__;
  assign new_new_n22770__ = ~new_new_n22739__ & po001;
  assign new_new_n22771__ = ~pi124 & ~po001;
  assign new_new_n22772__ = ~new_new_n22770__ & ~new_new_n22771__;
  assign new_new_n22773__ = new_new_n22760__ & ~new_new_n22772__;
  assign new_new_n22774__ = ~new_new_n22760__ & new_new_n22772__;
  assign new_new_n22775__ = ~new_new_n22773__ & ~new_new_n22774__;
  assign new_new_n22776__ = pi125 & ~new_new_n22775__;
  assign new_new_n22777__ = ~pi125 & new_new_n22775__;
  assign new_new_n22778__ = ~new_new_n22737__ & po001;
  assign new_new_n22779__ = pi123 & ~po001;
  assign new_new_n22780__ = ~new_new_n22778__ & ~new_new_n22779__;
  assign new_new_n22781__ = ~new_new_n22059__ & ~new_new_n22060__;
  assign new_new_n22782__ = ~new_new_n22780__ & new_new_n22781__;
  assign new_new_n22783__ = new_new_n22780__ & ~new_new_n22781__;
  assign new_new_n22784__ = ~new_new_n22782__ & ~new_new_n22783__;
  assign new_new_n22785__ = ~pi124 & ~new_new_n22784__;
  assign new_new_n22786__ = pi124 & new_new_n22784__;
  assign new_new_n22787__ = ~new_new_n22735__ & po001;
  assign new_new_n22788__ = pi122 & ~po001;
  assign new_new_n22789__ = ~new_new_n22787__ & ~new_new_n22788__;
  assign new_new_n22790__ = ~new_new_n22068__ & ~new_new_n22069__;
  assign new_new_n22791__ = ~new_new_n22789__ & new_new_n22790__;
  assign new_new_n22792__ = new_new_n22789__ & ~new_new_n22790__;
  assign new_new_n22793__ = ~new_new_n22791__ & ~new_new_n22792__;
  assign new_new_n22794__ = ~pi123 & ~new_new_n22793__;
  assign new_new_n22795__ = pi123 & new_new_n22793__;
  assign new_new_n22796__ = pi121 & ~new_new_n22733__;
  assign new_new_n22797__ = ~pi121 & new_new_n22733__;
  assign new_new_n22798__ = ~new_new_n22796__ & ~new_new_n22797__;
  assign new_new_n22799__ = po001 & new_new_n22798__;
  assign new_new_n22800__ = new_new_n22076__ & new_new_n22799__;
  assign new_new_n22801__ = ~new_new_n22076__ & ~new_new_n22799__;
  assign new_new_n22802__ = ~new_new_n22800__ & ~new_new_n22801__;
  assign new_new_n22803__ = ~pi122 & new_new_n22802__;
  assign new_new_n22804__ = pi122 & ~new_new_n22802__;
  assign new_new_n22805__ = ~new_new_n22731__ & po001;
  assign new_new_n22806__ = pi120 & ~po001;
  assign new_new_n22807__ = ~new_new_n22805__ & ~new_new_n22806__;
  assign new_new_n22808__ = ~new_new_n22086__ & ~new_new_n22087__;
  assign new_new_n22809__ = ~new_new_n22807__ & new_new_n22808__;
  assign new_new_n22810__ = new_new_n22807__ & ~new_new_n22808__;
  assign new_new_n22811__ = ~new_new_n22809__ & ~new_new_n22810__;
  assign new_new_n22812__ = ~pi121 & ~new_new_n22811__;
  assign new_new_n22813__ = pi121 & new_new_n22811__;
  assign new_new_n22814__ = ~new_new_n22095__ & ~new_new_n22096__;
  assign new_new_n22815__ = ~new_new_n22729__ & po001;
  assign new_new_n22816__ = ~pi119 & ~po001;
  assign new_new_n22817__ = ~new_new_n22815__ & ~new_new_n22816__;
  assign new_new_n22818__ = new_new_n22814__ & ~new_new_n22817__;
  assign new_new_n22819__ = ~new_new_n22814__ & new_new_n22817__;
  assign new_new_n22820__ = ~new_new_n22818__ & ~new_new_n22819__;
  assign new_new_n22821__ = pi120 & ~new_new_n22820__;
  assign new_new_n22822__ = ~pi120 & new_new_n22820__;
  assign new_new_n22823__ = ~new_new_n22104__ & ~new_new_n22105__;
  assign new_new_n22824__ = ~new_new_n22727__ & po001;
  assign new_new_n22825__ = pi118 & ~po001;
  assign new_new_n22826__ = ~new_new_n22824__ & ~new_new_n22825__;
  assign new_new_n22827__ = new_new_n22823__ & ~new_new_n22826__;
  assign new_new_n22828__ = ~new_new_n22823__ & new_new_n22826__;
  assign new_new_n22829__ = ~new_new_n22827__ & ~new_new_n22828__;
  assign new_new_n22830__ = ~pi119 & ~new_new_n22829__;
  assign new_new_n22831__ = pi119 & new_new_n22829__;
  assign new_new_n22832__ = ~new_new_n22113__ & ~new_new_n22114__;
  assign new_new_n22833__ = new_new_n22725__ & po001;
  assign new_new_n22834__ = ~pi117 & ~po001;
  assign new_new_n22835__ = ~new_new_n22833__ & ~new_new_n22834__;
  assign new_new_n22836__ = ~new_new_n22832__ & ~new_new_n22835__;
  assign new_new_n22837__ = new_new_n22832__ & new_new_n22835__;
  assign new_new_n22838__ = ~new_new_n22836__ & ~new_new_n22837__;
  assign new_new_n22839__ = ~pi118 & ~new_new_n22838__;
  assign new_new_n22840__ = pi118 & new_new_n22838__;
  assign new_new_n22841__ = pi116 & ~new_new_n22723__;
  assign new_new_n22842__ = ~pi116 & new_new_n22723__;
  assign new_new_n22843__ = ~new_new_n22841__ & ~new_new_n22842__;
  assign new_new_n22844__ = po001 & new_new_n22843__;
  assign new_new_n22845__ = new_new_n22121__ & new_new_n22844__;
  assign new_new_n22846__ = ~new_new_n22121__ & ~new_new_n22844__;
  assign new_new_n22847__ = ~new_new_n22845__ & ~new_new_n22846__;
  assign new_new_n22848__ = pi117 & ~new_new_n22847__;
  assign new_new_n22849__ = ~pi117 & new_new_n22847__;
  assign new_new_n22850__ = ~new_new_n22721__ & po001;
  assign new_new_n22851__ = pi115 & ~po001;
  assign new_new_n22852__ = ~new_new_n22850__ & ~new_new_n22851__;
  assign new_new_n22853__ = ~new_new_n22131__ & ~new_new_n22132__;
  assign new_new_n22854__ = ~new_new_n22852__ & new_new_n22853__;
  assign new_new_n22855__ = new_new_n22852__ & ~new_new_n22853__;
  assign new_new_n22856__ = ~new_new_n22854__ & ~new_new_n22855__;
  assign new_new_n22857__ = pi116 & new_new_n22856__;
  assign new_new_n22858__ = ~pi116 & ~new_new_n22856__;
  assign new_new_n22859__ = ~new_new_n22140__ & ~new_new_n22141__;
  assign new_new_n22860__ = ~new_new_n22719__ & po001;
  assign new_new_n22861__ = ~pi114 & ~po001;
  assign new_new_n22862__ = ~new_new_n22860__ & ~new_new_n22861__;
  assign new_new_n22863__ = new_new_n22859__ & ~new_new_n22862__;
  assign new_new_n22864__ = ~new_new_n22859__ & new_new_n22862__;
  assign new_new_n22865__ = ~new_new_n22863__ & ~new_new_n22864__;
  assign new_new_n22866__ = pi115 & ~new_new_n22865__;
  assign new_new_n22867__ = ~pi115 & new_new_n22865__;
  assign new_new_n22868__ = ~pi113 & ~new_new_n22717__;
  assign new_new_n22869__ = pi113 & new_new_n22717__;
  assign new_new_n22870__ = ~new_new_n22868__ & ~new_new_n22869__;
  assign new_new_n22871__ = po001 & new_new_n22870__;
  assign new_new_n22872__ = new_new_n22148__ & new_new_n22871__;
  assign new_new_n22873__ = ~new_new_n22148__ & ~new_new_n22871__;
  assign new_new_n22874__ = ~new_new_n22872__ & ~new_new_n22873__;
  assign new_new_n22875__ = ~pi114 & ~new_new_n22874__;
  assign new_new_n22876__ = pi114 & new_new_n22874__;
  assign new_new_n22877__ = ~new_new_n22715__ & po001;
  assign new_new_n22878__ = pi112 & ~po001;
  assign new_new_n22879__ = ~new_new_n22877__ & ~new_new_n22878__;
  assign new_new_n22880__ = ~new_new_n22158__ & ~new_new_n22159__;
  assign new_new_n22881__ = ~new_new_n22879__ & new_new_n22880__;
  assign new_new_n22882__ = new_new_n22879__ & ~new_new_n22880__;
  assign new_new_n22883__ = ~new_new_n22881__ & ~new_new_n22882__;
  assign new_new_n22884__ = ~pi113 & ~new_new_n22883__;
  assign new_new_n22885__ = pi113 & new_new_n22883__;
  assign new_new_n22886__ = ~new_new_n22167__ & ~new_new_n22168__;
  assign new_new_n22887__ = ~new_new_n22713__ & po001;
  assign new_new_n22888__ = pi111 & ~po001;
  assign new_new_n22889__ = ~new_new_n22887__ & ~new_new_n22888__;
  assign new_new_n22890__ = new_new_n22886__ & ~new_new_n22889__;
  assign new_new_n22891__ = ~new_new_n22886__ & new_new_n22889__;
  assign new_new_n22892__ = ~new_new_n22890__ & ~new_new_n22891__;
  assign new_new_n22893__ = pi112 & new_new_n22892__;
  assign new_new_n22894__ = ~pi112 & ~new_new_n22892__;
  assign new_new_n22895__ = ~new_new_n22176__ & ~new_new_n22177__;
  assign new_new_n22896__ = ~new_new_n22711__ & po001;
  assign new_new_n22897__ = ~pi110 & ~po001;
  assign new_new_n22898__ = ~new_new_n22896__ & ~new_new_n22897__;
  assign new_new_n22899__ = new_new_n22895__ & ~new_new_n22898__;
  assign new_new_n22900__ = ~new_new_n22895__ & new_new_n22898__;
  assign new_new_n22901__ = ~new_new_n22899__ & ~new_new_n22900__;
  assign new_new_n22902__ = pi111 & ~new_new_n22901__;
  assign new_new_n22903__ = ~pi111 & new_new_n22901__;
  assign new_new_n22904__ = ~new_new_n22709__ & po001;
  assign new_new_n22905__ = pi109 & ~po001;
  assign new_new_n22906__ = ~new_new_n22904__ & ~new_new_n22905__;
  assign new_new_n22907__ = ~new_new_n22185__ & ~new_new_n22186__;
  assign new_new_n22908__ = ~new_new_n22906__ & new_new_n22907__;
  assign new_new_n22909__ = new_new_n22906__ & ~new_new_n22907__;
  assign new_new_n22910__ = ~new_new_n22908__ & ~new_new_n22909__;
  assign new_new_n22911__ = ~pi110 & ~new_new_n22910__;
  assign new_new_n22912__ = pi110 & new_new_n22910__;
  assign new_new_n22913__ = ~new_new_n22707__ & po001;
  assign new_new_n22914__ = pi108 & ~po001;
  assign new_new_n22915__ = ~new_new_n22913__ & ~new_new_n22914__;
  assign new_new_n22916__ = ~new_new_n22194__ & ~new_new_n22195__;
  assign new_new_n22917__ = ~new_new_n22915__ & new_new_n22916__;
  assign new_new_n22918__ = new_new_n22915__ & ~new_new_n22916__;
  assign new_new_n22919__ = ~new_new_n22917__ & ~new_new_n22918__;
  assign new_new_n22920__ = ~pi109 & ~new_new_n22919__;
  assign new_new_n22921__ = pi109 & new_new_n22919__;
  assign new_new_n22922__ = ~new_new_n22203__ & ~new_new_n22204__;
  assign new_new_n22923__ = ~new_new_n22705__ & po001;
  assign new_new_n22924__ = ~pi107 & ~po001;
  assign new_new_n22925__ = ~new_new_n22923__ & ~new_new_n22924__;
  assign new_new_n22926__ = new_new_n22922__ & ~new_new_n22925__;
  assign new_new_n22927__ = ~new_new_n22922__ & new_new_n22925__;
  assign new_new_n22928__ = ~new_new_n22926__ & ~new_new_n22927__;
  assign new_new_n22929__ = ~pi108 & new_new_n22928__;
  assign new_new_n22930__ = pi108 & ~new_new_n22928__;
  assign new_new_n22931__ = ~new_new_n22212__ & ~new_new_n22213__;
  assign new_new_n22932__ = ~new_new_n22703__ & po001;
  assign new_new_n22933__ = pi106 & ~po001;
  assign new_new_n22934__ = ~new_new_n22932__ & ~new_new_n22933__;
  assign new_new_n22935__ = new_new_n22931__ & ~new_new_n22934__;
  assign new_new_n22936__ = ~new_new_n22931__ & new_new_n22934__;
  assign new_new_n22937__ = ~new_new_n22935__ & ~new_new_n22936__;
  assign new_new_n22938__ = ~pi107 & ~new_new_n22937__;
  assign new_new_n22939__ = pi107 & new_new_n22937__;
  assign new_new_n22940__ = ~new_new_n22221__ & ~new_new_n22222__;
  assign new_new_n22941__ = ~new_new_n22701__ & po001;
  assign new_new_n22942__ = ~pi105 & ~po001;
  assign new_new_n22943__ = ~new_new_n22941__ & ~new_new_n22942__;
  assign new_new_n22944__ = new_new_n22940__ & ~new_new_n22943__;
  assign new_new_n22945__ = ~new_new_n22940__ & new_new_n22943__;
  assign new_new_n22946__ = ~new_new_n22944__ & ~new_new_n22945__;
  assign new_new_n22947__ = ~pi106 & new_new_n22946__;
  assign new_new_n22948__ = pi106 & ~new_new_n22946__;
  assign new_new_n22949__ = ~new_new_n22230__ & ~new_new_n22231__;
  assign new_new_n22950__ = ~new_new_n22699__ & po001;
  assign new_new_n22951__ = ~pi104 & ~po001;
  assign new_new_n22952__ = ~new_new_n22950__ & ~new_new_n22951__;
  assign new_new_n22953__ = new_new_n22949__ & ~new_new_n22952__;
  assign new_new_n22954__ = ~new_new_n22949__ & new_new_n22952__;
  assign new_new_n22955__ = ~new_new_n22953__ & ~new_new_n22954__;
  assign new_new_n22956__ = ~pi105 & new_new_n22955__;
  assign new_new_n22957__ = pi105 & ~new_new_n22955__;
  assign new_new_n22958__ = ~new_new_n22239__ & ~new_new_n22240__;
  assign new_new_n22959__ = ~new_new_n22697__ & po001;
  assign new_new_n22960__ = ~pi103 & ~po001;
  assign new_new_n22961__ = ~new_new_n22959__ & ~new_new_n22960__;
  assign new_new_n22962__ = new_new_n22958__ & ~new_new_n22961__;
  assign new_new_n22963__ = ~new_new_n22958__ & new_new_n22961__;
  assign new_new_n22964__ = ~new_new_n22962__ & ~new_new_n22963__;
  assign new_new_n22965__ = ~pi104 & new_new_n22964__;
  assign new_new_n22966__ = pi104 & ~new_new_n22964__;
  assign new_new_n22967__ = ~new_new_n22248__ & ~new_new_n22249__;
  assign new_new_n22968__ = ~new_new_n22695__ & po001;
  assign new_new_n22969__ = ~pi102 & ~po001;
  assign new_new_n22970__ = ~new_new_n22968__ & ~new_new_n22969__;
  assign new_new_n22971__ = new_new_n22967__ & new_new_n22970__;
  assign new_new_n22972__ = ~new_new_n22967__ & ~new_new_n22970__;
  assign new_new_n22973__ = ~new_new_n22971__ & ~new_new_n22972__;
  assign new_new_n22974__ = ~pi103 & ~new_new_n22973__;
  assign new_new_n22975__ = pi103 & new_new_n22973__;
  assign new_new_n22976__ = ~pi101 & ~new_new_n22693__;
  assign new_new_n22977__ = pi101 & new_new_n22693__;
  assign new_new_n22978__ = ~new_new_n22976__ & ~new_new_n22977__;
  assign new_new_n22979__ = po001 & new_new_n22978__;
  assign new_new_n22980__ = new_new_n22256__ & new_new_n22979__;
  assign new_new_n22981__ = ~new_new_n22256__ & ~new_new_n22979__;
  assign new_new_n22982__ = ~new_new_n22980__ & ~new_new_n22981__;
  assign new_new_n22983__ = ~pi102 & ~new_new_n22982__;
  assign new_new_n22984__ = pi102 & new_new_n22982__;
  assign new_new_n22985__ = new_new_n22691__ & po001;
  assign new_new_n22986__ = ~pi100 & ~po001;
  assign new_new_n22987__ = ~new_new_n22985__ & ~new_new_n22986__;
  assign new_new_n22988__ = ~new_new_n22266__ & ~new_new_n22267__;
  assign new_new_n22989__ = ~new_new_n22987__ & ~new_new_n22988__;
  assign new_new_n22990__ = new_new_n22987__ & new_new_n22988__;
  assign new_new_n22991__ = ~new_new_n22989__ & ~new_new_n22990__;
  assign new_new_n22992__ = ~pi101 & ~new_new_n22991__;
  assign new_new_n22993__ = pi101 & new_new_n22991__;
  assign new_new_n22994__ = pi099 & ~new_new_n22689__;
  assign new_new_n22995__ = ~pi099 & new_new_n22689__;
  assign new_new_n22996__ = ~new_new_n22994__ & ~new_new_n22995__;
  assign new_new_n22997__ = po001 & new_new_n22996__;
  assign new_new_n22998__ = new_new_n22274__ & new_new_n22997__;
  assign new_new_n22999__ = ~new_new_n22274__ & ~new_new_n22997__;
  assign new_new_n23000__ = ~new_new_n22998__ & ~new_new_n22999__;
  assign new_new_n23001__ = pi100 & ~new_new_n23000__;
  assign new_new_n23002__ = ~pi100 & new_new_n23000__;
  assign new_new_n23003__ = ~new_new_n22284__ & ~new_new_n22285__;
  assign new_new_n23004__ = ~new_new_n22687__ & po001;
  assign new_new_n23005__ = ~pi098 & ~po001;
  assign new_new_n23006__ = ~new_new_n23004__ & ~new_new_n23005__;
  assign new_new_n23007__ = new_new_n23003__ & ~new_new_n23006__;
  assign new_new_n23008__ = ~new_new_n23003__ & new_new_n23006__;
  assign new_new_n23009__ = ~new_new_n23007__ & ~new_new_n23008__;
  assign new_new_n23010__ = ~pi099 & new_new_n23009__;
  assign new_new_n23011__ = pi099 & ~new_new_n23009__;
  assign new_new_n23012__ = ~pi097 & ~new_new_n22685__;
  assign new_new_n23013__ = pi097 & new_new_n22685__;
  assign new_new_n23014__ = ~new_new_n23012__ & ~new_new_n23013__;
  assign new_new_n23015__ = po001 & new_new_n23014__;
  assign new_new_n23016__ = new_new_n22292__ & new_new_n23015__;
  assign new_new_n23017__ = ~new_new_n22292__ & ~new_new_n23015__;
  assign new_new_n23018__ = ~new_new_n23016__ & ~new_new_n23017__;
  assign new_new_n23019__ = ~pi098 & ~new_new_n23018__;
  assign new_new_n23020__ = pi098 & new_new_n23018__;
  assign new_new_n23021__ = ~pi096 & ~new_new_n22683__;
  assign new_new_n23022__ = pi096 & new_new_n22683__;
  assign new_new_n23023__ = ~new_new_n23021__ & ~new_new_n23022__;
  assign new_new_n23024__ = po001 & new_new_n23023__;
  assign new_new_n23025__ = new_new_n22301__ & new_new_n23024__;
  assign new_new_n23026__ = ~new_new_n22301__ & ~new_new_n23024__;
  assign new_new_n23027__ = ~new_new_n23025__ & ~new_new_n23026__;
  assign new_new_n23028__ = ~pi097 & ~new_new_n23027__;
  assign new_new_n23029__ = pi097 & new_new_n23027__;
  assign new_new_n23030__ = ~new_new_n22311__ & ~new_new_n22312__;
  assign new_new_n23031__ = ~new_new_n22681__ & po001;
  assign new_new_n23032__ = ~pi095 & ~po001;
  assign new_new_n23033__ = ~new_new_n23031__ & ~new_new_n23032__;
  assign new_new_n23034__ = new_new_n23030__ & ~new_new_n23033__;
  assign new_new_n23035__ = ~new_new_n23030__ & new_new_n23033__;
  assign new_new_n23036__ = ~new_new_n23034__ & ~new_new_n23035__;
  assign new_new_n23037__ = ~pi096 & new_new_n23036__;
  assign new_new_n23038__ = pi096 & ~new_new_n23036__;
  assign new_new_n23039__ = ~pi094 & ~new_new_n22679__;
  assign new_new_n23040__ = pi094 & new_new_n22679__;
  assign new_new_n23041__ = ~new_new_n23039__ & ~new_new_n23040__;
  assign new_new_n23042__ = po001 & new_new_n23041__;
  assign new_new_n23043__ = new_new_n22319__ & new_new_n23042__;
  assign new_new_n23044__ = ~new_new_n22319__ & ~new_new_n23042__;
  assign new_new_n23045__ = ~new_new_n23043__ & ~new_new_n23044__;
  assign new_new_n23046__ = ~pi095 & ~new_new_n23045__;
  assign new_new_n23047__ = pi095 & new_new_n23045__;
  assign new_new_n23048__ = ~pi093 & ~new_new_n22677__;
  assign new_new_n23049__ = pi093 & new_new_n22677__;
  assign new_new_n23050__ = ~new_new_n23048__ & ~new_new_n23049__;
  assign new_new_n23051__ = po001 & new_new_n23050__;
  assign new_new_n23052__ = new_new_n22328__ & new_new_n23051__;
  assign new_new_n23053__ = ~new_new_n22328__ & ~new_new_n23051__;
  assign new_new_n23054__ = ~new_new_n23052__ & ~new_new_n23053__;
  assign new_new_n23055__ = ~pi094 & ~new_new_n23054__;
  assign new_new_n23056__ = pi094 & new_new_n23054__;
  assign new_new_n23057__ = ~new_new_n22675__ & po001;
  assign new_new_n23058__ = pi092 & ~po001;
  assign new_new_n23059__ = ~new_new_n23057__ & ~new_new_n23058__;
  assign new_new_n23060__ = ~new_new_n22338__ & ~new_new_n22339__;
  assign new_new_n23061__ = ~new_new_n23059__ & new_new_n23060__;
  assign new_new_n23062__ = new_new_n23059__ & ~new_new_n23060__;
  assign new_new_n23063__ = ~new_new_n23061__ & ~new_new_n23062__;
  assign new_new_n23064__ = ~pi093 & ~new_new_n23063__;
  assign new_new_n23065__ = pi093 & new_new_n23063__;
  assign new_new_n23066__ = ~new_new_n22347__ & ~new_new_n22348__;
  assign new_new_n23067__ = pi091 & ~po001;
  assign new_new_n23068__ = ~new_new_n22673__ & po001;
  assign new_new_n23069__ = ~new_new_n23067__ & ~new_new_n23068__;
  assign new_new_n23070__ = new_new_n23066__ & new_new_n23069__;
  assign new_new_n23071__ = ~new_new_n23066__ & ~new_new_n23069__;
  assign new_new_n23072__ = ~new_new_n23070__ & ~new_new_n23071__;
  assign new_new_n23073__ = ~pi092 & new_new_n23072__;
  assign new_new_n23074__ = pi092 & ~new_new_n23072__;
  assign new_new_n23075__ = ~new_new_n22671__ & po001;
  assign new_new_n23076__ = pi090 & ~po001;
  assign new_new_n23077__ = ~new_new_n23075__ & ~new_new_n23076__;
  assign new_new_n23078__ = ~new_new_n22356__ & ~new_new_n22357__;
  assign new_new_n23079__ = ~new_new_n23077__ & new_new_n23078__;
  assign new_new_n23080__ = new_new_n23077__ & ~new_new_n23078__;
  assign new_new_n23081__ = ~new_new_n23079__ & ~new_new_n23080__;
  assign new_new_n23082__ = ~pi091 & ~new_new_n23081__;
  assign new_new_n23083__ = pi091 & new_new_n23081__;
  assign new_new_n23084__ = pi089 & ~new_new_n22669__;
  assign new_new_n23085__ = ~pi089 & new_new_n22669__;
  assign new_new_n23086__ = ~new_new_n23084__ & ~new_new_n23085__;
  assign new_new_n23087__ = po001 & new_new_n23086__;
  assign new_new_n23088__ = new_new_n22364__ & new_new_n23087__;
  assign new_new_n23089__ = ~new_new_n22364__ & ~new_new_n23087__;
  assign new_new_n23090__ = ~new_new_n23088__ & ~new_new_n23089__;
  assign new_new_n23091__ = pi090 & ~new_new_n23090__;
  assign new_new_n23092__ = ~pi090 & new_new_n23090__;
  assign new_new_n23093__ = ~new_new_n22667__ & po001;
  assign new_new_n23094__ = pi088 & ~po001;
  assign new_new_n23095__ = ~new_new_n23093__ & ~new_new_n23094__;
  assign new_new_n23096__ = ~new_new_n22374__ & ~new_new_n22375__;
  assign new_new_n23097__ = ~new_new_n23095__ & new_new_n23096__;
  assign new_new_n23098__ = new_new_n23095__ & ~new_new_n23096__;
  assign new_new_n23099__ = ~new_new_n23097__ & ~new_new_n23098__;
  assign new_new_n23100__ = ~pi089 & ~new_new_n23099__;
  assign new_new_n23101__ = pi089 & new_new_n23099__;
  assign new_new_n23102__ = ~new_new_n22383__ & ~new_new_n22384__;
  assign new_new_n23103__ = new_new_n22665__ & po001;
  assign new_new_n23104__ = ~pi087 & ~po001;
  assign new_new_n23105__ = ~new_new_n23103__ & ~new_new_n23104__;
  assign new_new_n23106__ = ~new_new_n23102__ & ~new_new_n23105__;
  assign new_new_n23107__ = new_new_n23102__ & new_new_n23105__;
  assign new_new_n23108__ = ~new_new_n23106__ & ~new_new_n23107__;
  assign new_new_n23109__ = pi088 & new_new_n23108__;
  assign new_new_n23110__ = ~pi088 & ~new_new_n23108__;
  assign new_new_n23111__ = pi086 & ~new_new_n22663__;
  assign new_new_n23112__ = ~pi086 & new_new_n22663__;
  assign new_new_n23113__ = ~new_new_n23111__ & ~new_new_n23112__;
  assign new_new_n23114__ = po001 & new_new_n23113__;
  assign new_new_n23115__ = ~new_new_n22391__ & ~new_new_n23114__;
  assign new_new_n23116__ = new_new_n22391__ & new_new_n23114__;
  assign new_new_n23117__ = ~new_new_n23115__ & ~new_new_n23116__;
  assign new_new_n23118__ = pi087 & ~new_new_n23117__;
  assign new_new_n23119__ = ~pi087 & new_new_n23117__;
  assign new_new_n23120__ = ~new_new_n22401__ & ~new_new_n22402__;
  assign new_new_n23121__ = ~new_new_n22661__ & po001;
  assign new_new_n23122__ = ~pi085 & ~po001;
  assign new_new_n23123__ = ~new_new_n23121__ & ~new_new_n23122__;
  assign new_new_n23124__ = new_new_n23120__ & ~new_new_n23123__;
  assign new_new_n23125__ = ~new_new_n23120__ & new_new_n23123__;
  assign new_new_n23126__ = ~new_new_n23124__ & ~new_new_n23125__;
  assign new_new_n23127__ = pi086 & ~new_new_n23126__;
  assign new_new_n23128__ = ~pi086 & new_new_n23126__;
  assign new_new_n23129__ = ~new_new_n22659__ & po001;
  assign new_new_n23130__ = pi084 & ~po001;
  assign new_new_n23131__ = ~new_new_n23129__ & ~new_new_n23130__;
  assign new_new_n23132__ = ~new_new_n22410__ & ~new_new_n22411__;
  assign new_new_n23133__ = ~new_new_n23131__ & new_new_n23132__;
  assign new_new_n23134__ = new_new_n23131__ & ~new_new_n23132__;
  assign new_new_n23135__ = ~new_new_n23133__ & ~new_new_n23134__;
  assign new_new_n23136__ = ~pi085 & ~new_new_n23135__;
  assign new_new_n23137__ = pi085 & new_new_n23135__;
  assign new_new_n23138__ = pi083 & ~new_new_n22657__;
  assign new_new_n23139__ = ~pi083 & new_new_n22657__;
  assign new_new_n23140__ = ~new_new_n23138__ & ~new_new_n23139__;
  assign new_new_n23141__ = po001 & new_new_n23140__;
  assign new_new_n23142__ = new_new_n22418__ & new_new_n23141__;
  assign new_new_n23143__ = ~new_new_n22418__ & ~new_new_n23141__;
  assign new_new_n23144__ = ~new_new_n23142__ & ~new_new_n23143__;
  assign new_new_n23145__ = pi084 & ~new_new_n23144__;
  assign new_new_n23146__ = ~pi084 & new_new_n23144__;
  assign new_new_n23147__ = ~new_new_n22428__ & ~new_new_n22429__;
  assign new_new_n23148__ = ~new_new_n22655__ & po001;
  assign new_new_n23149__ = ~pi082 & ~po001;
  assign new_new_n23150__ = ~new_new_n23148__ & ~new_new_n23149__;
  assign new_new_n23151__ = new_new_n23147__ & ~new_new_n23150__;
  assign new_new_n23152__ = ~new_new_n23147__ & new_new_n23150__;
  assign new_new_n23153__ = ~new_new_n23151__ & ~new_new_n23152__;
  assign new_new_n23154__ = pi083 & ~new_new_n23153__;
  assign new_new_n23155__ = ~pi083 & new_new_n23153__;
  assign new_new_n23156__ = ~pi081 & ~new_new_n22653__;
  assign new_new_n23157__ = pi081 & new_new_n22653__;
  assign new_new_n23158__ = ~new_new_n23156__ & ~new_new_n23157__;
  assign new_new_n23159__ = po001 & new_new_n23158__;
  assign new_new_n23160__ = new_new_n22436__ & new_new_n23159__;
  assign new_new_n23161__ = ~new_new_n22436__ & ~new_new_n23159__;
  assign new_new_n23162__ = ~new_new_n23160__ & ~new_new_n23161__;
  assign new_new_n23163__ = ~pi082 & ~new_new_n23162__;
  assign new_new_n23164__ = pi082 & new_new_n23162__;
  assign new_new_n23165__ = ~pi080 & ~new_new_n22651__;
  assign new_new_n23166__ = pi080 & new_new_n22651__;
  assign new_new_n23167__ = ~new_new_n23165__ & ~new_new_n23166__;
  assign new_new_n23168__ = po001 & new_new_n23167__;
  assign new_new_n23169__ = new_new_n22445__ & new_new_n23168__;
  assign new_new_n23170__ = ~new_new_n22445__ & ~new_new_n23168__;
  assign new_new_n23171__ = ~new_new_n23169__ & ~new_new_n23170__;
  assign new_new_n23172__ = ~pi081 & ~new_new_n23171__;
  assign new_new_n23173__ = pi081 & new_new_n23171__;
  assign new_new_n23174__ = ~pi079 & ~new_new_n22649__;
  assign new_new_n23175__ = pi079 & new_new_n22649__;
  assign new_new_n23176__ = ~new_new_n23174__ & ~new_new_n23175__;
  assign new_new_n23177__ = po001 & new_new_n23176__;
  assign new_new_n23178__ = new_new_n22454__ & new_new_n23177__;
  assign new_new_n23179__ = ~new_new_n22454__ & ~new_new_n23177__;
  assign new_new_n23180__ = ~new_new_n23178__ & ~new_new_n23179__;
  assign new_new_n23181__ = ~pi080 & ~new_new_n23180__;
  assign new_new_n23182__ = pi080 & new_new_n23180__;
  assign new_new_n23183__ = ~pi078 & ~new_new_n22647__;
  assign new_new_n23184__ = pi078 & new_new_n22647__;
  assign new_new_n23185__ = ~new_new_n23183__ & ~new_new_n23184__;
  assign new_new_n23186__ = po001 & new_new_n23185__;
  assign new_new_n23187__ = new_new_n22463__ & new_new_n23186__;
  assign new_new_n23188__ = ~new_new_n22463__ & ~new_new_n23186__;
  assign new_new_n23189__ = ~new_new_n23187__ & ~new_new_n23188__;
  assign new_new_n23190__ = ~pi079 & ~new_new_n23189__;
  assign new_new_n23191__ = pi079 & new_new_n23189__;
  assign new_new_n23192__ = ~pi077 & ~new_new_n22645__;
  assign new_new_n23193__ = pi077 & new_new_n22645__;
  assign new_new_n23194__ = ~new_new_n23192__ & ~new_new_n23193__;
  assign new_new_n23195__ = po001 & new_new_n23194__;
  assign new_new_n23196__ = new_new_n22472__ & new_new_n23195__;
  assign new_new_n23197__ = ~new_new_n22472__ & ~new_new_n23195__;
  assign new_new_n23198__ = ~new_new_n23196__ & ~new_new_n23197__;
  assign new_new_n23199__ = ~pi078 & ~new_new_n23198__;
  assign new_new_n23200__ = pi078 & new_new_n23198__;
  assign new_new_n23201__ = ~new_new_n22643__ & po001;
  assign new_new_n23202__ = pi076 & ~po001;
  assign new_new_n23203__ = ~new_new_n23201__ & ~new_new_n23202__;
  assign new_new_n23204__ = ~new_new_n22482__ & ~new_new_n22483__;
  assign new_new_n23205__ = ~new_new_n23203__ & new_new_n23204__;
  assign new_new_n23206__ = new_new_n23203__ & ~new_new_n23204__;
  assign new_new_n23207__ = ~new_new_n23205__ & ~new_new_n23206__;
  assign new_new_n23208__ = ~pi077 & ~new_new_n23207__;
  assign new_new_n23209__ = pi077 & new_new_n23207__;
  assign new_new_n23210__ = ~new_new_n22491__ & ~new_new_n22492__;
  assign new_new_n23211__ = ~new_new_n22641__ & po001;
  assign new_new_n23212__ = ~pi075 & ~po001;
  assign new_new_n23213__ = ~new_new_n23211__ & ~new_new_n23212__;
  assign new_new_n23214__ = new_new_n23210__ & ~new_new_n23213__;
  assign new_new_n23215__ = ~new_new_n23210__ & new_new_n23213__;
  assign new_new_n23216__ = ~new_new_n23214__ & ~new_new_n23215__;
  assign new_new_n23217__ = ~pi076 & new_new_n23216__;
  assign new_new_n23218__ = pi076 & ~new_new_n23216__;
  assign new_new_n23219__ = ~new_new_n22500__ & ~new_new_n22501__;
  assign new_new_n23220__ = ~new_new_n22639__ & po001;
  assign new_new_n23221__ = ~pi074 & ~po001;
  assign new_new_n23222__ = ~new_new_n23220__ & ~new_new_n23221__;
  assign new_new_n23223__ = new_new_n23219__ & ~new_new_n23222__;
  assign new_new_n23224__ = ~new_new_n23219__ & new_new_n23222__;
  assign new_new_n23225__ = ~new_new_n23223__ & ~new_new_n23224__;
  assign new_new_n23226__ = ~pi075 & new_new_n23225__;
  assign new_new_n23227__ = pi075 & ~new_new_n23225__;
  assign new_new_n23228__ = ~new_new_n22507__ & ~new_new_n22508__;
  assign new_new_n23229__ = ~new_new_n22637__ & po001;
  assign new_new_n23230__ = ~pi073 & ~po001;
  assign new_new_n23231__ = ~new_new_n23229__ & ~new_new_n23230__;
  assign new_new_n23232__ = ~new_new_n23228__ & ~new_new_n23231__;
  assign new_new_n23233__ = new_new_n23228__ & new_new_n23231__;
  assign new_new_n23234__ = ~new_new_n23232__ & ~new_new_n23233__;
  assign new_new_n23235__ = ~pi074 & ~new_new_n23234__;
  assign new_new_n23236__ = pi074 & new_new_n23234__;
  assign new_new_n23237__ = ~new_new_n22516__ & ~new_new_n22517__;
  assign new_new_n23238__ = ~new_new_n22635__ & po001;
  assign new_new_n23239__ = ~pi072 & ~po001;
  assign new_new_n23240__ = ~new_new_n23238__ & ~new_new_n23239__;
  assign new_new_n23241__ = ~new_new_n23237__ & ~new_new_n23240__;
  assign new_new_n23242__ = new_new_n23237__ & new_new_n23240__;
  assign new_new_n23243__ = ~new_new_n23241__ & ~new_new_n23242__;
  assign new_new_n23244__ = ~pi073 & ~new_new_n23243__;
  assign new_new_n23245__ = pi073 & new_new_n23243__;
  assign new_new_n23246__ = new_new_n22633__ & po001;
  assign new_new_n23247__ = ~pi071 & ~po001;
  assign new_new_n23248__ = ~new_new_n23246__ & ~new_new_n23247__;
  assign new_new_n23249__ = ~new_new_n22525__ & ~new_new_n22526__;
  assign new_new_n23250__ = ~new_new_n23248__ & ~new_new_n23249__;
  assign new_new_n23251__ = new_new_n23248__ & new_new_n23249__;
  assign new_new_n23252__ = ~new_new_n23250__ & ~new_new_n23251__;
  assign new_new_n23253__ = pi072 & new_new_n23252__;
  assign new_new_n23254__ = ~pi072 & ~new_new_n23252__;
  assign new_new_n23255__ = pi070 & ~new_new_n22631__;
  assign new_new_n23256__ = ~pi070 & new_new_n22631__;
  assign new_new_n23257__ = ~new_new_n23255__ & ~new_new_n23256__;
  assign new_new_n23258__ = po001 & new_new_n23257__;
  assign new_new_n23259__ = ~new_new_n22533__ & ~new_new_n23258__;
  assign new_new_n23260__ = new_new_n22533__ & new_new_n23258__;
  assign new_new_n23261__ = ~new_new_n23259__ & ~new_new_n23260__;
  assign new_new_n23262__ = pi071 & ~new_new_n23261__;
  assign new_new_n23263__ = ~pi071 & new_new_n23261__;
  assign new_new_n23264__ = ~new_new_n22629__ & po001;
  assign new_new_n23265__ = pi069 & ~po001;
  assign new_new_n23266__ = ~new_new_n23264__ & ~new_new_n23265__;
  assign new_new_n23267__ = ~new_new_n22541__ & ~new_new_n22542__;
  assign new_new_n23268__ = ~new_new_n23266__ & new_new_n23267__;
  assign new_new_n23269__ = new_new_n23266__ & ~new_new_n23267__;
  assign new_new_n23270__ = ~new_new_n23268__ & ~new_new_n23269__;
  assign new_new_n23271__ = pi070 & new_new_n23270__;
  assign new_new_n23272__ = ~pi070 & ~new_new_n23270__;
  assign new_new_n23273__ = ~new_new_n22627__ & po001;
  assign new_new_n23274__ = pi068 & ~po001;
  assign new_new_n23275__ = ~new_new_n23273__ & ~new_new_n23274__;
  assign new_new_n23276__ = ~new_new_n22550__ & ~new_new_n22551__;
  assign new_new_n23277__ = ~new_new_n23275__ & new_new_n23276__;
  assign new_new_n23278__ = new_new_n23275__ & ~new_new_n23276__;
  assign new_new_n23279__ = ~new_new_n23277__ & ~new_new_n23278__;
  assign new_new_n23280__ = pi069 & new_new_n23279__;
  assign new_new_n23281__ = ~pi069 & ~new_new_n23279__;
  assign new_new_n23282__ = ~new_new_n22563__ & ~new_new_n22564__;
  assign new_new_n23283__ = po001 & new_new_n23282__;
  assign new_new_n23284__ = new_new_n22582__ & new_new_n23283__;
  assign new_new_n23285__ = ~new_new_n22582__ & ~new_new_n23283__;
  assign new_new_n23286__ = ~new_new_n23284__ & ~new_new_n23285__;
  assign new_new_n23287__ = pi067 & ~new_new_n23286__;
  assign new_new_n23288__ = ~pi067 & new_new_n23286__;
  assign new_new_n23289__ = pi001 & po001;
  assign new_new_n23290__ = pi000 & ~pi065;
  assign new_new_n23291__ = new_new_n23289__ & ~new_new_n23290__;
  assign new_new_n23292__ = ~pi001 & ~po001;
  assign new_new_n23293__ = ~pi065 & ~new_new_n23292__;
  assign new_new_n23294__ = ~pi000 & ~new_new_n23293__;
  assign new_new_n23295__ = ~new_new_n23291__ & ~new_new_n23294__;
  assign new_new_n23296__ = pi064 & ~new_new_n23295__;
  assign new_new_n23297__ = pi064 & po001;
  assign new_new_n23298__ = pi065 & ~new_new_n23297__;
  assign new_new_n23299__ = ~pi001 & new_new_n23298__;
  assign new_new_n23300__ = ~new_new_n23296__ & ~new_new_n23299__;
  assign new_new_n23301__ = pi066 & ~new_new_n23300__;
  assign new_new_n23302__ = ~pi066 & new_new_n23300__;
  assign new_new_n23303__ = pi065 & po001;
  assign new_new_n23304__ = ~new_new_n22560__ & ~new_new_n23303__;
  assign new_new_n23305__ = pi001 & ~new_new_n22574__;
  assign new_new_n23306__ = pi064 & ~new_new_n23305__;
  assign new_new_n23307__ = ~new_new_n23304__ & ~new_new_n23306__;
  assign new_new_n23308__ = ~pi065 & po001;
  assign new_new_n23309__ = ~po002 & ~new_new_n23308__;
  assign new_new_n23310__ = po002 & new_new_n23308__;
  assign new_new_n23311__ = pi064 & ~new_new_n23289__;
  assign new_new_n23312__ = ~new_new_n23309__ & new_new_n23311__;
  assign new_new_n23313__ = ~new_new_n23310__ & new_new_n23312__;
  assign new_new_n23314__ = ~new_new_n23307__ & ~new_new_n23313__;
  assign new_new_n23315__ = pi002 & ~new_new_n23314__;
  assign new_new_n23316__ = ~new_new_n332__ & po001;
  assign new_new_n23317__ = ~new_new_n22560__ & ~new_new_n23316__;
  assign new_new_n23318__ = ~new_new_n22566__ & ~new_new_n22574__;
  assign new_new_n23319__ = pi001 & ~new_new_n23318__;
  assign new_new_n23320__ = ~new_new_n23298__ & new_new_n23319__;
  assign new_new_n23321__ = ~pi065 & ~po001;
  assign new_new_n23322__ = ~pi001 & ~new_new_n403__;
  assign new_new_n23323__ = new_new_n23318__ & new_new_n23322__;
  assign new_new_n23324__ = ~new_new_n23321__ & new_new_n23323__;
  assign new_new_n23325__ = ~new_new_n23317__ & ~new_new_n23324__;
  assign new_new_n23326__ = ~new_new_n23320__ & new_new_n23325__;
  assign new_new_n23327__ = ~pi002 & ~new_new_n23326__;
  assign new_new_n23328__ = ~new_new_n23315__ & ~new_new_n23327__;
  assign new_new_n23329__ = ~new_new_n23302__ & ~new_new_n23328__;
  assign new_new_n23330__ = ~new_new_n23301__ & ~new_new_n23329__;
  assign new_new_n23331__ = ~new_new_n23288__ & ~new_new_n23330__;
  assign new_new_n23332__ = ~new_new_n23287__ & ~new_new_n23331__;
  assign new_new_n23333__ = pi068 & ~new_new_n23332__;
  assign new_new_n23334__ = ~pi068 & new_new_n23332__;
  assign new_new_n23335__ = ~new_new_n22585__ & ~new_new_n22586__;
  assign new_new_n23336__ = po001 & new_new_n23335__;
  assign new_new_n23337__ = new_new_n22625__ & new_new_n23336__;
  assign new_new_n23338__ = ~new_new_n22625__ & ~new_new_n23336__;
  assign new_new_n23339__ = ~new_new_n23337__ & ~new_new_n23338__;
  assign new_new_n23340__ = ~new_new_n23334__ & ~new_new_n23339__;
  assign new_new_n23341__ = ~new_new_n23333__ & ~new_new_n23340__;
  assign new_new_n23342__ = ~new_new_n23281__ & ~new_new_n23341__;
  assign new_new_n23343__ = ~new_new_n23280__ & ~new_new_n23342__;
  assign new_new_n23344__ = ~new_new_n23272__ & ~new_new_n23343__;
  assign new_new_n23345__ = ~new_new_n23271__ & ~new_new_n23344__;
  assign new_new_n23346__ = ~new_new_n23263__ & ~new_new_n23345__;
  assign new_new_n23347__ = ~new_new_n23262__ & ~new_new_n23346__;
  assign new_new_n23348__ = ~new_new_n23254__ & ~new_new_n23347__;
  assign new_new_n23349__ = ~new_new_n23253__ & ~new_new_n23348__;
  assign new_new_n23350__ = ~new_new_n23245__ & new_new_n23349__;
  assign new_new_n23351__ = ~new_new_n23244__ & ~new_new_n23350__;
  assign new_new_n23352__ = ~new_new_n23236__ & ~new_new_n23351__;
  assign new_new_n23353__ = ~new_new_n23235__ & ~new_new_n23352__;
  assign new_new_n23354__ = ~new_new_n23227__ & ~new_new_n23353__;
  assign new_new_n23355__ = ~new_new_n23226__ & ~new_new_n23354__;
  assign new_new_n23356__ = ~new_new_n23218__ & ~new_new_n23355__;
  assign new_new_n23357__ = ~new_new_n23217__ & ~new_new_n23356__;
  assign new_new_n23358__ = ~new_new_n23209__ & ~new_new_n23357__;
  assign new_new_n23359__ = ~new_new_n23208__ & ~new_new_n23358__;
  assign new_new_n23360__ = ~new_new_n23200__ & ~new_new_n23359__;
  assign new_new_n23361__ = ~new_new_n23199__ & ~new_new_n23360__;
  assign new_new_n23362__ = ~new_new_n23191__ & ~new_new_n23361__;
  assign new_new_n23363__ = ~new_new_n23190__ & ~new_new_n23362__;
  assign new_new_n23364__ = ~new_new_n23182__ & ~new_new_n23363__;
  assign new_new_n23365__ = ~new_new_n23181__ & ~new_new_n23364__;
  assign new_new_n23366__ = ~new_new_n23173__ & ~new_new_n23365__;
  assign new_new_n23367__ = ~new_new_n23172__ & ~new_new_n23366__;
  assign new_new_n23368__ = ~new_new_n23164__ & ~new_new_n23367__;
  assign new_new_n23369__ = ~new_new_n23163__ & ~new_new_n23368__;
  assign new_new_n23370__ = ~new_new_n23155__ & new_new_n23369__;
  assign new_new_n23371__ = ~new_new_n23154__ & ~new_new_n23370__;
  assign new_new_n23372__ = ~new_new_n23146__ & ~new_new_n23371__;
  assign new_new_n23373__ = ~new_new_n23145__ & ~new_new_n23372__;
  assign new_new_n23374__ = ~new_new_n23137__ & new_new_n23373__;
  assign new_new_n23375__ = ~new_new_n23136__ & ~new_new_n23374__;
  assign new_new_n23376__ = ~new_new_n23128__ & new_new_n23375__;
  assign new_new_n23377__ = ~new_new_n23127__ & ~new_new_n23376__;
  assign new_new_n23378__ = ~new_new_n23119__ & ~new_new_n23377__;
  assign new_new_n23379__ = ~new_new_n23118__ & ~new_new_n23378__;
  assign new_new_n23380__ = ~new_new_n23110__ & ~new_new_n23379__;
  assign new_new_n23381__ = ~new_new_n23109__ & ~new_new_n23380__;
  assign new_new_n23382__ = ~new_new_n23101__ & new_new_n23381__;
  assign new_new_n23383__ = ~new_new_n23100__ & ~new_new_n23382__;
  assign new_new_n23384__ = ~new_new_n23092__ & new_new_n23383__;
  assign new_new_n23385__ = ~new_new_n23091__ & ~new_new_n23384__;
  assign new_new_n23386__ = ~new_new_n23083__ & new_new_n23385__;
  assign new_new_n23387__ = ~new_new_n23082__ & ~new_new_n23386__;
  assign new_new_n23388__ = ~new_new_n23074__ & ~new_new_n23387__;
  assign new_new_n23389__ = ~new_new_n23073__ & ~new_new_n23388__;
  assign new_new_n23390__ = ~new_new_n23065__ & ~new_new_n23389__;
  assign new_new_n23391__ = ~new_new_n23064__ & ~new_new_n23390__;
  assign new_new_n23392__ = ~new_new_n23056__ & ~new_new_n23391__;
  assign new_new_n23393__ = ~new_new_n23055__ & ~new_new_n23392__;
  assign new_new_n23394__ = ~new_new_n23047__ & ~new_new_n23393__;
  assign new_new_n23395__ = ~new_new_n23046__ & ~new_new_n23394__;
  assign new_new_n23396__ = ~new_new_n23038__ & ~new_new_n23395__;
  assign new_new_n23397__ = ~new_new_n23037__ & ~new_new_n23396__;
  assign new_new_n23398__ = ~new_new_n23029__ & ~new_new_n23397__;
  assign new_new_n23399__ = ~new_new_n23028__ & ~new_new_n23398__;
  assign new_new_n23400__ = ~new_new_n23020__ & ~new_new_n23399__;
  assign new_new_n23401__ = ~new_new_n23019__ & ~new_new_n23400__;
  assign new_new_n23402__ = ~new_new_n23011__ & ~new_new_n23401__;
  assign new_new_n23403__ = ~new_new_n23010__ & ~new_new_n23402__;
  assign new_new_n23404__ = ~new_new_n23002__ & new_new_n23403__;
  assign new_new_n23405__ = ~new_new_n23001__ & ~new_new_n23404__;
  assign new_new_n23406__ = ~new_new_n22993__ & new_new_n23405__;
  assign new_new_n23407__ = ~new_new_n22992__ & ~new_new_n23406__;
  assign new_new_n23408__ = ~new_new_n22984__ & ~new_new_n23407__;
  assign new_new_n23409__ = ~new_new_n22983__ & ~new_new_n23408__;
  assign new_new_n23410__ = ~new_new_n22975__ & ~new_new_n23409__;
  assign new_new_n23411__ = ~new_new_n22974__ & ~new_new_n23410__;
  assign new_new_n23412__ = ~new_new_n22966__ & ~new_new_n23411__;
  assign new_new_n23413__ = ~new_new_n22965__ & ~new_new_n23412__;
  assign new_new_n23414__ = ~new_new_n22957__ & ~new_new_n23413__;
  assign new_new_n23415__ = ~new_new_n22956__ & ~new_new_n23414__;
  assign new_new_n23416__ = ~new_new_n22948__ & ~new_new_n23415__;
  assign new_new_n23417__ = ~new_new_n22947__ & ~new_new_n23416__;
  assign new_new_n23418__ = ~new_new_n22939__ & ~new_new_n23417__;
  assign new_new_n23419__ = ~new_new_n22938__ & ~new_new_n23418__;
  assign new_new_n23420__ = ~new_new_n22930__ & ~new_new_n23419__;
  assign new_new_n23421__ = ~new_new_n22929__ & ~new_new_n23420__;
  assign new_new_n23422__ = ~new_new_n22921__ & ~new_new_n23421__;
  assign new_new_n23423__ = ~new_new_n22920__ & ~new_new_n23422__;
  assign new_new_n23424__ = ~new_new_n22912__ & ~new_new_n23423__;
  assign new_new_n23425__ = ~new_new_n22911__ & ~new_new_n23424__;
  assign new_new_n23426__ = ~new_new_n22903__ & new_new_n23425__;
  assign new_new_n23427__ = ~new_new_n22902__ & ~new_new_n23426__;
  assign new_new_n23428__ = ~new_new_n22894__ & ~new_new_n23427__;
  assign new_new_n23429__ = ~new_new_n22893__ & ~new_new_n23428__;
  assign new_new_n23430__ = ~new_new_n22885__ & new_new_n23429__;
  assign new_new_n23431__ = ~new_new_n22884__ & ~new_new_n23430__;
  assign new_new_n23432__ = ~new_new_n22876__ & ~new_new_n23431__;
  assign new_new_n23433__ = ~new_new_n22875__ & ~new_new_n23432__;
  assign new_new_n23434__ = ~new_new_n22867__ & new_new_n23433__;
  assign new_new_n23435__ = ~new_new_n22866__ & ~new_new_n23434__;
  assign new_new_n23436__ = ~new_new_n22858__ & ~new_new_n23435__;
  assign new_new_n23437__ = ~new_new_n22857__ & ~new_new_n23436__;
  assign new_new_n23438__ = ~new_new_n22849__ & ~new_new_n23437__;
  assign new_new_n23439__ = ~new_new_n22848__ & ~new_new_n23438__;
  assign new_new_n23440__ = ~new_new_n22840__ & new_new_n23439__;
  assign new_new_n23441__ = ~new_new_n22839__ & ~new_new_n23440__;
  assign new_new_n23442__ = ~new_new_n22831__ & ~new_new_n23441__;
  assign new_new_n23443__ = ~new_new_n22830__ & ~new_new_n23442__;
  assign new_new_n23444__ = ~new_new_n22822__ & new_new_n23443__;
  assign new_new_n23445__ = ~new_new_n22821__ & ~new_new_n23444__;
  assign new_new_n23446__ = ~new_new_n22813__ & new_new_n23445__;
  assign new_new_n23447__ = ~new_new_n22812__ & ~new_new_n23446__;
  assign new_new_n23448__ = ~new_new_n22804__ & ~new_new_n23447__;
  assign new_new_n23449__ = ~new_new_n22803__ & ~new_new_n23448__;
  assign new_new_n23450__ = ~new_new_n22795__ & ~new_new_n23449__;
  assign new_new_n23451__ = ~new_new_n22794__ & ~new_new_n23450__;
  assign new_new_n23452__ = ~new_new_n22786__ & ~new_new_n23451__;
  assign new_new_n23453__ = ~new_new_n22785__ & ~new_new_n23452__;
  assign new_new_n23454__ = ~new_new_n22777__ & new_new_n23453__;
  assign new_new_n23455__ = ~new_new_n22776__ & ~new_new_n23454__;
  assign new_new_n23456__ = ~new_new_n22759__ & ~new_new_n23455__;
  assign new_new_n23457__ = ~new_new_n22758__ & ~new_new_n23456__;
  assign new_new_n23458__ = ~new_new_n20019__ & new_new_n23457__;
  assign new_new_n23459__ = ~new_new_n22765__ & ~new_new_n22767__;
  assign new_new_n23460__ = ~pi127 & ~new_new_n23459__;
  assign new_new_n23461__ = new_new_n22753__ & new_new_n23460__;
  assign po000 = new_new_n23458__ | new_new_n23461__;
  assign po062 = new_new_n322__ & ~new_new_n333__;
  assign new_new_n23464__ = ~pi063 & pi064;
  assign new_new_n23465__ = ~pi065 & new_new_n319__;
  assign new_new_n23466__ = ~new_new_n23464__ & new_new_n23465__;
  assign po063 = new_new_n315__ & new_new_n23466__;
  assign new_new_n23468__ = pi064 & po000;
  assign new_new_n23469__ = ~pi000 & ~new_new_n23468__;
  assign new_new_n23470__ = pi000 & new_new_n23468__;
  assign po064 = ~new_new_n23469__ & ~new_new_n23470__;
  assign new_new_n23472__ = pi065 & po000;
  assign new_new_n23473__ = ~new_new_n23297__ & ~new_new_n23472__;
  assign new_new_n23474__ = ~new_new_n23468__ & new_new_n23473__;
  assign new_new_n23475__ = po001 & ~po000;
  assign new_new_n23476__ = ~new_new_n426__ & ~po001;
  assign new_new_n23477__ = ~pi000 & ~new_new_n23303__;
  assign new_new_n23478__ = ~new_new_n23476__ & new_new_n23477__;
  assign new_new_n23479__ = ~new_new_n23475__ & new_new_n23478__;
  assign new_new_n23480__ = po001 & ~new_new_n23472__;
  assign new_new_n23481__ = pi000 & ~new_new_n23298__;
  assign new_new_n23482__ = ~new_new_n23480__ & new_new_n23481__;
  assign new_new_n23483__ = ~new_new_n23474__ & ~new_new_n23479__;
  assign new_new_n23484__ = ~new_new_n23482__ & new_new_n23483__;
  assign new_new_n23485__ = pi001 & ~new_new_n23484__;
  assign new_new_n23486__ = new_new_n23321__ & po000;
  assign new_new_n23487__ = ~new_new_n23303__ & ~new_new_n23486__;
  assign new_new_n23488__ = ~pi000 & ~new_new_n23487__;
  assign new_new_n23489__ = ~new_new_n23475__ & ~new_new_n23488__;
  assign new_new_n23490__ = pi064 & ~new_new_n23489__;
  assign new_new_n23491__ = pi000 & ~new_new_n23303__;
  assign new_new_n23492__ = pi064 & ~new_new_n23491__;
  assign new_new_n23493__ = ~new_new_n23473__ & ~new_new_n23492__;
  assign new_new_n23494__ = ~new_new_n23490__ & ~new_new_n23493__;
  assign new_new_n23495__ = ~pi001 & ~new_new_n23494__;
  assign po065 = new_new_n23485__ | new_new_n23495__;
  assign new_new_n23497__ = ~new_new_n23301__ & ~new_new_n23302__;
  assign new_new_n23498__ = po000 & new_new_n23497__;
  assign new_new_n23499__ = new_new_n23328__ & ~new_new_n23498__;
  assign new_new_n23500__ = ~new_new_n23328__ & new_new_n23498__;
  assign po066 = new_new_n23499__ | new_new_n23500__;
  assign new_new_n23502__ = pi067 & ~new_new_n23330__;
  assign new_new_n23503__ = ~pi067 & new_new_n23330__;
  assign new_new_n23504__ = ~new_new_n23502__ & ~new_new_n23503__;
  assign new_new_n23505__ = po000 & new_new_n23504__;
  assign new_new_n23506__ = new_new_n23286__ & new_new_n23505__;
  assign new_new_n23507__ = ~new_new_n23286__ & ~new_new_n23505__;
  assign po067 = ~new_new_n23506__ & ~new_new_n23507__;
  assign new_new_n23509__ = ~new_new_n23333__ & ~new_new_n23334__;
  assign new_new_n23510__ = po000 & new_new_n23509__;
  assign new_new_n23511__ = new_new_n23339__ & ~new_new_n23510__;
  assign new_new_n23512__ = ~new_new_n23339__ & new_new_n23510__;
  assign po068 = new_new_n23511__ | new_new_n23512__;
  assign new_new_n23514__ = new_new_n23341__ & po000;
  assign new_new_n23515__ = ~pi069 & ~po000;
  assign new_new_n23516__ = ~new_new_n23514__ & ~new_new_n23515__;
  assign new_new_n23517__ = ~new_new_n23280__ & ~new_new_n23281__;
  assign new_new_n23518__ = ~new_new_n23516__ & ~new_new_n23517__;
  assign new_new_n23519__ = new_new_n23516__ & new_new_n23517__;
  assign po069 = new_new_n23518__ | new_new_n23519__;
  assign new_new_n23521__ = new_new_n23343__ & po000;
  assign new_new_n23522__ = ~pi070 & ~po000;
  assign new_new_n23523__ = ~new_new_n23521__ & ~new_new_n23522__;
  assign new_new_n23524__ = ~new_new_n23271__ & ~new_new_n23272__;
  assign new_new_n23525__ = ~new_new_n23523__ & ~new_new_n23524__;
  assign new_new_n23526__ = new_new_n23523__ & new_new_n23524__;
  assign po070 = new_new_n23525__ | new_new_n23526__;
  assign new_new_n23528__ = ~new_new_n23262__ & ~new_new_n23263__;
  assign new_new_n23529__ = ~pi071 & ~po000;
  assign new_new_n23530__ = new_new_n23345__ & po000;
  assign new_new_n23531__ = ~new_new_n23529__ & ~new_new_n23530__;
  assign new_new_n23532__ = new_new_n23528__ & ~new_new_n23531__;
  assign new_new_n23533__ = ~new_new_n23528__ & new_new_n23531__;
  assign po071 = ~new_new_n23532__ & ~new_new_n23533__;
  assign new_new_n23535__ = ~new_new_n23253__ & ~new_new_n23254__;
  assign new_new_n23536__ = ~pi072 & ~po000;
  assign new_new_n23537__ = new_new_n23347__ & po000;
  assign new_new_n23538__ = ~new_new_n23536__ & ~new_new_n23537__;
  assign new_new_n23539__ = new_new_n23535__ & ~new_new_n23538__;
  assign new_new_n23540__ = ~new_new_n23535__ & new_new_n23538__;
  assign po072 = ~new_new_n23539__ & ~new_new_n23540__;
  assign new_new_n23542__ = ~new_new_n23244__ & ~new_new_n23245__;
  assign new_new_n23543__ = new_new_n23349__ & po000;
  assign new_new_n23544__ = ~pi073 & ~po000;
  assign new_new_n23545__ = ~new_new_n23543__ & ~new_new_n23544__;
  assign new_new_n23546__ = ~new_new_n23542__ & ~new_new_n23545__;
  assign new_new_n23547__ = new_new_n23542__ & new_new_n23545__;
  assign po073 = new_new_n23546__ | new_new_n23547__;
  assign new_new_n23549__ = ~pi074 & ~new_new_n23351__;
  assign new_new_n23550__ = pi074 & new_new_n23351__;
  assign new_new_n23551__ = ~new_new_n23549__ & ~new_new_n23550__;
  assign new_new_n23552__ = po000 & new_new_n23551__;
  assign new_new_n23553__ = ~new_new_n23234__ & new_new_n23552__;
  assign new_new_n23554__ = new_new_n23234__ & ~new_new_n23552__;
  assign po074 = ~new_new_n23553__ & ~new_new_n23554__;
  assign new_new_n23556__ = ~new_new_n23226__ & ~new_new_n23227__;
  assign new_new_n23557__ = ~pi075 & ~po000;
  assign new_new_n23558__ = ~new_new_n23353__ & po000;
  assign new_new_n23559__ = ~new_new_n23557__ & ~new_new_n23558__;
  assign new_new_n23560__ = new_new_n23556__ & ~new_new_n23559__;
  assign new_new_n23561__ = ~new_new_n23556__ & new_new_n23559__;
  assign po075 = ~new_new_n23560__ & ~new_new_n23561__;
  assign new_new_n23563__ = ~new_new_n23217__ & ~new_new_n23218__;
  assign new_new_n23564__ = ~pi076 & ~po000;
  assign new_new_n23565__ = ~new_new_n23355__ & po000;
  assign new_new_n23566__ = ~new_new_n23564__ & ~new_new_n23565__;
  assign new_new_n23567__ = new_new_n23563__ & ~new_new_n23566__;
  assign new_new_n23568__ = ~new_new_n23563__ & new_new_n23566__;
  assign po076 = ~new_new_n23567__ & ~new_new_n23568__;
  assign new_new_n23570__ = ~pi077 & ~new_new_n23357__;
  assign new_new_n23571__ = pi077 & new_new_n23357__;
  assign new_new_n23572__ = ~new_new_n23570__ & ~new_new_n23571__;
  assign new_new_n23573__ = po000 & new_new_n23572__;
  assign new_new_n23574__ = new_new_n23207__ & new_new_n23573__;
  assign new_new_n23575__ = ~new_new_n23207__ & ~new_new_n23573__;
  assign po077 = new_new_n23574__ | new_new_n23575__;
  assign new_new_n23577__ = ~pi078 & ~new_new_n23359__;
  assign new_new_n23578__ = pi078 & new_new_n23359__;
  assign new_new_n23579__ = ~new_new_n23577__ & ~new_new_n23578__;
  assign new_new_n23580__ = po000 & new_new_n23579__;
  assign new_new_n23581__ = new_new_n23198__ & new_new_n23580__;
  assign new_new_n23582__ = ~new_new_n23198__ & ~new_new_n23580__;
  assign po078 = new_new_n23581__ | new_new_n23582__;
  assign new_new_n23584__ = ~new_new_n23190__ & ~new_new_n23191__;
  assign new_new_n23585__ = ~pi079 & ~po000;
  assign new_new_n23586__ = ~new_new_n23361__ & po000;
  assign new_new_n23587__ = ~new_new_n23585__ & ~new_new_n23586__;
  assign new_new_n23588__ = new_new_n23584__ & ~new_new_n23587__;
  assign new_new_n23589__ = ~new_new_n23584__ & new_new_n23587__;
  assign po079 = ~new_new_n23588__ & ~new_new_n23589__;
  assign new_new_n23591__ = ~pi080 & ~new_new_n23363__;
  assign new_new_n23592__ = pi080 & new_new_n23363__;
  assign new_new_n23593__ = ~new_new_n23591__ & ~new_new_n23592__;
  assign new_new_n23594__ = po000 & new_new_n23593__;
  assign new_new_n23595__ = new_new_n23180__ & new_new_n23594__;
  assign new_new_n23596__ = ~new_new_n23180__ & ~new_new_n23594__;
  assign po080 = new_new_n23595__ | new_new_n23596__;
  assign new_new_n23598__ = ~new_new_n23172__ & ~new_new_n23173__;
  assign new_new_n23599__ = ~pi081 & ~po000;
  assign new_new_n23600__ = ~new_new_n23365__ & po000;
  assign new_new_n23601__ = ~new_new_n23599__ & ~new_new_n23600__;
  assign new_new_n23602__ = new_new_n23598__ & ~new_new_n23601__;
  assign new_new_n23603__ = ~new_new_n23598__ & new_new_n23601__;
  assign po081 = ~new_new_n23602__ & ~new_new_n23603__;
  assign new_new_n23605__ = ~pi082 & ~new_new_n23367__;
  assign new_new_n23606__ = pi082 & new_new_n23367__;
  assign new_new_n23607__ = ~new_new_n23605__ & ~new_new_n23606__;
  assign new_new_n23608__ = po000 & new_new_n23607__;
  assign new_new_n23609__ = ~new_new_n23162__ & ~new_new_n23608__;
  assign new_new_n23610__ = new_new_n23162__ & new_new_n23608__;
  assign po082 = new_new_n23609__ | new_new_n23610__;
  assign new_new_n23612__ = ~new_new_n23154__ & ~new_new_n23155__;
  assign new_new_n23613__ = ~pi083 & ~po000;
  assign new_new_n23614__ = ~new_new_n23369__ & po000;
  assign new_new_n23615__ = ~new_new_n23613__ & ~new_new_n23614__;
  assign new_new_n23616__ = new_new_n23612__ & ~new_new_n23615__;
  assign new_new_n23617__ = ~new_new_n23612__ & new_new_n23615__;
  assign po083 = ~new_new_n23616__ & ~new_new_n23617__;
  assign new_new_n23619__ = pi084 & ~new_new_n23371__;
  assign new_new_n23620__ = ~pi084 & new_new_n23371__;
  assign new_new_n23621__ = ~new_new_n23619__ & ~new_new_n23620__;
  assign new_new_n23622__ = po000 & new_new_n23621__;
  assign new_new_n23623__ = new_new_n23144__ & ~new_new_n23622__;
  assign new_new_n23624__ = ~new_new_n23144__ & new_new_n23622__;
  assign po084 = new_new_n23623__ | new_new_n23624__;
  assign new_new_n23626__ = ~new_new_n23136__ & ~new_new_n23137__;
  assign new_new_n23627__ = new_new_n23373__ & po000;
  assign new_new_n23628__ = ~pi085 & ~po000;
  assign new_new_n23629__ = ~new_new_n23627__ & ~new_new_n23628__;
  assign new_new_n23630__ = ~new_new_n23626__ & ~new_new_n23629__;
  assign new_new_n23631__ = new_new_n23626__ & new_new_n23629__;
  assign po085 = new_new_n23630__ | new_new_n23631__;
  assign new_new_n23633__ = ~new_new_n23127__ & ~new_new_n23128__;
  assign new_new_n23634__ = ~pi086 & ~po000;
  assign new_new_n23635__ = ~new_new_n23375__ & po000;
  assign new_new_n23636__ = ~new_new_n23634__ & ~new_new_n23635__;
  assign new_new_n23637__ = new_new_n23633__ & ~new_new_n23636__;
  assign new_new_n23638__ = ~new_new_n23633__ & new_new_n23636__;
  assign po086 = ~new_new_n23637__ & ~new_new_n23638__;
  assign new_new_n23640__ = ~new_new_n23118__ & ~new_new_n23119__;
  assign new_new_n23641__ = new_new_n23377__ & po000;
  assign new_new_n23642__ = ~pi087 & ~po000;
  assign new_new_n23643__ = ~new_new_n23641__ & ~new_new_n23642__;
  assign new_new_n23644__ = new_new_n23640__ & new_new_n23643__;
  assign new_new_n23645__ = ~new_new_n23640__ & ~new_new_n23643__;
  assign po087 = new_new_n23644__ | new_new_n23645__;
  assign new_new_n23647__ = ~new_new_n23109__ & ~new_new_n23110__;
  assign new_new_n23648__ = ~pi088 & ~po000;
  assign new_new_n23649__ = new_new_n23379__ & po000;
  assign new_new_n23650__ = ~new_new_n23648__ & ~new_new_n23649__;
  assign new_new_n23651__ = new_new_n23647__ & ~new_new_n23650__;
  assign new_new_n23652__ = ~new_new_n23647__ & new_new_n23650__;
  assign po088 = ~new_new_n23651__ & ~new_new_n23652__;
  assign new_new_n23654__ = ~new_new_n23100__ & ~new_new_n23101__;
  assign new_new_n23655__ = ~pi089 & ~po000;
  assign new_new_n23656__ = new_new_n23381__ & po000;
  assign new_new_n23657__ = ~new_new_n23655__ & ~new_new_n23656__;
  assign new_new_n23658__ = new_new_n23654__ & ~new_new_n23657__;
  assign new_new_n23659__ = ~new_new_n23654__ & new_new_n23657__;
  assign po089 = ~new_new_n23658__ & ~new_new_n23659__;
  assign new_new_n23661__ = ~new_new_n23091__ & ~new_new_n23092__;
  assign new_new_n23662__ = ~pi090 & ~po000;
  assign new_new_n23663__ = ~new_new_n23383__ & po000;
  assign new_new_n23664__ = ~new_new_n23662__ & ~new_new_n23663__;
  assign new_new_n23665__ = new_new_n23661__ & ~new_new_n23664__;
  assign new_new_n23666__ = ~new_new_n23661__ & new_new_n23664__;
  assign po090 = ~new_new_n23665__ & ~new_new_n23666__;
  assign new_new_n23668__ = ~new_new_n23082__ & ~new_new_n23083__;
  assign new_new_n23669__ = ~pi091 & ~po000;
  assign new_new_n23670__ = new_new_n23385__ & po000;
  assign new_new_n23671__ = ~new_new_n23669__ & ~new_new_n23670__;
  assign new_new_n23672__ = new_new_n23668__ & ~new_new_n23671__;
  assign new_new_n23673__ = ~new_new_n23668__ & new_new_n23671__;
  assign po091 = ~new_new_n23672__ & ~new_new_n23673__;
  assign new_new_n23675__ = ~new_new_n23073__ & ~new_new_n23074__;
  assign new_new_n23676__ = ~pi092 & ~po000;
  assign new_new_n23677__ = ~new_new_n23387__ & po000;
  assign new_new_n23678__ = ~new_new_n23676__ & ~new_new_n23677__;
  assign new_new_n23679__ = new_new_n23675__ & ~new_new_n23678__;
  assign new_new_n23680__ = ~new_new_n23675__ & new_new_n23678__;
  assign po092 = ~new_new_n23679__ & ~new_new_n23680__;
  assign new_new_n23682__ = ~new_new_n23064__ & ~new_new_n23065__;
  assign new_new_n23683__ = ~pi093 & ~po000;
  assign new_new_n23684__ = ~new_new_n23389__ & po000;
  assign new_new_n23685__ = ~new_new_n23683__ & ~new_new_n23684__;
  assign new_new_n23686__ = new_new_n23682__ & ~new_new_n23685__;
  assign new_new_n23687__ = ~new_new_n23682__ & new_new_n23685__;
  assign po093 = ~new_new_n23686__ & ~new_new_n23687__;
  assign new_new_n23689__ = ~pi094 & ~new_new_n23391__;
  assign new_new_n23690__ = pi094 & new_new_n23391__;
  assign new_new_n23691__ = ~new_new_n23689__ & ~new_new_n23690__;
  assign new_new_n23692__ = po000 & new_new_n23691__;
  assign new_new_n23693__ = new_new_n23054__ & new_new_n23692__;
  assign new_new_n23694__ = ~new_new_n23054__ & ~new_new_n23692__;
  assign po094 = new_new_n23693__ | new_new_n23694__;
  assign new_new_n23696__ = ~new_new_n23046__ & ~new_new_n23047__;
  assign new_new_n23697__ = ~pi095 & ~po000;
  assign new_new_n23698__ = ~new_new_n23393__ & po000;
  assign new_new_n23699__ = ~new_new_n23697__ & ~new_new_n23698__;
  assign new_new_n23700__ = new_new_n23696__ & ~new_new_n23699__;
  assign new_new_n23701__ = ~new_new_n23696__ & new_new_n23699__;
  assign po095 = ~new_new_n23700__ & ~new_new_n23701__;
  assign new_new_n23703__ = ~new_new_n23037__ & ~new_new_n23038__;
  assign new_new_n23704__ = ~pi096 & ~po000;
  assign new_new_n23705__ = ~new_new_n23395__ & po000;
  assign new_new_n23706__ = ~new_new_n23704__ & ~new_new_n23705__;
  assign new_new_n23707__ = new_new_n23703__ & ~new_new_n23706__;
  assign new_new_n23708__ = ~new_new_n23703__ & new_new_n23706__;
  assign po096 = ~new_new_n23707__ & ~new_new_n23708__;
  assign new_new_n23710__ = ~pi097 & ~new_new_n23397__;
  assign new_new_n23711__ = pi097 & new_new_n23397__;
  assign new_new_n23712__ = ~new_new_n23710__ & ~new_new_n23711__;
  assign new_new_n23713__ = po000 & new_new_n23712__;
  assign new_new_n23714__ = new_new_n23027__ & new_new_n23713__;
  assign new_new_n23715__ = ~new_new_n23027__ & ~new_new_n23713__;
  assign po097 = new_new_n23714__ | new_new_n23715__;
  assign new_new_n23717__ = ~pi098 & ~new_new_n23399__;
  assign new_new_n23718__ = pi098 & new_new_n23399__;
  assign new_new_n23719__ = ~new_new_n23717__ & ~new_new_n23718__;
  assign new_new_n23720__ = po000 & new_new_n23719__;
  assign new_new_n23721__ = ~new_new_n23018__ & ~new_new_n23720__;
  assign new_new_n23722__ = new_new_n23018__ & new_new_n23720__;
  assign po098 = new_new_n23721__ | new_new_n23722__;
  assign new_new_n23724__ = ~new_new_n23010__ & ~new_new_n23011__;
  assign new_new_n23725__ = ~pi099 & ~po000;
  assign new_new_n23726__ = ~new_new_n23401__ & po000;
  assign new_new_n23727__ = ~new_new_n23725__ & ~new_new_n23726__;
  assign new_new_n23728__ = new_new_n23724__ & ~new_new_n23727__;
  assign new_new_n23729__ = ~new_new_n23724__ & new_new_n23727__;
  assign po099 = ~new_new_n23728__ & ~new_new_n23729__;
  assign new_new_n23731__ = ~new_new_n23001__ & ~new_new_n23002__;
  assign new_new_n23732__ = ~pi100 & ~po000;
  assign new_new_n23733__ = ~new_new_n23403__ & po000;
  assign new_new_n23734__ = ~new_new_n23732__ & ~new_new_n23733__;
  assign new_new_n23735__ = new_new_n23731__ & ~new_new_n23734__;
  assign new_new_n23736__ = ~new_new_n23731__ & new_new_n23734__;
  assign po100 = ~new_new_n23735__ & ~new_new_n23736__;
  assign new_new_n23738__ = new_new_n23405__ & po000;
  assign new_new_n23739__ = ~pi101 & ~po000;
  assign new_new_n23740__ = ~new_new_n23738__ & ~new_new_n23739__;
  assign new_new_n23741__ = ~new_new_n22992__ & ~new_new_n22993__;
  assign new_new_n23742__ = ~new_new_n23740__ & ~new_new_n23741__;
  assign new_new_n23743__ = new_new_n23740__ & new_new_n23741__;
  assign po101 = new_new_n23742__ | new_new_n23743__;
  assign new_new_n23745__ = ~pi102 & ~new_new_n23407__;
  assign new_new_n23746__ = pi102 & new_new_n23407__;
  assign new_new_n23747__ = ~new_new_n23745__ & ~new_new_n23746__;
  assign new_new_n23748__ = po000 & new_new_n23747__;
  assign new_new_n23749__ = ~new_new_n22982__ & ~new_new_n23748__;
  assign new_new_n23750__ = new_new_n22982__ & new_new_n23748__;
  assign po102 = new_new_n23749__ | new_new_n23750__;
  assign new_new_n23752__ = ~new_new_n22974__ & ~new_new_n22975__;
  assign new_new_n23753__ = ~new_new_n23409__ & po000;
  assign new_new_n23754__ = ~pi103 & ~po000;
  assign new_new_n23755__ = ~new_new_n23753__ & ~new_new_n23754__;
  assign new_new_n23756__ = ~new_new_n23752__ & ~new_new_n23755__;
  assign new_new_n23757__ = new_new_n23752__ & new_new_n23755__;
  assign po103 = new_new_n23756__ | new_new_n23757__;
  assign new_new_n23759__ = new_new_n23411__ & po000;
  assign new_new_n23760__ = pi104 & ~po000;
  assign new_new_n23761__ = ~new_new_n23759__ & ~new_new_n23760__;
  assign new_new_n23762__ = ~new_new_n22965__ & ~new_new_n22966__;
  assign new_new_n23763__ = ~new_new_n23761__ & ~new_new_n23762__;
  assign new_new_n23764__ = new_new_n23761__ & new_new_n23762__;
  assign po104 = ~new_new_n23763__ & ~new_new_n23764__;
  assign new_new_n23766__ = new_new_n23413__ & po000;
  assign new_new_n23767__ = pi105 & ~po000;
  assign new_new_n23768__ = ~new_new_n23766__ & ~new_new_n23767__;
  assign new_new_n23769__ = ~new_new_n22956__ & ~new_new_n22957__;
  assign new_new_n23770__ = ~new_new_n23768__ & ~new_new_n23769__;
  assign new_new_n23771__ = new_new_n23768__ & new_new_n23769__;
  assign po105 = ~new_new_n23770__ & ~new_new_n23771__;
  assign new_new_n23773__ = new_new_n23415__ & po000;
  assign new_new_n23774__ = pi106 & ~po000;
  assign new_new_n23775__ = ~new_new_n23773__ & ~new_new_n23774__;
  assign new_new_n23776__ = ~new_new_n22947__ & ~new_new_n22948__;
  assign new_new_n23777__ = ~new_new_n23775__ & ~new_new_n23776__;
  assign new_new_n23778__ = new_new_n23775__ & new_new_n23776__;
  assign po106 = ~new_new_n23777__ & ~new_new_n23778__;
  assign new_new_n23780__ = ~new_new_n22938__ & ~new_new_n22939__;
  assign new_new_n23781__ = ~new_new_n23417__ & po000;
  assign new_new_n23782__ = ~pi107 & ~po000;
  assign new_new_n23783__ = ~new_new_n23781__ & ~new_new_n23782__;
  assign new_new_n23784__ = ~new_new_n23780__ & ~new_new_n23783__;
  assign new_new_n23785__ = new_new_n23780__ & new_new_n23783__;
  assign po107 = new_new_n23784__ | new_new_n23785__;
  assign new_new_n23787__ = new_new_n23419__ & po000;
  assign new_new_n23788__ = pi108 & ~po000;
  assign new_new_n23789__ = ~new_new_n23787__ & ~new_new_n23788__;
  assign new_new_n23790__ = ~new_new_n22929__ & ~new_new_n22930__;
  assign new_new_n23791__ = ~new_new_n23789__ & ~new_new_n23790__;
  assign new_new_n23792__ = new_new_n23789__ & new_new_n23790__;
  assign po108 = ~new_new_n23791__ & ~new_new_n23792__;
  assign new_new_n23794__ = ~new_new_n22920__ & ~new_new_n22921__;
  assign new_new_n23795__ = ~new_new_n23421__ & po000;
  assign new_new_n23796__ = ~pi109 & ~po000;
  assign new_new_n23797__ = ~new_new_n23795__ & ~new_new_n23796__;
  assign new_new_n23798__ = ~new_new_n23794__ & ~new_new_n23797__;
  assign new_new_n23799__ = new_new_n23794__ & new_new_n23797__;
  assign po109 = new_new_n23798__ | new_new_n23799__;
  assign new_new_n23801__ = ~new_new_n22911__ & ~new_new_n22912__;
  assign new_new_n23802__ = ~new_new_n23423__ & po000;
  assign new_new_n23803__ = ~pi110 & ~po000;
  assign new_new_n23804__ = ~new_new_n23802__ & ~new_new_n23803__;
  assign new_new_n23805__ = ~new_new_n23801__ & ~new_new_n23804__;
  assign new_new_n23806__ = new_new_n23801__ & new_new_n23804__;
  assign po110 = new_new_n23805__ | new_new_n23806__;
  assign new_new_n23808__ = ~new_new_n22902__ & ~new_new_n22903__;
  assign new_new_n23809__ = ~pi111 & ~po000;
  assign new_new_n23810__ = ~new_new_n23425__ & po000;
  assign new_new_n23811__ = ~new_new_n23809__ & ~new_new_n23810__;
  assign new_new_n23812__ = new_new_n23808__ & ~new_new_n23811__;
  assign new_new_n23813__ = ~new_new_n23808__ & new_new_n23811__;
  assign po111 = ~new_new_n23812__ & ~new_new_n23813__;
  assign new_new_n23815__ = ~new_new_n22893__ & ~new_new_n22894__;
  assign new_new_n23816__ = ~pi112 & ~po000;
  assign new_new_n23817__ = new_new_n23427__ & po000;
  assign new_new_n23818__ = ~new_new_n23816__ & ~new_new_n23817__;
  assign new_new_n23819__ = new_new_n23815__ & ~new_new_n23818__;
  assign new_new_n23820__ = ~new_new_n23815__ & new_new_n23818__;
  assign po112 = ~new_new_n23819__ & ~new_new_n23820__;
  assign new_new_n23822__ = ~new_new_n22884__ & ~new_new_n22885__;
  assign new_new_n23823__ = new_new_n23429__ & po000;
  assign new_new_n23824__ = ~pi113 & ~po000;
  assign new_new_n23825__ = ~new_new_n23823__ & ~new_new_n23824__;
  assign new_new_n23826__ = ~new_new_n23822__ & ~new_new_n23825__;
  assign new_new_n23827__ = new_new_n23822__ & new_new_n23825__;
  assign po113 = new_new_n23826__ | new_new_n23827__;
  assign new_new_n23829__ = ~pi114 & ~new_new_n23431__;
  assign new_new_n23830__ = pi114 & new_new_n23431__;
  assign new_new_n23831__ = ~new_new_n23829__ & ~new_new_n23830__;
  assign new_new_n23832__ = po000 & new_new_n23831__;
  assign new_new_n23833__ = new_new_n22874__ & new_new_n23832__;
  assign new_new_n23834__ = ~new_new_n22874__ & ~new_new_n23832__;
  assign po114 = new_new_n23833__ | new_new_n23834__;
  assign new_new_n23836__ = ~new_new_n22866__ & ~new_new_n22867__;
  assign new_new_n23837__ = ~pi115 & ~po000;
  assign new_new_n23838__ = ~new_new_n23433__ & po000;
  assign new_new_n23839__ = ~new_new_n23837__ & ~new_new_n23838__;
  assign new_new_n23840__ = new_new_n23836__ & ~new_new_n23839__;
  assign new_new_n23841__ = ~new_new_n23836__ & new_new_n23839__;
  assign po115 = ~new_new_n23840__ & ~new_new_n23841__;
  assign new_new_n23843__ = ~new_new_n22857__ & ~new_new_n22858__;
  assign new_new_n23844__ = new_new_n23435__ & po000;
  assign new_new_n23845__ = ~pi116 & ~po000;
  assign new_new_n23846__ = ~new_new_n23844__ & ~new_new_n23845__;
  assign new_new_n23847__ = ~new_new_n23843__ & ~new_new_n23846__;
  assign new_new_n23848__ = new_new_n23843__ & new_new_n23846__;
  assign po116 = new_new_n23847__ | new_new_n23848__;
  assign new_new_n23850__ = ~new_new_n22848__ & ~new_new_n22849__;
  assign new_new_n23851__ = ~pi117 & ~po000;
  assign new_new_n23852__ = new_new_n23437__ & po000;
  assign new_new_n23853__ = ~new_new_n23851__ & ~new_new_n23852__;
  assign new_new_n23854__ = new_new_n23850__ & ~new_new_n23853__;
  assign new_new_n23855__ = ~new_new_n23850__ & new_new_n23853__;
  assign po117 = ~new_new_n23854__ & ~new_new_n23855__;
  assign new_new_n23857__ = new_new_n23439__ & po000;
  assign new_new_n23858__ = ~pi118 & ~po000;
  assign new_new_n23859__ = ~new_new_n23857__ & ~new_new_n23858__;
  assign new_new_n23860__ = ~new_new_n22839__ & ~new_new_n22840__;
  assign new_new_n23861__ = ~new_new_n23859__ & ~new_new_n23860__;
  assign new_new_n23862__ = new_new_n23859__ & new_new_n23860__;
  assign po118 = new_new_n23861__ | new_new_n23862__;
  assign new_new_n23864__ = ~new_new_n22830__ & ~new_new_n22831__;
  assign new_new_n23865__ = ~new_new_n23441__ & po000;
  assign new_new_n23866__ = ~pi119 & ~po000;
  assign new_new_n23867__ = ~new_new_n23865__ & ~new_new_n23866__;
  assign new_new_n23868__ = ~new_new_n23864__ & ~new_new_n23867__;
  assign new_new_n23869__ = new_new_n23864__ & new_new_n23867__;
  assign po119 = new_new_n23868__ | new_new_n23869__;
  assign new_new_n23871__ = ~new_new_n22821__ & ~new_new_n22822__;
  assign new_new_n23872__ = ~pi120 & ~po000;
  assign new_new_n23873__ = ~new_new_n23443__ & po000;
  assign new_new_n23874__ = ~new_new_n23872__ & ~new_new_n23873__;
  assign new_new_n23875__ = new_new_n23871__ & ~new_new_n23874__;
  assign new_new_n23876__ = ~new_new_n23871__ & new_new_n23874__;
  assign po120 = ~new_new_n23875__ & ~new_new_n23876__;
  assign new_new_n23878__ = ~new_new_n22812__ & ~new_new_n22813__;
  assign new_new_n23879__ = ~pi121 & ~po000;
  assign new_new_n23880__ = new_new_n23445__ & po000;
  assign new_new_n23881__ = ~new_new_n23879__ & ~new_new_n23880__;
  assign new_new_n23882__ = new_new_n23878__ & ~new_new_n23881__;
  assign new_new_n23883__ = ~new_new_n23878__ & new_new_n23881__;
  assign po121 = ~new_new_n23882__ & ~new_new_n23883__;
  assign new_new_n23885__ = ~new_new_n22803__ & ~new_new_n22804__;
  assign new_new_n23886__ = ~pi122 & ~po000;
  assign new_new_n23887__ = ~new_new_n23447__ & po000;
  assign new_new_n23888__ = ~new_new_n23886__ & ~new_new_n23887__;
  assign new_new_n23889__ = new_new_n23885__ & ~new_new_n23888__;
  assign new_new_n23890__ = ~new_new_n23885__ & new_new_n23888__;
  assign po122 = ~new_new_n23889__ & ~new_new_n23890__;
  assign new_new_n23892__ = ~pi123 & ~new_new_n23449__;
  assign new_new_n23893__ = pi123 & new_new_n23449__;
  assign new_new_n23894__ = ~new_new_n23892__ & ~new_new_n23893__;
  assign new_new_n23895__ = po000 & new_new_n23894__;
  assign new_new_n23896__ = new_new_n22793__ & new_new_n23895__;
  assign new_new_n23897__ = ~new_new_n22793__ & ~new_new_n23895__;
  assign po123 = new_new_n23896__ | new_new_n23897__;
  assign new_new_n23899__ = ~new_new_n22785__ & ~new_new_n22786__;
  assign new_new_n23900__ = ~pi124 & ~po000;
  assign new_new_n23901__ = ~new_new_n23451__ & po000;
  assign new_new_n23902__ = ~new_new_n23900__ & ~new_new_n23901__;
  assign new_new_n23903__ = new_new_n23899__ & ~new_new_n23902__;
  assign new_new_n23904__ = ~new_new_n23899__ & new_new_n23902__;
  assign po124 = ~new_new_n23903__ & ~new_new_n23904__;
  assign new_new_n23906__ = ~new_new_n22776__ & ~new_new_n22777__;
  assign new_new_n23907__ = ~pi125 & ~po000;
  assign new_new_n23908__ = ~new_new_n23453__ & po000;
  assign new_new_n23909__ = ~new_new_n23907__ & ~new_new_n23908__;
  assign new_new_n23910__ = new_new_n23906__ & ~new_new_n23909__;
  assign new_new_n23911__ = ~new_new_n23906__ & new_new_n23909__;
  assign po125 = ~new_new_n23910__ & ~new_new_n23911__;
  assign new_new_n23913__ = ~new_new_n22758__ & ~new_new_n22759__;
  assign new_new_n23914__ = ~pi126 & ~po000;
  assign new_new_n23915__ = new_new_n23455__ & po000;
  assign new_new_n23916__ = ~new_new_n23914__ & ~new_new_n23915__;
  assign new_new_n23917__ = new_new_n23913__ & ~new_new_n23916__;
  assign new_new_n23918__ = ~new_new_n23913__ & new_new_n23916__;
  assign po126 = ~new_new_n23917__ & ~new_new_n23918__;
  assign new_new_n23920__ = ~pi127 & ~new_new_n23457__;
  assign new_new_n23921__ = new_new_n23457__ & ~new_new_n23460__;
  assign new_new_n23922__ = new_new_n22753__ & ~new_new_n23920__;
  assign po127 = ~new_new_n23921__ & new_new_n23922__;
endmodule


