// Benchmark "max" written by ABC on Wed Jul 13 18:49:13 2022

module max ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279,
    pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289,
    pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299,
    pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309,
    pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319,
    pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329,
    pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339,
    pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349,
    pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359,
    pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369,
    pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378, pi379,
    pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388, pi389,
    pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398, pi399,
    pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408, pi409,
    pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418, pi419,
    pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429,
    pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439,
    pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449,
    pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458, pi459,
    pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468, pi469,
    pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478, pi479,
    pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488, pi489,
    pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498, pi499,
    pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508, pi509,
    pi510, pi511,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258,
    pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288,
    pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298,
    pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308,
    pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318,
    pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328,
    pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338,
    pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348,
    pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358,
    pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368,
    pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378,
    pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388,
    pi389, pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398,
    pi399, pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408,
    pi409, pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418,
    pi419, pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428,
    pi429, pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438,
    pi439, pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448,
    pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458,
    pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468,
    pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478,
    pi479, pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488,
    pi489, pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498,
    pi499, pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508,
    pi509, pi510, pi511;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129;
  wire new_new_n643__, new_new_n644__, new_new_n645__, new_new_n646__,
    new_new_n647__, new_new_n648__, new_new_n649__, new_new_n650__,
    new_new_n651__, new_new_n652__, new_new_n653__, new_new_n654__,
    new_new_n655__, new_new_n656__, new_new_n657__, new_new_n658__,
    new_new_n659__, new_new_n660__, new_new_n661__, new_new_n662__,
    new_new_n663__, new_new_n664__, new_new_n665__, new_new_n666__,
    new_new_n667__, new_new_n668__, new_new_n669__, new_new_n670__,
    new_new_n671__, new_new_n672__, new_new_n673__, new_new_n674__,
    new_new_n675__, new_new_n676__, new_new_n677__, new_new_n678__,
    new_new_n679__, new_new_n680__, new_new_n681__, new_new_n682__,
    new_new_n683__, new_new_n684__, new_new_n685__, new_new_n686__,
    new_new_n687__, new_new_n688__, new_new_n689__, new_new_n690__,
    new_new_n691__, new_new_n692__, new_new_n693__, new_new_n694__,
    new_new_n695__, new_new_n696__, new_new_n697__, new_new_n698__,
    new_new_n699__, new_new_n700__, new_new_n701__, new_new_n702__,
    new_new_n703__, new_new_n704__, new_new_n705__, new_new_n706__,
    new_new_n707__, new_new_n708__, new_new_n709__, new_new_n710__,
    new_new_n711__, new_new_n712__, new_new_n713__, new_new_n714__,
    new_new_n715__, new_new_n716__, new_new_n717__, new_new_n718__,
    new_new_n719__, new_new_n720__, new_new_n721__, new_new_n722__,
    new_new_n723__, new_new_n724__, new_new_n725__, new_new_n726__,
    new_new_n727__, new_new_n728__, new_new_n729__, new_new_n730__,
    new_new_n731__, new_new_n732__, new_new_n733__, new_new_n734__,
    new_new_n735__, new_new_n736__, new_new_n737__, new_new_n738__,
    new_new_n739__, new_new_n740__, new_new_n741__, new_new_n742__,
    new_new_n743__, new_new_n744__, new_new_n745__, new_new_n746__,
    new_new_n747__, new_new_n748__, new_new_n749__, new_new_n750__,
    new_new_n751__, new_new_n752__, new_new_n753__, new_new_n754__,
    new_new_n755__, new_new_n756__, new_new_n757__, new_new_n758__,
    new_new_n759__, new_new_n760__, new_new_n761__, new_new_n762__,
    new_new_n763__, new_new_n764__, new_new_n765__, new_new_n766__,
    new_new_n767__, new_new_n768__, new_new_n769__, new_new_n770__,
    new_new_n771__, new_new_n772__, new_new_n773__, new_new_n774__,
    new_new_n775__, new_new_n776__, new_new_n777__, new_new_n778__,
    new_new_n779__, new_new_n780__, new_new_n781__, new_new_n782__,
    new_new_n783__, new_new_n784__, new_new_n785__, new_new_n786__,
    new_new_n787__, new_new_n788__, new_new_n789__, new_new_n790__,
    new_new_n791__, new_new_n792__, new_new_n793__, new_new_n794__,
    new_new_n795__, new_new_n796__, new_new_n797__, new_new_n798__,
    new_new_n799__, new_new_n800__, new_new_n801__, new_new_n802__,
    new_new_n803__, new_new_n804__, new_new_n805__, new_new_n806__,
    new_new_n807__, new_new_n808__, new_new_n809__, new_new_n810__,
    new_new_n811__, new_new_n812__, new_new_n813__, new_new_n814__,
    new_new_n815__, new_new_n816__, new_new_n817__, new_new_n818__,
    new_new_n819__, new_new_n820__, new_new_n821__, new_new_n822__,
    new_new_n823__, new_new_n824__, new_new_n825__, new_new_n826__,
    new_new_n827__, new_new_n828__, new_new_n829__, new_new_n830__,
    new_new_n831__, new_new_n832__, new_new_n833__, new_new_n834__,
    new_new_n835__, new_new_n836__, new_new_n837__, new_new_n838__,
    new_new_n839__, new_new_n840__, new_new_n841__, new_new_n842__,
    new_new_n843__, new_new_n844__, new_new_n845__, new_new_n846__,
    new_new_n847__, new_new_n848__, new_new_n849__, new_new_n850__,
    new_new_n851__, new_new_n852__, new_new_n853__, new_new_n854__,
    new_new_n855__, new_new_n856__, new_new_n857__, new_new_n858__,
    new_new_n859__, new_new_n860__, new_new_n861__, new_new_n862__,
    new_new_n863__, new_new_n864__, new_new_n865__, new_new_n866__,
    new_new_n867__, new_new_n868__, new_new_n869__, new_new_n870__,
    new_new_n871__, new_new_n872__, new_new_n873__, new_new_n874__,
    new_new_n875__, new_new_n876__, new_new_n877__, new_new_n878__,
    new_new_n879__, new_new_n880__, new_new_n881__, new_new_n882__,
    new_new_n883__, new_new_n884__, new_new_n885__, new_new_n886__,
    new_new_n887__, new_new_n888__, new_new_n889__, new_new_n890__,
    new_new_n891__, new_new_n892__, new_new_n893__, new_new_n894__,
    new_new_n895__, new_new_n896__, new_new_n897__, new_new_n898__,
    new_new_n899__, new_new_n900__, new_new_n901__, new_new_n902__,
    new_new_n903__, new_new_n904__, new_new_n905__, new_new_n906__,
    new_new_n907__, new_new_n908__, new_new_n909__, new_new_n910__,
    new_new_n911__, new_new_n912__, new_new_n913__, new_new_n914__,
    new_new_n915__, new_new_n916__, new_new_n917__, new_new_n918__,
    new_new_n919__, new_new_n920__, new_new_n921__, new_new_n922__,
    new_new_n923__, new_new_n924__, new_new_n925__, new_new_n926__,
    new_new_n927__, new_new_n928__, new_new_n929__, new_new_n930__,
    new_new_n931__, new_new_n932__, new_new_n933__, new_new_n934__,
    new_new_n935__, new_new_n936__, new_new_n937__, new_new_n938__,
    new_new_n939__, new_new_n940__, new_new_n941__, new_new_n942__,
    new_new_n943__, new_new_n944__, new_new_n945__, new_new_n946__,
    new_new_n947__, new_new_n948__, new_new_n949__, new_new_n950__,
    new_new_n951__, new_new_n952__, new_new_n953__, new_new_n954__,
    new_new_n955__, new_new_n956__, new_new_n957__, new_new_n958__,
    new_new_n959__, new_new_n960__, new_new_n961__, new_new_n962__,
    new_new_n963__, new_new_n964__, new_new_n965__, new_new_n966__,
    new_new_n967__, new_new_n968__, new_new_n969__, new_new_n970__,
    new_new_n971__, new_new_n972__, new_new_n973__, new_new_n974__,
    new_new_n975__, new_new_n976__, new_new_n977__, new_new_n978__,
    new_new_n979__, new_new_n980__, new_new_n981__, new_new_n982__,
    new_new_n983__, new_new_n984__, new_new_n985__, new_new_n986__,
    new_new_n987__, new_new_n988__, new_new_n989__, new_new_n990__,
    new_new_n991__, new_new_n992__, new_new_n993__, new_new_n994__,
    new_new_n995__, new_new_n996__, new_new_n997__, new_new_n998__,
    new_new_n999__, new_new_n1000__, new_new_n1001__, new_new_n1002__,
    new_new_n1003__, new_new_n1004__, new_new_n1005__, new_new_n1006__,
    new_new_n1007__, new_new_n1008__, new_new_n1009__, new_new_n1010__,
    new_new_n1011__, new_new_n1012__, new_new_n1013__, new_new_n1014__,
    new_new_n1015__, new_new_n1016__, new_new_n1017__, new_new_n1018__,
    new_new_n1019__, new_new_n1020__, new_new_n1021__, new_new_n1022__,
    new_new_n1023__, new_new_n1024__, new_new_n1025__, new_new_n1026__,
    new_new_n1027__, new_new_n1028__, new_new_n1029__, new_new_n1030__,
    new_new_n1031__, new_new_n1032__, new_new_n1033__, new_new_n1034__,
    new_new_n1035__, new_new_n1036__, new_new_n1037__, new_new_n1038__,
    new_new_n1039__, new_new_n1040__, new_new_n1041__, new_new_n1042__,
    new_new_n1043__, new_new_n1044__, new_new_n1045__, new_new_n1046__,
    new_new_n1047__, new_new_n1048__, new_new_n1049__, new_new_n1050__,
    new_new_n1051__, new_new_n1052__, new_new_n1053__, new_new_n1054__,
    new_new_n1055__, new_new_n1056__, new_new_n1057__, new_new_n1058__,
    new_new_n1059__, new_new_n1060__, new_new_n1061__, new_new_n1062__,
    new_new_n1063__, new_new_n1064__, new_new_n1065__, new_new_n1066__,
    new_new_n1067__, new_new_n1068__, new_new_n1069__, new_new_n1070__,
    new_new_n1071__, new_new_n1072__, new_new_n1073__, new_new_n1074__,
    new_new_n1075__, new_new_n1076__, new_new_n1077__, new_new_n1078__,
    new_new_n1079__, new_new_n1080__, new_new_n1081__, new_new_n1082__,
    new_new_n1083__, new_new_n1084__, new_new_n1085__, new_new_n1086__,
    new_new_n1087__, new_new_n1088__, new_new_n1089__, new_new_n1090__,
    new_new_n1091__, new_new_n1092__, new_new_n1093__, new_new_n1094__,
    new_new_n1095__, new_new_n1096__, new_new_n1097__, new_new_n1098__,
    new_new_n1099__, new_new_n1100__, new_new_n1101__, new_new_n1102__,
    new_new_n1103__, new_new_n1104__, new_new_n1105__, new_new_n1106__,
    new_new_n1107__, new_new_n1108__, new_new_n1109__, new_new_n1110__,
    new_new_n1111__, new_new_n1112__, new_new_n1113__, new_new_n1114__,
    new_new_n1115__, new_new_n1116__, new_new_n1117__, new_new_n1118__,
    new_new_n1119__, new_new_n1120__, new_new_n1121__, new_new_n1122__,
    new_new_n1123__, new_new_n1124__, new_new_n1125__, new_new_n1126__,
    new_new_n1127__, new_new_n1128__, new_new_n1129__, new_new_n1130__,
    new_new_n1131__, new_new_n1132__, new_new_n1133__, new_new_n1134__,
    new_new_n1135__, new_new_n1136__, new_new_n1137__, new_new_n1138__,
    new_new_n1139__, new_new_n1140__, new_new_n1141__, new_new_n1142__,
    new_new_n1143__, new_new_n1144__, new_new_n1145__, new_new_n1146__,
    new_new_n1147__, new_new_n1148__, new_new_n1149__, new_new_n1150__,
    new_new_n1151__, new_new_n1152__, new_new_n1153__, new_new_n1154__,
    new_new_n1155__, new_new_n1156__, new_new_n1157__, new_new_n1158__,
    new_new_n1159__, new_new_n1160__, new_new_n1161__, new_new_n1162__,
    new_new_n1163__, new_new_n1164__, new_new_n1165__, new_new_n1166__,
    new_new_n1167__, new_new_n1168__, new_new_n1169__, new_new_n1170__,
    new_new_n1171__, new_new_n1172__, new_new_n1173__, new_new_n1174__,
    new_new_n1175__, new_new_n1176__, new_new_n1177__, new_new_n1178__,
    new_new_n1179__, new_new_n1180__, new_new_n1181__, new_new_n1182__,
    new_new_n1183__, new_new_n1184__, new_new_n1185__, new_new_n1186__,
    new_new_n1187__, new_new_n1188__, new_new_n1189__, new_new_n1190__,
    new_new_n1191__, new_new_n1192__, new_new_n1193__, new_new_n1194__,
    new_new_n1195__, new_new_n1196__, new_new_n1197__, new_new_n1198__,
    new_new_n1199__, new_new_n1200__, new_new_n1201__, new_new_n1202__,
    new_new_n1203__, new_new_n1204__, new_new_n1205__, new_new_n1206__,
    new_new_n1207__, new_new_n1208__, new_new_n1209__, new_new_n1210__,
    new_new_n1211__, new_new_n1212__, new_new_n1213__, new_new_n1214__,
    new_new_n1215__, new_new_n1216__, new_new_n1217__, new_new_n1218__,
    new_new_n1219__, new_new_n1220__, new_new_n1221__, new_new_n1222__,
    new_new_n1223__, new_new_n1224__, new_new_n1225__, new_new_n1226__,
    new_new_n1227__, new_new_n1228__, new_new_n1229__, new_new_n1230__,
    new_new_n1231__, new_new_n1232__, new_new_n1233__, new_new_n1234__,
    new_new_n1235__, new_new_n1236__, new_new_n1237__, new_new_n1238__,
    new_new_n1239__, new_new_n1240__, new_new_n1241__, new_new_n1242__,
    new_new_n1243__, new_new_n1244__, new_new_n1245__, new_new_n1246__,
    new_new_n1247__, new_new_n1248__, new_new_n1249__, new_new_n1250__,
    new_new_n1251__, new_new_n1252__, new_new_n1253__, new_new_n1254__,
    new_new_n1255__, new_new_n1256__, new_new_n1257__, new_new_n1258__,
    new_new_n1259__, new_new_n1260__, new_new_n1261__, new_new_n1262__,
    new_new_n1263__, new_new_n1264__, new_new_n1265__, new_new_n1266__,
    new_new_n1267__, new_new_n1268__, new_new_n1269__, new_new_n1270__,
    new_new_n1271__, new_new_n1272__, new_new_n1273__, new_new_n1274__,
    new_new_n1275__, new_new_n1276__, new_new_n1277__, new_new_n1278__,
    new_new_n1279__, new_new_n1280__, new_new_n1281__, new_new_n1282__,
    new_new_n1283__, new_new_n1284__, new_new_n1285__, new_new_n1286__,
    new_new_n1287__, new_new_n1288__, new_new_n1289__, new_new_n1290__,
    new_new_n1291__, new_new_n1292__, new_new_n1293__, new_new_n1294__,
    new_new_n1295__, new_new_n1296__, new_new_n1297__, new_new_n1298__,
    new_new_n1299__, new_new_n1300__, new_new_n1301__, new_new_n1302__,
    new_new_n1303__, new_new_n1304__, new_new_n1305__, new_new_n1306__,
    new_new_n1307__, new_new_n1308__, new_new_n1309__, new_new_n1310__,
    new_new_n1311__, new_new_n1312__, new_new_n1313__, new_new_n1314__,
    new_new_n1315__, new_new_n1316__, new_new_n1317__, new_new_n1318__,
    new_new_n1319__, new_new_n1320__, new_new_n1321__, new_new_n1322__,
    new_new_n1323__, new_new_n1324__, new_new_n1325__, new_new_n1326__,
    new_new_n1327__, new_new_n1328__, new_new_n1329__, new_new_n1330__,
    new_new_n1331__, new_new_n1332__, new_new_n1333__, new_new_n1334__,
    new_new_n1335__, new_new_n1336__, new_new_n1337__, new_new_n1338__,
    new_new_n1339__, new_new_n1340__, new_new_n1341__, new_new_n1342__,
    new_new_n1343__, new_new_n1344__, new_new_n1345__, new_new_n1346__,
    new_new_n1347__, new_new_n1348__, new_new_n1349__, new_new_n1350__,
    new_new_n1351__, new_new_n1352__, new_new_n1353__, new_new_n1354__,
    new_new_n1355__, new_new_n1356__, new_new_n1357__, new_new_n1358__,
    new_new_n1359__, new_new_n1360__, new_new_n1361__, new_new_n1362__,
    new_new_n1363__, new_new_n1364__, new_new_n1365__, new_new_n1366__,
    new_new_n1367__, new_new_n1368__, new_new_n1369__, new_new_n1370__,
    new_new_n1371__, new_new_n1372__, new_new_n1373__, new_new_n1374__,
    new_new_n1375__, new_new_n1376__, new_new_n1377__, new_new_n1378__,
    new_new_n1379__, new_new_n1380__, new_new_n1381__, new_new_n1382__,
    new_new_n1383__, new_new_n1384__, new_new_n1385__, new_new_n1386__,
    new_new_n1387__, new_new_n1388__, new_new_n1389__, new_new_n1390__,
    new_new_n1391__, new_new_n1392__, new_new_n1393__, new_new_n1394__,
    new_new_n1395__, new_new_n1396__, new_new_n1397__, new_new_n1398__,
    new_new_n1399__, new_new_n1400__, new_new_n1401__, new_new_n1402__,
    new_new_n1403__, new_new_n1404__, new_new_n1405__, new_new_n1406__,
    new_new_n1407__, new_new_n1408__, new_new_n1409__, new_new_n1410__,
    new_new_n1411__, new_new_n1412__, new_new_n1413__, new_new_n1414__,
    new_new_n1415__, new_new_n1416__, new_new_n1417__, new_new_n1418__,
    new_new_n1419__, new_new_n1420__, new_new_n1421__, new_new_n1422__,
    new_new_n1423__, new_new_n1424__, new_new_n1425__, new_new_n1426__,
    new_new_n1427__, new_new_n1428__, new_new_n1429__, new_new_n1430__,
    new_new_n1431__, new_new_n1432__, new_new_n1433__, new_new_n1434__,
    new_new_n1435__, new_new_n1436__, new_new_n1437__, new_new_n1438__,
    new_new_n1439__, new_new_n1440__, new_new_n1441__, new_new_n1442__,
    new_new_n1443__, new_new_n1444__, new_new_n1445__, new_new_n1446__,
    new_new_n1447__, new_new_n1448__, new_new_n1449__, new_new_n1450__,
    new_new_n1451__, new_new_n1452__, new_new_n1453__, new_new_n1454__,
    new_new_n1455__, new_new_n1456__, new_new_n1457__, new_new_n1458__,
    new_new_n1459__, new_new_n1460__, new_new_n1461__, new_new_n1462__,
    new_new_n1463__, new_new_n1464__, new_new_n1465__, new_new_n1466__,
    new_new_n1467__, new_new_n1468__, new_new_n1469__, new_new_n1470__,
    new_new_n1471__, new_new_n1472__, new_new_n1473__, new_new_n1474__,
    new_new_n1475__, new_new_n1476__, new_new_n1477__, new_new_n1478__,
    new_new_n1479__, new_new_n1480__, new_new_n1481__, new_new_n1482__,
    new_new_n1483__, new_new_n1484__, new_new_n1485__, new_new_n1486__,
    new_new_n1487__, new_new_n1488__, new_new_n1489__, new_new_n1490__,
    new_new_n1491__, new_new_n1492__, new_new_n1493__, new_new_n1494__,
    new_new_n1495__, new_new_n1496__, new_new_n1497__, new_new_n1498__,
    new_new_n1499__, new_new_n1500__, new_new_n1501__, new_new_n1502__,
    new_new_n1503__, new_new_n1504__, new_new_n1505__, new_new_n1506__,
    new_new_n1507__, new_new_n1508__, new_new_n1509__, new_new_n1510__,
    new_new_n1511__, new_new_n1512__, new_new_n1513__, new_new_n1514__,
    new_new_n1515__, new_new_n1516__, new_new_n1517__, new_new_n1518__,
    new_new_n1519__, new_new_n1520__, new_new_n1521__, new_new_n1522__,
    new_new_n1523__, new_new_n1524__, new_new_n1525__, new_new_n1526__,
    new_new_n1527__, new_new_n1528__, new_new_n1529__, new_new_n1530__,
    new_new_n1531__, new_new_n1532__, new_new_n1533__, new_new_n1534__,
    new_new_n1535__, new_new_n1536__, new_new_n1537__, new_new_n1538__,
    new_new_n1539__, new_new_n1540__, new_new_n1541__, new_new_n1542__,
    new_new_n1543__, new_new_n1544__, new_new_n1545__, new_new_n1546__,
    new_new_n1547__, new_new_n1548__, new_new_n1549__, new_new_n1550__,
    new_new_n1551__, new_new_n1552__, new_new_n1553__, new_new_n1554__,
    new_new_n1555__, new_new_n1556__, new_new_n1557__, new_new_n1558__,
    new_new_n1559__, new_new_n1560__, new_new_n1561__, new_new_n1562__,
    new_new_n1563__, new_new_n1564__, new_new_n1565__, new_new_n1566__,
    new_new_n1567__, new_new_n1568__, new_new_n1569__, new_new_n1570__,
    new_new_n1571__, new_new_n1572__, new_new_n1573__, new_new_n1574__,
    new_new_n1575__, new_new_n1576__, new_new_n1577__, new_new_n1578__,
    new_new_n1579__, new_new_n1580__, new_new_n1581__, new_new_n1582__,
    new_new_n1583__, new_new_n1584__, new_new_n1585__, new_new_n1586__,
    new_new_n1587__, new_new_n1588__, new_new_n1589__, new_new_n1590__,
    new_new_n1591__, new_new_n1592__, new_new_n1593__, new_new_n1594__,
    new_new_n1595__, new_new_n1596__, new_new_n1597__, new_new_n1598__,
    new_new_n1599__, new_new_n1600__, new_new_n1601__, new_new_n1602__,
    new_new_n1603__, new_new_n1604__, new_new_n1605__, new_new_n1606__,
    new_new_n1607__, new_new_n1608__, new_new_n1609__, new_new_n1610__,
    new_new_n1611__, new_new_n1612__, new_new_n1613__, new_new_n1614__,
    new_new_n1615__, new_new_n1616__, new_new_n1617__, new_new_n1618__,
    new_new_n1619__, new_new_n1620__, new_new_n1621__, new_new_n1622__,
    new_new_n1623__, new_new_n1624__, new_new_n1625__, new_new_n1626__,
    new_new_n1627__, new_new_n1628__, new_new_n1629__, new_new_n1630__,
    new_new_n1631__, new_new_n1632__, new_new_n1633__, new_new_n1634__,
    new_new_n1635__, new_new_n1636__, new_new_n1637__, new_new_n1638__,
    new_new_n1639__, new_new_n1640__, new_new_n1641__, new_new_n1642__,
    new_new_n1643__, new_new_n1644__, new_new_n1645__, new_new_n1646__,
    new_new_n1647__, new_new_n1648__, new_new_n1649__, new_new_n1650__,
    new_new_n1651__, new_new_n1652__, new_new_n1653__, new_new_n1654__,
    new_new_n1655__, new_new_n1656__, new_new_n1657__, new_new_n1658__,
    new_new_n1659__, new_new_n1660__, new_new_n1661__, new_new_n1662__,
    new_new_n1663__, new_new_n1664__, new_new_n1665__, new_new_n1666__,
    new_new_n1667__, new_new_n1668__, new_new_n1669__, new_new_n1670__,
    new_new_n1671__, new_new_n1672__, new_new_n1673__, new_new_n1674__,
    new_new_n1675__, new_new_n1676__, new_new_n1677__, new_new_n1678__,
    new_new_n1679__, new_new_n1680__, new_new_n1681__, new_new_n1682__,
    new_new_n1683__, new_new_n1684__, new_new_n1685__, new_new_n1686__,
    new_new_n1687__, new_new_n1688__, new_new_n1689__, new_new_n1690__,
    new_new_n1691__, new_new_n1692__, new_new_n1693__, new_new_n1694__,
    new_new_n1695__, new_new_n1696__, new_new_n1697__, new_new_n1698__,
    new_new_n1699__, new_new_n1700__, new_new_n1701__, new_new_n1702__,
    new_new_n1703__, new_new_n1704__, new_new_n1705__, new_new_n1706__,
    new_new_n1707__, new_new_n1708__, new_new_n1709__, new_new_n1710__,
    new_new_n1711__, new_new_n1712__, new_new_n1713__, new_new_n1714__,
    new_new_n1715__, new_new_n1716__, new_new_n1717__, new_new_n1718__,
    new_new_n1719__, new_new_n1720__, new_new_n1721__, new_new_n1722__,
    new_new_n1723__, new_new_n1724__, new_new_n1725__, new_new_n1726__,
    new_new_n1727__, new_new_n1728__, new_new_n1729__, new_new_n1730__,
    new_new_n1731__, new_new_n1732__, new_new_n1733__, new_new_n1734__,
    new_new_n1735__, new_new_n1736__, new_new_n1737__, new_new_n1738__,
    new_new_n1739__, new_new_n1740__, new_new_n1741__, new_new_n1742__,
    new_new_n1743__, new_new_n1744__, new_new_n1745__, new_new_n1746__,
    new_new_n1747__, new_new_n1748__, new_new_n1749__, new_new_n1750__,
    new_new_n1751__, new_new_n1752__, new_new_n1753__, new_new_n1754__,
    new_new_n1755__, new_new_n1756__, new_new_n1757__, new_new_n1758__,
    new_new_n1759__, new_new_n1760__, new_new_n1761__, new_new_n1762__,
    new_new_n1763__, new_new_n1764__, new_new_n1765__, new_new_n1766__,
    new_new_n1767__, new_new_n1768__, new_new_n1769__, new_new_n1770__,
    new_new_n1771__, new_new_n1772__, new_new_n1773__, new_new_n1774__,
    new_new_n1775__, new_new_n1776__, new_new_n1777__, new_new_n1778__,
    new_new_n1779__, new_new_n1780__, new_new_n1781__, new_new_n1782__,
    new_new_n1783__, new_new_n1784__, new_new_n1785__, new_new_n1786__,
    new_new_n1787__, new_new_n1788__, new_new_n1789__, new_new_n1790__,
    new_new_n1791__, new_new_n1792__, new_new_n1793__, new_new_n1794__,
    new_new_n1795__, new_new_n1796__, new_new_n1797__, new_new_n1798__,
    new_new_n1799__, new_new_n1800__, new_new_n1801__, new_new_n1802__,
    new_new_n1803__, new_new_n1804__, new_new_n1805__, new_new_n1806__,
    new_new_n1807__, new_new_n1808__, new_new_n1809__, new_new_n1810__,
    new_new_n1811__, new_new_n1812__, new_new_n1813__, new_new_n1814__,
    new_new_n1815__, new_new_n1816__, new_new_n1817__, new_new_n1818__,
    new_new_n1819__, new_new_n1820__, new_new_n1821__, new_new_n1822__,
    new_new_n1823__, new_new_n1824__, new_new_n1825__, new_new_n1826__,
    new_new_n1827__, new_new_n1828__, new_new_n1829__, new_new_n1830__,
    new_new_n1831__, new_new_n1832__, new_new_n1833__, new_new_n1834__,
    new_new_n1835__, new_new_n1836__, new_new_n1837__, new_new_n1838__,
    new_new_n1839__, new_new_n1840__, new_new_n1841__, new_new_n1842__,
    new_new_n1843__, new_new_n1844__, new_new_n1845__, new_new_n1846__,
    new_new_n1847__, new_new_n1848__, new_new_n1849__, new_new_n1850__,
    new_new_n1851__, new_new_n1852__, new_new_n1853__, new_new_n1854__,
    new_new_n1855__, new_new_n1856__, new_new_n1857__, new_new_n1858__,
    new_new_n1859__, new_new_n1860__, new_new_n1861__, new_new_n1862__,
    new_new_n1863__, new_new_n1864__, new_new_n1865__, new_new_n1866__,
    new_new_n1867__, new_new_n1868__, new_new_n1869__, new_new_n1870__,
    new_new_n1871__, new_new_n1872__, new_new_n1873__, new_new_n1874__,
    new_new_n1875__, new_new_n1876__, new_new_n1877__, new_new_n1878__,
    new_new_n1879__, new_new_n1880__, new_new_n1881__, new_new_n1882__,
    new_new_n1883__, new_new_n1884__, new_new_n1885__, new_new_n1886__,
    new_new_n1887__, new_new_n1888__, new_new_n1889__, new_new_n1890__,
    new_new_n1891__, new_new_n1892__, new_new_n1893__, new_new_n1894__,
    new_new_n1895__, new_new_n1896__, new_new_n1897__, new_new_n1898__,
    new_new_n1899__, new_new_n1900__, new_new_n1901__, new_new_n1902__,
    new_new_n1903__, new_new_n1904__, new_new_n1905__, new_new_n1906__,
    new_new_n1907__, new_new_n1908__, new_new_n1909__, new_new_n1910__,
    new_new_n1911__, new_new_n1912__, new_new_n1913__, new_new_n1914__,
    new_new_n1915__, new_new_n1916__, new_new_n1917__, new_new_n1918__,
    new_new_n1919__, new_new_n1920__, new_new_n1921__, new_new_n1922__,
    new_new_n1923__, new_new_n1924__, new_new_n1925__, new_new_n1926__,
    new_new_n1927__, new_new_n1928__, new_new_n1929__, new_new_n1930__,
    new_new_n1931__, new_new_n1932__, new_new_n1933__, new_new_n1934__,
    new_new_n1935__, new_new_n1936__, new_new_n1937__, new_new_n1938__,
    new_new_n1939__, new_new_n1940__, new_new_n1941__, new_new_n1942__,
    new_new_n1943__, new_new_n1944__, new_new_n1945__, new_new_n1946__,
    new_new_n1947__, new_new_n1948__, new_new_n1949__, new_new_n1950__,
    new_new_n1951__, new_new_n1952__, new_new_n1953__, new_new_n1954__,
    new_new_n1955__, new_new_n1956__, new_new_n1957__, new_new_n1958__,
    new_new_n1959__, new_new_n1960__, new_new_n1961__, new_new_n1962__,
    new_new_n1963__, new_new_n1964__, new_new_n1965__, new_new_n1966__,
    new_new_n1967__, new_new_n1968__, new_new_n1969__, new_new_n1970__,
    new_new_n1971__, new_new_n1972__, new_new_n1973__, new_new_n1974__,
    new_new_n1975__, new_new_n1976__, new_new_n1977__, new_new_n1978__,
    new_new_n1979__, new_new_n1980__, new_new_n1981__, new_new_n1982__,
    new_new_n1983__, new_new_n1984__, new_new_n1985__, new_new_n1986__,
    new_new_n1987__, new_new_n1988__, new_new_n1989__, new_new_n1990__,
    new_new_n1991__, new_new_n1992__, new_new_n1993__, new_new_n1994__,
    new_new_n1995__, new_new_n1996__, new_new_n1997__, new_new_n1998__,
    new_new_n1999__, new_new_n2000__, new_new_n2001__, new_new_n2002__,
    new_new_n2003__, new_new_n2004__, new_new_n2005__, new_new_n2006__,
    new_new_n2007__, new_new_n2008__, new_new_n2009__, new_new_n2010__,
    new_new_n2011__, new_new_n2012__, new_new_n2013__, new_new_n2014__,
    new_new_n2015__, new_new_n2016__, new_new_n2017__, new_new_n2018__,
    new_new_n2019__, new_new_n2020__, new_new_n2021__, new_new_n2022__,
    new_new_n2023__, new_new_n2024__, new_new_n2025__, new_new_n2026__,
    new_new_n2027__, new_new_n2028__, new_new_n2029__, new_new_n2030__,
    new_new_n2031__, new_new_n2032__, new_new_n2033__, new_new_n2034__,
    new_new_n2035__, new_new_n2036__, new_new_n2037__, new_new_n2038__,
    new_new_n2039__, new_new_n2040__, new_new_n2041__, new_new_n2042__,
    new_new_n2043__, new_new_n2044__, new_new_n2045__, new_new_n2046__,
    new_new_n2047__, new_new_n2048__, new_new_n2049__, new_new_n2050__,
    new_new_n2051__, new_new_n2052__, new_new_n2053__, new_new_n2054__,
    new_new_n2055__, new_new_n2056__, new_new_n2057__, new_new_n2058__,
    new_new_n2059__, new_new_n2060__, new_new_n2061__, new_new_n2062__,
    new_new_n2063__, new_new_n2064__, new_new_n2065__, new_new_n2066__,
    new_new_n2067__, new_new_n2068__, new_new_n2069__, new_new_n2070__,
    new_new_n2071__, new_new_n2072__, new_new_n2073__, new_new_n2074__,
    new_new_n2075__, new_new_n2076__, new_new_n2077__, new_new_n2078__,
    new_new_n2079__, new_new_n2080__, new_new_n2081__, new_new_n2082__,
    new_new_n2083__, new_new_n2084__, new_new_n2085__, new_new_n2086__,
    new_new_n2087__, new_new_n2088__, new_new_n2089__, new_new_n2090__,
    new_new_n2091__, new_new_n2092__, new_new_n2093__, new_new_n2094__,
    new_new_n2095__, new_new_n2096__, new_new_n2097__, new_new_n2098__,
    new_new_n2099__, new_new_n2100__, new_new_n2101__, new_new_n2102__,
    new_new_n2103__, new_new_n2104__, new_new_n2105__, new_new_n2106__,
    new_new_n2107__, new_new_n2108__, new_new_n2109__, new_new_n2110__,
    new_new_n2111__, new_new_n2112__, new_new_n2113__, new_new_n2114__,
    new_new_n2115__, new_new_n2116__, new_new_n2117__, new_new_n2118__,
    new_new_n2119__, new_new_n2120__, new_new_n2121__, new_new_n2122__,
    new_new_n2123__, new_new_n2124__, new_new_n2125__, new_new_n2126__,
    new_new_n2127__, new_new_n2128__, new_new_n2129__, new_new_n2130__,
    new_new_n2131__, new_new_n2132__, new_new_n2133__, new_new_n2134__,
    new_new_n2135__, new_new_n2136__, new_new_n2137__, new_new_n2138__,
    new_new_n2139__, new_new_n2140__, new_new_n2141__, new_new_n2142__,
    new_new_n2143__, new_new_n2144__, new_new_n2145__, new_new_n2146__,
    new_new_n2147__, new_new_n2148__, new_new_n2149__, new_new_n2150__,
    new_new_n2151__, new_new_n2152__, new_new_n2153__, new_new_n2154__,
    new_new_n2155__, new_new_n2156__, new_new_n2157__, new_new_n2158__,
    new_new_n2159__, new_new_n2160__, new_new_n2161__, new_new_n2162__,
    new_new_n2163__, new_new_n2164__, new_new_n2165__, new_new_n2166__,
    new_new_n2167__, new_new_n2168__, new_new_n2169__, new_new_n2170__,
    new_new_n2171__, new_new_n2172__, new_new_n2173__, new_new_n2174__,
    new_new_n2175__, new_new_n2176__, new_new_n2177__, new_new_n2178__,
    new_new_n2179__, new_new_n2180__, new_new_n2181__, new_new_n2182__,
    new_new_n2183__, new_new_n2184__, new_new_n2185__, new_new_n2186__,
    new_new_n2187__, new_new_n2188__, new_new_n2189__, new_new_n2190__,
    new_new_n2191__, new_new_n2192__, new_new_n2193__, new_new_n2194__,
    new_new_n2195__, new_new_n2196__, new_new_n2197__, new_new_n2198__,
    new_new_n2199__, new_new_n2200__, new_new_n2201__, new_new_n2202__,
    new_new_n2203__, new_new_n2204__, new_new_n2205__, new_new_n2206__,
    new_new_n2207__, new_new_n2208__, new_new_n2209__, new_new_n2210__,
    new_new_n2211__, new_new_n2212__, new_new_n2213__, new_new_n2214__,
    new_new_n2215__, new_new_n2216__, new_new_n2217__, new_new_n2218__,
    new_new_n2219__, new_new_n2220__, new_new_n2221__, new_new_n2222__,
    new_new_n2223__, new_new_n2224__, new_new_n2225__, new_new_n2226__,
    new_new_n2227__, new_new_n2228__, new_new_n2229__, new_new_n2230__,
    new_new_n2231__, new_new_n2232__, new_new_n2233__, new_new_n2234__,
    new_new_n2235__, new_new_n2236__, new_new_n2237__, new_new_n2238__,
    new_new_n2239__, new_new_n2240__, new_new_n2241__, new_new_n2242__,
    new_new_n2243__, new_new_n2244__, new_new_n2245__, new_new_n2246__,
    new_new_n2247__, new_new_n2248__, new_new_n2249__, new_new_n2250__,
    new_new_n2251__, new_new_n2252__, new_new_n2253__, new_new_n2254__,
    new_new_n2255__, new_new_n2256__, new_new_n2257__, new_new_n2258__,
    new_new_n2259__, new_new_n2260__, new_new_n2261__, new_new_n2262__,
    new_new_n2263__, new_new_n2264__, new_new_n2265__, new_new_n2266__,
    new_new_n2267__, new_new_n2268__, new_new_n2269__, new_new_n2270__,
    new_new_n2271__, new_new_n2272__, new_new_n2273__, new_new_n2274__,
    new_new_n2275__, new_new_n2276__, new_new_n2277__, new_new_n2278__,
    new_new_n2279__, new_new_n2280__, new_new_n2281__, new_new_n2282__,
    new_new_n2283__, new_new_n2284__, new_new_n2285__, new_new_n2286__,
    new_new_n2287__, new_new_n2288__, new_new_n2289__, new_new_n2290__,
    new_new_n2291__, new_new_n2292__, new_new_n2293__, new_new_n2294__,
    new_new_n2295__, new_new_n2296__, new_new_n2297__, new_new_n2298__,
    new_new_n2299__, new_new_n2300__, new_new_n2301__, new_new_n2302__,
    new_new_n2303__, new_new_n2304__, new_new_n2305__, new_new_n2306__,
    new_new_n2307__, new_new_n2308__, new_new_n2309__, new_new_n2310__,
    new_new_n2311__, new_new_n2312__, new_new_n2313__, new_new_n2314__,
    new_new_n2315__, new_new_n2316__, new_new_n2317__, new_new_n2318__,
    new_new_n2319__, new_new_n2320__, new_new_n2321__, new_new_n2322__,
    new_new_n2323__, new_new_n2324__, new_new_n2325__, new_new_n2326__,
    new_new_n2327__, new_new_n2328__, new_new_n2329__, new_new_n2330__,
    new_new_n2331__, new_new_n2332__, new_new_n2333__, new_new_n2334__,
    new_new_n2335__, new_new_n2336__, new_new_n2337__, new_new_n2338__,
    new_new_n2339__, new_new_n2340__, new_new_n2341__, new_new_n2342__,
    new_new_n2343__, new_new_n2344__, new_new_n2345__, new_new_n2346__,
    new_new_n2347__, new_new_n2348__, new_new_n2349__, new_new_n2350__,
    new_new_n2351__, new_new_n2352__, new_new_n2353__, new_new_n2354__,
    new_new_n2355__, new_new_n2356__, new_new_n2357__, new_new_n2358__,
    new_new_n2359__, new_new_n2360__, new_new_n2361__, new_new_n2362__,
    new_new_n2363__, new_new_n2364__, new_new_n2365__, new_new_n2366__,
    new_new_n2367__, new_new_n2368__, new_new_n2369__, new_new_n2370__,
    new_new_n2371__, new_new_n2372__, new_new_n2373__, new_new_n2374__,
    new_new_n2375__, new_new_n2376__, new_new_n2377__, new_new_n2378__,
    new_new_n2379__, new_new_n2380__, new_new_n2381__, new_new_n2382__,
    new_new_n2383__, new_new_n2384__, new_new_n2385__, new_new_n2386__,
    new_new_n2387__, new_new_n2388__, new_new_n2389__, new_new_n2390__,
    new_new_n2391__, new_new_n2392__, new_new_n2393__, new_new_n2394__,
    new_new_n2395__, new_new_n2396__, new_new_n2397__, new_new_n2398__,
    new_new_n2399__, new_new_n2400__, new_new_n2401__, new_new_n2402__,
    new_new_n2403__, new_new_n2404__, new_new_n2405__, new_new_n2406__,
    new_new_n2407__, new_new_n2408__, new_new_n2409__, new_new_n2410__,
    new_new_n2411__, new_new_n2412__, new_new_n2413__, new_new_n2414__,
    new_new_n2415__, new_new_n2416__, new_new_n2417__, new_new_n2418__,
    new_new_n2419__, new_new_n2420__, new_new_n2421__, new_new_n2422__,
    new_new_n2423__, new_new_n2424__, new_new_n2425__, new_new_n2426__,
    new_new_n2427__, new_new_n2428__, new_new_n2429__, new_new_n2430__,
    new_new_n2431__, new_new_n2432__, new_new_n2433__, new_new_n2434__,
    new_new_n2435__, new_new_n2436__, new_new_n2437__, new_new_n2438__,
    new_new_n2439__, new_new_n2440__, new_new_n2441__, new_new_n2442__,
    new_new_n2443__, new_new_n2444__, new_new_n2445__, new_new_n2446__,
    new_new_n2447__, new_new_n2448__, new_new_n2449__, new_new_n2450__,
    new_new_n2451__, new_new_n2452__, new_new_n2453__, new_new_n2454__,
    new_new_n2455__, new_new_n2456__, new_new_n2457__, new_new_n2458__,
    new_new_n2459__, new_new_n2460__, new_new_n2461__, new_new_n2462__,
    new_new_n2463__, new_new_n2464__, new_new_n2465__, new_new_n2466__,
    new_new_n2467__, new_new_n2468__, new_new_n2469__, new_new_n2470__,
    new_new_n2471__, new_new_n2472__, new_new_n2473__, new_new_n2474__,
    new_new_n2475__, new_new_n2476__, new_new_n2477__, new_new_n2478__,
    new_new_n2479__, new_new_n2480__, new_new_n2481__, new_new_n2482__,
    new_new_n2483__, new_new_n2484__, new_new_n2485__, new_new_n2486__,
    new_new_n2487__, new_new_n2488__, new_new_n2489__, new_new_n2490__,
    new_new_n2491__, new_new_n2492__, new_new_n2493__, new_new_n2494__,
    new_new_n2495__, new_new_n2496__, new_new_n2497__, new_new_n2498__,
    new_new_n2499__, new_new_n2500__, new_new_n2501__, new_new_n2502__,
    new_new_n2503__, new_new_n2504__, new_new_n2505__, new_new_n2506__,
    new_new_n2507__, new_new_n2508__, new_new_n2509__, new_new_n2510__,
    new_new_n2511__, new_new_n2512__, new_new_n2513__, new_new_n2514__,
    new_new_n2515__, new_new_n2516__, new_new_n2517__, new_new_n2518__,
    new_new_n2519__, new_new_n2520__, new_new_n2521__, new_new_n2522__,
    new_new_n2523__, new_new_n2524__, new_new_n2525__, new_new_n2526__,
    new_new_n2527__, new_new_n2528__, new_new_n2529__, new_new_n2530__,
    new_new_n2531__, new_new_n2532__, new_new_n2533__, new_new_n2534__,
    new_new_n2535__, new_new_n2536__, new_new_n2537__, new_new_n2538__,
    new_new_n2539__, new_new_n2540__, new_new_n2541__, new_new_n2542__,
    new_new_n2543__, new_new_n2544__, new_new_n2545__, new_new_n2546__,
    new_new_n2547__, new_new_n2548__, new_new_n2549__, new_new_n2550__,
    new_new_n2551__, new_new_n2552__, new_new_n2553__, new_new_n2554__,
    new_new_n2555__, new_new_n2556__, new_new_n2557__, new_new_n2558__,
    new_new_n2559__, new_new_n2560__, new_new_n2561__, new_new_n2562__,
    new_new_n2563__, new_new_n2564__, new_new_n2565__, new_new_n2566__,
    new_new_n2567__, new_new_n2568__, new_new_n2569__, new_new_n2570__,
    new_new_n2571__, new_new_n2572__, new_new_n2573__, new_new_n2574__,
    new_new_n2575__, new_new_n2576__, new_new_n2577__, new_new_n2578__,
    new_new_n2579__, new_new_n2580__, new_new_n2581__, new_new_n2582__,
    new_new_n2583__, new_new_n2584__, new_new_n2585__, new_new_n2586__,
    new_new_n2587__, new_new_n2588__, new_new_n2589__, new_new_n2590__,
    new_new_n2591__, new_new_n2592__, new_new_n2593__, new_new_n2594__,
    new_new_n2595__, new_new_n2596__, new_new_n2597__, new_new_n2598__,
    new_new_n2599__, new_new_n2600__, new_new_n2601__, new_new_n2602__,
    new_new_n2603__, new_new_n2604__, new_new_n2605__, new_new_n2606__,
    new_new_n2607__, new_new_n2608__, new_new_n2609__, new_new_n2610__,
    new_new_n2611__, new_new_n2612__, new_new_n2613__, new_new_n2614__,
    new_new_n2615__, new_new_n2616__, new_new_n2617__, new_new_n2618__,
    new_new_n2619__, new_new_n2620__, new_new_n2621__, new_new_n2622__,
    new_new_n2623__, new_new_n2624__, new_new_n2625__, new_new_n2626__,
    new_new_n2627__, new_new_n2628__, new_new_n2629__, new_new_n2630__,
    new_new_n2631__, new_new_n2632__, new_new_n2633__, new_new_n2634__,
    new_new_n2635__, new_new_n2636__, new_new_n2637__, new_new_n2638__,
    new_new_n2639__, new_new_n2640__, new_new_n2641__, new_new_n2642__,
    new_new_n2643__, new_new_n2644__, new_new_n2645__, new_new_n2646__,
    new_new_n2647__, new_new_n2648__, new_new_n2649__, new_new_n2650__,
    new_new_n2651__, new_new_n2652__, new_new_n2653__, new_new_n2654__,
    new_new_n2655__, new_new_n2656__, new_new_n2657__, new_new_n2658__,
    new_new_n2659__, new_new_n2660__, new_new_n2661__, new_new_n2662__,
    new_new_n2663__, new_new_n2664__, new_new_n2665__, new_new_n2666__,
    new_new_n2667__, new_new_n2668__, new_new_n2669__, new_new_n2670__,
    new_new_n2671__, new_new_n2672__, new_new_n2673__, new_new_n2674__,
    new_new_n2675__, new_new_n2676__, new_new_n2677__, new_new_n2678__,
    new_new_n2679__, new_new_n2680__, new_new_n2681__, new_new_n2682__,
    new_new_n2683__, new_new_n2684__, new_new_n2685__, new_new_n2686__,
    new_new_n2687__, new_new_n2688__, new_new_n2689__, new_new_n2690__,
    new_new_n2691__, new_new_n2692__, new_new_n2693__, new_new_n2694__,
    new_new_n2695__, new_new_n2696__, new_new_n2697__, new_new_n2698__,
    new_new_n2699__, new_new_n2700__, new_new_n2701__, new_new_n2702__,
    new_new_n2703__, new_new_n2704__, new_new_n2705__, new_new_n2706__,
    new_new_n2707__, new_new_n2708__, new_new_n2709__, new_new_n2710__,
    new_new_n2711__, new_new_n2712__, new_new_n2713__, new_new_n2714__,
    new_new_n2715__, new_new_n2716__, new_new_n2717__, new_new_n2718__,
    new_new_n2719__, new_new_n2720__, new_new_n2721__, new_new_n2722__,
    new_new_n2723__, new_new_n2724__, new_new_n2725__, new_new_n2726__,
    new_new_n2727__, new_new_n2728__, new_new_n2729__, new_new_n2730__,
    new_new_n2731__, new_new_n2732__, new_new_n2733__, new_new_n2734__,
    new_new_n2735__, new_new_n2736__, new_new_n2737__, new_new_n2738__,
    new_new_n2739__, new_new_n2740__, new_new_n2741__, new_new_n2742__,
    new_new_n2743__, new_new_n2744__, new_new_n2745__, new_new_n2746__,
    new_new_n2747__, new_new_n2748__, new_new_n2749__, new_new_n2750__,
    new_new_n2751__, new_new_n2752__, new_new_n2753__, new_new_n2754__,
    new_new_n2755__, new_new_n2756__, new_new_n2757__, new_new_n2758__,
    new_new_n2759__, new_new_n2760__, new_new_n2761__, new_new_n2762__,
    new_new_n2763__, new_new_n2764__, new_new_n2765__, new_new_n2766__,
    new_new_n2767__, new_new_n2768__, new_new_n2769__, new_new_n2770__,
    new_new_n2771__, new_new_n2772__, new_new_n2773__, new_new_n2774__,
    new_new_n2775__, new_new_n2776__, new_new_n2777__, new_new_n2778__,
    new_new_n2779__, new_new_n2780__, new_new_n2781__, new_new_n2782__,
    new_new_n2783__, new_new_n2784__, new_new_n2785__, new_new_n2786__,
    new_new_n2787__, new_new_n2788__, new_new_n2789__, new_new_n2790__,
    new_new_n2791__, new_new_n2792__, new_new_n2793__, new_new_n2794__,
    new_new_n2795__, new_new_n2796__, new_new_n2797__, new_new_n2798__,
    new_new_n2799__, new_new_n2800__, new_new_n2801__, new_new_n2802__,
    new_new_n2803__, new_new_n2804__, new_new_n2805__, new_new_n2806__,
    new_new_n2807__, new_new_n2808__, new_new_n2809__, new_new_n2810__,
    new_new_n2811__, new_new_n2812__, new_new_n2813__, new_new_n2814__,
    new_new_n2815__, new_new_n2816__, new_new_n2817__, new_new_n2818__,
    new_new_n2819__, new_new_n2820__, new_new_n2821__, new_new_n2822__,
    new_new_n2823__, new_new_n2824__, new_new_n2825__, new_new_n2826__,
    new_new_n2827__, new_new_n2828__, new_new_n2829__, new_new_n2830__,
    new_new_n2831__, new_new_n2832__, new_new_n2833__, new_new_n2834__,
    new_new_n2835__, new_new_n2836__, new_new_n2837__, new_new_n2838__,
    new_new_n2839__, new_new_n2840__, new_new_n2841__, new_new_n2842__,
    new_new_n2843__, new_new_n2844__, new_new_n2845__, new_new_n2846__,
    new_new_n2847__, new_new_n2848__, new_new_n2849__, new_new_n2850__,
    new_new_n2851__, new_new_n2852__, new_new_n2853__, new_new_n2854__,
    new_new_n2855__, new_new_n2856__, new_new_n2857__, new_new_n2858__,
    new_new_n2859__, new_new_n2860__, new_new_n2861__, new_new_n2862__,
    new_new_n2863__, new_new_n2864__, new_new_n2865__, new_new_n2866__,
    new_new_n2867__, new_new_n2868__, new_new_n2869__, new_new_n2870__,
    new_new_n2871__, new_new_n2872__, new_new_n2873__, new_new_n2874__,
    new_new_n2875__, new_new_n2876__, new_new_n2877__, new_new_n2878__,
    new_new_n2879__, new_new_n2880__, new_new_n2881__, new_new_n2882__,
    new_new_n2883__, new_new_n2884__, new_new_n2885__, new_new_n2886__,
    new_new_n2887__, new_new_n2888__, new_new_n2889__, new_new_n2890__,
    new_new_n2891__, new_new_n2892__, new_new_n2893__, new_new_n2894__,
    new_new_n2895__, new_new_n2896__, new_new_n2897__, new_new_n2898__,
    new_new_n2899__, new_new_n2900__, new_new_n2901__, new_new_n2902__,
    new_new_n2903__, new_new_n2904__, new_new_n2905__, new_new_n2906__,
    new_new_n2907__, new_new_n2908__, new_new_n2909__, new_new_n2910__,
    new_new_n2911__, new_new_n2912__, new_new_n2913__, new_new_n2914__,
    new_new_n2915__, new_new_n2916__, new_new_n2917__, new_new_n2918__,
    new_new_n2919__, new_new_n2920__, new_new_n2921__, new_new_n2922__,
    new_new_n2923__, new_new_n2924__, new_new_n2925__, new_new_n2926__,
    new_new_n2927__, new_new_n2928__, new_new_n2929__, new_new_n2930__,
    new_new_n2931__, new_new_n2932__, new_new_n2933__, new_new_n2934__,
    new_new_n2935__, new_new_n2936__, new_new_n2937__, new_new_n2938__,
    new_new_n2939__, new_new_n2940__, new_new_n2941__, new_new_n2942__,
    new_new_n2944__, new_new_n2945__, new_new_n2947__, new_new_n2948__,
    new_new_n2950__, new_new_n2951__, new_new_n2953__, new_new_n2954__,
    new_new_n2956__, new_new_n2957__, new_new_n2959__, new_new_n2960__,
    new_new_n2962__, new_new_n2963__, new_new_n2965__, new_new_n2966__,
    new_new_n2968__, new_new_n2969__, new_new_n2971__, new_new_n2972__,
    new_new_n2974__, new_new_n2975__, new_new_n2977__, new_new_n2978__,
    new_new_n2980__, new_new_n2981__, new_new_n2983__, new_new_n2984__,
    new_new_n2986__, new_new_n2987__, new_new_n2989__, new_new_n2990__,
    new_new_n2992__, new_new_n2993__, new_new_n2995__, new_new_n2996__,
    new_new_n2998__, new_new_n2999__, new_new_n3001__, new_new_n3002__,
    new_new_n3004__, new_new_n3005__, new_new_n3007__, new_new_n3008__,
    new_new_n3010__, new_new_n3011__, new_new_n3013__, new_new_n3014__,
    new_new_n3016__, new_new_n3017__, new_new_n3019__, new_new_n3020__,
    new_new_n3022__, new_new_n3023__, new_new_n3025__, new_new_n3026__,
    new_new_n3028__, new_new_n3029__, new_new_n3031__, new_new_n3032__,
    new_new_n3034__, new_new_n3035__, new_new_n3037__, new_new_n3038__,
    new_new_n3040__, new_new_n3041__, new_new_n3043__, new_new_n3044__,
    new_new_n3046__, new_new_n3047__, new_new_n3049__, new_new_n3050__,
    new_new_n3052__, new_new_n3053__, new_new_n3055__, new_new_n3056__,
    new_new_n3058__, new_new_n3059__, new_new_n3061__, new_new_n3062__,
    new_new_n3064__, new_new_n3065__, new_new_n3067__, new_new_n3068__,
    new_new_n3070__, new_new_n3071__, new_new_n3073__, new_new_n3074__,
    new_new_n3076__, new_new_n3077__, new_new_n3079__, new_new_n3080__,
    new_new_n3082__, new_new_n3083__, new_new_n3085__, new_new_n3086__,
    new_new_n3088__, new_new_n3089__, new_new_n3091__, new_new_n3092__,
    new_new_n3094__, new_new_n3095__, new_new_n3097__, new_new_n3098__,
    new_new_n3100__, new_new_n3101__, new_new_n3103__, new_new_n3104__,
    new_new_n3106__, new_new_n3107__, new_new_n3109__, new_new_n3110__,
    new_new_n3112__, new_new_n3113__, new_new_n3115__, new_new_n3116__,
    new_new_n3118__, new_new_n3119__, new_new_n3121__, new_new_n3122__,
    new_new_n3124__, new_new_n3125__, new_new_n3127__, new_new_n3128__,
    new_new_n3130__, new_new_n3131__, new_new_n3133__, new_new_n3134__,
    new_new_n3136__, new_new_n3137__, new_new_n3139__, new_new_n3140__,
    new_new_n3142__, new_new_n3143__, new_new_n3145__, new_new_n3146__,
    new_new_n3148__, new_new_n3149__, new_new_n3151__, new_new_n3152__,
    new_new_n3154__, new_new_n3155__, new_new_n3157__, new_new_n3158__,
    new_new_n3160__, new_new_n3161__, new_new_n3163__, new_new_n3164__,
    new_new_n3166__, new_new_n3167__, new_new_n3169__, new_new_n3170__,
    new_new_n3172__, new_new_n3173__, new_new_n3175__, new_new_n3176__,
    new_new_n3178__, new_new_n3179__, new_new_n3181__, new_new_n3182__,
    new_new_n3184__, new_new_n3185__, new_new_n3187__, new_new_n3188__,
    new_new_n3190__, new_new_n3191__, new_new_n3193__, new_new_n3194__,
    new_new_n3196__, new_new_n3197__, new_new_n3199__, new_new_n3200__,
    new_new_n3202__, new_new_n3203__, new_new_n3205__, new_new_n3206__,
    new_new_n3208__, new_new_n3209__, new_new_n3211__, new_new_n3212__,
    new_new_n3214__, new_new_n3215__, new_new_n3217__, new_new_n3218__,
    new_new_n3220__, new_new_n3221__, new_new_n3223__, new_new_n3224__,
    new_new_n3226__, new_new_n3227__, new_new_n3229__, new_new_n3230__,
    new_new_n3232__, new_new_n3233__, new_new_n3235__, new_new_n3236__,
    new_new_n3238__, new_new_n3239__, new_new_n3241__, new_new_n3242__,
    new_new_n3244__, new_new_n3245__, new_new_n3247__, new_new_n3248__,
    new_new_n3250__, new_new_n3251__, new_new_n3253__, new_new_n3254__,
    new_new_n3256__, new_new_n3257__, new_new_n3259__, new_new_n3260__,
    new_new_n3262__, new_new_n3263__, new_new_n3265__, new_new_n3266__,
    new_new_n3268__, new_new_n3269__, new_new_n3271__, new_new_n3272__,
    new_new_n3274__, new_new_n3275__, new_new_n3277__, new_new_n3278__,
    new_new_n3280__, new_new_n3281__, new_new_n3283__, new_new_n3284__,
    new_new_n3286__, new_new_n3287__, new_new_n3289__, new_new_n3290__,
    new_new_n3292__, new_new_n3293__, new_new_n3295__, new_new_n3296__,
    new_new_n3298__, new_new_n3299__, new_new_n3301__, new_new_n3302__,
    new_new_n3304__, new_new_n3305__, new_new_n3307__, new_new_n3308__,
    new_new_n3310__, new_new_n3311__, new_new_n3313__, new_new_n3314__,
    new_new_n3316__, new_new_n3317__, new_new_n3319__, new_new_n3320__,
    new_new_n3322__, new_new_n3323__, new_new_n3326__, new_new_n3327__;
  assign new_new_n643__ = pi122 & ~pi250;
  assign new_new_n644__ = pi123 & ~pi251;
  assign new_new_n645__ = ~pi122 & pi250;
  assign new_new_n646__ = pi121 & ~pi249;
  assign new_new_n647__ = ~pi121 & pi249;
  assign new_new_n648__ = pi120 & ~pi248;
  assign new_new_n649__ = ~pi120 & pi248;
  assign new_new_n650__ = ~pi119 & pi247;
  assign new_new_n651__ = pi117 & ~pi245;
  assign new_new_n652__ = ~pi116 & pi244;
  assign new_new_n653__ = pi114 & ~pi242;
  assign new_new_n654__ = ~pi113 & pi241;
  assign new_new_n655__ = ~pi110 & pi238;
  assign new_new_n656__ = pi109 & ~pi237;
  assign new_new_n657__ = pi106 & ~pi234;
  assign new_new_n658__ = ~pi105 & pi233;
  assign new_new_n659__ = ~pi102 & pi230;
  assign new_new_n660__ = pi101 & ~pi229;
  assign new_new_n661__ = pi098 & ~pi226;
  assign new_new_n662__ = ~pi097 & pi225;
  assign new_new_n663__ = pi095 & ~pi223;
  assign new_new_n664__ = ~pi094 & pi222;
  assign new_new_n665__ = ~pi093 & pi221;
  assign new_new_n666__ = pi092 & ~pi220;
  assign new_new_n667__ = pi091 & ~pi219;
  assign new_new_n668__ = ~pi090 & pi218;
  assign new_new_n669__ = ~pi088 & pi216;
  assign new_new_n670__ = ~pi089 & pi217;
  assign new_new_n671__ = pi087 & ~pi215;
  assign new_new_n672__ = pi088 & ~pi216;
  assign new_new_n673__ = ~pi087 & pi215;
  assign new_new_n674__ = pi086 & ~pi214;
  assign new_new_n675__ = ~pi086 & pi214;
  assign new_new_n676__ = pi085 & ~pi213;
  assign new_new_n677__ = ~pi085 & pi213;
  assign new_new_n678__ = pi084 & ~pi212;
  assign new_new_n679__ = ~pi084 & pi212;
  assign new_new_n680__ = pi083 & ~pi211;
  assign new_new_n681__ = ~pi083 & pi211;
  assign new_new_n682__ = pi082 & ~pi210;
  assign new_new_n683__ = ~pi082 & pi210;
  assign new_new_n684__ = pi081 & ~pi209;
  assign new_new_n685__ = ~pi081 & pi209;
  assign new_new_n686__ = pi080 & ~pi208;
  assign new_new_n687__ = ~pi080 & pi208;
  assign new_new_n688__ = ~pi079 & pi207;
  assign new_new_n689__ = pi078 & ~pi206;
  assign new_new_n690__ = pi079 & ~pi207;
  assign new_new_n691__ = ~pi077 & pi205;
  assign new_new_n692__ = ~pi078 & pi206;
  assign new_new_n693__ = pi077 & ~pi205;
  assign new_new_n694__ = ~pi076 & pi204;
  assign new_new_n695__ = pi076 & ~pi204;
  assign new_new_n696__ = ~pi075 & pi203;
  assign new_new_n697__ = pi075 & ~pi203;
  assign new_new_n698__ = ~pi074 & pi202;
  assign new_new_n699__ = pi074 & ~pi202;
  assign new_new_n700__ = ~pi073 & pi201;
  assign new_new_n701__ = pi073 & ~pi201;
  assign new_new_n702__ = ~pi072 & pi200;
  assign new_new_n703__ = pi072 & ~pi200;
  assign new_new_n704__ = ~pi071 & pi199;
  assign new_new_n705__ = pi067 & ~pi195;
  assign new_new_n706__ = ~pi066 & pi194;
  assign new_new_n707__ = pi065 & ~pi193;
  assign new_new_n708__ = pi066 & ~pi194;
  assign new_new_n709__ = ~pi064 & pi192;
  assign new_new_n710__ = ~pi065 & pi193;
  assign new_new_n711__ = pi064 & ~pi192;
  assign new_new_n712__ = ~pi063 & pi191;
  assign new_new_n713__ = pi057 & ~pi185;
  assign new_new_n714__ = ~pi056 & pi184;
  assign new_new_n715__ = ~pi054 & pi182;
  assign new_new_n716__ = ~pi055 & pi183;
  assign new_new_n717__ = pi053 & ~pi181;
  assign new_new_n718__ = pi054 & ~pi182;
  assign new_new_n719__ = ~pi053 & pi181;
  assign new_new_n720__ = pi052 & ~pi180;
  assign new_new_n721__ = ~pi052 & pi180;
  assign new_new_n722__ = pi051 & ~pi179;
  assign new_new_n723__ = ~pi051 & pi179;
  assign new_new_n724__ = pi050 & ~pi178;
  assign new_new_n725__ = ~pi050 & pi178;
  assign new_new_n726__ = ~pi049 & pi177;
  assign new_new_n727__ = pi039 & ~pi167;
  assign new_new_n728__ = ~pi038 & pi166;
  assign new_new_n729__ = pi035 & ~pi163;
  assign new_new_n730__ = pi036 & ~pi164;
  assign new_new_n731__ = ~pi034 & pi162;
  assign new_new_n732__ = ~pi035 & pi163;
  assign new_new_n733__ = pi034 & ~pi162;
  assign new_new_n734__ = ~pi033 & pi161;
  assign new_new_n735__ = pi033 & ~pi161;
  assign new_new_n736__ = pi032 & ~pi160;
  assign new_new_n737__ = ~pi030 & pi158;
  assign new_new_n738__ = pi029 & ~pi157;
  assign new_new_n739__ = ~pi027 & pi155;
  assign new_new_n740__ = pi026 & ~pi154;
  assign new_new_n741__ = ~pi023 & pi151;
  assign new_new_n742__ = ~pi024 & pi152;
  assign new_new_n743__ = pi022 & ~pi150;
  assign new_new_n744__ = pi023 & ~pi151;
  assign new_new_n745__ = ~pi022 & pi150;
  assign new_new_n746__ = pi021 & ~pi149;
  assign new_new_n747__ = ~pi021 & pi149;
  assign new_new_n748__ = pi020 & ~pi148;
  assign new_new_n749__ = ~pi020 & pi148;
  assign new_new_n750__ = pi019 & ~pi147;
  assign new_new_n751__ = ~pi019 & pi147;
  assign new_new_n752__ = ~pi018 & pi146;
  assign new_new_n753__ = pi016 & ~pi144;
  assign new_new_n754__ = ~pi015 & pi143;
  assign new_new_n755__ = ~pi014 & pi142;
  assign new_new_n756__ = pi013 & ~pi141;
  assign new_new_n757__ = pi012 & ~pi140;
  assign new_new_n758__ = ~pi011 & pi139;
  assign new_new_n759__ = ~pi009 & pi137;
  assign new_new_n760__ = ~pi010 & pi138;
  assign new_new_n761__ = pi008 & ~pi136;
  assign new_new_n762__ = pi009 & ~pi137;
  assign new_new_n763__ = ~pi008 & pi136;
  assign new_new_n764__ = pi007 & ~pi135;
  assign new_new_n765__ = ~pi007 & pi135;
  assign new_new_n766__ = ~pi006 & pi134;
  assign new_new_n767__ = pi006 & ~pi134;
  assign new_new_n768__ = pi005 & ~pi133;
  assign new_new_n769__ = ~pi004 & pi132;
  assign new_new_n770__ = ~pi005 & pi133;
  assign new_new_n771__ = pi004 & ~pi132;
  assign new_new_n772__ = ~pi003 & pi131;
  assign new_new_n773__ = pi002 & ~pi130;
  assign new_new_n774__ = pi003 & ~pi131;
  assign new_new_n775__ = ~pi002 & pi130;
  assign new_new_n776__ = ~pi001 & pi129;
  assign new_new_n777__ = pi000 & ~pi128;
  assign new_new_n778__ = ~new_new_n776__ & new_new_n777__;
  assign new_new_n779__ = pi001 & ~pi129;
  assign new_new_n780__ = ~new_new_n778__ & ~new_new_n779__;
  assign new_new_n781__ = ~new_new_n775__ & ~new_new_n780__;
  assign new_new_n782__ = ~new_new_n773__ & ~new_new_n774__;
  assign new_new_n783__ = ~new_new_n781__ & new_new_n782__;
  assign new_new_n784__ = ~new_new_n772__ & ~new_new_n783__;
  assign new_new_n785__ = ~new_new_n771__ & ~new_new_n784__;
  assign new_new_n786__ = ~new_new_n769__ & ~new_new_n770__;
  assign new_new_n787__ = ~new_new_n785__ & new_new_n786__;
  assign new_new_n788__ = ~new_new_n767__ & ~new_new_n768__;
  assign new_new_n789__ = ~new_new_n787__ & new_new_n788__;
  assign new_new_n790__ = ~new_new_n765__ & ~new_new_n766__;
  assign new_new_n791__ = ~new_new_n789__ & new_new_n790__;
  assign new_new_n792__ = ~new_new_n764__ & ~new_new_n791__;
  assign new_new_n793__ = ~new_new_n763__ & ~new_new_n792__;
  assign new_new_n794__ = ~new_new_n761__ & ~new_new_n762__;
  assign new_new_n795__ = ~new_new_n793__ & new_new_n794__;
  assign new_new_n796__ = ~new_new_n759__ & ~new_new_n760__;
  assign new_new_n797__ = ~new_new_n795__ & new_new_n796__;
  assign new_new_n798__ = pi010 & ~pi138;
  assign new_new_n799__ = pi011 & ~pi139;
  assign new_new_n800__ = ~new_new_n798__ & ~new_new_n799__;
  assign new_new_n801__ = ~new_new_n797__ & new_new_n800__;
  assign new_new_n802__ = ~new_new_n758__ & ~new_new_n801__;
  assign new_new_n803__ = ~new_new_n757__ & ~new_new_n802__;
  assign new_new_n804__ = ~pi012 & pi140;
  assign new_new_n805__ = ~pi013 & pi141;
  assign new_new_n806__ = ~new_new_n804__ & ~new_new_n805__;
  assign new_new_n807__ = ~new_new_n803__ & new_new_n806__;
  assign new_new_n808__ = ~new_new_n756__ & ~new_new_n807__;
  assign new_new_n809__ = ~new_new_n755__ & ~new_new_n808__;
  assign new_new_n810__ = pi014 & ~pi142;
  assign new_new_n811__ = pi015 & ~pi143;
  assign new_new_n812__ = ~new_new_n810__ & ~new_new_n811__;
  assign new_new_n813__ = ~new_new_n809__ & new_new_n812__;
  assign new_new_n814__ = ~new_new_n754__ & ~new_new_n813__;
  assign new_new_n815__ = ~new_new_n753__ & ~new_new_n814__;
  assign new_new_n816__ = ~pi016 & pi144;
  assign new_new_n817__ = ~pi017 & pi145;
  assign new_new_n818__ = ~new_new_n816__ & ~new_new_n817__;
  assign new_new_n819__ = ~new_new_n815__ & new_new_n818__;
  assign new_new_n820__ = pi018 & ~pi146;
  assign new_new_n821__ = pi017 & ~pi145;
  assign new_new_n822__ = ~new_new_n820__ & ~new_new_n821__;
  assign new_new_n823__ = ~new_new_n819__ & new_new_n822__;
  assign new_new_n824__ = ~new_new_n751__ & ~new_new_n752__;
  assign new_new_n825__ = ~new_new_n823__ & new_new_n824__;
  assign new_new_n826__ = ~new_new_n750__ & ~new_new_n825__;
  assign new_new_n827__ = ~new_new_n749__ & ~new_new_n826__;
  assign new_new_n828__ = ~new_new_n748__ & ~new_new_n827__;
  assign new_new_n829__ = ~new_new_n747__ & ~new_new_n828__;
  assign new_new_n830__ = ~new_new_n746__ & ~new_new_n829__;
  assign new_new_n831__ = ~new_new_n745__ & ~new_new_n830__;
  assign new_new_n832__ = ~new_new_n743__ & ~new_new_n744__;
  assign new_new_n833__ = ~new_new_n831__ & new_new_n832__;
  assign new_new_n834__ = ~new_new_n741__ & ~new_new_n742__;
  assign new_new_n835__ = ~new_new_n833__ & new_new_n834__;
  assign new_new_n836__ = pi024 & ~pi152;
  assign new_new_n837__ = pi025 & ~pi153;
  assign new_new_n838__ = ~new_new_n836__ & ~new_new_n837__;
  assign new_new_n839__ = ~new_new_n835__ & new_new_n838__;
  assign new_new_n840__ = ~pi026 & pi154;
  assign new_new_n841__ = ~pi025 & pi153;
  assign new_new_n842__ = ~new_new_n840__ & ~new_new_n841__;
  assign new_new_n843__ = ~new_new_n839__ & new_new_n842__;
  assign new_new_n844__ = ~new_new_n740__ & ~new_new_n843__;
  assign new_new_n845__ = ~new_new_n739__ & ~new_new_n844__;
  assign new_new_n846__ = pi027 & ~pi155;
  assign new_new_n847__ = pi028 & ~pi156;
  assign new_new_n848__ = ~new_new_n846__ & ~new_new_n847__;
  assign new_new_n849__ = ~new_new_n845__ & new_new_n848__;
  assign new_new_n850__ = ~pi028 & pi156;
  assign new_new_n851__ = ~pi029 & pi157;
  assign new_new_n852__ = ~new_new_n850__ & ~new_new_n851__;
  assign new_new_n853__ = ~new_new_n849__ & new_new_n852__;
  assign new_new_n854__ = ~new_new_n738__ & ~new_new_n853__;
  assign new_new_n855__ = ~new_new_n737__ & ~new_new_n854__;
  assign new_new_n856__ = pi030 & ~pi158;
  assign new_new_n857__ = pi031 & ~pi159;
  assign new_new_n858__ = ~new_new_n856__ & ~new_new_n857__;
  assign new_new_n859__ = ~new_new_n855__ & new_new_n858__;
  assign new_new_n860__ = ~pi032 & pi160;
  assign new_new_n861__ = ~pi031 & pi159;
  assign new_new_n862__ = ~new_new_n860__ & ~new_new_n861__;
  assign new_new_n863__ = ~new_new_n859__ & new_new_n862__;
  assign new_new_n864__ = ~new_new_n735__ & ~new_new_n736__;
  assign new_new_n865__ = ~new_new_n863__ & new_new_n864__;
  assign new_new_n866__ = ~new_new_n734__ & ~new_new_n865__;
  assign new_new_n867__ = ~new_new_n733__ & ~new_new_n866__;
  assign new_new_n868__ = ~new_new_n731__ & ~new_new_n732__;
  assign new_new_n869__ = ~new_new_n867__ & new_new_n868__;
  assign new_new_n870__ = ~new_new_n729__ & ~new_new_n730__;
  assign new_new_n871__ = ~new_new_n869__ & new_new_n870__;
  assign new_new_n872__ = ~pi036 & pi164;
  assign new_new_n873__ = ~pi037 & pi165;
  assign new_new_n874__ = ~new_new_n872__ & ~new_new_n873__;
  assign new_new_n875__ = ~new_new_n871__ & new_new_n874__;
  assign new_new_n876__ = pi038 & ~pi166;
  assign new_new_n877__ = pi037 & ~pi165;
  assign new_new_n878__ = ~new_new_n876__ & ~new_new_n877__;
  assign new_new_n879__ = ~new_new_n875__ & new_new_n878__;
  assign new_new_n880__ = ~new_new_n728__ & ~new_new_n879__;
  assign new_new_n881__ = ~new_new_n727__ & ~new_new_n880__;
  assign new_new_n882__ = ~pi040 & pi168;
  assign new_new_n883__ = ~pi042 & pi170;
  assign new_new_n884__ = ~pi041 & pi169;
  assign new_new_n885__ = ~new_new_n883__ & ~new_new_n884__;
  assign new_new_n886__ = ~pi039 & pi167;
  assign new_new_n887__ = ~new_new_n882__ & ~new_new_n886__;
  assign new_new_n888__ = new_new_n885__ & new_new_n887__;
  assign new_new_n889__ = ~new_new_n881__ & new_new_n888__;
  assign new_new_n890__ = pi042 & ~pi170;
  assign new_new_n891__ = pi040 & ~pi168;
  assign new_new_n892__ = pi041 & ~pi169;
  assign new_new_n893__ = ~new_new_n891__ & ~new_new_n892__;
  assign new_new_n894__ = new_new_n885__ & ~new_new_n893__;
  assign new_new_n895__ = pi043 & ~pi171;
  assign new_new_n896__ = ~new_new_n890__ & ~new_new_n895__;
  assign new_new_n897__ = ~new_new_n894__ & new_new_n896__;
  assign new_new_n898__ = ~new_new_n889__ & new_new_n897__;
  assign new_new_n899__ = ~pi044 & pi172;
  assign new_new_n900__ = ~pi046 & pi174;
  assign new_new_n901__ = ~pi045 & pi173;
  assign new_new_n902__ = ~new_new_n900__ & ~new_new_n901__;
  assign new_new_n903__ = ~pi043 & pi171;
  assign new_new_n904__ = ~new_new_n899__ & ~new_new_n903__;
  assign new_new_n905__ = new_new_n902__ & new_new_n904__;
  assign new_new_n906__ = ~new_new_n898__ & new_new_n905__;
  assign new_new_n907__ = pi046 & ~pi174;
  assign new_new_n908__ = pi044 & ~pi172;
  assign new_new_n909__ = pi045 & ~pi173;
  assign new_new_n910__ = ~new_new_n908__ & ~new_new_n909__;
  assign new_new_n911__ = new_new_n902__ & ~new_new_n910__;
  assign new_new_n912__ = pi047 & ~pi175;
  assign new_new_n913__ = ~new_new_n907__ & ~new_new_n912__;
  assign new_new_n914__ = ~new_new_n911__ & new_new_n913__;
  assign new_new_n915__ = ~new_new_n906__ & new_new_n914__;
  assign new_new_n916__ = ~pi047 & pi175;
  assign new_new_n917__ = ~pi048 & pi176;
  assign new_new_n918__ = ~new_new_n916__ & ~new_new_n917__;
  assign new_new_n919__ = ~new_new_n915__ & new_new_n918__;
  assign new_new_n920__ = pi049 & ~pi177;
  assign new_new_n921__ = pi048 & ~pi176;
  assign new_new_n922__ = ~new_new_n920__ & ~new_new_n921__;
  assign new_new_n923__ = ~new_new_n919__ & new_new_n922__;
  assign new_new_n924__ = ~new_new_n725__ & ~new_new_n726__;
  assign new_new_n925__ = ~new_new_n923__ & new_new_n924__;
  assign new_new_n926__ = ~new_new_n724__ & ~new_new_n925__;
  assign new_new_n927__ = ~new_new_n723__ & ~new_new_n926__;
  assign new_new_n928__ = ~new_new_n722__ & ~new_new_n927__;
  assign new_new_n929__ = ~new_new_n721__ & ~new_new_n928__;
  assign new_new_n930__ = ~new_new_n720__ & ~new_new_n929__;
  assign new_new_n931__ = ~new_new_n719__ & ~new_new_n930__;
  assign new_new_n932__ = ~new_new_n717__ & ~new_new_n718__;
  assign new_new_n933__ = ~new_new_n931__ & new_new_n932__;
  assign new_new_n934__ = ~new_new_n715__ & ~new_new_n716__;
  assign new_new_n935__ = ~new_new_n933__ & new_new_n934__;
  assign new_new_n936__ = pi055 & ~pi183;
  assign new_new_n937__ = pi056 & ~pi184;
  assign new_new_n938__ = ~new_new_n936__ & ~new_new_n937__;
  assign new_new_n939__ = ~new_new_n935__ & new_new_n938__;
  assign new_new_n940__ = ~new_new_n714__ & ~new_new_n939__;
  assign new_new_n941__ = ~new_new_n713__ & ~new_new_n940__;
  assign new_new_n942__ = ~pi057 & pi185;
  assign new_new_n943__ = ~pi058 & pi186;
  assign new_new_n944__ = ~new_new_n942__ & ~new_new_n943__;
  assign new_new_n945__ = ~new_new_n941__ & new_new_n944__;
  assign new_new_n946__ = pi059 & ~pi187;
  assign new_new_n947__ = pi058 & ~pi186;
  assign new_new_n948__ = ~new_new_n946__ & ~new_new_n947__;
  assign new_new_n949__ = ~new_new_n945__ & new_new_n948__;
  assign new_new_n950__ = ~pi060 & pi188;
  assign new_new_n951__ = ~pi062 & pi190;
  assign new_new_n952__ = ~pi061 & pi189;
  assign new_new_n953__ = ~new_new_n951__ & ~new_new_n952__;
  assign new_new_n954__ = ~pi059 & pi187;
  assign new_new_n955__ = ~new_new_n950__ & ~new_new_n954__;
  assign new_new_n956__ = new_new_n953__ & new_new_n955__;
  assign new_new_n957__ = ~new_new_n949__ & new_new_n956__;
  assign new_new_n958__ = pi062 & ~pi190;
  assign new_new_n959__ = pi060 & ~pi188;
  assign new_new_n960__ = pi061 & ~pi189;
  assign new_new_n961__ = ~new_new_n959__ & ~new_new_n960__;
  assign new_new_n962__ = new_new_n953__ & ~new_new_n961__;
  assign new_new_n963__ = pi063 & ~pi191;
  assign new_new_n964__ = ~new_new_n958__ & ~new_new_n963__;
  assign new_new_n965__ = ~new_new_n962__ & new_new_n964__;
  assign new_new_n966__ = ~new_new_n957__ & new_new_n965__;
  assign new_new_n967__ = ~new_new_n712__ & ~new_new_n966__;
  assign new_new_n968__ = ~new_new_n711__ & ~new_new_n967__;
  assign new_new_n969__ = ~new_new_n709__ & ~new_new_n710__;
  assign new_new_n970__ = ~new_new_n968__ & new_new_n969__;
  assign new_new_n971__ = ~new_new_n707__ & ~new_new_n708__;
  assign new_new_n972__ = ~new_new_n970__ & new_new_n971__;
  assign new_new_n973__ = ~new_new_n706__ & ~new_new_n972__;
  assign new_new_n974__ = ~new_new_n705__ & ~new_new_n973__;
  assign new_new_n975__ = ~pi068 & pi196;
  assign new_new_n976__ = ~pi070 & pi198;
  assign new_new_n977__ = ~pi069 & pi197;
  assign new_new_n978__ = ~new_new_n976__ & ~new_new_n977__;
  assign new_new_n979__ = ~pi067 & pi195;
  assign new_new_n980__ = ~new_new_n975__ & ~new_new_n979__;
  assign new_new_n981__ = new_new_n978__ & new_new_n980__;
  assign new_new_n982__ = ~new_new_n974__ & new_new_n981__;
  assign new_new_n983__ = pi070 & ~pi198;
  assign new_new_n984__ = pi068 & ~pi196;
  assign new_new_n985__ = pi069 & ~pi197;
  assign new_new_n986__ = ~new_new_n984__ & ~new_new_n985__;
  assign new_new_n987__ = new_new_n978__ & ~new_new_n986__;
  assign new_new_n988__ = pi071 & ~pi199;
  assign new_new_n989__ = ~new_new_n983__ & ~new_new_n988__;
  assign new_new_n990__ = ~new_new_n987__ & new_new_n989__;
  assign new_new_n991__ = ~new_new_n982__ & new_new_n990__;
  assign new_new_n992__ = ~new_new_n704__ & ~new_new_n991__;
  assign new_new_n993__ = ~new_new_n703__ & ~new_new_n992__;
  assign new_new_n994__ = ~new_new_n702__ & ~new_new_n993__;
  assign new_new_n995__ = ~new_new_n701__ & ~new_new_n994__;
  assign new_new_n996__ = ~new_new_n700__ & ~new_new_n995__;
  assign new_new_n997__ = ~new_new_n699__ & ~new_new_n996__;
  assign new_new_n998__ = ~new_new_n698__ & ~new_new_n997__;
  assign new_new_n999__ = ~new_new_n697__ & ~new_new_n998__;
  assign new_new_n1000__ = ~new_new_n696__ & ~new_new_n999__;
  assign new_new_n1001__ = ~new_new_n695__ & ~new_new_n1000__;
  assign new_new_n1002__ = ~new_new_n694__ & ~new_new_n1001__;
  assign new_new_n1003__ = ~new_new_n693__ & ~new_new_n1002__;
  assign new_new_n1004__ = ~new_new_n691__ & ~new_new_n692__;
  assign new_new_n1005__ = ~new_new_n1003__ & new_new_n1004__;
  assign new_new_n1006__ = ~new_new_n689__ & ~new_new_n690__;
  assign new_new_n1007__ = ~new_new_n1005__ & new_new_n1006__;
  assign new_new_n1008__ = ~new_new_n687__ & ~new_new_n688__;
  assign new_new_n1009__ = ~new_new_n1007__ & new_new_n1008__;
  assign new_new_n1010__ = ~new_new_n686__ & ~new_new_n1009__;
  assign new_new_n1011__ = ~new_new_n685__ & ~new_new_n1010__;
  assign new_new_n1012__ = ~new_new_n684__ & ~new_new_n1011__;
  assign new_new_n1013__ = ~new_new_n683__ & ~new_new_n1012__;
  assign new_new_n1014__ = ~new_new_n682__ & ~new_new_n1013__;
  assign new_new_n1015__ = ~new_new_n681__ & ~new_new_n1014__;
  assign new_new_n1016__ = ~new_new_n680__ & ~new_new_n1015__;
  assign new_new_n1017__ = ~new_new_n679__ & ~new_new_n1016__;
  assign new_new_n1018__ = ~new_new_n678__ & ~new_new_n1017__;
  assign new_new_n1019__ = ~new_new_n677__ & ~new_new_n1018__;
  assign new_new_n1020__ = ~new_new_n676__ & ~new_new_n1019__;
  assign new_new_n1021__ = ~new_new_n675__ & ~new_new_n1020__;
  assign new_new_n1022__ = ~new_new_n674__ & ~new_new_n1021__;
  assign new_new_n1023__ = ~new_new_n673__ & ~new_new_n1022__;
  assign new_new_n1024__ = ~new_new_n671__ & ~new_new_n672__;
  assign new_new_n1025__ = ~new_new_n1023__ & new_new_n1024__;
  assign new_new_n1026__ = ~new_new_n669__ & ~new_new_n670__;
  assign new_new_n1027__ = ~new_new_n1025__ & new_new_n1026__;
  assign new_new_n1028__ = pi089 & ~pi217;
  assign new_new_n1029__ = pi090 & ~pi218;
  assign new_new_n1030__ = ~new_new_n1028__ & ~new_new_n1029__;
  assign new_new_n1031__ = ~new_new_n1027__ & new_new_n1030__;
  assign new_new_n1032__ = ~new_new_n668__ & ~new_new_n1031__;
  assign new_new_n1033__ = ~new_new_n667__ & ~new_new_n1032__;
  assign new_new_n1034__ = ~pi091 & pi219;
  assign new_new_n1035__ = ~pi092 & pi220;
  assign new_new_n1036__ = ~new_new_n1034__ & ~new_new_n1035__;
  assign new_new_n1037__ = ~new_new_n1033__ & new_new_n1036__;
  assign new_new_n1038__ = ~new_new_n666__ & ~new_new_n1037__;
  assign new_new_n1039__ = ~new_new_n665__ & ~new_new_n1038__;
  assign new_new_n1040__ = pi093 & ~pi221;
  assign new_new_n1041__ = pi094 & ~pi222;
  assign new_new_n1042__ = ~new_new_n1040__ & ~new_new_n1041__;
  assign new_new_n1043__ = ~new_new_n1039__ & new_new_n1042__;
  assign new_new_n1044__ = ~new_new_n664__ & ~new_new_n1043__;
  assign new_new_n1045__ = ~new_new_n663__ & ~new_new_n1044__;
  assign new_new_n1046__ = ~pi095 & pi223;
  assign new_new_n1047__ = ~pi096 & pi224;
  assign new_new_n1048__ = ~new_new_n1046__ & ~new_new_n1047__;
  assign new_new_n1049__ = ~new_new_n1045__ & new_new_n1048__;
  assign new_new_n1050__ = pi097 & ~pi225;
  assign new_new_n1051__ = pi096 & ~pi224;
  assign new_new_n1052__ = ~new_new_n1050__ & ~new_new_n1051__;
  assign new_new_n1053__ = ~new_new_n1049__ & new_new_n1052__;
  assign new_new_n1054__ = ~new_new_n662__ & ~new_new_n1053__;
  assign new_new_n1055__ = ~new_new_n661__ & ~new_new_n1054__;
  assign new_new_n1056__ = ~pi098 & pi226;
  assign new_new_n1057__ = ~pi099 & pi227;
  assign new_new_n1058__ = ~new_new_n1056__ & ~new_new_n1057__;
  assign new_new_n1059__ = ~new_new_n1055__ & new_new_n1058__;
  assign new_new_n1060__ = pi099 & ~pi227;
  assign new_new_n1061__ = pi100 & ~pi228;
  assign new_new_n1062__ = ~new_new_n1060__ & ~new_new_n1061__;
  assign new_new_n1063__ = ~new_new_n1059__ & new_new_n1062__;
  assign new_new_n1064__ = ~pi101 & pi229;
  assign new_new_n1065__ = ~pi100 & pi228;
  assign new_new_n1066__ = ~new_new_n1064__ & ~new_new_n1065__;
  assign new_new_n1067__ = ~new_new_n1063__ & new_new_n1066__;
  assign new_new_n1068__ = ~new_new_n660__ & ~new_new_n1067__;
  assign new_new_n1069__ = ~new_new_n659__ & ~new_new_n1068__;
  assign new_new_n1070__ = pi102 & ~pi230;
  assign new_new_n1071__ = pi103 & ~pi231;
  assign new_new_n1072__ = ~new_new_n1070__ & ~new_new_n1071__;
  assign new_new_n1073__ = ~new_new_n1069__ & new_new_n1072__;
  assign new_new_n1074__ = ~pi103 & pi231;
  assign new_new_n1075__ = ~pi104 & pi232;
  assign new_new_n1076__ = ~new_new_n1074__ & ~new_new_n1075__;
  assign new_new_n1077__ = ~new_new_n1073__ & new_new_n1076__;
  assign new_new_n1078__ = pi105 & ~pi233;
  assign new_new_n1079__ = pi104 & ~pi232;
  assign new_new_n1080__ = ~new_new_n1078__ & ~new_new_n1079__;
  assign new_new_n1081__ = ~new_new_n1077__ & new_new_n1080__;
  assign new_new_n1082__ = ~new_new_n658__ & ~new_new_n1081__;
  assign new_new_n1083__ = ~new_new_n657__ & ~new_new_n1082__;
  assign new_new_n1084__ = ~pi106 & pi234;
  assign new_new_n1085__ = ~pi107 & pi235;
  assign new_new_n1086__ = ~new_new_n1084__ & ~new_new_n1085__;
  assign new_new_n1087__ = ~new_new_n1083__ & new_new_n1086__;
  assign new_new_n1088__ = pi107 & ~pi235;
  assign new_new_n1089__ = pi108 & ~pi236;
  assign new_new_n1090__ = ~new_new_n1088__ & ~new_new_n1089__;
  assign new_new_n1091__ = ~new_new_n1087__ & new_new_n1090__;
  assign new_new_n1092__ = ~pi109 & pi237;
  assign new_new_n1093__ = ~pi108 & pi236;
  assign new_new_n1094__ = ~new_new_n1092__ & ~new_new_n1093__;
  assign new_new_n1095__ = ~new_new_n1091__ & new_new_n1094__;
  assign new_new_n1096__ = ~new_new_n656__ & ~new_new_n1095__;
  assign new_new_n1097__ = ~new_new_n655__ & ~new_new_n1096__;
  assign new_new_n1098__ = pi110 & ~pi238;
  assign new_new_n1099__ = pi111 & ~pi239;
  assign new_new_n1100__ = ~new_new_n1098__ & ~new_new_n1099__;
  assign new_new_n1101__ = ~new_new_n1097__ & new_new_n1100__;
  assign new_new_n1102__ = ~pi111 & pi239;
  assign new_new_n1103__ = ~pi112 & pi240;
  assign new_new_n1104__ = ~new_new_n1102__ & ~new_new_n1103__;
  assign new_new_n1105__ = ~new_new_n1101__ & new_new_n1104__;
  assign new_new_n1106__ = pi113 & ~pi241;
  assign new_new_n1107__ = pi112 & ~pi240;
  assign new_new_n1108__ = ~new_new_n1106__ & ~new_new_n1107__;
  assign new_new_n1109__ = ~new_new_n1105__ & new_new_n1108__;
  assign new_new_n1110__ = ~new_new_n654__ & ~new_new_n1109__;
  assign new_new_n1111__ = ~new_new_n653__ & ~new_new_n1110__;
  assign new_new_n1112__ = ~pi114 & pi242;
  assign new_new_n1113__ = ~pi115 & pi243;
  assign new_new_n1114__ = ~new_new_n1112__ & ~new_new_n1113__;
  assign new_new_n1115__ = ~new_new_n1111__ & new_new_n1114__;
  assign new_new_n1116__ = pi115 & ~pi243;
  assign new_new_n1117__ = pi116 & ~pi244;
  assign new_new_n1118__ = ~new_new_n1116__ & ~new_new_n1117__;
  assign new_new_n1119__ = ~new_new_n1115__ & new_new_n1118__;
  assign new_new_n1120__ = ~new_new_n652__ & ~new_new_n1119__;
  assign new_new_n1121__ = ~new_new_n651__ & ~new_new_n1120__;
  assign new_new_n1122__ = ~pi117 & pi245;
  assign new_new_n1123__ = ~pi118 & pi246;
  assign new_new_n1124__ = ~new_new_n1122__ & ~new_new_n1123__;
  assign new_new_n1125__ = ~new_new_n1121__ & new_new_n1124__;
  assign new_new_n1126__ = pi119 & ~pi247;
  assign new_new_n1127__ = pi118 & ~pi246;
  assign new_new_n1128__ = ~new_new_n1126__ & ~new_new_n1127__;
  assign new_new_n1129__ = ~new_new_n1125__ & new_new_n1128__;
  assign new_new_n1130__ = ~new_new_n649__ & ~new_new_n650__;
  assign new_new_n1131__ = ~new_new_n1129__ & new_new_n1130__;
  assign new_new_n1132__ = ~new_new_n648__ & ~new_new_n1131__;
  assign new_new_n1133__ = ~new_new_n647__ & ~new_new_n1132__;
  assign new_new_n1134__ = ~new_new_n646__ & ~new_new_n1133__;
  assign new_new_n1135__ = ~new_new_n645__ & ~new_new_n1134__;
  assign new_new_n1136__ = ~new_new_n643__ & ~new_new_n644__;
  assign new_new_n1137__ = ~new_new_n1135__ & new_new_n1136__;
  assign new_new_n1138__ = ~pi124 & pi252;
  assign new_new_n1139__ = ~pi126 & pi254;
  assign new_new_n1140__ = ~pi125 & pi253;
  assign new_new_n1141__ = ~new_new_n1139__ & ~new_new_n1140__;
  assign new_new_n1142__ = ~pi123 & pi251;
  assign new_new_n1143__ = ~new_new_n1138__ & ~new_new_n1142__;
  assign new_new_n1144__ = new_new_n1141__ & new_new_n1143__;
  assign new_new_n1145__ = ~new_new_n1137__ & new_new_n1144__;
  assign new_new_n1146__ = pi126 & ~pi254;
  assign new_new_n1147__ = pi124 & ~pi252;
  assign new_new_n1148__ = pi125 & ~pi253;
  assign new_new_n1149__ = ~new_new_n1147__ & ~new_new_n1148__;
  assign new_new_n1150__ = new_new_n1141__ & ~new_new_n1149__;
  assign new_new_n1151__ = ~new_new_n1146__ & ~new_new_n1150__;
  assign new_new_n1152__ = ~new_new_n1145__ & new_new_n1151__;
  assign new_new_n1153__ = pi127 & ~pi255;
  assign new_new_n1154__ = ~new_new_n1152__ & ~new_new_n1153__;
  assign new_new_n1155__ = ~pi127 & pi255;
  assign new_new_n1156__ = ~new_new_n1154__ & ~new_new_n1155__;
  assign new_new_n1157__ = pi000 & ~new_new_n1156__;
  assign new_new_n1158__ = pi128 & new_new_n1156__;
  assign new_new_n1159__ = ~new_new_n1157__ & ~new_new_n1158__;
  assign new_new_n1160__ = pi383 & pi511;
  assign new_new_n1161__ = pi378 & ~pi506;
  assign new_new_n1162__ = pi379 & ~pi507;
  assign new_new_n1163__ = ~pi377 & pi505;
  assign new_new_n1164__ = ~pi378 & pi506;
  assign new_new_n1165__ = pi377 & ~pi505;
  assign new_new_n1166__ = ~pi376 & pi504;
  assign new_new_n1167__ = pi376 & ~pi504;
  assign new_new_n1168__ = ~pi375 & pi503;
  assign new_new_n1169__ = pi375 & ~pi503;
  assign new_new_n1170__ = ~pi374 & pi502;
  assign new_new_n1171__ = pi374 & ~pi502;
  assign new_new_n1172__ = ~pi373 & pi501;
  assign new_new_n1173__ = pi373 & ~pi501;
  assign new_new_n1174__ = pi372 & ~pi500;
  assign new_new_n1175__ = ~pi369 & pi497;
  assign new_new_n1176__ = ~pi370 & pi498;
  assign new_new_n1177__ = pi368 & ~pi496;
  assign new_new_n1178__ = pi369 & ~pi497;
  assign new_new_n1179__ = ~pi368 & pi496;
  assign new_new_n1180__ = pi367 & ~pi495;
  assign new_new_n1181__ = ~pi367 & pi495;
  assign new_new_n1182__ = ~pi366 & pi494;
  assign new_new_n1183__ = pi364 & ~pi492;
  assign new_new_n1184__ = ~pi363 & pi491;
  assign new_new_n1185__ = ~pi362 & pi490;
  assign new_new_n1186__ = pi361 & ~pi489;
  assign new_new_n1187__ = pi360 & ~pi488;
  assign new_new_n1188__ = ~pi359 & pi487;
  assign new_new_n1189__ = ~pi357 & pi485;
  assign new_new_n1190__ = ~pi358 & pi486;
  assign new_new_n1191__ = pi356 & ~pi484;
  assign new_new_n1192__ = pi357 & ~pi485;
  assign new_new_n1193__ = ~pi356 & pi484;
  assign new_new_n1194__ = pi355 & ~pi483;
  assign new_new_n1195__ = ~pi355 & pi483;
  assign new_new_n1196__ = ~pi354 & pi482;
  assign new_new_n1197__ = pi351 & ~pi479;
  assign new_new_n1198__ = pi352 & ~pi480;
  assign new_new_n1199__ = ~pi350 & pi478;
  assign new_new_n1200__ = ~pi351 & pi479;
  assign new_new_n1201__ = pi350 & ~pi478;
  assign new_new_n1202__ = ~pi349 & pi477;
  assign new_new_n1203__ = pi349 & ~pi477;
  assign new_new_n1204__ = pi348 & ~pi476;
  assign new_new_n1205__ = ~pi346 & pi474;
  assign new_new_n1206__ = pi345 & ~pi473;
  assign new_new_n1207__ = pi344 & ~pi472;
  assign new_new_n1208__ = ~pi343 & pi471;
  assign new_new_n1209__ = ~pi341 & pi469;
  assign new_new_n1210__ = ~pi342 & pi470;
  assign new_new_n1211__ = pi340 & ~pi468;
  assign new_new_n1212__ = pi341 & ~pi469;
  assign new_new_n1213__ = ~pi340 & pi468;
  assign new_new_n1214__ = pi339 & ~pi467;
  assign new_new_n1215__ = ~pi339 & pi467;
  assign new_new_n1216__ = ~pi338 & pi466;
  assign new_new_n1217__ = ~pi335 & pi463;
  assign new_new_n1218__ = pi334 & ~pi462;
  assign new_new_n1219__ = ~pi332 & pi460;
  assign new_new_n1220__ = pi331 & ~pi459;
  assign new_new_n1221__ = ~pi329 & pi457;
  assign new_new_n1222__ = pi328 & ~pi456;
  assign new_new_n1223__ = pi321 & ~pi449;
  assign new_new_n1224__ = ~pi320 & pi448;
  assign new_new_n1225__ = pi314 & ~pi442;
  assign new_new_n1226__ = pi315 & ~pi443;
  assign new_new_n1227__ = ~pi314 & pi442;
  assign new_new_n1228__ = pi313 & ~pi441;
  assign new_new_n1229__ = ~pi313 & pi441;
  assign new_new_n1230__ = ~pi312 & pi440;
  assign new_new_n1231__ = pi311 & ~pi439;
  assign new_new_n1232__ = pi312 & ~pi440;
  assign new_new_n1233__ = ~pi310 & pi438;
  assign new_new_n1234__ = ~pi311 & pi439;
  assign new_new_n1235__ = pi310 & ~pi438;
  assign new_new_n1236__ = ~pi309 & pi437;
  assign new_new_n1237__ = pi309 & ~pi437;
  assign new_new_n1238__ = ~pi308 & pi436;
  assign new_new_n1239__ = pi308 & ~pi436;
  assign new_new_n1240__ = ~pi307 & pi435;
  assign new_new_n1241__ = pi307 & ~pi435;
  assign new_new_n1242__ = ~pi306 & pi434;
  assign new_new_n1243__ = pi306 & ~pi434;
  assign new_new_n1244__ = ~pi305 & pi433;
  assign new_new_n1245__ = pi305 & ~pi433;
  assign new_new_n1246__ = ~pi304 & pi432;
  assign new_new_n1247__ = pi304 & ~pi432;
  assign new_new_n1248__ = ~pi303 & pi431;
  assign new_new_n1249__ = ~pi294 & pi422;
  assign new_new_n1250__ = pi293 & ~pi421;
  assign new_new_n1251__ = pi292 & ~pi420;
  assign new_new_n1252__ = ~pi291 & pi419;
  assign new_new_n1253__ = ~pi289 & pi417;
  assign new_new_n1254__ = ~pi290 & pi418;
  assign new_new_n1255__ = pi288 & ~pi416;
  assign new_new_n1256__ = pi289 & ~pi417;
  assign new_new_n1257__ = ~pi288 & pi416;
  assign new_new_n1258__ = pi287 & ~pi415;
  assign new_new_n1259__ = ~pi287 & pi415;
  assign new_new_n1260__ = ~pi286 & pi414;
  assign new_new_n1261__ = ~pi283 & pi411;
  assign new_new_n1262__ = pi282 & ~pi410;
  assign new_new_n1263__ = ~pi279 & pi407;
  assign new_new_n1264__ = ~pi280 & pi408;
  assign new_new_n1265__ = pi278 & ~pi406;
  assign new_new_n1266__ = pi279 & ~pi407;
  assign new_new_n1267__ = ~pi278 & pi406;
  assign new_new_n1268__ = pi277 & ~pi405;
  assign new_new_n1269__ = ~pi277 & pi405;
  assign new_new_n1270__ = pi276 & ~pi404;
  assign new_new_n1271__ = ~pi276 & pi404;
  assign new_new_n1272__ = pi275 & ~pi403;
  assign new_new_n1273__ = ~pi275 & pi403;
  assign new_new_n1274__ = ~pi274 & pi402;
  assign new_new_n1275__ = ~pi273 & pi401;
  assign new_new_n1276__ = pi272 & ~pi400;
  assign new_new_n1277__ = pi271 & ~pi399;
  assign new_new_n1278__ = ~pi270 & pi398;
  assign new_new_n1279__ = ~pi269 & pi397;
  assign new_new_n1280__ = pi268 & ~pi396;
  assign new_new_n1281__ = pi267 & ~pi395;
  assign new_new_n1282__ = ~pi266 & pi394;
  assign new_new_n1283__ = pi265 & ~pi393;
  assign new_new_n1284__ = pi266 & ~pi394;
  assign new_new_n1285__ = ~pi264 & pi392;
  assign new_new_n1286__ = ~pi265 & pi393;
  assign new_new_n1287__ = pi264 & ~pi392;
  assign new_new_n1288__ = ~pi263 & pi391;
  assign new_new_n1289__ = pi263 & ~pi391;
  assign new_new_n1290__ = ~pi262 & pi390;
  assign new_new_n1291__ = pi262 & ~pi390;
  assign new_new_n1292__ = ~pi261 & pi389;
  assign new_new_n1293__ = pi261 & ~pi389;
  assign new_new_n1294__ = ~pi260 & pi388;
  assign new_new_n1295__ = pi260 & ~pi388;
  assign new_new_n1296__ = ~pi259 & pi387;
  assign new_new_n1297__ = pi259 & ~pi387;
  assign new_new_n1298__ = pi258 & ~pi386;
  assign new_new_n1299__ = pi256 & ~pi384;
  assign new_new_n1300__ = pi257 & ~pi385;
  assign new_new_n1301__ = ~new_new_n1299__ & ~new_new_n1300__;
  assign new_new_n1302__ = ~pi257 & pi385;
  assign new_new_n1303__ = ~pi258 & pi386;
  assign new_new_n1304__ = ~new_new_n1302__ & ~new_new_n1303__;
  assign new_new_n1305__ = ~new_new_n1301__ & new_new_n1304__;
  assign new_new_n1306__ = ~new_new_n1297__ & ~new_new_n1298__;
  assign new_new_n1307__ = ~new_new_n1305__ & new_new_n1306__;
  assign new_new_n1308__ = ~new_new_n1296__ & ~new_new_n1307__;
  assign new_new_n1309__ = ~new_new_n1295__ & ~new_new_n1308__;
  assign new_new_n1310__ = ~new_new_n1294__ & ~new_new_n1309__;
  assign new_new_n1311__ = ~new_new_n1293__ & ~new_new_n1310__;
  assign new_new_n1312__ = ~new_new_n1292__ & ~new_new_n1311__;
  assign new_new_n1313__ = ~new_new_n1291__ & ~new_new_n1312__;
  assign new_new_n1314__ = ~new_new_n1290__ & ~new_new_n1313__;
  assign new_new_n1315__ = ~new_new_n1289__ & ~new_new_n1314__;
  assign new_new_n1316__ = ~new_new_n1288__ & ~new_new_n1315__;
  assign new_new_n1317__ = ~new_new_n1287__ & ~new_new_n1316__;
  assign new_new_n1318__ = ~new_new_n1285__ & ~new_new_n1286__;
  assign new_new_n1319__ = ~new_new_n1317__ & new_new_n1318__;
  assign new_new_n1320__ = ~new_new_n1283__ & ~new_new_n1284__;
  assign new_new_n1321__ = ~new_new_n1319__ & new_new_n1320__;
  assign new_new_n1322__ = ~new_new_n1282__ & ~new_new_n1321__;
  assign new_new_n1323__ = ~new_new_n1281__ & ~new_new_n1322__;
  assign new_new_n1324__ = ~pi267 & pi395;
  assign new_new_n1325__ = ~pi268 & pi396;
  assign new_new_n1326__ = ~new_new_n1324__ & ~new_new_n1325__;
  assign new_new_n1327__ = ~new_new_n1323__ & new_new_n1326__;
  assign new_new_n1328__ = ~new_new_n1280__ & ~new_new_n1327__;
  assign new_new_n1329__ = ~new_new_n1279__ & ~new_new_n1328__;
  assign new_new_n1330__ = pi269 & ~pi397;
  assign new_new_n1331__ = pi270 & ~pi398;
  assign new_new_n1332__ = ~new_new_n1330__ & ~new_new_n1331__;
  assign new_new_n1333__ = ~new_new_n1329__ & new_new_n1332__;
  assign new_new_n1334__ = ~new_new_n1278__ & ~new_new_n1333__;
  assign new_new_n1335__ = ~new_new_n1277__ & ~new_new_n1334__;
  assign new_new_n1336__ = ~pi271 & pi399;
  assign new_new_n1337__ = ~pi272 & pi400;
  assign new_new_n1338__ = ~new_new_n1336__ & ~new_new_n1337__;
  assign new_new_n1339__ = ~new_new_n1335__ & new_new_n1338__;
  assign new_new_n1340__ = ~new_new_n1276__ & ~new_new_n1339__;
  assign new_new_n1341__ = ~new_new_n1275__ & ~new_new_n1340__;
  assign new_new_n1342__ = pi273 & ~pi401;
  assign new_new_n1343__ = pi274 & ~pi402;
  assign new_new_n1344__ = ~new_new_n1342__ & ~new_new_n1343__;
  assign new_new_n1345__ = ~new_new_n1341__ & new_new_n1344__;
  assign new_new_n1346__ = ~new_new_n1273__ & ~new_new_n1274__;
  assign new_new_n1347__ = ~new_new_n1345__ & new_new_n1346__;
  assign new_new_n1348__ = ~new_new_n1272__ & ~new_new_n1347__;
  assign new_new_n1349__ = ~new_new_n1271__ & ~new_new_n1348__;
  assign new_new_n1350__ = ~new_new_n1270__ & ~new_new_n1349__;
  assign new_new_n1351__ = ~new_new_n1269__ & ~new_new_n1350__;
  assign new_new_n1352__ = ~new_new_n1268__ & ~new_new_n1351__;
  assign new_new_n1353__ = ~new_new_n1267__ & ~new_new_n1352__;
  assign new_new_n1354__ = ~new_new_n1265__ & ~new_new_n1266__;
  assign new_new_n1355__ = ~new_new_n1353__ & new_new_n1354__;
  assign new_new_n1356__ = ~new_new_n1263__ & ~new_new_n1264__;
  assign new_new_n1357__ = ~new_new_n1355__ & new_new_n1356__;
  assign new_new_n1358__ = pi280 & ~pi408;
  assign new_new_n1359__ = pi281 & ~pi409;
  assign new_new_n1360__ = ~new_new_n1358__ & ~new_new_n1359__;
  assign new_new_n1361__ = ~new_new_n1357__ & new_new_n1360__;
  assign new_new_n1362__ = ~pi282 & pi410;
  assign new_new_n1363__ = ~pi281 & pi409;
  assign new_new_n1364__ = ~new_new_n1362__ & ~new_new_n1363__;
  assign new_new_n1365__ = ~new_new_n1361__ & new_new_n1364__;
  assign new_new_n1366__ = ~new_new_n1262__ & ~new_new_n1365__;
  assign new_new_n1367__ = ~new_new_n1261__ & ~new_new_n1366__;
  assign new_new_n1368__ = pi283 & ~pi411;
  assign new_new_n1369__ = pi284 & ~pi412;
  assign new_new_n1370__ = ~new_new_n1368__ & ~new_new_n1369__;
  assign new_new_n1371__ = ~new_new_n1367__ & new_new_n1370__;
  assign new_new_n1372__ = ~pi284 & pi412;
  assign new_new_n1373__ = ~pi285 & pi413;
  assign new_new_n1374__ = ~new_new_n1372__ & ~new_new_n1373__;
  assign new_new_n1375__ = ~new_new_n1371__ & new_new_n1374__;
  assign new_new_n1376__ = pi286 & ~pi414;
  assign new_new_n1377__ = pi285 & ~pi413;
  assign new_new_n1378__ = ~new_new_n1376__ & ~new_new_n1377__;
  assign new_new_n1379__ = ~new_new_n1375__ & new_new_n1378__;
  assign new_new_n1380__ = ~new_new_n1259__ & ~new_new_n1260__;
  assign new_new_n1381__ = ~new_new_n1379__ & new_new_n1380__;
  assign new_new_n1382__ = ~new_new_n1258__ & ~new_new_n1381__;
  assign new_new_n1383__ = ~new_new_n1257__ & ~new_new_n1382__;
  assign new_new_n1384__ = ~new_new_n1255__ & ~new_new_n1256__;
  assign new_new_n1385__ = ~new_new_n1383__ & new_new_n1384__;
  assign new_new_n1386__ = ~new_new_n1253__ & ~new_new_n1254__;
  assign new_new_n1387__ = ~new_new_n1385__ & new_new_n1386__;
  assign new_new_n1388__ = pi290 & ~pi418;
  assign new_new_n1389__ = pi291 & ~pi419;
  assign new_new_n1390__ = ~new_new_n1388__ & ~new_new_n1389__;
  assign new_new_n1391__ = ~new_new_n1387__ & new_new_n1390__;
  assign new_new_n1392__ = ~new_new_n1252__ & ~new_new_n1391__;
  assign new_new_n1393__ = ~new_new_n1251__ & ~new_new_n1392__;
  assign new_new_n1394__ = ~pi292 & pi420;
  assign new_new_n1395__ = ~pi293 & pi421;
  assign new_new_n1396__ = ~new_new_n1394__ & ~new_new_n1395__;
  assign new_new_n1397__ = ~new_new_n1393__ & new_new_n1396__;
  assign new_new_n1398__ = ~new_new_n1250__ & ~new_new_n1397__;
  assign new_new_n1399__ = ~new_new_n1249__ & ~new_new_n1398__;
  assign new_new_n1400__ = pi294 & ~pi422;
  assign new_new_n1401__ = pi295 & ~pi423;
  assign new_new_n1402__ = ~new_new_n1400__ & ~new_new_n1401__;
  assign new_new_n1403__ = ~new_new_n1399__ & new_new_n1402__;
  assign new_new_n1404__ = ~pi296 & pi424;
  assign new_new_n1405__ = ~pi298 & pi426;
  assign new_new_n1406__ = ~pi297 & pi425;
  assign new_new_n1407__ = ~new_new_n1405__ & ~new_new_n1406__;
  assign new_new_n1408__ = ~pi295 & pi423;
  assign new_new_n1409__ = ~new_new_n1404__ & ~new_new_n1408__;
  assign new_new_n1410__ = new_new_n1407__ & new_new_n1409__;
  assign new_new_n1411__ = ~new_new_n1403__ & new_new_n1410__;
  assign new_new_n1412__ = pi298 & ~pi426;
  assign new_new_n1413__ = pi296 & ~pi424;
  assign new_new_n1414__ = pi297 & ~pi425;
  assign new_new_n1415__ = ~new_new_n1413__ & ~new_new_n1414__;
  assign new_new_n1416__ = new_new_n1407__ & ~new_new_n1415__;
  assign new_new_n1417__ = pi299 & ~pi427;
  assign new_new_n1418__ = ~new_new_n1412__ & ~new_new_n1417__;
  assign new_new_n1419__ = ~new_new_n1416__ & new_new_n1418__;
  assign new_new_n1420__ = ~new_new_n1411__ & new_new_n1419__;
  assign new_new_n1421__ = ~pi299 & pi427;
  assign new_new_n1422__ = ~pi302 & pi430;
  assign new_new_n1423__ = ~pi301 & pi429;
  assign new_new_n1424__ = ~new_new_n1422__ & ~new_new_n1423__;
  assign new_new_n1425__ = ~pi300 & pi428;
  assign new_new_n1426__ = ~new_new_n1421__ & ~new_new_n1425__;
  assign new_new_n1427__ = new_new_n1424__ & new_new_n1426__;
  assign new_new_n1428__ = ~new_new_n1420__ & new_new_n1427__;
  assign new_new_n1429__ = pi302 & ~pi430;
  assign new_new_n1430__ = pi300 & ~pi428;
  assign new_new_n1431__ = pi301 & ~pi429;
  assign new_new_n1432__ = ~new_new_n1430__ & ~new_new_n1431__;
  assign new_new_n1433__ = new_new_n1424__ & ~new_new_n1432__;
  assign new_new_n1434__ = pi303 & ~pi431;
  assign new_new_n1435__ = ~new_new_n1429__ & ~new_new_n1434__;
  assign new_new_n1436__ = ~new_new_n1433__ & new_new_n1435__;
  assign new_new_n1437__ = ~new_new_n1428__ & new_new_n1436__;
  assign new_new_n1438__ = ~new_new_n1248__ & ~new_new_n1437__;
  assign new_new_n1439__ = ~new_new_n1247__ & ~new_new_n1438__;
  assign new_new_n1440__ = ~new_new_n1246__ & ~new_new_n1439__;
  assign new_new_n1441__ = ~new_new_n1245__ & ~new_new_n1440__;
  assign new_new_n1442__ = ~new_new_n1244__ & ~new_new_n1441__;
  assign new_new_n1443__ = ~new_new_n1243__ & ~new_new_n1442__;
  assign new_new_n1444__ = ~new_new_n1242__ & ~new_new_n1443__;
  assign new_new_n1445__ = ~new_new_n1241__ & ~new_new_n1444__;
  assign new_new_n1446__ = ~new_new_n1240__ & ~new_new_n1445__;
  assign new_new_n1447__ = ~new_new_n1239__ & ~new_new_n1446__;
  assign new_new_n1448__ = ~new_new_n1238__ & ~new_new_n1447__;
  assign new_new_n1449__ = ~new_new_n1237__ & ~new_new_n1448__;
  assign new_new_n1450__ = ~new_new_n1236__ & ~new_new_n1449__;
  assign new_new_n1451__ = ~new_new_n1235__ & ~new_new_n1450__;
  assign new_new_n1452__ = ~new_new_n1233__ & ~new_new_n1234__;
  assign new_new_n1453__ = ~new_new_n1451__ & new_new_n1452__;
  assign new_new_n1454__ = ~new_new_n1231__ & ~new_new_n1232__;
  assign new_new_n1455__ = ~new_new_n1453__ & new_new_n1454__;
  assign new_new_n1456__ = ~new_new_n1229__ & ~new_new_n1230__;
  assign new_new_n1457__ = ~new_new_n1455__ & new_new_n1456__;
  assign new_new_n1458__ = ~new_new_n1228__ & ~new_new_n1457__;
  assign new_new_n1459__ = ~new_new_n1227__ & ~new_new_n1458__;
  assign new_new_n1460__ = ~new_new_n1225__ & ~new_new_n1226__;
  assign new_new_n1461__ = ~new_new_n1459__ & new_new_n1460__;
  assign new_new_n1462__ = ~pi316 & pi444;
  assign new_new_n1463__ = ~pi318 & pi446;
  assign new_new_n1464__ = ~pi317 & pi445;
  assign new_new_n1465__ = ~new_new_n1463__ & ~new_new_n1464__;
  assign new_new_n1466__ = ~pi315 & pi443;
  assign new_new_n1467__ = ~new_new_n1462__ & ~new_new_n1466__;
  assign new_new_n1468__ = new_new_n1465__ & new_new_n1467__;
  assign new_new_n1469__ = ~new_new_n1461__ & new_new_n1468__;
  assign new_new_n1470__ = pi318 & ~pi446;
  assign new_new_n1471__ = pi316 & ~pi444;
  assign new_new_n1472__ = pi317 & ~pi445;
  assign new_new_n1473__ = ~new_new_n1471__ & ~new_new_n1472__;
  assign new_new_n1474__ = new_new_n1465__ & ~new_new_n1473__;
  assign new_new_n1475__ = ~new_new_n1470__ & ~new_new_n1474__;
  assign new_new_n1476__ = ~new_new_n1469__ & new_new_n1475__;
  assign new_new_n1477__ = ~pi319 & pi447;
  assign new_new_n1478__ = ~new_new_n1476__ & ~new_new_n1477__;
  assign new_new_n1479__ = pi319 & ~pi447;
  assign new_new_n1480__ = pi320 & ~pi448;
  assign new_new_n1481__ = ~new_new_n1479__ & ~new_new_n1480__;
  assign new_new_n1482__ = ~new_new_n1478__ & new_new_n1481__;
  assign new_new_n1483__ = ~new_new_n1224__ & ~new_new_n1482__;
  assign new_new_n1484__ = ~new_new_n1223__ & ~new_new_n1483__;
  assign new_new_n1485__ = ~pi321 & pi449;
  assign new_new_n1486__ = ~pi322 & pi450;
  assign new_new_n1487__ = ~new_new_n1485__ & ~new_new_n1486__;
  assign new_new_n1488__ = ~new_new_n1484__ & new_new_n1487__;
  assign new_new_n1489__ = pi322 & ~pi450;
  assign new_new_n1490__ = pi323 & ~pi451;
  assign new_new_n1491__ = ~new_new_n1489__ & ~new_new_n1490__;
  assign new_new_n1492__ = ~new_new_n1488__ & new_new_n1491__;
  assign new_new_n1493__ = ~pi324 & pi452;
  assign new_new_n1494__ = ~pi326 & pi454;
  assign new_new_n1495__ = ~pi325 & pi453;
  assign new_new_n1496__ = ~new_new_n1494__ & ~new_new_n1495__;
  assign new_new_n1497__ = ~pi323 & pi451;
  assign new_new_n1498__ = ~new_new_n1493__ & ~new_new_n1497__;
  assign new_new_n1499__ = new_new_n1496__ & new_new_n1498__;
  assign new_new_n1500__ = ~new_new_n1492__ & new_new_n1499__;
  assign new_new_n1501__ = pi326 & ~pi454;
  assign new_new_n1502__ = pi324 & ~pi452;
  assign new_new_n1503__ = pi325 & ~pi453;
  assign new_new_n1504__ = ~new_new_n1502__ & ~new_new_n1503__;
  assign new_new_n1505__ = new_new_n1496__ & ~new_new_n1504__;
  assign new_new_n1506__ = pi327 & ~pi455;
  assign new_new_n1507__ = ~new_new_n1501__ & ~new_new_n1506__;
  assign new_new_n1508__ = ~new_new_n1505__ & new_new_n1507__;
  assign new_new_n1509__ = ~new_new_n1500__ & new_new_n1508__;
  assign new_new_n1510__ = ~pi327 & pi455;
  assign new_new_n1511__ = ~pi328 & pi456;
  assign new_new_n1512__ = ~new_new_n1510__ & ~new_new_n1511__;
  assign new_new_n1513__ = ~new_new_n1509__ & new_new_n1512__;
  assign new_new_n1514__ = ~new_new_n1222__ & ~new_new_n1513__;
  assign new_new_n1515__ = ~new_new_n1221__ & ~new_new_n1514__;
  assign new_new_n1516__ = pi329 & ~pi457;
  assign new_new_n1517__ = pi330 & ~pi458;
  assign new_new_n1518__ = ~new_new_n1516__ & ~new_new_n1517__;
  assign new_new_n1519__ = ~new_new_n1515__ & new_new_n1518__;
  assign new_new_n1520__ = ~pi330 & pi458;
  assign new_new_n1521__ = ~pi331 & pi459;
  assign new_new_n1522__ = ~new_new_n1520__ & ~new_new_n1521__;
  assign new_new_n1523__ = ~new_new_n1519__ & new_new_n1522__;
  assign new_new_n1524__ = ~new_new_n1220__ & ~new_new_n1523__;
  assign new_new_n1525__ = ~new_new_n1219__ & ~new_new_n1524__;
  assign new_new_n1526__ = pi332 & ~pi460;
  assign new_new_n1527__ = pi333 & ~pi461;
  assign new_new_n1528__ = ~new_new_n1526__ & ~new_new_n1527__;
  assign new_new_n1529__ = ~new_new_n1525__ & new_new_n1528__;
  assign new_new_n1530__ = ~pi334 & pi462;
  assign new_new_n1531__ = ~pi333 & pi461;
  assign new_new_n1532__ = ~new_new_n1530__ & ~new_new_n1531__;
  assign new_new_n1533__ = ~new_new_n1529__ & new_new_n1532__;
  assign new_new_n1534__ = ~new_new_n1218__ & ~new_new_n1533__;
  assign new_new_n1535__ = ~new_new_n1217__ & ~new_new_n1534__;
  assign new_new_n1536__ = pi335 & ~pi463;
  assign new_new_n1537__ = pi336 & ~pi464;
  assign new_new_n1538__ = ~new_new_n1536__ & ~new_new_n1537__;
  assign new_new_n1539__ = ~new_new_n1535__ & new_new_n1538__;
  assign new_new_n1540__ = ~pi336 & pi464;
  assign new_new_n1541__ = ~pi337 & pi465;
  assign new_new_n1542__ = ~new_new_n1540__ & ~new_new_n1541__;
  assign new_new_n1543__ = ~new_new_n1539__ & new_new_n1542__;
  assign new_new_n1544__ = pi338 & ~pi466;
  assign new_new_n1545__ = pi337 & ~pi465;
  assign new_new_n1546__ = ~new_new_n1544__ & ~new_new_n1545__;
  assign new_new_n1547__ = ~new_new_n1543__ & new_new_n1546__;
  assign new_new_n1548__ = ~new_new_n1215__ & ~new_new_n1216__;
  assign new_new_n1549__ = ~new_new_n1547__ & new_new_n1548__;
  assign new_new_n1550__ = ~new_new_n1214__ & ~new_new_n1549__;
  assign new_new_n1551__ = ~new_new_n1213__ & ~new_new_n1550__;
  assign new_new_n1552__ = ~new_new_n1211__ & ~new_new_n1212__;
  assign new_new_n1553__ = ~new_new_n1551__ & new_new_n1552__;
  assign new_new_n1554__ = ~new_new_n1209__ & ~new_new_n1210__;
  assign new_new_n1555__ = ~new_new_n1553__ & new_new_n1554__;
  assign new_new_n1556__ = pi342 & ~pi470;
  assign new_new_n1557__ = pi343 & ~pi471;
  assign new_new_n1558__ = ~new_new_n1556__ & ~new_new_n1557__;
  assign new_new_n1559__ = ~new_new_n1555__ & new_new_n1558__;
  assign new_new_n1560__ = ~new_new_n1208__ & ~new_new_n1559__;
  assign new_new_n1561__ = ~new_new_n1207__ & ~new_new_n1560__;
  assign new_new_n1562__ = ~pi344 & pi472;
  assign new_new_n1563__ = ~pi345 & pi473;
  assign new_new_n1564__ = ~new_new_n1562__ & ~new_new_n1563__;
  assign new_new_n1565__ = ~new_new_n1561__ & new_new_n1564__;
  assign new_new_n1566__ = ~new_new_n1206__ & ~new_new_n1565__;
  assign new_new_n1567__ = ~new_new_n1205__ & ~new_new_n1566__;
  assign new_new_n1568__ = pi346 & ~pi474;
  assign new_new_n1569__ = pi347 & ~pi475;
  assign new_new_n1570__ = ~new_new_n1568__ & ~new_new_n1569__;
  assign new_new_n1571__ = ~new_new_n1567__ & new_new_n1570__;
  assign new_new_n1572__ = ~pi348 & pi476;
  assign new_new_n1573__ = ~pi347 & pi475;
  assign new_new_n1574__ = ~new_new_n1572__ & ~new_new_n1573__;
  assign new_new_n1575__ = ~new_new_n1571__ & new_new_n1574__;
  assign new_new_n1576__ = ~new_new_n1203__ & ~new_new_n1204__;
  assign new_new_n1577__ = ~new_new_n1575__ & new_new_n1576__;
  assign new_new_n1578__ = ~new_new_n1202__ & ~new_new_n1577__;
  assign new_new_n1579__ = ~new_new_n1201__ & ~new_new_n1578__;
  assign new_new_n1580__ = ~new_new_n1199__ & ~new_new_n1200__;
  assign new_new_n1581__ = ~new_new_n1579__ & new_new_n1580__;
  assign new_new_n1582__ = ~new_new_n1197__ & ~new_new_n1198__;
  assign new_new_n1583__ = ~new_new_n1581__ & new_new_n1582__;
  assign new_new_n1584__ = ~pi352 & pi480;
  assign new_new_n1585__ = ~pi353 & pi481;
  assign new_new_n1586__ = ~new_new_n1584__ & ~new_new_n1585__;
  assign new_new_n1587__ = ~new_new_n1583__ & new_new_n1586__;
  assign new_new_n1588__ = pi354 & ~pi482;
  assign new_new_n1589__ = pi353 & ~pi481;
  assign new_new_n1590__ = ~new_new_n1588__ & ~new_new_n1589__;
  assign new_new_n1591__ = ~new_new_n1587__ & new_new_n1590__;
  assign new_new_n1592__ = ~new_new_n1195__ & ~new_new_n1196__;
  assign new_new_n1593__ = ~new_new_n1591__ & new_new_n1592__;
  assign new_new_n1594__ = ~new_new_n1194__ & ~new_new_n1593__;
  assign new_new_n1595__ = ~new_new_n1193__ & ~new_new_n1594__;
  assign new_new_n1596__ = ~new_new_n1191__ & ~new_new_n1192__;
  assign new_new_n1597__ = ~new_new_n1595__ & new_new_n1596__;
  assign new_new_n1598__ = ~new_new_n1189__ & ~new_new_n1190__;
  assign new_new_n1599__ = ~new_new_n1597__ & new_new_n1598__;
  assign new_new_n1600__ = pi358 & ~pi486;
  assign new_new_n1601__ = pi359 & ~pi487;
  assign new_new_n1602__ = ~new_new_n1600__ & ~new_new_n1601__;
  assign new_new_n1603__ = ~new_new_n1599__ & new_new_n1602__;
  assign new_new_n1604__ = ~new_new_n1188__ & ~new_new_n1603__;
  assign new_new_n1605__ = ~new_new_n1187__ & ~new_new_n1604__;
  assign new_new_n1606__ = ~pi360 & pi488;
  assign new_new_n1607__ = ~pi361 & pi489;
  assign new_new_n1608__ = ~new_new_n1606__ & ~new_new_n1607__;
  assign new_new_n1609__ = ~new_new_n1605__ & new_new_n1608__;
  assign new_new_n1610__ = ~new_new_n1186__ & ~new_new_n1609__;
  assign new_new_n1611__ = ~new_new_n1185__ & ~new_new_n1610__;
  assign new_new_n1612__ = pi362 & ~pi490;
  assign new_new_n1613__ = pi363 & ~pi491;
  assign new_new_n1614__ = ~new_new_n1612__ & ~new_new_n1613__;
  assign new_new_n1615__ = ~new_new_n1611__ & new_new_n1614__;
  assign new_new_n1616__ = ~new_new_n1184__ & ~new_new_n1615__;
  assign new_new_n1617__ = ~new_new_n1183__ & ~new_new_n1616__;
  assign new_new_n1618__ = ~pi364 & pi492;
  assign new_new_n1619__ = ~pi365 & pi493;
  assign new_new_n1620__ = ~new_new_n1618__ & ~new_new_n1619__;
  assign new_new_n1621__ = ~new_new_n1617__ & new_new_n1620__;
  assign new_new_n1622__ = pi366 & ~pi494;
  assign new_new_n1623__ = pi365 & ~pi493;
  assign new_new_n1624__ = ~new_new_n1622__ & ~new_new_n1623__;
  assign new_new_n1625__ = ~new_new_n1621__ & new_new_n1624__;
  assign new_new_n1626__ = ~new_new_n1181__ & ~new_new_n1182__;
  assign new_new_n1627__ = ~new_new_n1625__ & new_new_n1626__;
  assign new_new_n1628__ = ~new_new_n1180__ & ~new_new_n1627__;
  assign new_new_n1629__ = ~new_new_n1179__ & ~new_new_n1628__;
  assign new_new_n1630__ = ~new_new_n1177__ & ~new_new_n1178__;
  assign new_new_n1631__ = ~new_new_n1629__ & new_new_n1630__;
  assign new_new_n1632__ = ~new_new_n1175__ & ~new_new_n1176__;
  assign new_new_n1633__ = ~new_new_n1631__ & new_new_n1632__;
  assign new_new_n1634__ = pi370 & ~pi498;
  assign new_new_n1635__ = pi371 & ~pi499;
  assign new_new_n1636__ = ~new_new_n1634__ & ~new_new_n1635__;
  assign new_new_n1637__ = ~new_new_n1633__ & new_new_n1636__;
  assign new_new_n1638__ = ~pi372 & pi500;
  assign new_new_n1639__ = ~pi371 & pi499;
  assign new_new_n1640__ = ~new_new_n1638__ & ~new_new_n1639__;
  assign new_new_n1641__ = ~new_new_n1637__ & new_new_n1640__;
  assign new_new_n1642__ = ~new_new_n1173__ & ~new_new_n1174__;
  assign new_new_n1643__ = ~new_new_n1641__ & new_new_n1642__;
  assign new_new_n1644__ = ~new_new_n1172__ & ~new_new_n1643__;
  assign new_new_n1645__ = ~new_new_n1171__ & ~new_new_n1644__;
  assign new_new_n1646__ = ~new_new_n1170__ & ~new_new_n1645__;
  assign new_new_n1647__ = ~new_new_n1169__ & ~new_new_n1646__;
  assign new_new_n1648__ = ~new_new_n1168__ & ~new_new_n1647__;
  assign new_new_n1649__ = ~new_new_n1167__ & ~new_new_n1648__;
  assign new_new_n1650__ = ~new_new_n1166__ & ~new_new_n1649__;
  assign new_new_n1651__ = ~new_new_n1165__ & ~new_new_n1650__;
  assign new_new_n1652__ = ~new_new_n1163__ & ~new_new_n1164__;
  assign new_new_n1653__ = ~new_new_n1651__ & new_new_n1652__;
  assign new_new_n1654__ = ~new_new_n1161__ & ~new_new_n1162__;
  assign new_new_n1655__ = ~new_new_n1653__ & new_new_n1654__;
  assign new_new_n1656__ = ~pi380 & pi508;
  assign new_new_n1657__ = ~pi382 & pi510;
  assign new_new_n1658__ = ~pi381 & pi509;
  assign new_new_n1659__ = ~new_new_n1657__ & ~new_new_n1658__;
  assign new_new_n1660__ = ~pi379 & pi507;
  assign new_new_n1661__ = ~new_new_n1656__ & ~new_new_n1660__;
  assign new_new_n1662__ = new_new_n1659__ & new_new_n1661__;
  assign new_new_n1663__ = ~new_new_n1655__ & new_new_n1662__;
  assign new_new_n1664__ = pi382 & ~pi510;
  assign new_new_n1665__ = pi380 & ~pi508;
  assign new_new_n1666__ = pi381 & ~pi509;
  assign new_new_n1667__ = ~new_new_n1665__ & ~new_new_n1666__;
  assign new_new_n1668__ = new_new_n1659__ & ~new_new_n1667__;
  assign new_new_n1669__ = ~new_new_n1664__ & ~new_new_n1668__;
  assign new_new_n1670__ = ~new_new_n1663__ & new_new_n1669__;
  assign new_new_n1671__ = pi383 & ~pi511;
  assign new_new_n1672__ = ~new_new_n1670__ & ~new_new_n1671__;
  assign new_new_n1673__ = ~pi383 & pi511;
  assign new_new_n1674__ = ~new_new_n1672__ & ~new_new_n1673__;
  assign new_new_n1675__ = pi373 & ~new_new_n1674__;
  assign new_new_n1676__ = pi501 & new_new_n1674__;
  assign new_new_n1677__ = ~new_new_n1675__ & ~new_new_n1676__;
  assign new_new_n1678__ = pi372 & ~new_new_n1674__;
  assign new_new_n1679__ = pi500 & new_new_n1674__;
  assign new_new_n1680__ = ~new_new_n1678__ & ~new_new_n1679__;
  assign new_new_n1681__ = pi371 & ~new_new_n1674__;
  assign new_new_n1682__ = pi499 & new_new_n1674__;
  assign new_new_n1683__ = ~new_new_n1681__ & ~new_new_n1682__;
  assign new_new_n1684__ = pi370 & ~new_new_n1674__;
  assign new_new_n1685__ = pi498 & new_new_n1674__;
  assign new_new_n1686__ = ~new_new_n1684__ & ~new_new_n1685__;
  assign new_new_n1687__ = pi369 & ~new_new_n1674__;
  assign new_new_n1688__ = pi497 & new_new_n1674__;
  assign new_new_n1689__ = ~new_new_n1687__ & ~new_new_n1688__;
  assign new_new_n1690__ = pi368 & ~new_new_n1674__;
  assign new_new_n1691__ = pi496 & new_new_n1674__;
  assign new_new_n1692__ = ~new_new_n1690__ & ~new_new_n1691__;
  assign new_new_n1693__ = pi366 & ~new_new_n1674__;
  assign new_new_n1694__ = pi494 & new_new_n1674__;
  assign new_new_n1695__ = ~new_new_n1693__ & ~new_new_n1694__;
  assign new_new_n1696__ = pi365 & ~new_new_n1674__;
  assign new_new_n1697__ = pi493 & new_new_n1674__;
  assign new_new_n1698__ = ~new_new_n1696__ & ~new_new_n1697__;
  assign new_new_n1699__ = pi363 & ~new_new_n1674__;
  assign new_new_n1700__ = pi491 & new_new_n1674__;
  assign new_new_n1701__ = ~new_new_n1699__ & ~new_new_n1700__;
  assign new_new_n1702__ = pi362 & ~new_new_n1674__;
  assign new_new_n1703__ = pi490 & new_new_n1674__;
  assign new_new_n1704__ = ~new_new_n1702__ & ~new_new_n1703__;
  assign new_new_n1705__ = pi359 & ~new_new_n1674__;
  assign new_new_n1706__ = pi487 & new_new_n1674__;
  assign new_new_n1707__ = ~new_new_n1705__ & ~new_new_n1706__;
  assign new_new_n1708__ = pi358 & ~new_new_n1674__;
  assign new_new_n1709__ = pi486 & new_new_n1674__;
  assign new_new_n1710__ = ~new_new_n1708__ & ~new_new_n1709__;
  assign new_new_n1711__ = pi357 & ~new_new_n1674__;
  assign new_new_n1712__ = pi485 & new_new_n1674__;
  assign new_new_n1713__ = ~new_new_n1711__ & ~new_new_n1712__;
  assign new_new_n1714__ = pi356 & ~new_new_n1674__;
  assign new_new_n1715__ = pi484 & new_new_n1674__;
  assign new_new_n1716__ = ~new_new_n1714__ & ~new_new_n1715__;
  assign new_new_n1717__ = pi354 & ~new_new_n1674__;
  assign new_new_n1718__ = pi482 & new_new_n1674__;
  assign new_new_n1719__ = ~new_new_n1717__ & ~new_new_n1718__;
  assign new_new_n1720__ = pi351 & ~new_new_n1674__;
  assign new_new_n1721__ = pi479 & new_new_n1674__;
  assign new_new_n1722__ = ~new_new_n1720__ & ~new_new_n1721__;
  assign new_new_n1723__ = pi350 & ~new_new_n1674__;
  assign new_new_n1724__ = pi478 & new_new_n1674__;
  assign new_new_n1725__ = ~new_new_n1723__ & ~new_new_n1724__;
  assign new_new_n1726__ = pi349 & ~new_new_n1674__;
  assign new_new_n1727__ = pi477 & new_new_n1674__;
  assign new_new_n1728__ = ~new_new_n1726__ & ~new_new_n1727__;
  assign new_new_n1729__ = pi348 & ~new_new_n1674__;
  assign new_new_n1730__ = pi476 & new_new_n1674__;
  assign new_new_n1731__ = ~new_new_n1729__ & ~new_new_n1730__;
  assign new_new_n1732__ = pi347 & ~new_new_n1674__;
  assign new_new_n1733__ = pi475 & new_new_n1674__;
  assign new_new_n1734__ = ~new_new_n1732__ & ~new_new_n1733__;
  assign new_new_n1735__ = pi089 & ~new_new_n1156__;
  assign new_new_n1736__ = pi217 & new_new_n1156__;
  assign new_new_n1737__ = ~new_new_n1735__ & ~new_new_n1736__;
  assign new_new_n1738__ = pi088 & ~new_new_n1156__;
  assign new_new_n1739__ = pi216 & new_new_n1156__;
  assign new_new_n1740__ = ~new_new_n1738__ & ~new_new_n1739__;
  assign new_new_n1741__ = pi087 & ~new_new_n1156__;
  assign new_new_n1742__ = pi215 & new_new_n1156__;
  assign new_new_n1743__ = ~new_new_n1741__ & ~new_new_n1742__;
  assign new_new_n1744__ = pi086 & ~new_new_n1156__;
  assign new_new_n1745__ = pi214 & new_new_n1156__;
  assign new_new_n1746__ = ~new_new_n1744__ & ~new_new_n1745__;
  assign new_new_n1747__ = pi340 & ~new_new_n1674__;
  assign new_new_n1748__ = pi468 & new_new_n1674__;
  assign new_new_n1749__ = ~new_new_n1747__ & ~new_new_n1748__;
  assign new_new_n1750__ = pi081 & ~new_new_n1156__;
  assign new_new_n1751__ = pi209 & new_new_n1156__;
  assign new_new_n1752__ = ~new_new_n1750__ & ~new_new_n1751__;
  assign new_new_n1753__ = pi080 & ~new_new_n1156__;
  assign new_new_n1754__ = pi208 & new_new_n1156__;
  assign new_new_n1755__ = ~new_new_n1753__ & ~new_new_n1754__;
  assign new_new_n1756__ = pi079 & ~new_new_n1156__;
  assign new_new_n1757__ = pi207 & new_new_n1156__;
  assign new_new_n1758__ = ~new_new_n1756__ & ~new_new_n1757__;
  assign new_new_n1759__ = pi078 & ~new_new_n1156__;
  assign new_new_n1760__ = pi206 & new_new_n1156__;
  assign new_new_n1761__ = ~new_new_n1759__ & ~new_new_n1760__;
  assign new_new_n1762__ = pi077 & ~new_new_n1156__;
  assign new_new_n1763__ = pi205 & new_new_n1156__;
  assign new_new_n1764__ = ~new_new_n1762__ & ~new_new_n1763__;
  assign new_new_n1765__ = pi076 & ~new_new_n1156__;
  assign new_new_n1766__ = pi204 & new_new_n1156__;
  assign new_new_n1767__ = ~new_new_n1765__ & ~new_new_n1766__;
  assign new_new_n1768__ = pi075 & ~new_new_n1156__;
  assign new_new_n1769__ = pi203 & new_new_n1156__;
  assign new_new_n1770__ = ~new_new_n1768__ & ~new_new_n1769__;
  assign new_new_n1771__ = pi328 & ~new_new_n1674__;
  assign new_new_n1772__ = pi456 & new_new_n1674__;
  assign new_new_n1773__ = ~new_new_n1771__ & ~new_new_n1772__;
  assign new_new_n1774__ = pi326 & ~new_new_n1674__;
  assign new_new_n1775__ = pi454 & new_new_n1674__;
  assign new_new_n1776__ = ~new_new_n1774__ & ~new_new_n1775__;
  assign new_new_n1777__ = pi323 & ~new_new_n1674__;
  assign new_new_n1778__ = pi451 & new_new_n1674__;
  assign new_new_n1779__ = ~new_new_n1777__ & ~new_new_n1778__;
  assign new_new_n1780__ = pi322 & ~new_new_n1674__;
  assign new_new_n1781__ = pi450 & new_new_n1674__;
  assign new_new_n1782__ = ~new_new_n1780__ & ~new_new_n1781__;
  assign new_new_n1783__ = pi061 & ~new_new_n1156__;
  assign new_new_n1784__ = pi189 & new_new_n1156__;
  assign new_new_n1785__ = ~new_new_n1783__ & ~new_new_n1784__;
  assign new_new_n1786__ = pi058 & ~new_new_n1156__;
  assign new_new_n1787__ = pi186 & new_new_n1156__;
  assign new_new_n1788__ = ~new_new_n1786__ & ~new_new_n1787__;
  assign new_new_n1789__ = pi053 & ~new_new_n1156__;
  assign new_new_n1790__ = pi181 & new_new_n1156__;
  assign new_new_n1791__ = ~new_new_n1789__ & ~new_new_n1790__;
  assign new_new_n1792__ = pi052 & ~new_new_n1156__;
  assign new_new_n1793__ = pi180 & new_new_n1156__;
  assign new_new_n1794__ = ~new_new_n1792__ & ~new_new_n1793__;
  assign new_new_n1795__ = pi051 & ~new_new_n1156__;
  assign new_new_n1796__ = pi179 & new_new_n1156__;
  assign new_new_n1797__ = ~new_new_n1795__ & ~new_new_n1796__;
  assign new_new_n1798__ = pi304 & ~new_new_n1674__;
  assign new_new_n1799__ = pi432 & new_new_n1674__;
  assign new_new_n1800__ = ~new_new_n1798__ & ~new_new_n1799__;
  assign new_new_n1801__ = pi303 & ~new_new_n1674__;
  assign new_new_n1802__ = pi431 & new_new_n1674__;
  assign new_new_n1803__ = ~new_new_n1801__ & ~new_new_n1802__;
  assign new_new_n1804__ = pi045 & ~new_new_n1156__;
  assign new_new_n1805__ = pi173 & new_new_n1156__;
  assign new_new_n1806__ = ~new_new_n1804__ & ~new_new_n1805__;
  assign new_new_n1807__ = pi043 & ~new_new_n1156__;
  assign new_new_n1808__ = pi171 & new_new_n1156__;
  assign new_new_n1809__ = ~new_new_n1807__ & ~new_new_n1808__;
  assign new_new_n1810__ = pi291 & ~new_new_n1674__;
  assign new_new_n1811__ = pi419 & new_new_n1674__;
  assign new_new_n1812__ = ~new_new_n1810__ & ~new_new_n1811__;
  assign new_new_n1813__ = pi033 & ~new_new_n1156__;
  assign new_new_n1814__ = pi161 & new_new_n1156__;
  assign new_new_n1815__ = ~new_new_n1813__ & ~new_new_n1814__;
  assign new_new_n1816__ = pi285 & ~new_new_n1674__;
  assign new_new_n1817__ = pi413 & new_new_n1674__;
  assign new_new_n1818__ = ~new_new_n1816__ & ~new_new_n1817__;
  assign new_new_n1819__ = pi284 & ~new_new_n1674__;
  assign new_new_n1820__ = pi412 & new_new_n1674__;
  assign new_new_n1821__ = ~new_new_n1819__ & ~new_new_n1820__;
  assign new_new_n1822__ = pi026 & ~new_new_n1156__;
  assign new_new_n1823__ = pi154 & new_new_n1156__;
  assign new_new_n1824__ = ~new_new_n1822__ & ~new_new_n1823__;
  assign new_new_n1825__ = pi280 & ~new_new_n1674__;
  assign new_new_n1826__ = pi408 & new_new_n1674__;
  assign new_new_n1827__ = ~new_new_n1825__ & ~new_new_n1826__;
  assign new_new_n1828__ = pi279 & ~new_new_n1674__;
  assign new_new_n1829__ = pi407 & new_new_n1674__;
  assign new_new_n1830__ = ~new_new_n1828__ & ~new_new_n1829__;
  assign new_new_n1831__ = pi278 & ~new_new_n1674__;
  assign new_new_n1832__ = pi406 & new_new_n1674__;
  assign new_new_n1833__ = ~new_new_n1831__ & ~new_new_n1832__;
  assign new_new_n1834__ = pi277 & ~new_new_n1674__;
  assign new_new_n1835__ = pi405 & new_new_n1674__;
  assign new_new_n1836__ = ~new_new_n1834__ & ~new_new_n1835__;
  assign new_new_n1837__ = pi272 & ~new_new_n1674__;
  assign new_new_n1838__ = pi400 & new_new_n1674__;
  assign new_new_n1839__ = ~new_new_n1837__ & ~new_new_n1838__;
  assign new_new_n1840__ = pi271 & ~new_new_n1674__;
  assign new_new_n1841__ = pi399 & new_new_n1674__;
  assign new_new_n1842__ = ~new_new_n1840__ & ~new_new_n1841__;
  assign new_new_n1843__ = pi010 & ~new_new_n1156__;
  assign new_new_n1844__ = pi138 & new_new_n1156__;
  assign new_new_n1845__ = ~new_new_n1843__ & ~new_new_n1844__;
  assign new_new_n1846__ = pi009 & ~new_new_n1156__;
  assign new_new_n1847__ = pi137 & new_new_n1156__;
  assign new_new_n1848__ = ~new_new_n1846__ & ~new_new_n1847__;
  assign new_new_n1849__ = pi007 & ~new_new_n1156__;
  assign new_new_n1850__ = pi135 & new_new_n1156__;
  assign new_new_n1851__ = ~new_new_n1849__ & ~new_new_n1850__;
  assign new_new_n1852__ = pi006 & ~new_new_n1156__;
  assign new_new_n1853__ = pi134 & new_new_n1156__;
  assign new_new_n1854__ = ~new_new_n1852__ & ~new_new_n1853__;
  assign new_new_n1855__ = pi260 & ~new_new_n1674__;
  assign new_new_n1856__ = pi388 & new_new_n1674__;
  assign new_new_n1857__ = ~new_new_n1855__ & ~new_new_n1856__;
  assign new_new_n1858__ = pi259 & ~new_new_n1674__;
  assign new_new_n1859__ = pi387 & new_new_n1674__;
  assign new_new_n1860__ = ~new_new_n1858__ & ~new_new_n1859__;
  assign new_new_n1861__ = pi258 & ~new_new_n1674__;
  assign new_new_n1862__ = pi386 & new_new_n1674__;
  assign new_new_n1863__ = ~new_new_n1861__ & ~new_new_n1862__;
  assign new_new_n1864__ = pi257 & ~new_new_n1674__;
  assign new_new_n1865__ = pi385 & new_new_n1674__;
  assign new_new_n1866__ = ~new_new_n1864__ & ~new_new_n1865__;
  assign new_new_n1867__ = pi256 & ~new_new_n1674__;
  assign new_new_n1868__ = pi384 & new_new_n1674__;
  assign new_new_n1869__ = ~new_new_n1867__ & ~new_new_n1868__;
  assign new_new_n1870__ = ~new_new_n1159__ & new_new_n1869__;
  assign new_new_n1871__ = pi001 & ~new_new_n1156__;
  assign new_new_n1872__ = pi129 & new_new_n1156__;
  assign new_new_n1873__ = ~new_new_n1871__ & ~new_new_n1872__;
  assign new_new_n1874__ = ~new_new_n1870__ & new_new_n1873__;
  assign new_new_n1875__ = new_new_n1866__ & ~new_new_n1874__;
  assign new_new_n1876__ = new_new_n1870__ & ~new_new_n1873__;
  assign new_new_n1877__ = ~new_new_n1875__ & ~new_new_n1876__;
  assign new_new_n1878__ = pi002 & ~new_new_n1156__;
  assign new_new_n1879__ = pi130 & new_new_n1156__;
  assign new_new_n1880__ = ~new_new_n1878__ & ~new_new_n1879__;
  assign new_new_n1881__ = new_new_n1877__ & new_new_n1880__;
  assign new_new_n1882__ = new_new_n1863__ & ~new_new_n1881__;
  assign new_new_n1883__ = ~new_new_n1877__ & ~new_new_n1880__;
  assign new_new_n1884__ = ~new_new_n1882__ & ~new_new_n1883__;
  assign new_new_n1885__ = pi003 & ~new_new_n1156__;
  assign new_new_n1886__ = pi131 & new_new_n1156__;
  assign new_new_n1887__ = ~new_new_n1885__ & ~new_new_n1886__;
  assign new_new_n1888__ = new_new_n1884__ & new_new_n1887__;
  assign new_new_n1889__ = new_new_n1860__ & ~new_new_n1888__;
  assign new_new_n1890__ = ~new_new_n1884__ & ~new_new_n1887__;
  assign new_new_n1891__ = ~new_new_n1889__ & ~new_new_n1890__;
  assign new_new_n1892__ = pi004 & ~new_new_n1156__;
  assign new_new_n1893__ = pi132 & new_new_n1156__;
  assign new_new_n1894__ = ~new_new_n1892__ & ~new_new_n1893__;
  assign new_new_n1895__ = new_new_n1891__ & new_new_n1894__;
  assign new_new_n1896__ = new_new_n1857__ & ~new_new_n1895__;
  assign new_new_n1897__ = ~new_new_n1891__ & ~new_new_n1894__;
  assign new_new_n1898__ = ~new_new_n1896__ & ~new_new_n1897__;
  assign new_new_n1899__ = pi261 & ~new_new_n1674__;
  assign new_new_n1900__ = pi389 & new_new_n1674__;
  assign new_new_n1901__ = ~new_new_n1899__ & ~new_new_n1900__;
  assign new_new_n1902__ = ~new_new_n1898__ & new_new_n1901__;
  assign new_new_n1903__ = new_new_n1898__ & ~new_new_n1901__;
  assign new_new_n1904__ = pi005 & ~new_new_n1156__;
  assign new_new_n1905__ = pi133 & new_new_n1156__;
  assign new_new_n1906__ = ~new_new_n1904__ & ~new_new_n1905__;
  assign new_new_n1907__ = ~new_new_n1903__ & ~new_new_n1906__;
  assign new_new_n1908__ = ~new_new_n1902__ & ~new_new_n1907__;
  assign new_new_n1909__ = pi262 & ~new_new_n1674__;
  assign new_new_n1910__ = pi390 & new_new_n1674__;
  assign new_new_n1911__ = ~new_new_n1909__ & ~new_new_n1910__;
  assign new_new_n1912__ = ~new_new_n1908__ & new_new_n1911__;
  assign new_new_n1913__ = new_new_n1854__ & ~new_new_n1912__;
  assign new_new_n1914__ = new_new_n1908__ & ~new_new_n1911__;
  assign new_new_n1915__ = ~new_new_n1913__ & ~new_new_n1914__;
  assign new_new_n1916__ = pi263 & ~new_new_n1674__;
  assign new_new_n1917__ = pi391 & new_new_n1674__;
  assign new_new_n1918__ = ~new_new_n1916__ & ~new_new_n1917__;
  assign new_new_n1919__ = new_new_n1915__ & new_new_n1918__;
  assign new_new_n1920__ = new_new_n1851__ & ~new_new_n1919__;
  assign new_new_n1921__ = ~new_new_n1915__ & ~new_new_n1918__;
  assign new_new_n1922__ = ~new_new_n1920__ & ~new_new_n1921__;
  assign new_new_n1923__ = pi264 & ~new_new_n1674__;
  assign new_new_n1924__ = pi392 & new_new_n1674__;
  assign new_new_n1925__ = ~new_new_n1923__ & ~new_new_n1924__;
  assign new_new_n1926__ = new_new_n1922__ & new_new_n1925__;
  assign new_new_n1927__ = ~new_new_n1922__ & ~new_new_n1925__;
  assign new_new_n1928__ = pi008 & ~new_new_n1156__;
  assign new_new_n1929__ = pi136 & new_new_n1156__;
  assign new_new_n1930__ = ~new_new_n1928__ & ~new_new_n1929__;
  assign new_new_n1931__ = ~new_new_n1927__ & ~new_new_n1930__;
  assign new_new_n1932__ = ~new_new_n1926__ & ~new_new_n1931__;
  assign new_new_n1933__ = pi265 & ~new_new_n1674__;
  assign new_new_n1934__ = pi393 & new_new_n1674__;
  assign new_new_n1935__ = ~new_new_n1933__ & ~new_new_n1934__;
  assign new_new_n1936__ = ~new_new_n1932__ & new_new_n1935__;
  assign new_new_n1937__ = new_new_n1848__ & ~new_new_n1936__;
  assign new_new_n1938__ = new_new_n1932__ & ~new_new_n1935__;
  assign new_new_n1939__ = ~new_new_n1937__ & ~new_new_n1938__;
  assign new_new_n1940__ = pi266 & ~new_new_n1674__;
  assign new_new_n1941__ = pi394 & new_new_n1674__;
  assign new_new_n1942__ = ~new_new_n1940__ & ~new_new_n1941__;
  assign new_new_n1943__ = new_new_n1939__ & new_new_n1942__;
  assign new_new_n1944__ = new_new_n1845__ & ~new_new_n1943__;
  assign new_new_n1945__ = ~new_new_n1939__ & ~new_new_n1942__;
  assign new_new_n1946__ = ~new_new_n1944__ & ~new_new_n1945__;
  assign new_new_n1947__ = pi267 & ~new_new_n1674__;
  assign new_new_n1948__ = pi395 & new_new_n1674__;
  assign new_new_n1949__ = ~new_new_n1947__ & ~new_new_n1948__;
  assign new_new_n1950__ = new_new_n1946__ & new_new_n1949__;
  assign new_new_n1951__ = ~new_new_n1946__ & ~new_new_n1949__;
  assign new_new_n1952__ = pi011 & ~new_new_n1156__;
  assign new_new_n1953__ = pi139 & new_new_n1156__;
  assign new_new_n1954__ = ~new_new_n1952__ & ~new_new_n1953__;
  assign new_new_n1955__ = ~new_new_n1951__ & ~new_new_n1954__;
  assign new_new_n1956__ = ~new_new_n1950__ & ~new_new_n1955__;
  assign new_new_n1957__ = pi012 & ~new_new_n1156__;
  assign new_new_n1958__ = pi140 & new_new_n1156__;
  assign new_new_n1959__ = ~new_new_n1957__ & ~new_new_n1958__;
  assign new_new_n1960__ = new_new_n1956__ & new_new_n1959__;
  assign new_new_n1961__ = ~new_new_n1956__ & ~new_new_n1959__;
  assign new_new_n1962__ = pi268 & ~new_new_n1674__;
  assign new_new_n1963__ = pi396 & new_new_n1674__;
  assign new_new_n1964__ = ~new_new_n1962__ & ~new_new_n1963__;
  assign new_new_n1965__ = ~new_new_n1961__ & ~new_new_n1964__;
  assign new_new_n1966__ = ~new_new_n1960__ & ~new_new_n1965__;
  assign new_new_n1967__ = pi013 & ~new_new_n1156__;
  assign new_new_n1968__ = pi141 & new_new_n1156__;
  assign new_new_n1969__ = ~new_new_n1967__ & ~new_new_n1968__;
  assign new_new_n1970__ = ~new_new_n1966__ & new_new_n1969__;
  assign new_new_n1971__ = new_new_n1966__ & ~new_new_n1969__;
  assign new_new_n1972__ = pi269 & ~new_new_n1674__;
  assign new_new_n1973__ = pi397 & new_new_n1674__;
  assign new_new_n1974__ = ~new_new_n1972__ & ~new_new_n1973__;
  assign new_new_n1975__ = ~new_new_n1971__ & ~new_new_n1974__;
  assign new_new_n1976__ = ~new_new_n1970__ & ~new_new_n1975__;
  assign new_new_n1977__ = pi014 & ~new_new_n1156__;
  assign new_new_n1978__ = pi142 & new_new_n1156__;
  assign new_new_n1979__ = ~new_new_n1977__ & ~new_new_n1978__;
  assign new_new_n1980__ = ~new_new_n1976__ & new_new_n1979__;
  assign new_new_n1981__ = new_new_n1976__ & ~new_new_n1979__;
  assign new_new_n1982__ = pi270 & ~new_new_n1674__;
  assign new_new_n1983__ = pi398 & new_new_n1674__;
  assign new_new_n1984__ = ~new_new_n1982__ & ~new_new_n1983__;
  assign new_new_n1985__ = ~new_new_n1981__ & ~new_new_n1984__;
  assign new_new_n1986__ = ~new_new_n1980__ & ~new_new_n1985__;
  assign new_new_n1987__ = pi015 & ~new_new_n1156__;
  assign new_new_n1988__ = pi143 & new_new_n1156__;
  assign new_new_n1989__ = ~new_new_n1987__ & ~new_new_n1988__;
  assign new_new_n1990__ = ~new_new_n1986__ & new_new_n1989__;
  assign new_new_n1991__ = new_new_n1842__ & ~new_new_n1990__;
  assign new_new_n1992__ = new_new_n1986__ & ~new_new_n1989__;
  assign new_new_n1993__ = ~new_new_n1991__ & ~new_new_n1992__;
  assign new_new_n1994__ = pi016 & ~new_new_n1156__;
  assign new_new_n1995__ = pi144 & new_new_n1156__;
  assign new_new_n1996__ = ~new_new_n1994__ & ~new_new_n1995__;
  assign new_new_n1997__ = new_new_n1993__ & new_new_n1996__;
  assign new_new_n1998__ = new_new_n1839__ & ~new_new_n1997__;
  assign new_new_n1999__ = ~new_new_n1993__ & ~new_new_n1996__;
  assign new_new_n2000__ = ~new_new_n1998__ & ~new_new_n1999__;
  assign new_new_n2001__ = pi017 & ~new_new_n1156__;
  assign new_new_n2002__ = pi145 & new_new_n1156__;
  assign new_new_n2003__ = ~new_new_n2001__ & ~new_new_n2002__;
  assign new_new_n2004__ = new_new_n2000__ & new_new_n2003__;
  assign new_new_n2005__ = ~new_new_n2000__ & ~new_new_n2003__;
  assign new_new_n2006__ = pi273 & ~new_new_n1674__;
  assign new_new_n2007__ = pi401 & new_new_n1674__;
  assign new_new_n2008__ = ~new_new_n2006__ & ~new_new_n2007__;
  assign new_new_n2009__ = ~new_new_n2005__ & ~new_new_n2008__;
  assign new_new_n2010__ = ~new_new_n2004__ & ~new_new_n2009__;
  assign new_new_n2011__ = pi018 & ~new_new_n1156__;
  assign new_new_n2012__ = pi146 & new_new_n1156__;
  assign new_new_n2013__ = ~new_new_n2011__ & ~new_new_n2012__;
  assign new_new_n2014__ = ~new_new_n2010__ & new_new_n2013__;
  assign new_new_n2015__ = new_new_n2010__ & ~new_new_n2013__;
  assign new_new_n2016__ = pi274 & ~new_new_n1674__;
  assign new_new_n2017__ = pi402 & new_new_n1674__;
  assign new_new_n2018__ = ~new_new_n2016__ & ~new_new_n2017__;
  assign new_new_n2019__ = ~new_new_n2015__ & ~new_new_n2018__;
  assign new_new_n2020__ = ~new_new_n2014__ & ~new_new_n2019__;
  assign new_new_n2021__ = pi019 & ~new_new_n1156__;
  assign new_new_n2022__ = pi147 & new_new_n1156__;
  assign new_new_n2023__ = ~new_new_n2021__ & ~new_new_n2022__;
  assign new_new_n2024__ = ~new_new_n2020__ & new_new_n2023__;
  assign new_new_n2025__ = new_new_n2020__ & ~new_new_n2023__;
  assign new_new_n2026__ = pi275 & ~new_new_n1674__;
  assign new_new_n2027__ = pi403 & new_new_n1674__;
  assign new_new_n2028__ = ~new_new_n2026__ & ~new_new_n2027__;
  assign new_new_n2029__ = ~new_new_n2025__ & ~new_new_n2028__;
  assign new_new_n2030__ = ~new_new_n2024__ & ~new_new_n2029__;
  assign new_new_n2031__ = pi020 & ~new_new_n1156__;
  assign new_new_n2032__ = pi148 & new_new_n1156__;
  assign new_new_n2033__ = ~new_new_n2031__ & ~new_new_n2032__;
  assign new_new_n2034__ = ~new_new_n2030__ & new_new_n2033__;
  assign new_new_n2035__ = new_new_n2030__ & ~new_new_n2033__;
  assign new_new_n2036__ = pi276 & ~new_new_n1674__;
  assign new_new_n2037__ = pi404 & new_new_n1674__;
  assign new_new_n2038__ = ~new_new_n2036__ & ~new_new_n2037__;
  assign new_new_n2039__ = ~new_new_n2035__ & ~new_new_n2038__;
  assign new_new_n2040__ = ~new_new_n2034__ & ~new_new_n2039__;
  assign new_new_n2041__ = pi021 & ~new_new_n1156__;
  assign new_new_n2042__ = pi149 & new_new_n1156__;
  assign new_new_n2043__ = ~new_new_n2041__ & ~new_new_n2042__;
  assign new_new_n2044__ = ~new_new_n2040__ & new_new_n2043__;
  assign new_new_n2045__ = new_new_n1836__ & ~new_new_n2044__;
  assign new_new_n2046__ = new_new_n2040__ & ~new_new_n2043__;
  assign new_new_n2047__ = ~new_new_n2045__ & ~new_new_n2046__;
  assign new_new_n2048__ = pi022 & ~new_new_n1156__;
  assign new_new_n2049__ = pi150 & new_new_n1156__;
  assign new_new_n2050__ = ~new_new_n2048__ & ~new_new_n2049__;
  assign new_new_n2051__ = new_new_n2047__ & new_new_n2050__;
  assign new_new_n2052__ = new_new_n1833__ & ~new_new_n2051__;
  assign new_new_n2053__ = ~new_new_n2047__ & ~new_new_n2050__;
  assign new_new_n2054__ = ~new_new_n2052__ & ~new_new_n2053__;
  assign new_new_n2055__ = pi023 & ~new_new_n1156__;
  assign new_new_n2056__ = pi151 & new_new_n1156__;
  assign new_new_n2057__ = ~new_new_n2055__ & ~new_new_n2056__;
  assign new_new_n2058__ = new_new_n2054__ & new_new_n2057__;
  assign new_new_n2059__ = new_new_n1830__ & ~new_new_n2058__;
  assign new_new_n2060__ = ~new_new_n2054__ & ~new_new_n2057__;
  assign new_new_n2061__ = ~new_new_n2059__ & ~new_new_n2060__;
  assign new_new_n2062__ = pi024 & ~new_new_n1156__;
  assign new_new_n2063__ = pi152 & new_new_n1156__;
  assign new_new_n2064__ = ~new_new_n2062__ & ~new_new_n2063__;
  assign new_new_n2065__ = new_new_n2061__ & new_new_n2064__;
  assign new_new_n2066__ = new_new_n1827__ & ~new_new_n2065__;
  assign new_new_n2067__ = ~new_new_n2061__ & ~new_new_n2064__;
  assign new_new_n2068__ = ~new_new_n2066__ & ~new_new_n2067__;
  assign new_new_n2069__ = pi281 & ~new_new_n1674__;
  assign new_new_n2070__ = pi409 & new_new_n1674__;
  assign new_new_n2071__ = ~new_new_n2069__ & ~new_new_n2070__;
  assign new_new_n2072__ = ~new_new_n2068__ & new_new_n2071__;
  assign new_new_n2073__ = new_new_n2068__ & ~new_new_n2071__;
  assign new_new_n2074__ = pi025 & ~new_new_n1156__;
  assign new_new_n2075__ = pi153 & new_new_n1156__;
  assign new_new_n2076__ = ~new_new_n2074__ & ~new_new_n2075__;
  assign new_new_n2077__ = ~new_new_n2073__ & ~new_new_n2076__;
  assign new_new_n2078__ = ~new_new_n2072__ & ~new_new_n2077__;
  assign new_new_n2079__ = pi282 & ~new_new_n1674__;
  assign new_new_n2080__ = pi410 & new_new_n1674__;
  assign new_new_n2081__ = ~new_new_n2079__ & ~new_new_n2080__;
  assign new_new_n2082__ = ~new_new_n2078__ & new_new_n2081__;
  assign new_new_n2083__ = new_new_n1824__ & ~new_new_n2082__;
  assign new_new_n2084__ = new_new_n2078__ & ~new_new_n2081__;
  assign new_new_n2085__ = ~new_new_n2083__ & ~new_new_n2084__;
  assign new_new_n2086__ = pi027 & ~new_new_n1156__;
  assign new_new_n2087__ = pi155 & new_new_n1156__;
  assign new_new_n2088__ = ~new_new_n2086__ & ~new_new_n2087__;
  assign new_new_n2089__ = ~new_new_n2085__ & new_new_n2088__;
  assign new_new_n2090__ = new_new_n2085__ & ~new_new_n2088__;
  assign new_new_n2091__ = pi283 & ~new_new_n1674__;
  assign new_new_n2092__ = pi411 & new_new_n1674__;
  assign new_new_n2093__ = ~new_new_n2091__ & ~new_new_n2092__;
  assign new_new_n2094__ = ~new_new_n2090__ & ~new_new_n2093__;
  assign new_new_n2095__ = ~new_new_n2089__ & ~new_new_n2094__;
  assign new_new_n2096__ = pi028 & ~new_new_n1156__;
  assign new_new_n2097__ = pi156 & new_new_n1156__;
  assign new_new_n2098__ = ~new_new_n2096__ & ~new_new_n2097__;
  assign new_new_n2099__ = ~new_new_n2095__ & new_new_n2098__;
  assign new_new_n2100__ = new_new_n1821__ & ~new_new_n2099__;
  assign new_new_n2101__ = new_new_n2095__ & ~new_new_n2098__;
  assign new_new_n2102__ = ~new_new_n2100__ & ~new_new_n2101__;
  assign new_new_n2103__ = pi029 & ~new_new_n1156__;
  assign new_new_n2104__ = pi157 & new_new_n1156__;
  assign new_new_n2105__ = ~new_new_n2103__ & ~new_new_n2104__;
  assign new_new_n2106__ = new_new_n2102__ & new_new_n2105__;
  assign new_new_n2107__ = new_new_n1818__ & ~new_new_n2106__;
  assign new_new_n2108__ = ~new_new_n2102__ & ~new_new_n2105__;
  assign new_new_n2109__ = ~new_new_n2107__ & ~new_new_n2108__;
  assign new_new_n2110__ = pi030 & ~new_new_n1156__;
  assign new_new_n2111__ = pi158 & new_new_n1156__;
  assign new_new_n2112__ = ~new_new_n2110__ & ~new_new_n2111__;
  assign new_new_n2113__ = new_new_n2109__ & new_new_n2112__;
  assign new_new_n2114__ = ~new_new_n2109__ & ~new_new_n2112__;
  assign new_new_n2115__ = pi286 & ~new_new_n1674__;
  assign new_new_n2116__ = pi414 & new_new_n1674__;
  assign new_new_n2117__ = ~new_new_n2115__ & ~new_new_n2116__;
  assign new_new_n2118__ = ~new_new_n2114__ & ~new_new_n2117__;
  assign new_new_n2119__ = ~new_new_n2113__ & ~new_new_n2118__;
  assign new_new_n2120__ = pi287 & ~new_new_n1674__;
  assign new_new_n2121__ = pi415 & new_new_n1674__;
  assign new_new_n2122__ = ~new_new_n2120__ & ~new_new_n2121__;
  assign new_new_n2123__ = new_new_n2119__ & new_new_n2122__;
  assign new_new_n2124__ = ~new_new_n2119__ & ~new_new_n2122__;
  assign new_new_n2125__ = pi031 & ~new_new_n1156__;
  assign new_new_n2126__ = pi159 & new_new_n1156__;
  assign new_new_n2127__ = ~new_new_n2125__ & ~new_new_n2126__;
  assign new_new_n2128__ = ~new_new_n2124__ & ~new_new_n2127__;
  assign new_new_n2129__ = ~new_new_n2123__ & ~new_new_n2128__;
  assign new_new_n2130__ = pi288 & ~new_new_n1674__;
  assign new_new_n2131__ = pi416 & new_new_n1674__;
  assign new_new_n2132__ = ~new_new_n2130__ & ~new_new_n2131__;
  assign new_new_n2133__ = ~new_new_n2129__ & new_new_n2132__;
  assign new_new_n2134__ = new_new_n2129__ & ~new_new_n2132__;
  assign new_new_n2135__ = pi032 & ~new_new_n1156__;
  assign new_new_n2136__ = pi160 & new_new_n1156__;
  assign new_new_n2137__ = ~new_new_n2135__ & ~new_new_n2136__;
  assign new_new_n2138__ = ~new_new_n2134__ & ~new_new_n2137__;
  assign new_new_n2139__ = ~new_new_n2133__ & ~new_new_n2138__;
  assign new_new_n2140__ = pi289 & ~new_new_n1674__;
  assign new_new_n2141__ = pi417 & new_new_n1674__;
  assign new_new_n2142__ = ~new_new_n2140__ & ~new_new_n2141__;
  assign new_new_n2143__ = ~new_new_n2139__ & new_new_n2142__;
  assign new_new_n2144__ = new_new_n1815__ & ~new_new_n2143__;
  assign new_new_n2145__ = new_new_n2139__ & ~new_new_n2142__;
  assign new_new_n2146__ = ~new_new_n2144__ & ~new_new_n2145__;
  assign new_new_n2147__ = pi034 & ~new_new_n1156__;
  assign new_new_n2148__ = pi162 & new_new_n1156__;
  assign new_new_n2149__ = ~new_new_n2147__ & ~new_new_n2148__;
  assign new_new_n2150__ = ~new_new_n2146__ & new_new_n2149__;
  assign new_new_n2151__ = new_new_n2146__ & ~new_new_n2149__;
  assign new_new_n2152__ = pi290 & ~new_new_n1674__;
  assign new_new_n2153__ = pi418 & new_new_n1674__;
  assign new_new_n2154__ = ~new_new_n2152__ & ~new_new_n2153__;
  assign new_new_n2155__ = ~new_new_n2151__ & ~new_new_n2154__;
  assign new_new_n2156__ = ~new_new_n2150__ & ~new_new_n2155__;
  assign new_new_n2157__ = pi035 & ~new_new_n1156__;
  assign new_new_n2158__ = pi163 & new_new_n1156__;
  assign new_new_n2159__ = ~new_new_n2157__ & ~new_new_n2158__;
  assign new_new_n2160__ = ~new_new_n2156__ & new_new_n2159__;
  assign new_new_n2161__ = new_new_n1812__ & ~new_new_n2160__;
  assign new_new_n2162__ = new_new_n2156__ & ~new_new_n2159__;
  assign new_new_n2163__ = ~new_new_n2161__ & ~new_new_n2162__;
  assign new_new_n2164__ = pi036 & ~new_new_n1156__;
  assign new_new_n2165__ = pi164 & new_new_n1156__;
  assign new_new_n2166__ = ~new_new_n2164__ & ~new_new_n2165__;
  assign new_new_n2167__ = new_new_n2163__ & new_new_n2166__;
  assign new_new_n2168__ = ~new_new_n2163__ & ~new_new_n2166__;
  assign new_new_n2169__ = pi292 & ~new_new_n1674__;
  assign new_new_n2170__ = pi420 & new_new_n1674__;
  assign new_new_n2171__ = ~new_new_n2169__ & ~new_new_n2170__;
  assign new_new_n2172__ = ~new_new_n2168__ & ~new_new_n2171__;
  assign new_new_n2173__ = ~new_new_n2167__ & ~new_new_n2172__;
  assign new_new_n2174__ = pi037 & ~new_new_n1156__;
  assign new_new_n2175__ = pi165 & new_new_n1156__;
  assign new_new_n2176__ = ~new_new_n2174__ & ~new_new_n2175__;
  assign new_new_n2177__ = ~new_new_n2173__ & new_new_n2176__;
  assign new_new_n2178__ = new_new_n2173__ & ~new_new_n2176__;
  assign new_new_n2179__ = pi293 & ~new_new_n1674__;
  assign new_new_n2180__ = pi421 & new_new_n1674__;
  assign new_new_n2181__ = ~new_new_n2179__ & ~new_new_n2180__;
  assign new_new_n2182__ = ~new_new_n2178__ & ~new_new_n2181__;
  assign new_new_n2183__ = ~new_new_n2177__ & ~new_new_n2182__;
  assign new_new_n2184__ = pi294 & ~new_new_n1674__;
  assign new_new_n2185__ = pi422 & new_new_n1674__;
  assign new_new_n2186__ = ~new_new_n2184__ & ~new_new_n2185__;
  assign new_new_n2187__ = new_new_n2183__ & new_new_n2186__;
  assign new_new_n2188__ = ~new_new_n2183__ & ~new_new_n2186__;
  assign new_new_n2189__ = pi038 & ~new_new_n1156__;
  assign new_new_n2190__ = pi166 & new_new_n1156__;
  assign new_new_n2191__ = ~new_new_n2189__ & ~new_new_n2190__;
  assign new_new_n2192__ = ~new_new_n2188__ & ~new_new_n2191__;
  assign new_new_n2193__ = ~new_new_n2187__ & ~new_new_n2192__;
  assign new_new_n2194__ = pi295 & ~new_new_n1674__;
  assign new_new_n2195__ = pi423 & new_new_n1674__;
  assign new_new_n2196__ = ~new_new_n2194__ & ~new_new_n2195__;
  assign new_new_n2197__ = ~new_new_n2193__ & new_new_n2196__;
  assign new_new_n2198__ = new_new_n2193__ & ~new_new_n2196__;
  assign new_new_n2199__ = pi039 & ~new_new_n1156__;
  assign new_new_n2200__ = pi167 & new_new_n1156__;
  assign new_new_n2201__ = ~new_new_n2199__ & ~new_new_n2200__;
  assign new_new_n2202__ = ~new_new_n2198__ & ~new_new_n2201__;
  assign new_new_n2203__ = ~new_new_n2197__ & ~new_new_n2202__;
  assign new_new_n2204__ = pi040 & ~new_new_n1156__;
  assign new_new_n2205__ = pi168 & new_new_n1156__;
  assign new_new_n2206__ = ~new_new_n2204__ & ~new_new_n2205__;
  assign new_new_n2207__ = new_new_n2203__ & new_new_n2206__;
  assign new_new_n2208__ = ~new_new_n2203__ & ~new_new_n2206__;
  assign new_new_n2209__ = pi296 & ~new_new_n1674__;
  assign new_new_n2210__ = pi424 & new_new_n1674__;
  assign new_new_n2211__ = ~new_new_n2209__ & ~new_new_n2210__;
  assign new_new_n2212__ = ~new_new_n2208__ & ~new_new_n2211__;
  assign new_new_n2213__ = ~new_new_n2207__ & ~new_new_n2212__;
  assign new_new_n2214__ = pi297 & ~new_new_n1674__;
  assign new_new_n2215__ = pi425 & new_new_n1674__;
  assign new_new_n2216__ = ~new_new_n2214__ & ~new_new_n2215__;
  assign new_new_n2217__ = new_new_n2213__ & new_new_n2216__;
  assign new_new_n2218__ = ~new_new_n2213__ & ~new_new_n2216__;
  assign new_new_n2219__ = pi041 & ~new_new_n1156__;
  assign new_new_n2220__ = pi169 & new_new_n1156__;
  assign new_new_n2221__ = ~new_new_n2219__ & ~new_new_n2220__;
  assign new_new_n2222__ = ~new_new_n2218__ & ~new_new_n2221__;
  assign new_new_n2223__ = ~new_new_n2217__ & ~new_new_n2222__;
  assign new_new_n2224__ = pi298 & ~new_new_n1674__;
  assign new_new_n2225__ = pi426 & new_new_n1674__;
  assign new_new_n2226__ = ~new_new_n2224__ & ~new_new_n2225__;
  assign new_new_n2227__ = ~new_new_n2223__ & new_new_n2226__;
  assign new_new_n2228__ = new_new_n2223__ & ~new_new_n2226__;
  assign new_new_n2229__ = pi042 & ~new_new_n1156__;
  assign new_new_n2230__ = pi170 & new_new_n1156__;
  assign new_new_n2231__ = ~new_new_n2229__ & ~new_new_n2230__;
  assign new_new_n2232__ = ~new_new_n2228__ & ~new_new_n2231__;
  assign new_new_n2233__ = ~new_new_n2227__ & ~new_new_n2232__;
  assign new_new_n2234__ = pi299 & ~new_new_n1674__;
  assign new_new_n2235__ = pi427 & new_new_n1674__;
  assign new_new_n2236__ = ~new_new_n2234__ & ~new_new_n2235__;
  assign new_new_n2237__ = ~new_new_n2233__ & new_new_n2236__;
  assign new_new_n2238__ = new_new_n1809__ & ~new_new_n2237__;
  assign new_new_n2239__ = new_new_n2233__ & ~new_new_n2236__;
  assign new_new_n2240__ = ~new_new_n2238__ & ~new_new_n2239__;
  assign new_new_n2241__ = pi300 & ~new_new_n1674__;
  assign new_new_n2242__ = pi428 & new_new_n1674__;
  assign new_new_n2243__ = ~new_new_n2241__ & ~new_new_n2242__;
  assign new_new_n2244__ = new_new_n2240__ & new_new_n2243__;
  assign new_new_n2245__ = ~new_new_n2240__ & ~new_new_n2243__;
  assign new_new_n2246__ = pi044 & ~new_new_n1156__;
  assign new_new_n2247__ = pi172 & new_new_n1156__;
  assign new_new_n2248__ = ~new_new_n2246__ & ~new_new_n2247__;
  assign new_new_n2249__ = ~new_new_n2245__ & ~new_new_n2248__;
  assign new_new_n2250__ = ~new_new_n2244__ & ~new_new_n2249__;
  assign new_new_n2251__ = pi301 & ~new_new_n1674__;
  assign new_new_n2252__ = pi429 & new_new_n1674__;
  assign new_new_n2253__ = ~new_new_n2251__ & ~new_new_n2252__;
  assign new_new_n2254__ = ~new_new_n2250__ & new_new_n2253__;
  assign new_new_n2255__ = new_new_n1806__ & ~new_new_n2254__;
  assign new_new_n2256__ = new_new_n2250__ & ~new_new_n2253__;
  assign new_new_n2257__ = ~new_new_n2255__ & ~new_new_n2256__;
  assign new_new_n2258__ = pi046 & ~new_new_n1156__;
  assign new_new_n2259__ = pi174 & new_new_n1156__;
  assign new_new_n2260__ = ~new_new_n2258__ & ~new_new_n2259__;
  assign new_new_n2261__ = ~new_new_n2257__ & new_new_n2260__;
  assign new_new_n2262__ = new_new_n2257__ & ~new_new_n2260__;
  assign new_new_n2263__ = pi302 & ~new_new_n1674__;
  assign new_new_n2264__ = pi430 & new_new_n1674__;
  assign new_new_n2265__ = ~new_new_n2263__ & ~new_new_n2264__;
  assign new_new_n2266__ = ~new_new_n2262__ & ~new_new_n2265__;
  assign new_new_n2267__ = ~new_new_n2261__ & ~new_new_n2266__;
  assign new_new_n2268__ = pi047 & ~new_new_n1156__;
  assign new_new_n2269__ = pi175 & new_new_n1156__;
  assign new_new_n2270__ = ~new_new_n2268__ & ~new_new_n2269__;
  assign new_new_n2271__ = ~new_new_n2267__ & new_new_n2270__;
  assign new_new_n2272__ = new_new_n1803__ & ~new_new_n2271__;
  assign new_new_n2273__ = new_new_n2267__ & ~new_new_n2270__;
  assign new_new_n2274__ = ~new_new_n2272__ & ~new_new_n2273__;
  assign new_new_n2275__ = pi048 & ~new_new_n1156__;
  assign new_new_n2276__ = pi176 & new_new_n1156__;
  assign new_new_n2277__ = ~new_new_n2275__ & ~new_new_n2276__;
  assign new_new_n2278__ = new_new_n2274__ & new_new_n2277__;
  assign new_new_n2279__ = new_new_n1800__ & ~new_new_n2278__;
  assign new_new_n2280__ = ~new_new_n2274__ & ~new_new_n2277__;
  assign new_new_n2281__ = ~new_new_n2279__ & ~new_new_n2280__;
  assign new_new_n2282__ = pi049 & ~new_new_n1156__;
  assign new_new_n2283__ = pi177 & new_new_n1156__;
  assign new_new_n2284__ = ~new_new_n2282__ & ~new_new_n2283__;
  assign new_new_n2285__ = new_new_n2281__ & new_new_n2284__;
  assign new_new_n2286__ = ~new_new_n2281__ & ~new_new_n2284__;
  assign new_new_n2287__ = pi305 & ~new_new_n1674__;
  assign new_new_n2288__ = pi433 & new_new_n1674__;
  assign new_new_n2289__ = ~new_new_n2287__ & ~new_new_n2288__;
  assign new_new_n2290__ = ~new_new_n2286__ & ~new_new_n2289__;
  assign new_new_n2291__ = ~new_new_n2285__ & ~new_new_n2290__;
  assign new_new_n2292__ = pi306 & ~new_new_n1674__;
  assign new_new_n2293__ = pi434 & new_new_n1674__;
  assign new_new_n2294__ = ~new_new_n2292__ & ~new_new_n2293__;
  assign new_new_n2295__ = new_new_n2291__ & new_new_n2294__;
  assign new_new_n2296__ = ~new_new_n2291__ & ~new_new_n2294__;
  assign new_new_n2297__ = pi050 & ~new_new_n1156__;
  assign new_new_n2298__ = pi178 & new_new_n1156__;
  assign new_new_n2299__ = ~new_new_n2297__ & ~new_new_n2298__;
  assign new_new_n2300__ = ~new_new_n2296__ & ~new_new_n2299__;
  assign new_new_n2301__ = ~new_new_n2295__ & ~new_new_n2300__;
  assign new_new_n2302__ = pi307 & ~new_new_n1674__;
  assign new_new_n2303__ = pi435 & new_new_n1674__;
  assign new_new_n2304__ = ~new_new_n2302__ & ~new_new_n2303__;
  assign new_new_n2305__ = ~new_new_n2301__ & new_new_n2304__;
  assign new_new_n2306__ = new_new_n1797__ & ~new_new_n2305__;
  assign new_new_n2307__ = new_new_n2301__ & ~new_new_n2304__;
  assign new_new_n2308__ = ~new_new_n2306__ & ~new_new_n2307__;
  assign new_new_n2309__ = pi308 & ~new_new_n1674__;
  assign new_new_n2310__ = pi436 & new_new_n1674__;
  assign new_new_n2311__ = ~new_new_n2309__ & ~new_new_n2310__;
  assign new_new_n2312__ = new_new_n2308__ & new_new_n2311__;
  assign new_new_n2313__ = new_new_n1794__ & ~new_new_n2312__;
  assign new_new_n2314__ = ~new_new_n2308__ & ~new_new_n2311__;
  assign new_new_n2315__ = ~new_new_n2313__ & ~new_new_n2314__;
  assign new_new_n2316__ = pi309 & ~new_new_n1674__;
  assign new_new_n2317__ = pi437 & new_new_n1674__;
  assign new_new_n2318__ = ~new_new_n2316__ & ~new_new_n2317__;
  assign new_new_n2319__ = new_new_n2315__ & new_new_n2318__;
  assign new_new_n2320__ = new_new_n1791__ & ~new_new_n2319__;
  assign new_new_n2321__ = ~new_new_n2315__ & ~new_new_n2318__;
  assign new_new_n2322__ = ~new_new_n2320__ & ~new_new_n2321__;
  assign new_new_n2323__ = pi054 & ~new_new_n1156__;
  assign new_new_n2324__ = pi182 & new_new_n1156__;
  assign new_new_n2325__ = ~new_new_n2323__ & ~new_new_n2324__;
  assign new_new_n2326__ = ~new_new_n2322__ & new_new_n2325__;
  assign new_new_n2327__ = new_new_n2322__ & ~new_new_n2325__;
  assign new_new_n2328__ = pi310 & ~new_new_n1674__;
  assign new_new_n2329__ = pi438 & new_new_n1674__;
  assign new_new_n2330__ = ~new_new_n2328__ & ~new_new_n2329__;
  assign new_new_n2331__ = ~new_new_n2327__ & ~new_new_n2330__;
  assign new_new_n2332__ = ~new_new_n2326__ & ~new_new_n2331__;
  assign new_new_n2333__ = pi311 & ~new_new_n1674__;
  assign new_new_n2334__ = pi439 & new_new_n1674__;
  assign new_new_n2335__ = ~new_new_n2333__ & ~new_new_n2334__;
  assign new_new_n2336__ = new_new_n2332__ & new_new_n2335__;
  assign new_new_n2337__ = ~new_new_n2332__ & ~new_new_n2335__;
  assign new_new_n2338__ = pi055 & ~new_new_n1156__;
  assign new_new_n2339__ = pi183 & new_new_n1156__;
  assign new_new_n2340__ = ~new_new_n2338__ & ~new_new_n2339__;
  assign new_new_n2341__ = ~new_new_n2337__ & ~new_new_n2340__;
  assign new_new_n2342__ = ~new_new_n2336__ & ~new_new_n2341__;
  assign new_new_n2343__ = pi056 & ~new_new_n1156__;
  assign new_new_n2344__ = pi184 & new_new_n1156__;
  assign new_new_n2345__ = ~new_new_n2343__ & ~new_new_n2344__;
  assign new_new_n2346__ = new_new_n2342__ & new_new_n2345__;
  assign new_new_n2347__ = ~new_new_n2342__ & ~new_new_n2345__;
  assign new_new_n2348__ = pi312 & ~new_new_n1674__;
  assign new_new_n2349__ = pi440 & new_new_n1674__;
  assign new_new_n2350__ = ~new_new_n2348__ & ~new_new_n2349__;
  assign new_new_n2351__ = ~new_new_n2347__ & ~new_new_n2350__;
  assign new_new_n2352__ = ~new_new_n2346__ & ~new_new_n2351__;
  assign new_new_n2353__ = pi313 & ~new_new_n1674__;
  assign new_new_n2354__ = pi441 & new_new_n1674__;
  assign new_new_n2355__ = ~new_new_n2353__ & ~new_new_n2354__;
  assign new_new_n2356__ = new_new_n2352__ & new_new_n2355__;
  assign new_new_n2357__ = ~new_new_n2352__ & ~new_new_n2355__;
  assign new_new_n2358__ = pi057 & ~new_new_n1156__;
  assign new_new_n2359__ = pi185 & new_new_n1156__;
  assign new_new_n2360__ = ~new_new_n2358__ & ~new_new_n2359__;
  assign new_new_n2361__ = ~new_new_n2357__ & ~new_new_n2360__;
  assign new_new_n2362__ = ~new_new_n2356__ & ~new_new_n2361__;
  assign new_new_n2363__ = pi314 & ~new_new_n1674__;
  assign new_new_n2364__ = pi442 & new_new_n1674__;
  assign new_new_n2365__ = ~new_new_n2363__ & ~new_new_n2364__;
  assign new_new_n2366__ = ~new_new_n2362__ & new_new_n2365__;
  assign new_new_n2367__ = new_new_n1788__ & ~new_new_n2366__;
  assign new_new_n2368__ = new_new_n2362__ & ~new_new_n2365__;
  assign new_new_n2369__ = ~new_new_n2367__ & ~new_new_n2368__;
  assign new_new_n2370__ = pi315 & ~new_new_n1674__;
  assign new_new_n2371__ = pi443 & new_new_n1674__;
  assign new_new_n2372__ = ~new_new_n2370__ & ~new_new_n2371__;
  assign new_new_n2373__ = new_new_n2369__ & new_new_n2372__;
  assign new_new_n2374__ = ~new_new_n2369__ & ~new_new_n2372__;
  assign new_new_n2375__ = pi059 & ~new_new_n1156__;
  assign new_new_n2376__ = pi187 & new_new_n1156__;
  assign new_new_n2377__ = ~new_new_n2375__ & ~new_new_n2376__;
  assign new_new_n2378__ = ~new_new_n2374__ & ~new_new_n2377__;
  assign new_new_n2379__ = ~new_new_n2373__ & ~new_new_n2378__;
  assign new_new_n2380__ = pi316 & ~new_new_n1674__;
  assign new_new_n2381__ = pi444 & new_new_n1674__;
  assign new_new_n2382__ = ~new_new_n2380__ & ~new_new_n2381__;
  assign new_new_n2383__ = ~new_new_n2379__ & new_new_n2382__;
  assign new_new_n2384__ = new_new_n2379__ & ~new_new_n2382__;
  assign new_new_n2385__ = pi060 & ~new_new_n1156__;
  assign new_new_n2386__ = pi188 & new_new_n1156__;
  assign new_new_n2387__ = ~new_new_n2385__ & ~new_new_n2386__;
  assign new_new_n2388__ = ~new_new_n2384__ & ~new_new_n2387__;
  assign new_new_n2389__ = ~new_new_n2383__ & ~new_new_n2388__;
  assign new_new_n2390__ = pi317 & ~new_new_n1674__;
  assign new_new_n2391__ = pi445 & new_new_n1674__;
  assign new_new_n2392__ = ~new_new_n2390__ & ~new_new_n2391__;
  assign new_new_n2393__ = ~new_new_n2389__ & new_new_n2392__;
  assign new_new_n2394__ = new_new_n1785__ & ~new_new_n2393__;
  assign new_new_n2395__ = new_new_n2389__ & ~new_new_n2392__;
  assign new_new_n2396__ = ~new_new_n2394__ & ~new_new_n2395__;
  assign new_new_n2397__ = pi318 & ~new_new_n1674__;
  assign new_new_n2398__ = pi446 & new_new_n1674__;
  assign new_new_n2399__ = ~new_new_n2397__ & ~new_new_n2398__;
  assign new_new_n2400__ = new_new_n2396__ & new_new_n2399__;
  assign new_new_n2401__ = ~new_new_n2396__ & ~new_new_n2399__;
  assign new_new_n2402__ = pi062 & ~new_new_n1156__;
  assign new_new_n2403__ = pi190 & new_new_n1156__;
  assign new_new_n2404__ = ~new_new_n2402__ & ~new_new_n2403__;
  assign new_new_n2405__ = ~new_new_n2401__ & ~new_new_n2404__;
  assign new_new_n2406__ = ~new_new_n2400__ & ~new_new_n2405__;
  assign new_new_n2407__ = pi319 & ~new_new_n1674__;
  assign new_new_n2408__ = pi447 & new_new_n1674__;
  assign new_new_n2409__ = ~new_new_n2407__ & ~new_new_n2408__;
  assign new_new_n2410__ = ~new_new_n2406__ & new_new_n2409__;
  assign new_new_n2411__ = new_new_n2406__ & ~new_new_n2409__;
  assign new_new_n2412__ = pi063 & ~new_new_n1156__;
  assign new_new_n2413__ = pi191 & new_new_n1156__;
  assign new_new_n2414__ = ~new_new_n2412__ & ~new_new_n2413__;
  assign new_new_n2415__ = ~new_new_n2411__ & ~new_new_n2414__;
  assign new_new_n2416__ = ~new_new_n2410__ & ~new_new_n2415__;
  assign new_new_n2417__ = pi320 & ~new_new_n1674__;
  assign new_new_n2418__ = pi448 & new_new_n1674__;
  assign new_new_n2419__ = ~new_new_n2417__ & ~new_new_n2418__;
  assign new_new_n2420__ = ~new_new_n2416__ & new_new_n2419__;
  assign new_new_n2421__ = new_new_n2416__ & ~new_new_n2419__;
  assign new_new_n2422__ = pi064 & ~new_new_n1156__;
  assign new_new_n2423__ = pi192 & new_new_n1156__;
  assign new_new_n2424__ = ~new_new_n2422__ & ~new_new_n2423__;
  assign new_new_n2425__ = ~new_new_n2421__ & ~new_new_n2424__;
  assign new_new_n2426__ = ~new_new_n2420__ & ~new_new_n2425__;
  assign new_new_n2427__ = pi065 & ~new_new_n1156__;
  assign new_new_n2428__ = pi193 & new_new_n1156__;
  assign new_new_n2429__ = ~new_new_n2427__ & ~new_new_n2428__;
  assign new_new_n2430__ = new_new_n2426__ & new_new_n2429__;
  assign new_new_n2431__ = ~new_new_n2426__ & ~new_new_n2429__;
  assign new_new_n2432__ = pi321 & ~new_new_n1674__;
  assign new_new_n2433__ = pi449 & new_new_n1674__;
  assign new_new_n2434__ = ~new_new_n2432__ & ~new_new_n2433__;
  assign new_new_n2435__ = ~new_new_n2431__ & ~new_new_n2434__;
  assign new_new_n2436__ = ~new_new_n2430__ & ~new_new_n2435__;
  assign new_new_n2437__ = pi066 & ~new_new_n1156__;
  assign new_new_n2438__ = pi194 & new_new_n1156__;
  assign new_new_n2439__ = ~new_new_n2437__ & ~new_new_n2438__;
  assign new_new_n2440__ = ~new_new_n2436__ & new_new_n2439__;
  assign new_new_n2441__ = new_new_n1782__ & ~new_new_n2440__;
  assign new_new_n2442__ = new_new_n2436__ & ~new_new_n2439__;
  assign new_new_n2443__ = ~new_new_n2441__ & ~new_new_n2442__;
  assign new_new_n2444__ = pi067 & ~new_new_n1156__;
  assign new_new_n2445__ = pi195 & new_new_n1156__;
  assign new_new_n2446__ = ~new_new_n2444__ & ~new_new_n2445__;
  assign new_new_n2447__ = new_new_n2443__ & new_new_n2446__;
  assign new_new_n2448__ = new_new_n1779__ & ~new_new_n2447__;
  assign new_new_n2449__ = ~new_new_n2443__ & ~new_new_n2446__;
  assign new_new_n2450__ = ~new_new_n2448__ & ~new_new_n2449__;
  assign new_new_n2451__ = pi068 & ~new_new_n1156__;
  assign new_new_n2452__ = pi196 & new_new_n1156__;
  assign new_new_n2453__ = ~new_new_n2451__ & ~new_new_n2452__;
  assign new_new_n2454__ = new_new_n2450__ & new_new_n2453__;
  assign new_new_n2455__ = ~new_new_n2450__ & ~new_new_n2453__;
  assign new_new_n2456__ = pi324 & ~new_new_n1674__;
  assign new_new_n2457__ = pi452 & new_new_n1674__;
  assign new_new_n2458__ = ~new_new_n2456__ & ~new_new_n2457__;
  assign new_new_n2459__ = ~new_new_n2455__ & ~new_new_n2458__;
  assign new_new_n2460__ = ~new_new_n2454__ & ~new_new_n2459__;
  assign new_new_n2461__ = pi069 & ~new_new_n1156__;
  assign new_new_n2462__ = pi197 & new_new_n1156__;
  assign new_new_n2463__ = ~new_new_n2461__ & ~new_new_n2462__;
  assign new_new_n2464__ = ~new_new_n2460__ & new_new_n2463__;
  assign new_new_n2465__ = new_new_n2460__ & ~new_new_n2463__;
  assign new_new_n2466__ = pi325 & ~new_new_n1674__;
  assign new_new_n2467__ = pi453 & new_new_n1674__;
  assign new_new_n2468__ = ~new_new_n2466__ & ~new_new_n2467__;
  assign new_new_n2469__ = ~new_new_n2465__ & ~new_new_n2468__;
  assign new_new_n2470__ = ~new_new_n2464__ & ~new_new_n2469__;
  assign new_new_n2471__ = pi070 & ~new_new_n1156__;
  assign new_new_n2472__ = pi198 & new_new_n1156__;
  assign new_new_n2473__ = ~new_new_n2471__ & ~new_new_n2472__;
  assign new_new_n2474__ = ~new_new_n2470__ & new_new_n2473__;
  assign new_new_n2475__ = new_new_n1776__ & ~new_new_n2474__;
  assign new_new_n2476__ = new_new_n2470__ & ~new_new_n2473__;
  assign new_new_n2477__ = ~new_new_n2475__ & ~new_new_n2476__;
  assign new_new_n2478__ = pi071 & ~new_new_n1156__;
  assign new_new_n2479__ = pi199 & new_new_n1156__;
  assign new_new_n2480__ = ~new_new_n2478__ & ~new_new_n2479__;
  assign new_new_n2481__ = new_new_n2477__ & new_new_n2480__;
  assign new_new_n2482__ = ~new_new_n2477__ & ~new_new_n2480__;
  assign new_new_n2483__ = pi327 & ~new_new_n1674__;
  assign new_new_n2484__ = pi455 & new_new_n1674__;
  assign new_new_n2485__ = ~new_new_n2483__ & ~new_new_n2484__;
  assign new_new_n2486__ = ~new_new_n2482__ & ~new_new_n2485__;
  assign new_new_n2487__ = ~new_new_n2481__ & ~new_new_n2486__;
  assign new_new_n2488__ = pi072 & ~new_new_n1156__;
  assign new_new_n2489__ = pi200 & new_new_n1156__;
  assign new_new_n2490__ = ~new_new_n2488__ & ~new_new_n2489__;
  assign new_new_n2491__ = ~new_new_n2487__ & new_new_n2490__;
  assign new_new_n2492__ = new_new_n1773__ & ~new_new_n2491__;
  assign new_new_n2493__ = new_new_n2487__ & ~new_new_n2490__;
  assign new_new_n2494__ = ~new_new_n2492__ & ~new_new_n2493__;
  assign new_new_n2495__ = pi073 & ~new_new_n1156__;
  assign new_new_n2496__ = pi201 & new_new_n1156__;
  assign new_new_n2497__ = ~new_new_n2495__ & ~new_new_n2496__;
  assign new_new_n2498__ = new_new_n2494__ & new_new_n2497__;
  assign new_new_n2499__ = ~new_new_n2494__ & ~new_new_n2497__;
  assign new_new_n2500__ = pi329 & ~new_new_n1674__;
  assign new_new_n2501__ = pi457 & new_new_n1674__;
  assign new_new_n2502__ = ~new_new_n2500__ & ~new_new_n2501__;
  assign new_new_n2503__ = ~new_new_n2499__ & ~new_new_n2502__;
  assign new_new_n2504__ = ~new_new_n2498__ & ~new_new_n2503__;
  assign new_new_n2505__ = pi330 & ~new_new_n1674__;
  assign new_new_n2506__ = pi458 & new_new_n1674__;
  assign new_new_n2507__ = ~new_new_n2505__ & ~new_new_n2506__;
  assign new_new_n2508__ = new_new_n2504__ & new_new_n2507__;
  assign new_new_n2509__ = ~new_new_n2504__ & ~new_new_n2507__;
  assign new_new_n2510__ = pi074 & ~new_new_n1156__;
  assign new_new_n2511__ = pi202 & new_new_n1156__;
  assign new_new_n2512__ = ~new_new_n2510__ & ~new_new_n2511__;
  assign new_new_n2513__ = ~new_new_n2509__ & ~new_new_n2512__;
  assign new_new_n2514__ = ~new_new_n2508__ & ~new_new_n2513__;
  assign new_new_n2515__ = pi331 & ~new_new_n1674__;
  assign new_new_n2516__ = pi459 & new_new_n1674__;
  assign new_new_n2517__ = ~new_new_n2515__ & ~new_new_n2516__;
  assign new_new_n2518__ = ~new_new_n2514__ & new_new_n2517__;
  assign new_new_n2519__ = new_new_n1770__ & ~new_new_n2518__;
  assign new_new_n2520__ = new_new_n2514__ & ~new_new_n2517__;
  assign new_new_n2521__ = ~new_new_n2519__ & ~new_new_n2520__;
  assign new_new_n2522__ = pi332 & ~new_new_n1674__;
  assign new_new_n2523__ = pi460 & new_new_n1674__;
  assign new_new_n2524__ = ~new_new_n2522__ & ~new_new_n2523__;
  assign new_new_n2525__ = new_new_n2521__ & new_new_n2524__;
  assign new_new_n2526__ = new_new_n1767__ & ~new_new_n2525__;
  assign new_new_n2527__ = ~new_new_n2521__ & ~new_new_n2524__;
  assign new_new_n2528__ = ~new_new_n2526__ & ~new_new_n2527__;
  assign new_new_n2529__ = pi333 & ~new_new_n1674__;
  assign new_new_n2530__ = pi461 & new_new_n1674__;
  assign new_new_n2531__ = ~new_new_n2529__ & ~new_new_n2530__;
  assign new_new_n2532__ = new_new_n2528__ & new_new_n2531__;
  assign new_new_n2533__ = new_new_n1764__ & ~new_new_n2532__;
  assign new_new_n2534__ = ~new_new_n2528__ & ~new_new_n2531__;
  assign new_new_n2535__ = ~new_new_n2533__ & ~new_new_n2534__;
  assign new_new_n2536__ = pi334 & ~new_new_n1674__;
  assign new_new_n2537__ = pi462 & new_new_n1674__;
  assign new_new_n2538__ = ~new_new_n2536__ & ~new_new_n2537__;
  assign new_new_n2539__ = new_new_n2535__ & new_new_n2538__;
  assign new_new_n2540__ = new_new_n1761__ & ~new_new_n2539__;
  assign new_new_n2541__ = ~new_new_n2535__ & ~new_new_n2538__;
  assign new_new_n2542__ = ~new_new_n2540__ & ~new_new_n2541__;
  assign new_new_n2543__ = pi335 & ~new_new_n1674__;
  assign new_new_n2544__ = pi463 & new_new_n1674__;
  assign new_new_n2545__ = ~new_new_n2543__ & ~new_new_n2544__;
  assign new_new_n2546__ = new_new_n2542__ & new_new_n2545__;
  assign new_new_n2547__ = new_new_n1758__ & ~new_new_n2546__;
  assign new_new_n2548__ = ~new_new_n2542__ & ~new_new_n2545__;
  assign new_new_n2549__ = ~new_new_n2547__ & ~new_new_n2548__;
  assign new_new_n2550__ = pi336 & ~new_new_n1674__;
  assign new_new_n2551__ = pi464 & new_new_n1674__;
  assign new_new_n2552__ = ~new_new_n2550__ & ~new_new_n2551__;
  assign new_new_n2553__ = new_new_n2549__ & new_new_n2552__;
  assign new_new_n2554__ = new_new_n1755__ & ~new_new_n2553__;
  assign new_new_n2555__ = ~new_new_n2549__ & ~new_new_n2552__;
  assign new_new_n2556__ = ~new_new_n2554__ & ~new_new_n2555__;
  assign new_new_n2557__ = pi337 & ~new_new_n1674__;
  assign new_new_n2558__ = pi465 & new_new_n1674__;
  assign new_new_n2559__ = ~new_new_n2557__ & ~new_new_n2558__;
  assign new_new_n2560__ = new_new_n2556__ & new_new_n2559__;
  assign new_new_n2561__ = new_new_n1752__ & ~new_new_n2560__;
  assign new_new_n2562__ = ~new_new_n2556__ & ~new_new_n2559__;
  assign new_new_n2563__ = ~new_new_n2561__ & ~new_new_n2562__;
  assign new_new_n2564__ = pi338 & ~new_new_n1674__;
  assign new_new_n2565__ = pi466 & new_new_n1674__;
  assign new_new_n2566__ = ~new_new_n2564__ & ~new_new_n2565__;
  assign new_new_n2567__ = new_new_n2563__ & new_new_n2566__;
  assign new_new_n2568__ = ~new_new_n2563__ & ~new_new_n2566__;
  assign new_new_n2569__ = pi082 & ~new_new_n1156__;
  assign new_new_n2570__ = pi210 & new_new_n1156__;
  assign new_new_n2571__ = ~new_new_n2569__ & ~new_new_n2570__;
  assign new_new_n2572__ = ~new_new_n2568__ & ~new_new_n2571__;
  assign new_new_n2573__ = ~new_new_n2567__ & ~new_new_n2572__;
  assign new_new_n2574__ = pi083 & ~new_new_n1156__;
  assign new_new_n2575__ = pi211 & new_new_n1156__;
  assign new_new_n2576__ = ~new_new_n2574__ & ~new_new_n2575__;
  assign new_new_n2577__ = new_new_n2573__ & new_new_n2576__;
  assign new_new_n2578__ = ~new_new_n2573__ & ~new_new_n2576__;
  assign new_new_n2579__ = pi339 & ~new_new_n1674__;
  assign new_new_n2580__ = pi467 & new_new_n1674__;
  assign new_new_n2581__ = ~new_new_n2579__ & ~new_new_n2580__;
  assign new_new_n2582__ = ~new_new_n2578__ & ~new_new_n2581__;
  assign new_new_n2583__ = ~new_new_n2577__ & ~new_new_n2582__;
  assign new_new_n2584__ = pi084 & ~new_new_n1156__;
  assign new_new_n2585__ = pi212 & new_new_n1156__;
  assign new_new_n2586__ = ~new_new_n2584__ & ~new_new_n2585__;
  assign new_new_n2587__ = ~new_new_n2583__ & new_new_n2586__;
  assign new_new_n2588__ = new_new_n1749__ & ~new_new_n2587__;
  assign new_new_n2589__ = new_new_n2583__ & ~new_new_n2586__;
  assign new_new_n2590__ = ~new_new_n2588__ & ~new_new_n2589__;
  assign new_new_n2591__ = pi341 & ~new_new_n1674__;
  assign new_new_n2592__ = pi469 & new_new_n1674__;
  assign new_new_n2593__ = ~new_new_n2591__ & ~new_new_n2592__;
  assign new_new_n2594__ = ~new_new_n2590__ & new_new_n2593__;
  assign new_new_n2595__ = new_new_n2590__ & ~new_new_n2593__;
  assign new_new_n2596__ = pi085 & ~new_new_n1156__;
  assign new_new_n2597__ = pi213 & new_new_n1156__;
  assign new_new_n2598__ = ~new_new_n2596__ & ~new_new_n2597__;
  assign new_new_n2599__ = ~new_new_n2595__ & ~new_new_n2598__;
  assign new_new_n2600__ = ~new_new_n2594__ & ~new_new_n2599__;
  assign new_new_n2601__ = pi342 & ~new_new_n1674__;
  assign new_new_n2602__ = pi470 & new_new_n1674__;
  assign new_new_n2603__ = ~new_new_n2601__ & ~new_new_n2602__;
  assign new_new_n2604__ = ~new_new_n2600__ & new_new_n2603__;
  assign new_new_n2605__ = new_new_n1746__ & ~new_new_n2604__;
  assign new_new_n2606__ = new_new_n2600__ & ~new_new_n2603__;
  assign new_new_n2607__ = ~new_new_n2605__ & ~new_new_n2606__;
  assign new_new_n2608__ = pi343 & ~new_new_n1674__;
  assign new_new_n2609__ = pi471 & new_new_n1674__;
  assign new_new_n2610__ = ~new_new_n2608__ & ~new_new_n2609__;
  assign new_new_n2611__ = new_new_n2607__ & new_new_n2610__;
  assign new_new_n2612__ = new_new_n1743__ & ~new_new_n2611__;
  assign new_new_n2613__ = ~new_new_n2607__ & ~new_new_n2610__;
  assign new_new_n2614__ = ~new_new_n2612__ & ~new_new_n2613__;
  assign new_new_n2615__ = pi344 & ~new_new_n1674__;
  assign new_new_n2616__ = pi472 & new_new_n1674__;
  assign new_new_n2617__ = ~new_new_n2615__ & ~new_new_n2616__;
  assign new_new_n2618__ = new_new_n2614__ & new_new_n2617__;
  assign new_new_n2619__ = new_new_n1740__ & ~new_new_n2618__;
  assign new_new_n2620__ = ~new_new_n2614__ & ~new_new_n2617__;
  assign new_new_n2621__ = ~new_new_n2619__ & ~new_new_n2620__;
  assign new_new_n2622__ = pi345 & ~new_new_n1674__;
  assign new_new_n2623__ = pi473 & new_new_n1674__;
  assign new_new_n2624__ = ~new_new_n2622__ & ~new_new_n2623__;
  assign new_new_n2625__ = new_new_n2621__ & new_new_n2624__;
  assign new_new_n2626__ = new_new_n1737__ & ~new_new_n2625__;
  assign new_new_n2627__ = ~new_new_n2621__ & ~new_new_n2624__;
  assign new_new_n2628__ = ~new_new_n2626__ & ~new_new_n2627__;
  assign new_new_n2629__ = pi090 & ~new_new_n1156__;
  assign new_new_n2630__ = pi218 & new_new_n1156__;
  assign new_new_n2631__ = ~new_new_n2629__ & ~new_new_n2630__;
  assign new_new_n2632__ = ~new_new_n2628__ & new_new_n2631__;
  assign new_new_n2633__ = new_new_n2628__ & ~new_new_n2631__;
  assign new_new_n2634__ = pi346 & ~new_new_n1674__;
  assign new_new_n2635__ = pi474 & new_new_n1674__;
  assign new_new_n2636__ = ~new_new_n2634__ & ~new_new_n2635__;
  assign new_new_n2637__ = ~new_new_n2633__ & ~new_new_n2636__;
  assign new_new_n2638__ = ~new_new_n2632__ & ~new_new_n2637__;
  assign new_new_n2639__ = pi091 & ~new_new_n1156__;
  assign new_new_n2640__ = pi219 & new_new_n1156__;
  assign new_new_n2641__ = ~new_new_n2639__ & ~new_new_n2640__;
  assign new_new_n2642__ = ~new_new_n2638__ & new_new_n2641__;
  assign new_new_n2643__ = new_new_n1734__ & ~new_new_n2642__;
  assign new_new_n2644__ = new_new_n2638__ & ~new_new_n2641__;
  assign new_new_n2645__ = ~new_new_n2643__ & ~new_new_n2644__;
  assign new_new_n2646__ = pi092 & ~new_new_n1156__;
  assign new_new_n2647__ = pi220 & new_new_n1156__;
  assign new_new_n2648__ = ~new_new_n2646__ & ~new_new_n2647__;
  assign new_new_n2649__ = new_new_n2645__ & new_new_n2648__;
  assign new_new_n2650__ = new_new_n1731__ & ~new_new_n2649__;
  assign new_new_n2651__ = ~new_new_n2645__ & ~new_new_n2648__;
  assign new_new_n2652__ = ~new_new_n2650__ & ~new_new_n2651__;
  assign new_new_n2653__ = pi093 & ~new_new_n1156__;
  assign new_new_n2654__ = pi221 & new_new_n1156__;
  assign new_new_n2655__ = ~new_new_n2653__ & ~new_new_n2654__;
  assign new_new_n2656__ = new_new_n2652__ & new_new_n2655__;
  assign new_new_n2657__ = new_new_n1728__ & ~new_new_n2656__;
  assign new_new_n2658__ = ~new_new_n2652__ & ~new_new_n2655__;
  assign new_new_n2659__ = ~new_new_n2657__ & ~new_new_n2658__;
  assign new_new_n2660__ = pi094 & ~new_new_n1156__;
  assign new_new_n2661__ = pi222 & new_new_n1156__;
  assign new_new_n2662__ = ~new_new_n2660__ & ~new_new_n2661__;
  assign new_new_n2663__ = new_new_n2659__ & new_new_n2662__;
  assign new_new_n2664__ = new_new_n1725__ & ~new_new_n2663__;
  assign new_new_n2665__ = ~new_new_n2659__ & ~new_new_n2662__;
  assign new_new_n2666__ = ~new_new_n2664__ & ~new_new_n2665__;
  assign new_new_n2667__ = pi095 & ~new_new_n1156__;
  assign new_new_n2668__ = pi223 & new_new_n1156__;
  assign new_new_n2669__ = ~new_new_n2667__ & ~new_new_n2668__;
  assign new_new_n2670__ = new_new_n2666__ & new_new_n2669__;
  assign new_new_n2671__ = new_new_n1722__ & ~new_new_n2670__;
  assign new_new_n2672__ = ~new_new_n2666__ & ~new_new_n2669__;
  assign new_new_n2673__ = ~new_new_n2671__ & ~new_new_n2672__;
  assign new_new_n2674__ = pi096 & ~new_new_n1156__;
  assign new_new_n2675__ = pi224 & new_new_n1156__;
  assign new_new_n2676__ = ~new_new_n2674__ & ~new_new_n2675__;
  assign new_new_n2677__ = new_new_n2673__ & new_new_n2676__;
  assign new_new_n2678__ = ~new_new_n2673__ & ~new_new_n2676__;
  assign new_new_n2679__ = pi352 & ~new_new_n1674__;
  assign new_new_n2680__ = pi480 & new_new_n1674__;
  assign new_new_n2681__ = ~new_new_n2679__ & ~new_new_n2680__;
  assign new_new_n2682__ = ~new_new_n2678__ & ~new_new_n2681__;
  assign new_new_n2683__ = ~new_new_n2677__ & ~new_new_n2682__;
  assign new_new_n2684__ = pi097 & ~new_new_n1156__;
  assign new_new_n2685__ = pi225 & new_new_n1156__;
  assign new_new_n2686__ = ~new_new_n2684__ & ~new_new_n2685__;
  assign new_new_n2687__ = ~new_new_n2683__ & new_new_n2686__;
  assign new_new_n2688__ = new_new_n2683__ & ~new_new_n2686__;
  assign new_new_n2689__ = pi353 & ~new_new_n1674__;
  assign new_new_n2690__ = pi481 & new_new_n1674__;
  assign new_new_n2691__ = ~new_new_n2689__ & ~new_new_n2690__;
  assign new_new_n2692__ = ~new_new_n2688__ & ~new_new_n2691__;
  assign new_new_n2693__ = ~new_new_n2687__ & ~new_new_n2692__;
  assign new_new_n2694__ = pi098 & ~new_new_n1156__;
  assign new_new_n2695__ = pi226 & new_new_n1156__;
  assign new_new_n2696__ = ~new_new_n2694__ & ~new_new_n2695__;
  assign new_new_n2697__ = ~new_new_n2693__ & new_new_n2696__;
  assign new_new_n2698__ = new_new_n1719__ & ~new_new_n2697__;
  assign new_new_n2699__ = new_new_n2693__ & ~new_new_n2696__;
  assign new_new_n2700__ = ~new_new_n2698__ & ~new_new_n2699__;
  assign new_new_n2701__ = pi099 & ~new_new_n1156__;
  assign new_new_n2702__ = pi227 & new_new_n1156__;
  assign new_new_n2703__ = ~new_new_n2701__ & ~new_new_n2702__;
  assign new_new_n2704__ = new_new_n2700__ & new_new_n2703__;
  assign new_new_n2705__ = ~new_new_n2700__ & ~new_new_n2703__;
  assign new_new_n2706__ = pi355 & ~new_new_n1674__;
  assign new_new_n2707__ = pi483 & new_new_n1674__;
  assign new_new_n2708__ = ~new_new_n2706__ & ~new_new_n2707__;
  assign new_new_n2709__ = ~new_new_n2705__ & ~new_new_n2708__;
  assign new_new_n2710__ = ~new_new_n2704__ & ~new_new_n2709__;
  assign new_new_n2711__ = pi100 & ~new_new_n1156__;
  assign new_new_n2712__ = pi228 & new_new_n1156__;
  assign new_new_n2713__ = ~new_new_n2711__ & ~new_new_n2712__;
  assign new_new_n2714__ = ~new_new_n2710__ & new_new_n2713__;
  assign new_new_n2715__ = new_new_n1716__ & ~new_new_n2714__;
  assign new_new_n2716__ = new_new_n2710__ & ~new_new_n2713__;
  assign new_new_n2717__ = ~new_new_n2715__ & ~new_new_n2716__;
  assign new_new_n2718__ = pi101 & ~new_new_n1156__;
  assign new_new_n2719__ = pi229 & new_new_n1156__;
  assign new_new_n2720__ = ~new_new_n2718__ & ~new_new_n2719__;
  assign new_new_n2721__ = new_new_n2717__ & new_new_n2720__;
  assign new_new_n2722__ = new_new_n1713__ & ~new_new_n2721__;
  assign new_new_n2723__ = ~new_new_n2717__ & ~new_new_n2720__;
  assign new_new_n2724__ = ~new_new_n2722__ & ~new_new_n2723__;
  assign new_new_n2725__ = pi102 & ~new_new_n1156__;
  assign new_new_n2726__ = pi230 & new_new_n1156__;
  assign new_new_n2727__ = ~new_new_n2725__ & ~new_new_n2726__;
  assign new_new_n2728__ = new_new_n2724__ & new_new_n2727__;
  assign new_new_n2729__ = new_new_n1710__ & ~new_new_n2728__;
  assign new_new_n2730__ = ~new_new_n2724__ & ~new_new_n2727__;
  assign new_new_n2731__ = ~new_new_n2729__ & ~new_new_n2730__;
  assign new_new_n2732__ = pi103 & ~new_new_n1156__;
  assign new_new_n2733__ = pi231 & new_new_n1156__;
  assign new_new_n2734__ = ~new_new_n2732__ & ~new_new_n2733__;
  assign new_new_n2735__ = new_new_n2731__ & new_new_n2734__;
  assign new_new_n2736__ = new_new_n1707__ & ~new_new_n2735__;
  assign new_new_n2737__ = ~new_new_n2731__ & ~new_new_n2734__;
  assign new_new_n2738__ = ~new_new_n2736__ & ~new_new_n2737__;
  assign new_new_n2739__ = pi104 & ~new_new_n1156__;
  assign new_new_n2740__ = pi232 & new_new_n1156__;
  assign new_new_n2741__ = ~new_new_n2739__ & ~new_new_n2740__;
  assign new_new_n2742__ = new_new_n2738__ & new_new_n2741__;
  assign new_new_n2743__ = ~new_new_n2738__ & ~new_new_n2741__;
  assign new_new_n2744__ = pi360 & ~new_new_n1674__;
  assign new_new_n2745__ = pi488 & new_new_n1674__;
  assign new_new_n2746__ = ~new_new_n2744__ & ~new_new_n2745__;
  assign new_new_n2747__ = ~new_new_n2743__ & ~new_new_n2746__;
  assign new_new_n2748__ = ~new_new_n2742__ & ~new_new_n2747__;
  assign new_new_n2749__ = pi105 & ~new_new_n1156__;
  assign new_new_n2750__ = pi233 & new_new_n1156__;
  assign new_new_n2751__ = ~new_new_n2749__ & ~new_new_n2750__;
  assign new_new_n2752__ = ~new_new_n2748__ & new_new_n2751__;
  assign new_new_n2753__ = new_new_n2748__ & ~new_new_n2751__;
  assign new_new_n2754__ = pi361 & ~new_new_n1674__;
  assign new_new_n2755__ = pi489 & new_new_n1674__;
  assign new_new_n2756__ = ~new_new_n2754__ & ~new_new_n2755__;
  assign new_new_n2757__ = ~new_new_n2753__ & ~new_new_n2756__;
  assign new_new_n2758__ = ~new_new_n2752__ & ~new_new_n2757__;
  assign new_new_n2759__ = pi106 & ~new_new_n1156__;
  assign new_new_n2760__ = pi234 & new_new_n1156__;
  assign new_new_n2761__ = ~new_new_n2759__ & ~new_new_n2760__;
  assign new_new_n2762__ = ~new_new_n2758__ & new_new_n2761__;
  assign new_new_n2763__ = new_new_n1704__ & ~new_new_n2762__;
  assign new_new_n2764__ = new_new_n2758__ & ~new_new_n2761__;
  assign new_new_n2765__ = ~new_new_n2763__ & ~new_new_n2764__;
  assign new_new_n2766__ = pi107 & ~new_new_n1156__;
  assign new_new_n2767__ = pi235 & new_new_n1156__;
  assign new_new_n2768__ = ~new_new_n2766__ & ~new_new_n2767__;
  assign new_new_n2769__ = new_new_n2765__ & new_new_n2768__;
  assign new_new_n2770__ = new_new_n1701__ & ~new_new_n2769__;
  assign new_new_n2771__ = ~new_new_n2765__ & ~new_new_n2768__;
  assign new_new_n2772__ = ~new_new_n2770__ & ~new_new_n2771__;
  assign new_new_n2773__ = pi108 & ~new_new_n1156__;
  assign new_new_n2774__ = pi236 & new_new_n1156__;
  assign new_new_n2775__ = ~new_new_n2773__ & ~new_new_n2774__;
  assign new_new_n2776__ = new_new_n2772__ & new_new_n2775__;
  assign new_new_n2777__ = ~new_new_n2772__ & ~new_new_n2775__;
  assign new_new_n2778__ = pi364 & ~new_new_n1674__;
  assign new_new_n2779__ = pi492 & new_new_n1674__;
  assign new_new_n2780__ = ~new_new_n2778__ & ~new_new_n2779__;
  assign new_new_n2781__ = ~new_new_n2777__ & ~new_new_n2780__;
  assign new_new_n2782__ = ~new_new_n2776__ & ~new_new_n2781__;
  assign new_new_n2783__ = pi109 & ~new_new_n1156__;
  assign new_new_n2784__ = pi237 & new_new_n1156__;
  assign new_new_n2785__ = ~new_new_n2783__ & ~new_new_n2784__;
  assign new_new_n2786__ = ~new_new_n2782__ & new_new_n2785__;
  assign new_new_n2787__ = new_new_n1698__ & ~new_new_n2786__;
  assign new_new_n2788__ = new_new_n2782__ & ~new_new_n2785__;
  assign new_new_n2789__ = ~new_new_n2787__ & ~new_new_n2788__;
  assign new_new_n2790__ = pi110 & ~new_new_n1156__;
  assign new_new_n2791__ = pi238 & new_new_n1156__;
  assign new_new_n2792__ = ~new_new_n2790__ & ~new_new_n2791__;
  assign new_new_n2793__ = new_new_n2789__ & new_new_n2792__;
  assign new_new_n2794__ = new_new_n1695__ & ~new_new_n2793__;
  assign new_new_n2795__ = ~new_new_n2789__ & ~new_new_n2792__;
  assign new_new_n2796__ = ~new_new_n2794__ & ~new_new_n2795__;
  assign new_new_n2797__ = pi111 & ~new_new_n1156__;
  assign new_new_n2798__ = pi239 & new_new_n1156__;
  assign new_new_n2799__ = ~new_new_n2797__ & ~new_new_n2798__;
  assign new_new_n2800__ = new_new_n2796__ & new_new_n2799__;
  assign new_new_n2801__ = ~new_new_n2796__ & ~new_new_n2799__;
  assign new_new_n2802__ = pi367 & ~new_new_n1674__;
  assign new_new_n2803__ = pi495 & new_new_n1674__;
  assign new_new_n2804__ = ~new_new_n2802__ & ~new_new_n2803__;
  assign new_new_n2805__ = ~new_new_n2801__ & ~new_new_n2804__;
  assign new_new_n2806__ = ~new_new_n2800__ & ~new_new_n2805__;
  assign new_new_n2807__ = pi112 & ~new_new_n1156__;
  assign new_new_n2808__ = pi240 & new_new_n1156__;
  assign new_new_n2809__ = ~new_new_n2807__ & ~new_new_n2808__;
  assign new_new_n2810__ = ~new_new_n2806__ & new_new_n2809__;
  assign new_new_n2811__ = new_new_n1692__ & ~new_new_n2810__;
  assign new_new_n2812__ = new_new_n2806__ & ~new_new_n2809__;
  assign new_new_n2813__ = ~new_new_n2811__ & ~new_new_n2812__;
  assign new_new_n2814__ = pi113 & ~new_new_n1156__;
  assign new_new_n2815__ = pi241 & new_new_n1156__;
  assign new_new_n2816__ = ~new_new_n2814__ & ~new_new_n2815__;
  assign new_new_n2817__ = new_new_n2813__ & new_new_n2816__;
  assign new_new_n2818__ = new_new_n1689__ & ~new_new_n2817__;
  assign new_new_n2819__ = ~new_new_n2813__ & ~new_new_n2816__;
  assign new_new_n2820__ = ~new_new_n2818__ & ~new_new_n2819__;
  assign new_new_n2821__ = pi114 & ~new_new_n1156__;
  assign new_new_n2822__ = pi242 & new_new_n1156__;
  assign new_new_n2823__ = ~new_new_n2821__ & ~new_new_n2822__;
  assign new_new_n2824__ = new_new_n2820__ & new_new_n2823__;
  assign new_new_n2825__ = new_new_n1686__ & ~new_new_n2824__;
  assign new_new_n2826__ = ~new_new_n2820__ & ~new_new_n2823__;
  assign new_new_n2827__ = ~new_new_n2825__ & ~new_new_n2826__;
  assign new_new_n2828__ = pi115 & ~new_new_n1156__;
  assign new_new_n2829__ = pi243 & new_new_n1156__;
  assign new_new_n2830__ = ~new_new_n2828__ & ~new_new_n2829__;
  assign new_new_n2831__ = new_new_n2827__ & new_new_n2830__;
  assign new_new_n2832__ = new_new_n1683__ & ~new_new_n2831__;
  assign new_new_n2833__ = ~new_new_n2827__ & ~new_new_n2830__;
  assign new_new_n2834__ = ~new_new_n2832__ & ~new_new_n2833__;
  assign new_new_n2835__ = pi116 & ~new_new_n1156__;
  assign new_new_n2836__ = pi244 & new_new_n1156__;
  assign new_new_n2837__ = ~new_new_n2835__ & ~new_new_n2836__;
  assign new_new_n2838__ = new_new_n2834__ & new_new_n2837__;
  assign new_new_n2839__ = new_new_n1680__ & ~new_new_n2838__;
  assign new_new_n2840__ = ~new_new_n2834__ & ~new_new_n2837__;
  assign new_new_n2841__ = ~new_new_n2839__ & ~new_new_n2840__;
  assign new_new_n2842__ = pi117 & ~new_new_n1156__;
  assign new_new_n2843__ = pi245 & new_new_n1156__;
  assign new_new_n2844__ = ~new_new_n2842__ & ~new_new_n2843__;
  assign new_new_n2845__ = new_new_n2841__ & new_new_n2844__;
  assign new_new_n2846__ = new_new_n1677__ & ~new_new_n2845__;
  assign new_new_n2847__ = ~new_new_n2841__ & ~new_new_n2844__;
  assign new_new_n2848__ = ~new_new_n2846__ & ~new_new_n2847__;
  assign new_new_n2849__ = pi118 & ~new_new_n1156__;
  assign new_new_n2850__ = pi246 & new_new_n1156__;
  assign new_new_n2851__ = ~new_new_n2849__ & ~new_new_n2850__;
  assign new_new_n2852__ = new_new_n2848__ & new_new_n2851__;
  assign new_new_n2853__ = ~new_new_n2848__ & ~new_new_n2851__;
  assign new_new_n2854__ = pi374 & ~new_new_n1674__;
  assign new_new_n2855__ = pi502 & new_new_n1674__;
  assign new_new_n2856__ = ~new_new_n2854__ & ~new_new_n2855__;
  assign new_new_n2857__ = ~new_new_n2853__ & ~new_new_n2856__;
  assign new_new_n2858__ = ~new_new_n2852__ & ~new_new_n2857__;
  assign new_new_n2859__ = pi119 & ~new_new_n1156__;
  assign new_new_n2860__ = pi247 & new_new_n1156__;
  assign new_new_n2861__ = ~new_new_n2859__ & ~new_new_n2860__;
  assign new_new_n2862__ = ~new_new_n2858__ & new_new_n2861__;
  assign new_new_n2863__ = new_new_n2858__ & ~new_new_n2861__;
  assign new_new_n2864__ = pi375 & ~new_new_n1674__;
  assign new_new_n2865__ = pi503 & new_new_n1674__;
  assign new_new_n2866__ = ~new_new_n2864__ & ~new_new_n2865__;
  assign new_new_n2867__ = ~new_new_n2863__ & ~new_new_n2866__;
  assign new_new_n2868__ = ~new_new_n2862__ & ~new_new_n2867__;
  assign new_new_n2869__ = pi120 & ~new_new_n1156__;
  assign new_new_n2870__ = pi248 & new_new_n1156__;
  assign new_new_n2871__ = ~new_new_n2869__ & ~new_new_n2870__;
  assign new_new_n2872__ = ~new_new_n2868__ & new_new_n2871__;
  assign new_new_n2873__ = new_new_n2868__ & ~new_new_n2871__;
  assign new_new_n2874__ = pi376 & ~new_new_n1674__;
  assign new_new_n2875__ = pi504 & new_new_n1674__;
  assign new_new_n2876__ = ~new_new_n2874__ & ~new_new_n2875__;
  assign new_new_n2877__ = ~new_new_n2873__ & ~new_new_n2876__;
  assign new_new_n2878__ = ~new_new_n2872__ & ~new_new_n2877__;
  assign new_new_n2879__ = pi121 & ~new_new_n1156__;
  assign new_new_n2880__ = pi249 & new_new_n1156__;
  assign new_new_n2881__ = ~new_new_n2879__ & ~new_new_n2880__;
  assign new_new_n2882__ = ~new_new_n2878__ & new_new_n2881__;
  assign new_new_n2883__ = new_new_n2878__ & ~new_new_n2881__;
  assign new_new_n2884__ = pi377 & ~new_new_n1674__;
  assign new_new_n2885__ = pi505 & new_new_n1674__;
  assign new_new_n2886__ = ~new_new_n2884__ & ~new_new_n2885__;
  assign new_new_n2887__ = ~new_new_n2883__ & ~new_new_n2886__;
  assign new_new_n2888__ = ~new_new_n2882__ & ~new_new_n2887__;
  assign new_new_n2889__ = pi122 & ~new_new_n1156__;
  assign new_new_n2890__ = pi250 & new_new_n1156__;
  assign new_new_n2891__ = ~new_new_n2889__ & ~new_new_n2890__;
  assign new_new_n2892__ = ~new_new_n2888__ & new_new_n2891__;
  assign new_new_n2893__ = new_new_n2888__ & ~new_new_n2891__;
  assign new_new_n2894__ = pi378 & ~new_new_n1674__;
  assign new_new_n2895__ = pi506 & new_new_n1674__;
  assign new_new_n2896__ = ~new_new_n2894__ & ~new_new_n2895__;
  assign new_new_n2897__ = ~new_new_n2893__ & ~new_new_n2896__;
  assign new_new_n2898__ = ~new_new_n2892__ & ~new_new_n2897__;
  assign new_new_n2899__ = pi123 & ~new_new_n1156__;
  assign new_new_n2900__ = pi251 & new_new_n1156__;
  assign new_new_n2901__ = ~new_new_n2899__ & ~new_new_n2900__;
  assign new_new_n2902__ = ~new_new_n2898__ & new_new_n2901__;
  assign new_new_n2903__ = new_new_n2898__ & ~new_new_n2901__;
  assign new_new_n2904__ = pi379 & ~new_new_n1674__;
  assign new_new_n2905__ = pi507 & new_new_n1674__;
  assign new_new_n2906__ = ~new_new_n2904__ & ~new_new_n2905__;
  assign new_new_n2907__ = ~new_new_n2903__ & ~new_new_n2906__;
  assign new_new_n2908__ = ~new_new_n2902__ & ~new_new_n2907__;
  assign new_new_n2909__ = pi124 & ~new_new_n1156__;
  assign new_new_n2910__ = pi252 & new_new_n1156__;
  assign new_new_n2911__ = ~new_new_n2909__ & ~new_new_n2910__;
  assign new_new_n2912__ = ~new_new_n2908__ & new_new_n2911__;
  assign new_new_n2913__ = new_new_n2908__ & ~new_new_n2911__;
  assign new_new_n2914__ = pi380 & ~new_new_n1674__;
  assign new_new_n2915__ = pi508 & new_new_n1674__;
  assign new_new_n2916__ = ~new_new_n2914__ & ~new_new_n2915__;
  assign new_new_n2917__ = ~new_new_n2913__ & ~new_new_n2916__;
  assign new_new_n2918__ = ~new_new_n2912__ & ~new_new_n2917__;
  assign new_new_n2919__ = pi125 & ~new_new_n1156__;
  assign new_new_n2920__ = pi253 & new_new_n1156__;
  assign new_new_n2921__ = ~new_new_n2919__ & ~new_new_n2920__;
  assign new_new_n2922__ = ~new_new_n2918__ & new_new_n2921__;
  assign new_new_n2923__ = new_new_n2918__ & ~new_new_n2921__;
  assign new_new_n2924__ = pi381 & ~new_new_n1674__;
  assign new_new_n2925__ = pi509 & new_new_n1674__;
  assign new_new_n2926__ = ~new_new_n2924__ & ~new_new_n2925__;
  assign new_new_n2927__ = ~new_new_n2923__ & ~new_new_n2926__;
  assign new_new_n2928__ = ~new_new_n2922__ & ~new_new_n2927__;
  assign new_new_n2929__ = pi382 & ~new_new_n1674__;
  assign new_new_n2930__ = pi510 & new_new_n1674__;
  assign new_new_n2931__ = ~new_new_n2929__ & ~new_new_n2930__;
  assign new_new_n2932__ = new_new_n2928__ & new_new_n2931__;
  assign new_new_n2933__ = ~new_new_n2928__ & ~new_new_n2931__;
  assign new_new_n2934__ = pi126 & ~new_new_n1156__;
  assign new_new_n2935__ = pi254 & new_new_n1156__;
  assign new_new_n2936__ = ~new_new_n2934__ & ~new_new_n2935__;
  assign new_new_n2937__ = ~new_new_n2933__ & ~new_new_n2936__;
  assign new_new_n2938__ = ~new_new_n2932__ & ~new_new_n2937__;
  assign new_new_n2939__ = new_new_n1160__ & ~new_new_n2938__;
  assign new_new_n2940__ = pi127 & pi255;
  assign new_new_n2941__ = ~new_new_n1160__ & new_new_n2938__;
  assign new_new_n2942__ = ~new_new_n2940__ & ~new_new_n2941__;
  assign po129 = ~new_new_n2939__ & ~new_new_n2942__;
  assign new_new_n2944__ = ~new_new_n1159__ & ~po129;
  assign new_new_n2945__ = ~new_new_n1869__ & po129;
  assign po000 = new_new_n2944__ | new_new_n2945__;
  assign new_new_n2947__ = ~new_new_n1873__ & ~po129;
  assign new_new_n2948__ = ~new_new_n1866__ & po129;
  assign po001 = new_new_n2947__ | new_new_n2948__;
  assign new_new_n2950__ = ~new_new_n1880__ & ~po129;
  assign new_new_n2951__ = ~new_new_n1863__ & po129;
  assign po002 = new_new_n2950__ | new_new_n2951__;
  assign new_new_n2953__ = ~new_new_n1887__ & ~po129;
  assign new_new_n2954__ = ~new_new_n1860__ & po129;
  assign po003 = new_new_n2953__ | new_new_n2954__;
  assign new_new_n2956__ = ~new_new_n1894__ & ~po129;
  assign new_new_n2957__ = ~new_new_n1857__ & po129;
  assign po004 = new_new_n2956__ | new_new_n2957__;
  assign new_new_n2959__ = ~new_new_n1906__ & ~po129;
  assign new_new_n2960__ = ~new_new_n1901__ & po129;
  assign po005 = new_new_n2959__ | new_new_n2960__;
  assign new_new_n2962__ = ~new_new_n1854__ & ~po129;
  assign new_new_n2963__ = ~new_new_n1911__ & po129;
  assign po006 = new_new_n2962__ | new_new_n2963__;
  assign new_new_n2965__ = ~new_new_n1851__ & ~po129;
  assign new_new_n2966__ = ~new_new_n1918__ & po129;
  assign po007 = new_new_n2965__ | new_new_n2966__;
  assign new_new_n2968__ = ~new_new_n1930__ & ~po129;
  assign new_new_n2969__ = ~new_new_n1925__ & po129;
  assign po008 = new_new_n2968__ | new_new_n2969__;
  assign new_new_n2971__ = ~new_new_n1848__ & ~po129;
  assign new_new_n2972__ = ~new_new_n1935__ & po129;
  assign po009 = new_new_n2971__ | new_new_n2972__;
  assign new_new_n2974__ = ~new_new_n1845__ & ~po129;
  assign new_new_n2975__ = ~new_new_n1942__ & po129;
  assign po010 = new_new_n2974__ | new_new_n2975__;
  assign new_new_n2977__ = ~new_new_n1954__ & ~po129;
  assign new_new_n2978__ = ~new_new_n1949__ & po129;
  assign po011 = new_new_n2977__ | new_new_n2978__;
  assign new_new_n2980__ = ~new_new_n1959__ & ~po129;
  assign new_new_n2981__ = ~new_new_n1964__ & po129;
  assign po012 = new_new_n2980__ | new_new_n2981__;
  assign new_new_n2983__ = ~new_new_n1969__ & ~po129;
  assign new_new_n2984__ = ~new_new_n1974__ & po129;
  assign po013 = new_new_n2983__ | new_new_n2984__;
  assign new_new_n2986__ = ~new_new_n1979__ & ~po129;
  assign new_new_n2987__ = ~new_new_n1984__ & po129;
  assign po014 = new_new_n2986__ | new_new_n2987__;
  assign new_new_n2989__ = ~new_new_n1989__ & ~po129;
  assign new_new_n2990__ = ~new_new_n1842__ & po129;
  assign po015 = new_new_n2989__ | new_new_n2990__;
  assign new_new_n2992__ = ~new_new_n1996__ & ~po129;
  assign new_new_n2993__ = ~new_new_n1839__ & po129;
  assign po016 = new_new_n2992__ | new_new_n2993__;
  assign new_new_n2995__ = ~new_new_n2003__ & ~po129;
  assign new_new_n2996__ = ~new_new_n2008__ & po129;
  assign po017 = new_new_n2995__ | new_new_n2996__;
  assign new_new_n2998__ = ~new_new_n2013__ & ~po129;
  assign new_new_n2999__ = ~new_new_n2018__ & po129;
  assign po018 = new_new_n2998__ | new_new_n2999__;
  assign new_new_n3001__ = ~new_new_n2023__ & ~po129;
  assign new_new_n3002__ = ~new_new_n2028__ & po129;
  assign po019 = new_new_n3001__ | new_new_n3002__;
  assign new_new_n3004__ = ~new_new_n2033__ & ~po129;
  assign new_new_n3005__ = ~new_new_n2038__ & po129;
  assign po020 = new_new_n3004__ | new_new_n3005__;
  assign new_new_n3007__ = ~new_new_n2043__ & ~po129;
  assign new_new_n3008__ = ~new_new_n1836__ & po129;
  assign po021 = new_new_n3007__ | new_new_n3008__;
  assign new_new_n3010__ = ~new_new_n2050__ & ~po129;
  assign new_new_n3011__ = ~new_new_n1833__ & po129;
  assign po022 = new_new_n3010__ | new_new_n3011__;
  assign new_new_n3013__ = ~new_new_n2057__ & ~po129;
  assign new_new_n3014__ = ~new_new_n1830__ & po129;
  assign po023 = new_new_n3013__ | new_new_n3014__;
  assign new_new_n3016__ = ~new_new_n2064__ & ~po129;
  assign new_new_n3017__ = ~new_new_n1827__ & po129;
  assign po024 = new_new_n3016__ | new_new_n3017__;
  assign new_new_n3019__ = ~new_new_n2076__ & ~po129;
  assign new_new_n3020__ = ~new_new_n2071__ & po129;
  assign po025 = new_new_n3019__ | new_new_n3020__;
  assign new_new_n3022__ = ~new_new_n1824__ & ~po129;
  assign new_new_n3023__ = ~new_new_n2081__ & po129;
  assign po026 = new_new_n3022__ | new_new_n3023__;
  assign new_new_n3025__ = ~new_new_n2088__ & ~po129;
  assign new_new_n3026__ = ~new_new_n2093__ & po129;
  assign po027 = new_new_n3025__ | new_new_n3026__;
  assign new_new_n3028__ = ~new_new_n2098__ & ~po129;
  assign new_new_n3029__ = ~new_new_n1821__ & po129;
  assign po028 = new_new_n3028__ | new_new_n3029__;
  assign new_new_n3031__ = ~new_new_n2105__ & ~po129;
  assign new_new_n3032__ = ~new_new_n1818__ & po129;
  assign po029 = new_new_n3031__ | new_new_n3032__;
  assign new_new_n3034__ = ~new_new_n2112__ & ~po129;
  assign new_new_n3035__ = ~new_new_n2117__ & po129;
  assign po030 = new_new_n3034__ | new_new_n3035__;
  assign new_new_n3037__ = ~new_new_n2127__ & ~po129;
  assign new_new_n3038__ = ~new_new_n2122__ & po129;
  assign po031 = new_new_n3037__ | new_new_n3038__;
  assign new_new_n3040__ = ~new_new_n2137__ & ~po129;
  assign new_new_n3041__ = ~new_new_n2132__ & po129;
  assign po032 = new_new_n3040__ | new_new_n3041__;
  assign new_new_n3043__ = ~new_new_n1815__ & ~po129;
  assign new_new_n3044__ = ~new_new_n2142__ & po129;
  assign po033 = new_new_n3043__ | new_new_n3044__;
  assign new_new_n3046__ = ~new_new_n2149__ & ~po129;
  assign new_new_n3047__ = ~new_new_n2154__ & po129;
  assign po034 = new_new_n3046__ | new_new_n3047__;
  assign new_new_n3049__ = ~new_new_n2159__ & ~po129;
  assign new_new_n3050__ = ~new_new_n1812__ & po129;
  assign po035 = new_new_n3049__ | new_new_n3050__;
  assign new_new_n3052__ = ~new_new_n2166__ & ~po129;
  assign new_new_n3053__ = ~new_new_n2171__ & po129;
  assign po036 = new_new_n3052__ | new_new_n3053__;
  assign new_new_n3055__ = ~new_new_n2176__ & ~po129;
  assign new_new_n3056__ = ~new_new_n2181__ & po129;
  assign po037 = new_new_n3055__ | new_new_n3056__;
  assign new_new_n3058__ = ~new_new_n2191__ & ~po129;
  assign new_new_n3059__ = ~new_new_n2186__ & po129;
  assign po038 = new_new_n3058__ | new_new_n3059__;
  assign new_new_n3061__ = ~new_new_n2201__ & ~po129;
  assign new_new_n3062__ = ~new_new_n2196__ & po129;
  assign po039 = new_new_n3061__ | new_new_n3062__;
  assign new_new_n3064__ = ~new_new_n2206__ & ~po129;
  assign new_new_n3065__ = ~new_new_n2211__ & po129;
  assign po040 = new_new_n3064__ | new_new_n3065__;
  assign new_new_n3067__ = ~new_new_n2221__ & ~po129;
  assign new_new_n3068__ = ~new_new_n2216__ & po129;
  assign po041 = new_new_n3067__ | new_new_n3068__;
  assign new_new_n3070__ = ~new_new_n2231__ & ~po129;
  assign new_new_n3071__ = ~new_new_n2226__ & po129;
  assign po042 = new_new_n3070__ | new_new_n3071__;
  assign new_new_n3073__ = ~new_new_n1809__ & ~po129;
  assign new_new_n3074__ = ~new_new_n2236__ & po129;
  assign po043 = new_new_n3073__ | new_new_n3074__;
  assign new_new_n3076__ = ~new_new_n2248__ & ~po129;
  assign new_new_n3077__ = ~new_new_n2243__ & po129;
  assign po044 = new_new_n3076__ | new_new_n3077__;
  assign new_new_n3079__ = ~new_new_n1806__ & ~po129;
  assign new_new_n3080__ = ~new_new_n2253__ & po129;
  assign po045 = new_new_n3079__ | new_new_n3080__;
  assign new_new_n3082__ = ~new_new_n2260__ & ~po129;
  assign new_new_n3083__ = ~new_new_n2265__ & po129;
  assign po046 = new_new_n3082__ | new_new_n3083__;
  assign new_new_n3085__ = ~new_new_n2270__ & ~po129;
  assign new_new_n3086__ = ~new_new_n1803__ & po129;
  assign po047 = new_new_n3085__ | new_new_n3086__;
  assign new_new_n3088__ = ~new_new_n2277__ & ~po129;
  assign new_new_n3089__ = ~new_new_n1800__ & po129;
  assign po048 = new_new_n3088__ | new_new_n3089__;
  assign new_new_n3091__ = ~new_new_n2284__ & ~po129;
  assign new_new_n3092__ = ~new_new_n2289__ & po129;
  assign po049 = new_new_n3091__ | new_new_n3092__;
  assign new_new_n3094__ = ~new_new_n2299__ & ~po129;
  assign new_new_n3095__ = ~new_new_n2294__ & po129;
  assign po050 = new_new_n3094__ | new_new_n3095__;
  assign new_new_n3097__ = ~new_new_n1797__ & ~po129;
  assign new_new_n3098__ = ~new_new_n2304__ & po129;
  assign po051 = new_new_n3097__ | new_new_n3098__;
  assign new_new_n3100__ = ~new_new_n1794__ & ~po129;
  assign new_new_n3101__ = ~new_new_n2311__ & po129;
  assign po052 = new_new_n3100__ | new_new_n3101__;
  assign new_new_n3103__ = ~new_new_n1791__ & ~po129;
  assign new_new_n3104__ = ~new_new_n2318__ & po129;
  assign po053 = new_new_n3103__ | new_new_n3104__;
  assign new_new_n3106__ = ~new_new_n2325__ & ~po129;
  assign new_new_n3107__ = ~new_new_n2330__ & po129;
  assign po054 = new_new_n3106__ | new_new_n3107__;
  assign new_new_n3109__ = ~new_new_n2340__ & ~po129;
  assign new_new_n3110__ = ~new_new_n2335__ & po129;
  assign po055 = new_new_n3109__ | new_new_n3110__;
  assign new_new_n3112__ = ~new_new_n2345__ & ~po129;
  assign new_new_n3113__ = ~new_new_n2350__ & po129;
  assign po056 = new_new_n3112__ | new_new_n3113__;
  assign new_new_n3115__ = ~new_new_n2360__ & ~po129;
  assign new_new_n3116__ = ~new_new_n2355__ & po129;
  assign po057 = new_new_n3115__ | new_new_n3116__;
  assign new_new_n3118__ = ~new_new_n1788__ & ~po129;
  assign new_new_n3119__ = ~new_new_n2365__ & po129;
  assign po058 = new_new_n3118__ | new_new_n3119__;
  assign new_new_n3121__ = ~new_new_n2377__ & ~po129;
  assign new_new_n3122__ = ~new_new_n2372__ & po129;
  assign po059 = new_new_n3121__ | new_new_n3122__;
  assign new_new_n3124__ = ~new_new_n2387__ & ~po129;
  assign new_new_n3125__ = ~new_new_n2382__ & po129;
  assign po060 = new_new_n3124__ | new_new_n3125__;
  assign new_new_n3127__ = ~new_new_n1785__ & ~po129;
  assign new_new_n3128__ = ~new_new_n2392__ & po129;
  assign po061 = new_new_n3127__ | new_new_n3128__;
  assign new_new_n3130__ = ~new_new_n2404__ & ~po129;
  assign new_new_n3131__ = ~new_new_n2399__ & po129;
  assign po062 = new_new_n3130__ | new_new_n3131__;
  assign new_new_n3133__ = ~new_new_n2414__ & ~po129;
  assign new_new_n3134__ = ~new_new_n2409__ & po129;
  assign po063 = new_new_n3133__ | new_new_n3134__;
  assign new_new_n3136__ = ~new_new_n2424__ & ~po129;
  assign new_new_n3137__ = ~new_new_n2419__ & po129;
  assign po064 = new_new_n3136__ | new_new_n3137__;
  assign new_new_n3139__ = ~new_new_n2429__ & ~po129;
  assign new_new_n3140__ = ~new_new_n2434__ & po129;
  assign po065 = new_new_n3139__ | new_new_n3140__;
  assign new_new_n3142__ = ~new_new_n2439__ & ~po129;
  assign new_new_n3143__ = ~new_new_n1782__ & po129;
  assign po066 = new_new_n3142__ | new_new_n3143__;
  assign new_new_n3145__ = ~new_new_n2446__ & ~po129;
  assign new_new_n3146__ = ~new_new_n1779__ & po129;
  assign po067 = new_new_n3145__ | new_new_n3146__;
  assign new_new_n3148__ = ~new_new_n2453__ & ~po129;
  assign new_new_n3149__ = ~new_new_n2458__ & po129;
  assign po068 = new_new_n3148__ | new_new_n3149__;
  assign new_new_n3151__ = ~new_new_n2463__ & ~po129;
  assign new_new_n3152__ = ~new_new_n2468__ & po129;
  assign po069 = new_new_n3151__ | new_new_n3152__;
  assign new_new_n3154__ = ~new_new_n2473__ & ~po129;
  assign new_new_n3155__ = ~new_new_n1776__ & po129;
  assign po070 = new_new_n3154__ | new_new_n3155__;
  assign new_new_n3157__ = ~new_new_n2480__ & ~po129;
  assign new_new_n3158__ = ~new_new_n2485__ & po129;
  assign po071 = new_new_n3157__ | new_new_n3158__;
  assign new_new_n3160__ = ~new_new_n2490__ & ~po129;
  assign new_new_n3161__ = ~new_new_n1773__ & po129;
  assign po072 = new_new_n3160__ | new_new_n3161__;
  assign new_new_n3163__ = ~new_new_n2497__ & ~po129;
  assign new_new_n3164__ = ~new_new_n2502__ & po129;
  assign po073 = new_new_n3163__ | new_new_n3164__;
  assign new_new_n3166__ = ~new_new_n2512__ & ~po129;
  assign new_new_n3167__ = ~new_new_n2507__ & po129;
  assign po074 = new_new_n3166__ | new_new_n3167__;
  assign new_new_n3169__ = ~new_new_n1770__ & ~po129;
  assign new_new_n3170__ = ~new_new_n2517__ & po129;
  assign po075 = new_new_n3169__ | new_new_n3170__;
  assign new_new_n3172__ = ~new_new_n1767__ & ~po129;
  assign new_new_n3173__ = ~new_new_n2524__ & po129;
  assign po076 = new_new_n3172__ | new_new_n3173__;
  assign new_new_n3175__ = ~new_new_n1764__ & ~po129;
  assign new_new_n3176__ = ~new_new_n2531__ & po129;
  assign po077 = new_new_n3175__ | new_new_n3176__;
  assign new_new_n3178__ = ~new_new_n1761__ & ~po129;
  assign new_new_n3179__ = ~new_new_n2538__ & po129;
  assign po078 = new_new_n3178__ | new_new_n3179__;
  assign new_new_n3181__ = ~new_new_n1758__ & ~po129;
  assign new_new_n3182__ = ~new_new_n2545__ & po129;
  assign po079 = new_new_n3181__ | new_new_n3182__;
  assign new_new_n3184__ = ~new_new_n1755__ & ~po129;
  assign new_new_n3185__ = ~new_new_n2552__ & po129;
  assign po080 = new_new_n3184__ | new_new_n3185__;
  assign new_new_n3187__ = ~new_new_n1752__ & ~po129;
  assign new_new_n3188__ = ~new_new_n2559__ & po129;
  assign po081 = new_new_n3187__ | new_new_n3188__;
  assign new_new_n3190__ = ~new_new_n2571__ & ~po129;
  assign new_new_n3191__ = ~new_new_n2566__ & po129;
  assign po082 = new_new_n3190__ | new_new_n3191__;
  assign new_new_n3193__ = ~new_new_n2576__ & ~po129;
  assign new_new_n3194__ = ~new_new_n2581__ & po129;
  assign po083 = new_new_n3193__ | new_new_n3194__;
  assign new_new_n3196__ = ~new_new_n2586__ & ~po129;
  assign new_new_n3197__ = ~new_new_n1749__ & po129;
  assign po084 = new_new_n3196__ | new_new_n3197__;
  assign new_new_n3199__ = ~new_new_n2598__ & ~po129;
  assign new_new_n3200__ = ~new_new_n2593__ & po129;
  assign po085 = new_new_n3199__ | new_new_n3200__;
  assign new_new_n3202__ = ~new_new_n1746__ & ~po129;
  assign new_new_n3203__ = ~new_new_n2603__ & po129;
  assign po086 = new_new_n3202__ | new_new_n3203__;
  assign new_new_n3205__ = ~new_new_n1743__ & ~po129;
  assign new_new_n3206__ = ~new_new_n2610__ & po129;
  assign po087 = new_new_n3205__ | new_new_n3206__;
  assign new_new_n3208__ = ~new_new_n1740__ & ~po129;
  assign new_new_n3209__ = ~new_new_n2617__ & po129;
  assign po088 = new_new_n3208__ | new_new_n3209__;
  assign new_new_n3211__ = ~new_new_n1737__ & ~po129;
  assign new_new_n3212__ = ~new_new_n2624__ & po129;
  assign po089 = new_new_n3211__ | new_new_n3212__;
  assign new_new_n3214__ = ~new_new_n2631__ & ~po129;
  assign new_new_n3215__ = ~new_new_n2636__ & po129;
  assign po090 = new_new_n3214__ | new_new_n3215__;
  assign new_new_n3217__ = ~new_new_n2641__ & ~po129;
  assign new_new_n3218__ = ~new_new_n1734__ & po129;
  assign po091 = new_new_n3217__ | new_new_n3218__;
  assign new_new_n3220__ = ~new_new_n2648__ & ~po129;
  assign new_new_n3221__ = ~new_new_n1731__ & po129;
  assign po092 = new_new_n3220__ | new_new_n3221__;
  assign new_new_n3223__ = ~new_new_n2655__ & ~po129;
  assign new_new_n3224__ = ~new_new_n1728__ & po129;
  assign po093 = new_new_n3223__ | new_new_n3224__;
  assign new_new_n3226__ = ~new_new_n2662__ & ~po129;
  assign new_new_n3227__ = ~new_new_n1725__ & po129;
  assign po094 = new_new_n3226__ | new_new_n3227__;
  assign new_new_n3229__ = ~new_new_n2669__ & ~po129;
  assign new_new_n3230__ = ~new_new_n1722__ & po129;
  assign po095 = new_new_n3229__ | new_new_n3230__;
  assign new_new_n3232__ = ~new_new_n2676__ & ~po129;
  assign new_new_n3233__ = ~new_new_n2681__ & po129;
  assign po096 = new_new_n3232__ | new_new_n3233__;
  assign new_new_n3235__ = ~new_new_n2686__ & ~po129;
  assign new_new_n3236__ = ~new_new_n2691__ & po129;
  assign po097 = new_new_n3235__ | new_new_n3236__;
  assign new_new_n3238__ = ~new_new_n2696__ & ~po129;
  assign new_new_n3239__ = ~new_new_n1719__ & po129;
  assign po098 = new_new_n3238__ | new_new_n3239__;
  assign new_new_n3241__ = ~new_new_n2703__ & ~po129;
  assign new_new_n3242__ = ~new_new_n2708__ & po129;
  assign po099 = new_new_n3241__ | new_new_n3242__;
  assign new_new_n3244__ = ~new_new_n2713__ & ~po129;
  assign new_new_n3245__ = ~new_new_n1716__ & po129;
  assign po100 = new_new_n3244__ | new_new_n3245__;
  assign new_new_n3247__ = ~new_new_n2720__ & ~po129;
  assign new_new_n3248__ = ~new_new_n1713__ & po129;
  assign po101 = new_new_n3247__ | new_new_n3248__;
  assign new_new_n3250__ = ~new_new_n2727__ & ~po129;
  assign new_new_n3251__ = ~new_new_n1710__ & po129;
  assign po102 = new_new_n3250__ | new_new_n3251__;
  assign new_new_n3253__ = ~new_new_n2734__ & ~po129;
  assign new_new_n3254__ = ~new_new_n1707__ & po129;
  assign po103 = new_new_n3253__ | new_new_n3254__;
  assign new_new_n3256__ = ~new_new_n2741__ & ~po129;
  assign new_new_n3257__ = ~new_new_n2746__ & po129;
  assign po104 = new_new_n3256__ | new_new_n3257__;
  assign new_new_n3259__ = ~new_new_n2751__ & ~po129;
  assign new_new_n3260__ = ~new_new_n2756__ & po129;
  assign po105 = new_new_n3259__ | new_new_n3260__;
  assign new_new_n3262__ = ~new_new_n2761__ & ~po129;
  assign new_new_n3263__ = ~new_new_n1704__ & po129;
  assign po106 = new_new_n3262__ | new_new_n3263__;
  assign new_new_n3265__ = ~new_new_n2768__ & ~po129;
  assign new_new_n3266__ = ~new_new_n1701__ & po129;
  assign po107 = new_new_n3265__ | new_new_n3266__;
  assign new_new_n3268__ = ~new_new_n2775__ & ~po129;
  assign new_new_n3269__ = ~new_new_n2780__ & po129;
  assign po108 = new_new_n3268__ | new_new_n3269__;
  assign new_new_n3271__ = ~new_new_n2785__ & ~po129;
  assign new_new_n3272__ = ~new_new_n1698__ & po129;
  assign po109 = new_new_n3271__ | new_new_n3272__;
  assign new_new_n3274__ = ~new_new_n2792__ & ~po129;
  assign new_new_n3275__ = ~new_new_n1695__ & po129;
  assign po110 = new_new_n3274__ | new_new_n3275__;
  assign new_new_n3277__ = ~new_new_n2799__ & ~po129;
  assign new_new_n3278__ = ~new_new_n2804__ & po129;
  assign po111 = new_new_n3277__ | new_new_n3278__;
  assign new_new_n3280__ = ~new_new_n2809__ & ~po129;
  assign new_new_n3281__ = ~new_new_n1692__ & po129;
  assign po112 = new_new_n3280__ | new_new_n3281__;
  assign new_new_n3283__ = ~new_new_n2816__ & ~po129;
  assign new_new_n3284__ = ~new_new_n1689__ & po129;
  assign po113 = new_new_n3283__ | new_new_n3284__;
  assign new_new_n3286__ = ~new_new_n2823__ & ~po129;
  assign new_new_n3287__ = ~new_new_n1686__ & po129;
  assign po114 = new_new_n3286__ | new_new_n3287__;
  assign new_new_n3289__ = ~new_new_n2830__ & ~po129;
  assign new_new_n3290__ = ~new_new_n1683__ & po129;
  assign po115 = new_new_n3289__ | new_new_n3290__;
  assign new_new_n3292__ = ~new_new_n2837__ & ~po129;
  assign new_new_n3293__ = ~new_new_n1680__ & po129;
  assign po116 = new_new_n3292__ | new_new_n3293__;
  assign new_new_n3295__ = ~new_new_n2844__ & ~po129;
  assign new_new_n3296__ = ~new_new_n1677__ & po129;
  assign po117 = new_new_n3295__ | new_new_n3296__;
  assign new_new_n3298__ = ~new_new_n2851__ & ~po129;
  assign new_new_n3299__ = ~new_new_n2856__ & po129;
  assign po118 = new_new_n3298__ | new_new_n3299__;
  assign new_new_n3301__ = ~new_new_n2861__ & ~po129;
  assign new_new_n3302__ = ~new_new_n2866__ & po129;
  assign po119 = new_new_n3301__ | new_new_n3302__;
  assign new_new_n3304__ = ~new_new_n2871__ & ~po129;
  assign new_new_n3305__ = ~new_new_n2876__ & po129;
  assign po120 = new_new_n3304__ | new_new_n3305__;
  assign new_new_n3307__ = ~new_new_n2881__ & ~po129;
  assign new_new_n3308__ = ~new_new_n2886__ & po129;
  assign po121 = new_new_n3307__ | new_new_n3308__;
  assign new_new_n3310__ = ~new_new_n2891__ & ~po129;
  assign new_new_n3311__ = ~new_new_n2896__ & po129;
  assign po122 = new_new_n3310__ | new_new_n3311__;
  assign new_new_n3313__ = ~new_new_n2901__ & ~po129;
  assign new_new_n3314__ = ~new_new_n2906__ & po129;
  assign po123 = new_new_n3313__ | new_new_n3314__;
  assign new_new_n3316__ = ~new_new_n2911__ & ~po129;
  assign new_new_n3317__ = ~new_new_n2916__ & po129;
  assign po124 = new_new_n3316__ | new_new_n3317__;
  assign new_new_n3319__ = ~new_new_n2921__ & ~po129;
  assign new_new_n3320__ = ~new_new_n2926__ & po129;
  assign po125 = new_new_n3319__ | new_new_n3320__;
  assign new_new_n3322__ = ~new_new_n2936__ & ~po129;
  assign new_new_n3323__ = ~new_new_n2931__ & po129;
  assign po126 = new_new_n3322__ | new_new_n3323__;
  assign po127 = new_new_n1160__ & new_new_n2940__;
  assign new_new_n3326__ = ~new_new_n1674__ & po129;
  assign new_new_n3327__ = ~new_new_n1156__ & ~po129;
  assign po128 = ~new_new_n3326__ & ~new_new_n3327__;
endmodule


