// Benchmark "bar" written by ABC on Wed Jul 13 18:48:48 2022

module bar ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \shift[0] , \shift[1] , \shift[2] ,
    \shift[3] , \shift[4] , \shift[5] , \shift[6] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \shift[0] , \shift[1] ,
    \shift[2] , \shift[3] , \shift[4] , \shift[5] , \shift[6] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ;
  wire new_new_n264__, new_new_n265__, new_new_n266__, new_new_n267__,
    new_new_n268__, new_new_n269__, new_new_n270__, new_new_n271__,
    new_new_n272__, new_new_n273__, new_new_n274__, new_new_n275__,
    new_new_n276__, new_new_n277__, new_new_n278__, new_new_n279__,
    new_new_n280__, new_new_n281__, new_new_n282__, new_new_n283__,
    new_new_n284__, new_new_n285__, new_new_n286__, new_new_n287__,
    new_new_n288__, new_new_n289__, new_new_n290__, new_new_n291__,
    new_new_n292__, new_new_n293__, new_new_n294__, new_new_n295__,
    new_new_n296__, new_new_n297__, new_new_n298__, new_new_n299__,
    new_new_n300__, new_new_n301__, new_new_n302__, new_new_n303__,
    new_new_n304__, new_new_n305__, new_new_n306__, new_new_n307__,
    new_new_n308__, new_new_n309__, new_new_n310__, new_new_n311__,
    new_new_n312__, new_new_n313__, new_new_n314__, new_new_n315__,
    new_new_n316__, new_new_n317__, new_new_n318__, new_new_n319__,
    new_new_n320__, new_new_n321__, new_new_n322__, new_new_n323__,
    new_new_n324__, new_new_n325__, new_new_n326__, new_new_n327__,
    new_new_n328__, new_new_n329__, new_new_n330__, new_new_n331__,
    new_new_n332__, new_new_n333__, new_new_n334__, new_new_n335__,
    new_new_n336__, new_new_n337__, new_new_n338__, new_new_n339__,
    new_new_n340__, new_new_n341__, new_new_n342__, new_new_n343__,
    new_new_n344__, new_new_n345__, new_new_n346__, new_new_n347__,
    new_new_n348__, new_new_n349__, new_new_n350__, new_new_n351__,
    new_new_n352__, new_new_n353__, new_new_n354__, new_new_n355__,
    new_new_n356__, new_new_n357__, new_new_n358__, new_new_n359__,
    new_new_n360__, new_new_n361__, new_new_n362__, new_new_n363__,
    new_new_n364__, new_new_n365__, new_new_n366__, new_new_n367__,
    new_new_n368__, new_new_n369__, new_new_n370__, new_new_n371__,
    new_new_n372__, new_new_n373__, new_new_n374__, new_new_n375__,
    new_new_n376__, new_new_n377__, new_new_n378__, new_new_n379__,
    new_new_n380__, new_new_n381__, new_new_n382__, new_new_n383__,
    new_new_n384__, new_new_n385__, new_new_n386__, new_new_n387__,
    new_new_n388__, new_new_n389__, new_new_n390__, new_new_n391__,
    new_new_n392__, new_new_n393__, new_new_n394__, new_new_n395__,
    new_new_n396__, new_new_n397__, new_new_n398__, new_new_n399__,
    new_new_n400__, new_new_n401__, new_new_n402__, new_new_n403__,
    new_new_n404__, new_new_n405__, new_new_n406__, new_new_n407__,
    new_new_n408__, new_new_n409__, new_new_n410__, new_new_n411__,
    new_new_n412__, new_new_n413__, new_new_n414__, new_new_n415__,
    new_new_n416__, new_new_n417__, new_new_n418__, new_new_n419__,
    new_new_n420__, new_new_n421__, new_new_n422__, new_new_n423__,
    new_new_n424__, new_new_n425__, new_new_n426__, new_new_n427__,
    new_new_n428__, new_new_n429__, new_new_n430__, new_new_n431__,
    new_new_n432__, new_new_n433__, new_new_n434__, new_new_n435__,
    new_new_n436__, new_new_n437__, new_new_n438__, new_new_n439__,
    new_new_n440__, new_new_n441__, new_new_n442__, new_new_n443__,
    new_new_n444__, new_new_n445__, new_new_n446__, new_new_n447__,
    new_new_n448__, new_new_n449__, new_new_n450__, new_new_n451__,
    new_new_n452__, new_new_n453__, new_new_n454__, new_new_n455__,
    new_new_n456__, new_new_n457__, new_new_n458__, new_new_n459__,
    new_new_n460__, new_new_n461__, new_new_n462__, new_new_n463__,
    new_new_n464__, new_new_n465__, new_new_n466__, new_new_n467__,
    new_new_n468__, new_new_n469__, new_new_n470__, new_new_n471__,
    new_new_n472__, new_new_n473__, new_new_n474__, new_new_n475__,
    new_new_n476__, new_new_n477__, new_new_n478__, new_new_n479__,
    new_new_n480__, new_new_n481__, new_new_n482__, new_new_n483__,
    new_new_n484__, new_new_n485__, new_new_n486__, new_new_n487__,
    new_new_n488__, new_new_n489__, new_new_n490__, new_new_n491__,
    new_new_n492__, new_new_n493__, new_new_n494__, new_new_n495__,
    new_new_n496__, new_new_n497__, new_new_n498__, new_new_n499__,
    new_new_n500__, new_new_n501__, new_new_n502__, new_new_n503__,
    new_new_n504__, new_new_n505__, new_new_n506__, new_new_n507__,
    new_new_n508__, new_new_n509__, new_new_n510__, new_new_n511__,
    new_new_n512__, new_new_n513__, new_new_n514__, new_new_n515__,
    new_new_n516__, new_new_n517__, new_new_n518__, new_new_n519__,
    new_new_n520__, new_new_n521__, new_new_n522__, new_new_n523__,
    new_new_n524__, new_new_n525__, new_new_n526__, new_new_n527__,
    new_new_n528__, new_new_n529__, new_new_n530__, new_new_n531__,
    new_new_n532__, new_new_n533__, new_new_n534__, new_new_n535__,
    new_new_n536__, new_new_n537__, new_new_n538__, new_new_n539__,
    new_new_n540__, new_new_n541__, new_new_n542__, new_new_n543__,
    new_new_n544__, new_new_n545__, new_new_n546__, new_new_n547__,
    new_new_n548__, new_new_n549__, new_new_n550__, new_new_n551__,
    new_new_n552__, new_new_n553__, new_new_n554__, new_new_n555__,
    new_new_n556__, new_new_n557__, new_new_n558__, new_new_n559__,
    new_new_n560__, new_new_n561__, new_new_n562__, new_new_n563__,
    new_new_n564__, new_new_n565__, new_new_n566__, new_new_n567__,
    new_new_n568__, new_new_n569__, new_new_n570__, new_new_n571__,
    new_new_n572__, new_new_n573__, new_new_n574__, new_new_n575__,
    new_new_n576__, new_new_n577__, new_new_n578__, new_new_n579__,
    new_new_n580__, new_new_n581__, new_new_n582__, new_new_n583__,
    new_new_n584__, new_new_n585__, new_new_n586__, new_new_n587__,
    new_new_n588__, new_new_n589__, new_new_n590__, new_new_n591__,
    new_new_n592__, new_new_n593__, new_new_n594__, new_new_n595__,
    new_new_n596__, new_new_n597__, new_new_n598__, new_new_n599__,
    new_new_n600__, new_new_n601__, new_new_n602__, new_new_n603__,
    new_new_n604__, new_new_n605__, new_new_n606__, new_new_n607__,
    new_new_n608__, new_new_n609__, new_new_n610__, new_new_n611__,
    new_new_n612__, new_new_n613__, new_new_n614__, new_new_n615__,
    new_new_n616__, new_new_n617__, new_new_n618__, new_new_n619__,
    new_new_n620__, new_new_n621__, new_new_n622__, new_new_n623__,
    new_new_n624__, new_new_n625__, new_new_n626__, new_new_n627__,
    new_new_n628__, new_new_n629__, new_new_n630__, new_new_n631__,
    new_new_n632__, new_new_n633__, new_new_n634__, new_new_n635__,
    new_new_n636__, new_new_n637__, new_new_n638__, new_new_n639__,
    new_new_n640__, new_new_n641__, new_new_n642__, new_new_n643__,
    new_new_n645__, new_new_n646__, new_new_n647__, new_new_n648__,
    new_new_n649__, new_new_n650__, new_new_n651__, new_new_n652__,
    new_new_n653__, new_new_n654__, new_new_n655__, new_new_n656__,
    new_new_n657__, new_new_n658__, new_new_n659__, new_new_n660__,
    new_new_n661__, new_new_n662__, new_new_n663__, new_new_n664__,
    new_new_n665__, new_new_n666__, new_new_n667__, new_new_n668__,
    new_new_n669__, new_new_n670__, new_new_n671__, new_new_n672__,
    new_new_n673__, new_new_n674__, new_new_n675__, new_new_n676__,
    new_new_n677__, new_new_n678__, new_new_n679__, new_new_n680__,
    new_new_n681__, new_new_n682__, new_new_n683__, new_new_n684__,
    new_new_n685__, new_new_n686__, new_new_n687__, new_new_n688__,
    new_new_n689__, new_new_n690__, new_new_n691__, new_new_n692__,
    new_new_n693__, new_new_n694__, new_new_n695__, new_new_n696__,
    new_new_n697__, new_new_n698__, new_new_n699__, new_new_n700__,
    new_new_n701__, new_new_n702__, new_new_n703__, new_new_n704__,
    new_new_n705__, new_new_n706__, new_new_n707__, new_new_n708__,
    new_new_n709__, new_new_n710__, new_new_n711__, new_new_n712__,
    new_new_n713__, new_new_n714__, new_new_n715__, new_new_n716__,
    new_new_n717__, new_new_n718__, new_new_n719__, new_new_n720__,
    new_new_n721__, new_new_n722__, new_new_n723__, new_new_n724__,
    new_new_n725__, new_new_n726__, new_new_n727__, new_new_n728__,
    new_new_n729__, new_new_n730__, new_new_n731__, new_new_n732__,
    new_new_n733__, new_new_n734__, new_new_n735__, new_new_n736__,
    new_new_n737__, new_new_n738__, new_new_n739__, new_new_n740__,
    new_new_n741__, new_new_n742__, new_new_n743__, new_new_n744__,
    new_new_n745__, new_new_n746__, new_new_n747__, new_new_n748__,
    new_new_n749__, new_new_n750__, new_new_n751__, new_new_n752__,
    new_new_n753__, new_new_n754__, new_new_n755__, new_new_n756__,
    new_new_n757__, new_new_n758__, new_new_n759__, new_new_n760__,
    new_new_n761__, new_new_n762__, new_new_n763__, new_new_n764__,
    new_new_n765__, new_new_n766__, new_new_n767__, new_new_n768__,
    new_new_n769__, new_new_n770__, new_new_n771__, new_new_n772__,
    new_new_n773__, new_new_n774__, new_new_n775__, new_new_n776__,
    new_new_n777__, new_new_n778__, new_new_n779__, new_new_n780__,
    new_new_n781__, new_new_n782__, new_new_n783__, new_new_n784__,
    new_new_n785__, new_new_n786__, new_new_n787__, new_new_n788__,
    new_new_n789__, new_new_n790__, new_new_n791__, new_new_n792__,
    new_new_n793__, new_new_n794__, new_new_n795__, new_new_n796__,
    new_new_n797__, new_new_n798__, new_new_n799__, new_new_n800__,
    new_new_n801__, new_new_n802__, new_new_n803__, new_new_n804__,
    new_new_n805__, new_new_n806__, new_new_n807__, new_new_n808__,
    new_new_n809__, new_new_n810__, new_new_n811__, new_new_n812__,
    new_new_n813__, new_new_n814__, new_new_n815__, new_new_n816__,
    new_new_n817__, new_new_n818__, new_new_n819__, new_new_n820__,
    new_new_n821__, new_new_n822__, new_new_n823__, new_new_n824__,
    new_new_n825__, new_new_n826__, new_new_n827__, new_new_n828__,
    new_new_n829__, new_new_n830__, new_new_n831__, new_new_n832__,
    new_new_n833__, new_new_n834__, new_new_n835__, new_new_n836__,
    new_new_n837__, new_new_n838__, new_new_n839__, new_new_n840__,
    new_new_n841__, new_new_n842__, new_new_n843__, new_new_n844__,
    new_new_n845__, new_new_n846__, new_new_n847__, new_new_n848__,
    new_new_n849__, new_new_n850__, new_new_n851__, new_new_n852__,
    new_new_n853__, new_new_n854__, new_new_n855__, new_new_n856__,
    new_new_n857__, new_new_n858__, new_new_n859__, new_new_n860__,
    new_new_n861__, new_new_n862__, new_new_n863__, new_new_n864__,
    new_new_n865__, new_new_n866__, new_new_n867__, new_new_n868__,
    new_new_n869__, new_new_n870__, new_new_n871__, new_new_n872__,
    new_new_n873__, new_new_n874__, new_new_n875__, new_new_n876__,
    new_new_n877__, new_new_n878__, new_new_n879__, new_new_n880__,
    new_new_n881__, new_new_n882__, new_new_n883__, new_new_n884__,
    new_new_n885__, new_new_n886__, new_new_n887__, new_new_n888__,
    new_new_n889__, new_new_n890__, new_new_n891__, new_new_n892__,
    new_new_n893__, new_new_n894__, new_new_n895__, new_new_n896__,
    new_new_n897__, new_new_n898__, new_new_n899__, new_new_n900__,
    new_new_n901__, new_new_n902__, new_new_n903__, new_new_n904__,
    new_new_n905__, new_new_n906__, new_new_n907__, new_new_n908__,
    new_new_n909__, new_new_n910__, new_new_n911__, new_new_n912__,
    new_new_n913__, new_new_n914__, new_new_n915__, new_new_n916__,
    new_new_n917__, new_new_n918__, new_new_n919__, new_new_n920__,
    new_new_n921__, new_new_n922__, new_new_n923__, new_new_n924__,
    new_new_n925__, new_new_n926__, new_new_n927__, new_new_n928__,
    new_new_n930__, new_new_n931__, new_new_n932__, new_new_n933__,
    new_new_n934__, new_new_n935__, new_new_n936__, new_new_n937__,
    new_new_n938__, new_new_n939__, new_new_n940__, new_new_n941__,
    new_new_n942__, new_new_n943__, new_new_n944__, new_new_n945__,
    new_new_n946__, new_new_n947__, new_new_n948__, new_new_n949__,
    new_new_n950__, new_new_n951__, new_new_n952__, new_new_n953__,
    new_new_n954__, new_new_n955__, new_new_n956__, new_new_n957__,
    new_new_n958__, new_new_n959__, new_new_n960__, new_new_n961__,
    new_new_n962__, new_new_n963__, new_new_n964__, new_new_n965__,
    new_new_n966__, new_new_n967__, new_new_n968__, new_new_n969__,
    new_new_n970__, new_new_n971__, new_new_n972__, new_new_n973__,
    new_new_n974__, new_new_n975__, new_new_n976__, new_new_n977__,
    new_new_n978__, new_new_n979__, new_new_n980__, new_new_n981__,
    new_new_n982__, new_new_n983__, new_new_n984__, new_new_n985__,
    new_new_n986__, new_new_n987__, new_new_n988__, new_new_n989__,
    new_new_n990__, new_new_n991__, new_new_n992__, new_new_n993__,
    new_new_n994__, new_new_n995__, new_new_n996__, new_new_n997__,
    new_new_n998__, new_new_n999__, new_new_n1000__, new_new_n1001__,
    new_new_n1002__, new_new_n1003__, new_new_n1004__, new_new_n1005__,
    new_new_n1006__, new_new_n1007__, new_new_n1008__, new_new_n1009__,
    new_new_n1010__, new_new_n1011__, new_new_n1012__, new_new_n1013__,
    new_new_n1014__, new_new_n1015__, new_new_n1016__, new_new_n1017__,
    new_new_n1018__, new_new_n1019__, new_new_n1020__, new_new_n1021__,
    new_new_n1022__, new_new_n1023__, new_new_n1024__, new_new_n1025__,
    new_new_n1026__, new_new_n1027__, new_new_n1028__, new_new_n1029__,
    new_new_n1030__, new_new_n1031__, new_new_n1032__, new_new_n1033__,
    new_new_n1034__, new_new_n1035__, new_new_n1036__, new_new_n1037__,
    new_new_n1038__, new_new_n1039__, new_new_n1040__, new_new_n1041__,
    new_new_n1042__, new_new_n1043__, new_new_n1044__, new_new_n1045__,
    new_new_n1046__, new_new_n1047__, new_new_n1048__, new_new_n1049__,
    new_new_n1050__, new_new_n1051__, new_new_n1052__, new_new_n1053__,
    new_new_n1054__, new_new_n1055__, new_new_n1056__, new_new_n1057__,
    new_new_n1058__, new_new_n1059__, new_new_n1060__, new_new_n1061__,
    new_new_n1062__, new_new_n1063__, new_new_n1064__, new_new_n1065__,
    new_new_n1066__, new_new_n1067__, new_new_n1068__, new_new_n1069__,
    new_new_n1070__, new_new_n1071__, new_new_n1072__, new_new_n1073__,
    new_new_n1074__, new_new_n1075__, new_new_n1076__, new_new_n1077__,
    new_new_n1078__, new_new_n1079__, new_new_n1080__, new_new_n1081__,
    new_new_n1082__, new_new_n1083__, new_new_n1084__, new_new_n1085__,
    new_new_n1086__, new_new_n1087__, new_new_n1088__, new_new_n1089__,
    new_new_n1090__, new_new_n1091__, new_new_n1092__, new_new_n1093__,
    new_new_n1094__, new_new_n1095__, new_new_n1096__, new_new_n1097__,
    new_new_n1098__, new_new_n1099__, new_new_n1100__, new_new_n1101__,
    new_new_n1102__, new_new_n1103__, new_new_n1104__, new_new_n1105__,
    new_new_n1106__, new_new_n1107__, new_new_n1108__, new_new_n1109__,
    new_new_n1110__, new_new_n1111__, new_new_n1112__, new_new_n1113__,
    new_new_n1114__, new_new_n1115__, new_new_n1116__, new_new_n1117__,
    new_new_n1118__, new_new_n1119__, new_new_n1120__, new_new_n1121__,
    new_new_n1122__, new_new_n1123__, new_new_n1124__, new_new_n1125__,
    new_new_n1126__, new_new_n1127__, new_new_n1128__, new_new_n1129__,
    new_new_n1130__, new_new_n1131__, new_new_n1132__, new_new_n1133__,
    new_new_n1134__, new_new_n1135__, new_new_n1136__, new_new_n1137__,
    new_new_n1138__, new_new_n1139__, new_new_n1140__, new_new_n1141__,
    new_new_n1142__, new_new_n1143__, new_new_n1144__, new_new_n1145__,
    new_new_n1146__, new_new_n1147__, new_new_n1148__, new_new_n1149__,
    new_new_n1150__, new_new_n1151__, new_new_n1152__, new_new_n1153__,
    new_new_n1154__, new_new_n1155__, new_new_n1156__, new_new_n1157__,
    new_new_n1158__, new_new_n1159__, new_new_n1160__, new_new_n1161__,
    new_new_n1162__, new_new_n1163__, new_new_n1164__, new_new_n1165__,
    new_new_n1166__, new_new_n1167__, new_new_n1168__, new_new_n1169__,
    new_new_n1170__, new_new_n1171__, new_new_n1172__, new_new_n1173__,
    new_new_n1174__, new_new_n1175__, new_new_n1176__, new_new_n1177__,
    new_new_n1178__, new_new_n1179__, new_new_n1180__, new_new_n1181__,
    new_new_n1182__, new_new_n1183__, new_new_n1184__, new_new_n1185__,
    new_new_n1186__, new_new_n1187__, new_new_n1188__, new_new_n1189__,
    new_new_n1190__, new_new_n1191__, new_new_n1192__, new_new_n1193__,
    new_new_n1194__, new_new_n1195__, new_new_n1196__, new_new_n1197__,
    new_new_n1198__, new_new_n1199__, new_new_n1200__, new_new_n1201__,
    new_new_n1202__, new_new_n1203__, new_new_n1204__, new_new_n1205__,
    new_new_n1206__, new_new_n1207__, new_new_n1208__, new_new_n1209__,
    new_new_n1210__, new_new_n1211__, new_new_n1212__, new_new_n1213__,
    new_new_n1215__, new_new_n1216__, new_new_n1217__, new_new_n1218__,
    new_new_n1219__, new_new_n1220__, new_new_n1221__, new_new_n1222__,
    new_new_n1223__, new_new_n1224__, new_new_n1225__, new_new_n1226__,
    new_new_n1227__, new_new_n1228__, new_new_n1229__, new_new_n1230__,
    new_new_n1231__, new_new_n1232__, new_new_n1233__, new_new_n1234__,
    new_new_n1235__, new_new_n1236__, new_new_n1237__, new_new_n1238__,
    new_new_n1239__, new_new_n1240__, new_new_n1241__, new_new_n1242__,
    new_new_n1243__, new_new_n1244__, new_new_n1245__, new_new_n1246__,
    new_new_n1247__, new_new_n1248__, new_new_n1249__, new_new_n1250__,
    new_new_n1251__, new_new_n1252__, new_new_n1253__, new_new_n1254__,
    new_new_n1255__, new_new_n1256__, new_new_n1257__, new_new_n1258__,
    new_new_n1259__, new_new_n1260__, new_new_n1261__, new_new_n1262__,
    new_new_n1263__, new_new_n1264__, new_new_n1265__, new_new_n1266__,
    new_new_n1267__, new_new_n1268__, new_new_n1269__, new_new_n1270__,
    new_new_n1271__, new_new_n1272__, new_new_n1273__, new_new_n1274__,
    new_new_n1275__, new_new_n1276__, new_new_n1277__, new_new_n1278__,
    new_new_n1279__, new_new_n1280__, new_new_n1281__, new_new_n1282__,
    new_new_n1283__, new_new_n1284__, new_new_n1285__, new_new_n1286__,
    new_new_n1287__, new_new_n1288__, new_new_n1289__, new_new_n1290__,
    new_new_n1291__, new_new_n1292__, new_new_n1293__, new_new_n1294__,
    new_new_n1295__, new_new_n1296__, new_new_n1297__, new_new_n1298__,
    new_new_n1299__, new_new_n1300__, new_new_n1301__, new_new_n1302__,
    new_new_n1303__, new_new_n1304__, new_new_n1305__, new_new_n1306__,
    new_new_n1307__, new_new_n1308__, new_new_n1309__, new_new_n1310__,
    new_new_n1311__, new_new_n1312__, new_new_n1313__, new_new_n1314__,
    new_new_n1315__, new_new_n1316__, new_new_n1317__, new_new_n1318__,
    new_new_n1319__, new_new_n1320__, new_new_n1321__, new_new_n1322__,
    new_new_n1323__, new_new_n1324__, new_new_n1325__, new_new_n1326__,
    new_new_n1327__, new_new_n1328__, new_new_n1329__, new_new_n1330__,
    new_new_n1331__, new_new_n1332__, new_new_n1333__, new_new_n1334__,
    new_new_n1335__, new_new_n1336__, new_new_n1337__, new_new_n1338__,
    new_new_n1339__, new_new_n1340__, new_new_n1341__, new_new_n1342__,
    new_new_n1343__, new_new_n1344__, new_new_n1345__, new_new_n1346__,
    new_new_n1347__, new_new_n1348__, new_new_n1349__, new_new_n1350__,
    new_new_n1351__, new_new_n1352__, new_new_n1353__, new_new_n1354__,
    new_new_n1355__, new_new_n1356__, new_new_n1357__, new_new_n1358__,
    new_new_n1359__, new_new_n1360__, new_new_n1361__, new_new_n1362__,
    new_new_n1363__, new_new_n1364__, new_new_n1365__, new_new_n1366__,
    new_new_n1367__, new_new_n1368__, new_new_n1369__, new_new_n1370__,
    new_new_n1371__, new_new_n1372__, new_new_n1373__, new_new_n1374__,
    new_new_n1375__, new_new_n1376__, new_new_n1377__, new_new_n1378__,
    new_new_n1379__, new_new_n1380__, new_new_n1381__, new_new_n1382__,
    new_new_n1383__, new_new_n1384__, new_new_n1385__, new_new_n1386__,
    new_new_n1387__, new_new_n1388__, new_new_n1389__, new_new_n1390__,
    new_new_n1391__, new_new_n1392__, new_new_n1393__, new_new_n1394__,
    new_new_n1395__, new_new_n1396__, new_new_n1397__, new_new_n1398__,
    new_new_n1399__, new_new_n1400__, new_new_n1401__, new_new_n1402__,
    new_new_n1404__, new_new_n1405__, new_new_n1406__, new_new_n1407__,
    new_new_n1408__, new_new_n1409__, new_new_n1410__, new_new_n1411__,
    new_new_n1412__, new_new_n1413__, new_new_n1414__, new_new_n1415__,
    new_new_n1416__, new_new_n1417__, new_new_n1418__, new_new_n1419__,
    new_new_n1420__, new_new_n1421__, new_new_n1422__, new_new_n1423__,
    new_new_n1424__, new_new_n1425__, new_new_n1426__, new_new_n1427__,
    new_new_n1428__, new_new_n1429__, new_new_n1430__, new_new_n1431__,
    new_new_n1432__, new_new_n1433__, new_new_n1434__, new_new_n1435__,
    new_new_n1436__, new_new_n1437__, new_new_n1438__, new_new_n1439__,
    new_new_n1440__, new_new_n1441__, new_new_n1442__, new_new_n1443__,
    new_new_n1444__, new_new_n1445__, new_new_n1446__, new_new_n1447__,
    new_new_n1448__, new_new_n1449__, new_new_n1450__, new_new_n1451__,
    new_new_n1452__, new_new_n1453__, new_new_n1454__, new_new_n1455__,
    new_new_n1456__, new_new_n1457__, new_new_n1458__, new_new_n1459__,
    new_new_n1460__, new_new_n1461__, new_new_n1462__, new_new_n1463__,
    new_new_n1464__, new_new_n1465__, new_new_n1466__, new_new_n1467__,
    new_new_n1468__, new_new_n1469__, new_new_n1470__, new_new_n1471__,
    new_new_n1473__, new_new_n1474__, new_new_n1475__, new_new_n1476__,
    new_new_n1477__, new_new_n1478__, new_new_n1479__, new_new_n1480__,
    new_new_n1481__, new_new_n1482__, new_new_n1483__, new_new_n1484__,
    new_new_n1485__, new_new_n1486__, new_new_n1487__, new_new_n1488__,
    new_new_n1489__, new_new_n1490__, new_new_n1491__, new_new_n1492__,
    new_new_n1493__, new_new_n1494__, new_new_n1495__, new_new_n1496__,
    new_new_n1497__, new_new_n1498__, new_new_n1499__, new_new_n1500__,
    new_new_n1501__, new_new_n1502__, new_new_n1503__, new_new_n1504__,
    new_new_n1505__, new_new_n1506__, new_new_n1507__, new_new_n1508__,
    new_new_n1509__, new_new_n1510__, new_new_n1511__, new_new_n1512__,
    new_new_n1513__, new_new_n1514__, new_new_n1515__, new_new_n1516__,
    new_new_n1517__, new_new_n1518__, new_new_n1519__, new_new_n1520__,
    new_new_n1521__, new_new_n1522__, new_new_n1523__, new_new_n1524__,
    new_new_n1525__, new_new_n1526__, new_new_n1527__, new_new_n1528__,
    new_new_n1529__, new_new_n1530__, new_new_n1531__, new_new_n1532__,
    new_new_n1533__, new_new_n1534__, new_new_n1535__, new_new_n1536__,
    new_new_n1537__, new_new_n1538__, new_new_n1539__, new_new_n1540__,
    new_new_n1542__, new_new_n1543__, new_new_n1544__, new_new_n1545__,
    new_new_n1546__, new_new_n1547__, new_new_n1548__, new_new_n1549__,
    new_new_n1550__, new_new_n1551__, new_new_n1552__, new_new_n1553__,
    new_new_n1554__, new_new_n1555__, new_new_n1556__, new_new_n1557__,
    new_new_n1558__, new_new_n1559__, new_new_n1560__, new_new_n1561__,
    new_new_n1562__, new_new_n1563__, new_new_n1564__, new_new_n1565__,
    new_new_n1566__, new_new_n1567__, new_new_n1568__, new_new_n1569__,
    new_new_n1570__, new_new_n1571__, new_new_n1572__, new_new_n1573__,
    new_new_n1574__, new_new_n1575__, new_new_n1576__, new_new_n1577__,
    new_new_n1578__, new_new_n1579__, new_new_n1580__, new_new_n1581__,
    new_new_n1582__, new_new_n1583__, new_new_n1584__, new_new_n1585__,
    new_new_n1586__, new_new_n1587__, new_new_n1588__, new_new_n1589__,
    new_new_n1590__, new_new_n1591__, new_new_n1592__, new_new_n1593__,
    new_new_n1594__, new_new_n1595__, new_new_n1596__, new_new_n1597__,
    new_new_n1598__, new_new_n1599__, new_new_n1600__, new_new_n1601__,
    new_new_n1602__, new_new_n1603__, new_new_n1604__, new_new_n1605__,
    new_new_n1606__, new_new_n1607__, new_new_n1608__, new_new_n1609__,
    new_new_n1611__, new_new_n1612__, new_new_n1613__, new_new_n1614__,
    new_new_n1615__, new_new_n1616__, new_new_n1617__, new_new_n1618__,
    new_new_n1619__, new_new_n1620__, new_new_n1621__, new_new_n1622__,
    new_new_n1623__, new_new_n1624__, new_new_n1625__, new_new_n1626__,
    new_new_n1627__, new_new_n1628__, new_new_n1629__, new_new_n1630__,
    new_new_n1631__, new_new_n1632__, new_new_n1633__, new_new_n1634__,
    new_new_n1635__, new_new_n1636__, new_new_n1637__, new_new_n1638__,
    new_new_n1639__, new_new_n1640__, new_new_n1641__, new_new_n1642__,
    new_new_n1643__, new_new_n1644__, new_new_n1645__, new_new_n1646__,
    new_new_n1647__, new_new_n1648__, new_new_n1649__, new_new_n1650__,
    new_new_n1651__, new_new_n1652__, new_new_n1653__, new_new_n1654__,
    new_new_n1655__, new_new_n1656__, new_new_n1657__, new_new_n1658__,
    new_new_n1659__, new_new_n1660__, new_new_n1661__, new_new_n1662__,
    new_new_n1663__, new_new_n1664__, new_new_n1665__, new_new_n1666__,
    new_new_n1667__, new_new_n1668__, new_new_n1669__, new_new_n1670__,
    new_new_n1671__, new_new_n1672__, new_new_n1673__, new_new_n1674__,
    new_new_n1675__, new_new_n1676__, new_new_n1677__, new_new_n1678__,
    new_new_n1680__, new_new_n1681__, new_new_n1682__, new_new_n1683__,
    new_new_n1684__, new_new_n1685__, new_new_n1686__, new_new_n1687__,
    new_new_n1688__, new_new_n1689__, new_new_n1690__, new_new_n1691__,
    new_new_n1692__, new_new_n1693__, new_new_n1694__, new_new_n1695__,
    new_new_n1696__, new_new_n1697__, new_new_n1698__, new_new_n1699__,
    new_new_n1700__, new_new_n1701__, new_new_n1702__, new_new_n1703__,
    new_new_n1704__, new_new_n1705__, new_new_n1706__, new_new_n1707__,
    new_new_n1708__, new_new_n1709__, new_new_n1710__, new_new_n1711__,
    new_new_n1712__, new_new_n1713__, new_new_n1714__, new_new_n1715__,
    new_new_n1716__, new_new_n1717__, new_new_n1718__, new_new_n1719__,
    new_new_n1720__, new_new_n1721__, new_new_n1722__, new_new_n1723__,
    new_new_n1724__, new_new_n1725__, new_new_n1726__, new_new_n1727__,
    new_new_n1728__, new_new_n1729__, new_new_n1730__, new_new_n1731__,
    new_new_n1732__, new_new_n1733__, new_new_n1734__, new_new_n1735__,
    new_new_n1736__, new_new_n1737__, new_new_n1738__, new_new_n1739__,
    new_new_n1740__, new_new_n1741__, new_new_n1742__, new_new_n1743__,
    new_new_n1744__, new_new_n1745__, new_new_n1746__, new_new_n1747__,
    new_new_n1749__, new_new_n1750__, new_new_n1751__, new_new_n1752__,
    new_new_n1753__, new_new_n1754__, new_new_n1755__, new_new_n1756__,
    new_new_n1757__, new_new_n1758__, new_new_n1759__, new_new_n1760__,
    new_new_n1761__, new_new_n1762__, new_new_n1763__, new_new_n1764__,
    new_new_n1765__, new_new_n1766__, new_new_n1767__, new_new_n1768__,
    new_new_n1769__, new_new_n1770__, new_new_n1771__, new_new_n1772__,
    new_new_n1773__, new_new_n1774__, new_new_n1775__, new_new_n1776__,
    new_new_n1777__, new_new_n1778__, new_new_n1779__, new_new_n1780__,
    new_new_n1781__, new_new_n1782__, new_new_n1783__, new_new_n1784__,
    new_new_n1785__, new_new_n1786__, new_new_n1787__, new_new_n1788__,
    new_new_n1789__, new_new_n1790__, new_new_n1791__, new_new_n1792__,
    new_new_n1793__, new_new_n1794__, new_new_n1795__, new_new_n1796__,
    new_new_n1797__, new_new_n1798__, new_new_n1799__, new_new_n1800__,
    new_new_n1801__, new_new_n1802__, new_new_n1803__, new_new_n1804__,
    new_new_n1805__, new_new_n1806__, new_new_n1807__, new_new_n1808__,
    new_new_n1809__, new_new_n1810__, new_new_n1811__, new_new_n1812__,
    new_new_n1813__, new_new_n1814__, new_new_n1815__, new_new_n1816__,
    new_new_n1818__, new_new_n1819__, new_new_n1820__, new_new_n1821__,
    new_new_n1822__, new_new_n1823__, new_new_n1824__, new_new_n1825__,
    new_new_n1826__, new_new_n1827__, new_new_n1828__, new_new_n1829__,
    new_new_n1830__, new_new_n1831__, new_new_n1832__, new_new_n1833__,
    new_new_n1834__, new_new_n1835__, new_new_n1836__, new_new_n1837__,
    new_new_n1838__, new_new_n1839__, new_new_n1840__, new_new_n1841__,
    new_new_n1842__, new_new_n1843__, new_new_n1844__, new_new_n1845__,
    new_new_n1846__, new_new_n1847__, new_new_n1848__, new_new_n1849__,
    new_new_n1850__, new_new_n1851__, new_new_n1852__, new_new_n1853__,
    new_new_n1854__, new_new_n1855__, new_new_n1856__, new_new_n1857__,
    new_new_n1858__, new_new_n1859__, new_new_n1860__, new_new_n1861__,
    new_new_n1862__, new_new_n1863__, new_new_n1864__, new_new_n1865__,
    new_new_n1866__, new_new_n1867__, new_new_n1868__, new_new_n1869__,
    new_new_n1870__, new_new_n1871__, new_new_n1872__, new_new_n1873__,
    new_new_n1874__, new_new_n1875__, new_new_n1876__, new_new_n1877__,
    new_new_n1878__, new_new_n1879__, new_new_n1880__, new_new_n1881__,
    new_new_n1882__, new_new_n1883__, new_new_n1884__, new_new_n1885__,
    new_new_n1887__, new_new_n1888__, new_new_n1889__, new_new_n1890__,
    new_new_n1891__, new_new_n1892__, new_new_n1893__, new_new_n1894__,
    new_new_n1895__, new_new_n1896__, new_new_n1897__, new_new_n1898__,
    new_new_n1899__, new_new_n1900__, new_new_n1901__, new_new_n1902__,
    new_new_n1903__, new_new_n1904__, new_new_n1905__, new_new_n1906__,
    new_new_n1907__, new_new_n1908__, new_new_n1909__, new_new_n1910__,
    new_new_n1911__, new_new_n1912__, new_new_n1913__, new_new_n1914__,
    new_new_n1915__, new_new_n1916__, new_new_n1917__, new_new_n1918__,
    new_new_n1919__, new_new_n1920__, new_new_n1921__, new_new_n1922__,
    new_new_n1923__, new_new_n1924__, new_new_n1925__, new_new_n1926__,
    new_new_n1927__, new_new_n1928__, new_new_n1929__, new_new_n1930__,
    new_new_n1931__, new_new_n1932__, new_new_n1933__, new_new_n1934__,
    new_new_n1935__, new_new_n1936__, new_new_n1937__, new_new_n1938__,
    new_new_n1939__, new_new_n1940__, new_new_n1941__, new_new_n1942__,
    new_new_n1943__, new_new_n1944__, new_new_n1945__, new_new_n1946__,
    new_new_n1947__, new_new_n1948__, new_new_n1949__, new_new_n1950__,
    new_new_n1951__, new_new_n1952__, new_new_n1953__, new_new_n1954__,
    new_new_n1956__, new_new_n1957__, new_new_n1958__, new_new_n1959__,
    new_new_n1960__, new_new_n1961__, new_new_n1962__, new_new_n1963__,
    new_new_n1964__, new_new_n1965__, new_new_n1966__, new_new_n1967__,
    new_new_n1968__, new_new_n1969__, new_new_n1970__, new_new_n1971__,
    new_new_n1972__, new_new_n1973__, new_new_n1974__, new_new_n1975__,
    new_new_n1976__, new_new_n1977__, new_new_n1978__, new_new_n1979__,
    new_new_n1980__, new_new_n1981__, new_new_n1982__, new_new_n1983__,
    new_new_n1984__, new_new_n1985__, new_new_n1986__, new_new_n1987__,
    new_new_n1988__, new_new_n1989__, new_new_n1990__, new_new_n1991__,
    new_new_n1992__, new_new_n1993__, new_new_n1994__, new_new_n1995__,
    new_new_n1996__, new_new_n1997__, new_new_n1998__, new_new_n1999__,
    new_new_n2001__, new_new_n2002__, new_new_n2003__, new_new_n2004__,
    new_new_n2005__, new_new_n2006__, new_new_n2007__, new_new_n2008__,
    new_new_n2009__, new_new_n2010__, new_new_n2011__, new_new_n2012__,
    new_new_n2013__, new_new_n2014__, new_new_n2015__, new_new_n2016__,
    new_new_n2017__, new_new_n2018__, new_new_n2019__, new_new_n2020__,
    new_new_n2021__, new_new_n2022__, new_new_n2023__, new_new_n2024__,
    new_new_n2025__, new_new_n2026__, new_new_n2027__, new_new_n2028__,
    new_new_n2029__, new_new_n2030__, new_new_n2031__, new_new_n2032__,
    new_new_n2033__, new_new_n2034__, new_new_n2035__, new_new_n2036__,
    new_new_n2037__, new_new_n2038__, new_new_n2039__, new_new_n2040__,
    new_new_n2041__, new_new_n2042__, new_new_n2043__, new_new_n2044__,
    new_new_n2046__, new_new_n2047__, new_new_n2048__, new_new_n2049__,
    new_new_n2050__, new_new_n2051__, new_new_n2052__, new_new_n2053__,
    new_new_n2054__, new_new_n2055__, new_new_n2056__, new_new_n2057__,
    new_new_n2058__, new_new_n2059__, new_new_n2060__, new_new_n2061__,
    new_new_n2062__, new_new_n2063__, new_new_n2064__, new_new_n2065__,
    new_new_n2066__, new_new_n2067__, new_new_n2068__, new_new_n2069__,
    new_new_n2070__, new_new_n2071__, new_new_n2072__, new_new_n2073__,
    new_new_n2074__, new_new_n2075__, new_new_n2076__, new_new_n2077__,
    new_new_n2078__, new_new_n2079__, new_new_n2080__, new_new_n2081__,
    new_new_n2082__, new_new_n2083__, new_new_n2084__, new_new_n2085__,
    new_new_n2086__, new_new_n2087__, new_new_n2088__, new_new_n2089__,
    new_new_n2091__, new_new_n2092__, new_new_n2093__, new_new_n2094__,
    new_new_n2095__, new_new_n2096__, new_new_n2097__, new_new_n2098__,
    new_new_n2099__, new_new_n2100__, new_new_n2101__, new_new_n2102__,
    new_new_n2103__, new_new_n2104__, new_new_n2105__, new_new_n2106__,
    new_new_n2107__, new_new_n2108__, new_new_n2109__, new_new_n2110__,
    new_new_n2111__, new_new_n2112__, new_new_n2113__, new_new_n2114__,
    new_new_n2115__, new_new_n2116__, new_new_n2117__, new_new_n2118__,
    new_new_n2119__, new_new_n2120__, new_new_n2121__, new_new_n2122__,
    new_new_n2123__, new_new_n2124__, new_new_n2125__, new_new_n2126__,
    new_new_n2127__, new_new_n2128__, new_new_n2129__, new_new_n2130__,
    new_new_n2131__, new_new_n2132__, new_new_n2133__, new_new_n2134__,
    new_new_n2136__, new_new_n2137__, new_new_n2138__, new_new_n2139__,
    new_new_n2140__, new_new_n2141__, new_new_n2142__, new_new_n2143__,
    new_new_n2144__, new_new_n2145__, new_new_n2146__, new_new_n2147__,
    new_new_n2148__, new_new_n2149__, new_new_n2151__, new_new_n2152__,
    new_new_n2153__, new_new_n2154__, new_new_n2155__, new_new_n2156__,
    new_new_n2157__, new_new_n2158__, new_new_n2159__, new_new_n2160__,
    new_new_n2161__, new_new_n2162__, new_new_n2163__, new_new_n2164__,
    new_new_n2166__, new_new_n2167__, new_new_n2168__, new_new_n2169__,
    new_new_n2170__, new_new_n2171__, new_new_n2172__, new_new_n2173__,
    new_new_n2174__, new_new_n2175__, new_new_n2176__, new_new_n2177__,
    new_new_n2178__, new_new_n2179__, new_new_n2181__, new_new_n2182__,
    new_new_n2183__, new_new_n2184__, new_new_n2185__, new_new_n2186__,
    new_new_n2187__, new_new_n2188__, new_new_n2189__, new_new_n2190__,
    new_new_n2191__, new_new_n2192__, new_new_n2193__, new_new_n2194__,
    new_new_n2196__, new_new_n2197__, new_new_n2198__, new_new_n2199__,
    new_new_n2200__, new_new_n2201__, new_new_n2202__, new_new_n2203__,
    new_new_n2204__, new_new_n2205__, new_new_n2206__, new_new_n2207__,
    new_new_n2208__, new_new_n2209__, new_new_n2211__, new_new_n2212__,
    new_new_n2213__, new_new_n2214__, new_new_n2215__, new_new_n2216__,
    new_new_n2217__, new_new_n2218__, new_new_n2219__, new_new_n2220__,
    new_new_n2221__, new_new_n2222__, new_new_n2223__, new_new_n2224__,
    new_new_n2226__, new_new_n2227__, new_new_n2228__, new_new_n2229__,
    new_new_n2230__, new_new_n2231__, new_new_n2232__, new_new_n2233__,
    new_new_n2234__, new_new_n2235__, new_new_n2236__, new_new_n2237__,
    new_new_n2238__, new_new_n2239__, new_new_n2241__, new_new_n2242__,
    new_new_n2243__, new_new_n2244__, new_new_n2245__, new_new_n2246__,
    new_new_n2247__, new_new_n2248__, new_new_n2249__, new_new_n2250__,
    new_new_n2251__, new_new_n2252__, new_new_n2253__, new_new_n2254__,
    new_new_n2256__, new_new_n2257__, new_new_n2258__, new_new_n2259__,
    new_new_n2260__, new_new_n2261__, new_new_n2262__, new_new_n2263__,
    new_new_n2264__, new_new_n2265__, new_new_n2266__, new_new_n2267__,
    new_new_n2268__, new_new_n2269__, new_new_n2271__, new_new_n2272__,
    new_new_n2273__, new_new_n2274__, new_new_n2275__, new_new_n2276__,
    new_new_n2277__, new_new_n2278__, new_new_n2279__, new_new_n2280__,
    new_new_n2281__, new_new_n2282__, new_new_n2283__, new_new_n2284__,
    new_new_n2286__, new_new_n2287__, new_new_n2288__, new_new_n2289__,
    new_new_n2290__, new_new_n2291__, new_new_n2292__, new_new_n2293__,
    new_new_n2294__, new_new_n2295__, new_new_n2296__, new_new_n2297__,
    new_new_n2298__, new_new_n2299__, new_new_n2301__, new_new_n2302__,
    new_new_n2303__, new_new_n2304__, new_new_n2305__, new_new_n2306__,
    new_new_n2307__, new_new_n2308__, new_new_n2309__, new_new_n2310__,
    new_new_n2311__, new_new_n2312__, new_new_n2313__, new_new_n2314__,
    new_new_n2316__, new_new_n2317__, new_new_n2318__, new_new_n2319__,
    new_new_n2320__, new_new_n2321__, new_new_n2322__, new_new_n2323__,
    new_new_n2324__, new_new_n2325__, new_new_n2326__, new_new_n2327__,
    new_new_n2328__, new_new_n2329__, new_new_n2331__, new_new_n2332__,
    new_new_n2333__, new_new_n2334__, new_new_n2335__, new_new_n2336__,
    new_new_n2337__, new_new_n2338__, new_new_n2339__, new_new_n2340__,
    new_new_n2341__, new_new_n2342__, new_new_n2343__, new_new_n2344__,
    new_new_n2346__, new_new_n2347__, new_new_n2348__, new_new_n2349__,
    new_new_n2350__, new_new_n2351__, new_new_n2352__, new_new_n2353__,
    new_new_n2354__, new_new_n2355__, new_new_n2356__, new_new_n2357__,
    new_new_n2358__, new_new_n2359__, new_new_n2361__, new_new_n2362__,
    new_new_n2363__, new_new_n2364__, new_new_n2365__, new_new_n2366__,
    new_new_n2367__, new_new_n2368__, new_new_n2369__, new_new_n2370__,
    new_new_n2371__, new_new_n2372__, new_new_n2373__, new_new_n2374__,
    new_new_n2376__, new_new_n2377__, new_new_n2378__, new_new_n2379__,
    new_new_n2380__, new_new_n2381__, new_new_n2382__, new_new_n2383__,
    new_new_n2384__, new_new_n2385__, new_new_n2386__, new_new_n2387__,
    new_new_n2388__, new_new_n2389__, new_new_n2391__, new_new_n2392__,
    new_new_n2393__, new_new_n2394__, new_new_n2395__, new_new_n2396__,
    new_new_n2397__, new_new_n2398__, new_new_n2399__, new_new_n2400__,
    new_new_n2401__, new_new_n2402__, new_new_n2403__, new_new_n2404__,
    new_new_n2406__, new_new_n2407__, new_new_n2408__, new_new_n2409__,
    new_new_n2410__, new_new_n2411__, new_new_n2412__, new_new_n2413__,
    new_new_n2414__, new_new_n2415__, new_new_n2416__, new_new_n2417__,
    new_new_n2418__, new_new_n2419__, new_new_n2421__, new_new_n2422__,
    new_new_n2423__, new_new_n2424__, new_new_n2425__, new_new_n2426__,
    new_new_n2427__, new_new_n2428__, new_new_n2429__, new_new_n2430__,
    new_new_n2431__, new_new_n2432__, new_new_n2433__, new_new_n2434__,
    new_new_n2436__, new_new_n2437__, new_new_n2438__, new_new_n2439__,
    new_new_n2440__, new_new_n2441__, new_new_n2442__, new_new_n2443__,
    new_new_n2444__, new_new_n2445__, new_new_n2446__, new_new_n2447__,
    new_new_n2448__, new_new_n2449__, new_new_n2451__, new_new_n2452__,
    new_new_n2453__, new_new_n2454__, new_new_n2455__, new_new_n2456__,
    new_new_n2457__, new_new_n2458__, new_new_n2459__, new_new_n2460__,
    new_new_n2461__, new_new_n2462__, new_new_n2463__, new_new_n2464__,
    new_new_n2466__, new_new_n2467__, new_new_n2468__, new_new_n2469__,
    new_new_n2470__, new_new_n2471__, new_new_n2472__, new_new_n2473__,
    new_new_n2474__, new_new_n2475__, new_new_n2476__, new_new_n2477__,
    new_new_n2478__, new_new_n2479__, new_new_n2481__, new_new_n2482__,
    new_new_n2483__, new_new_n2484__, new_new_n2485__, new_new_n2486__,
    new_new_n2487__, new_new_n2488__, new_new_n2489__, new_new_n2490__,
    new_new_n2491__, new_new_n2492__, new_new_n2493__, new_new_n2494__,
    new_new_n2496__, new_new_n2497__, new_new_n2498__, new_new_n2499__,
    new_new_n2500__, new_new_n2501__, new_new_n2502__, new_new_n2503__,
    new_new_n2504__, new_new_n2505__, new_new_n2506__, new_new_n2507__,
    new_new_n2508__, new_new_n2509__, new_new_n2511__, new_new_n2512__,
    new_new_n2513__, new_new_n2514__, new_new_n2515__, new_new_n2516__,
    new_new_n2517__, new_new_n2518__, new_new_n2519__, new_new_n2520__,
    new_new_n2521__, new_new_n2522__, new_new_n2523__, new_new_n2524__,
    new_new_n2526__, new_new_n2527__, new_new_n2528__, new_new_n2529__,
    new_new_n2530__, new_new_n2531__, new_new_n2532__, new_new_n2533__,
    new_new_n2534__, new_new_n2535__, new_new_n2536__, new_new_n2537__,
    new_new_n2538__, new_new_n2539__, new_new_n2541__, new_new_n2542__,
    new_new_n2543__, new_new_n2544__, new_new_n2545__, new_new_n2546__,
    new_new_n2547__, new_new_n2548__, new_new_n2549__, new_new_n2550__,
    new_new_n2551__, new_new_n2552__, new_new_n2553__, new_new_n2554__,
    new_new_n2556__, new_new_n2557__, new_new_n2558__, new_new_n2559__,
    new_new_n2560__, new_new_n2561__, new_new_n2562__, new_new_n2563__,
    new_new_n2564__, new_new_n2565__, new_new_n2566__, new_new_n2567__,
    new_new_n2568__, new_new_n2569__, new_new_n2571__, new_new_n2572__,
    new_new_n2573__, new_new_n2574__, new_new_n2575__, new_new_n2576__,
    new_new_n2577__, new_new_n2578__, new_new_n2579__, new_new_n2580__,
    new_new_n2581__, new_new_n2582__, new_new_n2583__, new_new_n2584__,
    new_new_n2586__, new_new_n2587__, new_new_n2588__, new_new_n2589__,
    new_new_n2590__, new_new_n2591__, new_new_n2592__, new_new_n2593__,
    new_new_n2594__, new_new_n2595__, new_new_n2596__, new_new_n2597__,
    new_new_n2598__, new_new_n2599__, new_new_n2601__, new_new_n2602__,
    new_new_n2603__, new_new_n2604__, new_new_n2605__, new_new_n2606__,
    new_new_n2607__, new_new_n2608__, new_new_n2609__, new_new_n2610__,
    new_new_n2611__, new_new_n2612__, new_new_n2613__, new_new_n2614__,
    new_new_n2616__, new_new_n2617__, new_new_n2618__, new_new_n2619__,
    new_new_n2620__, new_new_n2621__, new_new_n2622__, new_new_n2623__,
    new_new_n2625__, new_new_n2626__, new_new_n2627__, new_new_n2628__,
    new_new_n2629__, new_new_n2630__, new_new_n2631__, new_new_n2632__,
    new_new_n2634__, new_new_n2635__, new_new_n2636__, new_new_n2637__,
    new_new_n2638__, new_new_n2639__, new_new_n2640__, new_new_n2641__,
    new_new_n2643__, new_new_n2644__, new_new_n2645__, new_new_n2646__,
    new_new_n2647__, new_new_n2648__, new_new_n2649__, new_new_n2650__,
    new_new_n2652__, new_new_n2653__, new_new_n2654__, new_new_n2655__,
    new_new_n2656__, new_new_n2657__, new_new_n2658__, new_new_n2659__,
    new_new_n2661__, new_new_n2662__, new_new_n2663__, new_new_n2664__,
    new_new_n2665__, new_new_n2666__, new_new_n2667__, new_new_n2668__,
    new_new_n2670__, new_new_n2671__, new_new_n2672__, new_new_n2673__,
    new_new_n2674__, new_new_n2675__, new_new_n2676__, new_new_n2677__,
    new_new_n2679__, new_new_n2680__, new_new_n2681__, new_new_n2682__,
    new_new_n2683__, new_new_n2684__, new_new_n2685__, new_new_n2686__,
    new_new_n2688__, new_new_n2689__, new_new_n2690__, new_new_n2691__,
    new_new_n2692__, new_new_n2693__, new_new_n2694__, new_new_n2695__,
    new_new_n2697__, new_new_n2698__, new_new_n2699__, new_new_n2700__,
    new_new_n2701__, new_new_n2702__, new_new_n2703__, new_new_n2704__,
    new_new_n2706__, new_new_n2707__, new_new_n2708__, new_new_n2709__,
    new_new_n2710__, new_new_n2711__, new_new_n2712__, new_new_n2713__,
    new_new_n2715__, new_new_n2716__, new_new_n2717__, new_new_n2718__,
    new_new_n2719__, new_new_n2720__, new_new_n2721__, new_new_n2722__,
    new_new_n2724__, new_new_n2725__, new_new_n2726__, new_new_n2727__,
    new_new_n2728__, new_new_n2729__, new_new_n2730__, new_new_n2731__,
    new_new_n2733__, new_new_n2734__, new_new_n2735__, new_new_n2736__,
    new_new_n2737__, new_new_n2738__, new_new_n2739__, new_new_n2740__,
    new_new_n2742__, new_new_n2743__, new_new_n2744__, new_new_n2745__,
    new_new_n2746__, new_new_n2747__, new_new_n2748__, new_new_n2749__,
    new_new_n2751__, new_new_n2752__, new_new_n2753__, new_new_n2754__,
    new_new_n2755__, new_new_n2756__, new_new_n2757__, new_new_n2758__,
    new_new_n2760__, new_new_n2761__, new_new_n2763__, new_new_n2764__,
    new_new_n2766__, new_new_n2767__, new_new_n2769__, new_new_n2770__,
    new_new_n2772__, new_new_n2773__, new_new_n2775__, new_new_n2776__,
    new_new_n2778__, new_new_n2779__, new_new_n2781__, new_new_n2782__,
    new_new_n2784__, new_new_n2785__, new_new_n2787__, new_new_n2788__,
    new_new_n2790__, new_new_n2791__, new_new_n2793__, new_new_n2794__,
    new_new_n2796__, new_new_n2797__, new_new_n2799__, new_new_n2800__,
    new_new_n2802__, new_new_n2803__, new_new_n2805__, new_new_n2806__,
    new_new_n2808__, new_new_n2809__, new_new_n2811__, new_new_n2812__,
    new_new_n2814__, new_new_n2815__, new_new_n2817__, new_new_n2818__,
    new_new_n2820__, new_new_n2821__, new_new_n2823__, new_new_n2824__,
    new_new_n2826__, new_new_n2827__, new_new_n2829__, new_new_n2830__,
    new_new_n2832__, new_new_n2833__, new_new_n2835__, new_new_n2836__,
    new_new_n2838__, new_new_n2839__, new_new_n2841__, new_new_n2842__,
    new_new_n2844__, new_new_n2845__, new_new_n2847__, new_new_n2848__,
    new_new_n2850__, new_new_n2851__, new_new_n2853__, new_new_n2854__,
    new_new_n2856__, new_new_n2857__, new_new_n2859__, new_new_n2860__,
    new_new_n2862__, new_new_n2863__, new_new_n2865__, new_new_n2866__,
    new_new_n2868__, new_new_n2869__, new_new_n2871__, new_new_n2872__,
    new_new_n2874__, new_new_n2875__, new_new_n2877__, new_new_n2878__,
    new_new_n2880__, new_new_n2881__, new_new_n2883__, new_new_n2884__,
    new_new_n2886__, new_new_n2887__, new_new_n2889__, new_new_n2890__,
    new_new_n2892__, new_new_n2893__, new_new_n2895__, new_new_n2896__,
    new_new_n2898__, new_new_n2899__, new_new_n2901__, new_new_n2902__,
    new_new_n2904__, new_new_n2905__, new_new_n2907__, new_new_n2908__,
    new_new_n2910__, new_new_n2911__, new_new_n2913__, new_new_n2914__,
    new_new_n2916__, new_new_n2917__, new_new_n2919__, new_new_n2920__,
    new_new_n2922__, new_new_n2923__, new_new_n2925__, new_new_n2926__,
    new_new_n2928__, new_new_n2929__, new_new_n2931__, new_new_n2932__,
    new_new_n2934__, new_new_n2935__, new_new_n2937__, new_new_n2938__,
    new_new_n2940__, new_new_n2941__, new_new_n2943__, new_new_n2944__,
    new_new_n2946__, new_new_n2947__, new_new_n2949__, new_new_n2950__;
  assign new_new_n264__ = ~\a[1]  & \shift[1] ;
  assign new_new_n265__ = ~\a[3]  & ~\shift[1] ;
  assign new_new_n266__ = ~new_new_n264__ & ~new_new_n265__;
  assign new_new_n267__ = \shift[0]  & ~new_new_n266__;
  assign new_new_n268__ = ~\a[4]  & ~\shift[1] ;
  assign new_new_n269__ = ~\a[2]  & \shift[1] ;
  assign new_new_n270__ = ~new_new_n268__ & ~new_new_n269__;
  assign new_new_n271__ = ~\shift[0]  & ~new_new_n270__;
  assign new_new_n272__ = ~new_new_n267__ & ~new_new_n271__;
  assign new_new_n273__ = \shift[3]  & ~new_new_n272__;
  assign new_new_n274__ = ~\a[9]  & \shift[1] ;
  assign new_new_n275__ = ~\a[11]  & ~\shift[1] ;
  assign new_new_n276__ = ~new_new_n274__ & ~new_new_n275__;
  assign new_new_n277__ = \shift[0]  & ~new_new_n276__;
  assign new_new_n278__ = ~\a[12]  & ~\shift[1] ;
  assign new_new_n279__ = ~\a[10]  & \shift[1] ;
  assign new_new_n280__ = ~new_new_n278__ & ~new_new_n279__;
  assign new_new_n281__ = ~\shift[0]  & ~new_new_n280__;
  assign new_new_n282__ = ~new_new_n277__ & ~new_new_n281__;
  assign new_new_n283__ = ~\shift[3]  & ~new_new_n282__;
  assign new_new_n284__ = ~new_new_n273__ & ~new_new_n283__;
  assign new_new_n285__ = \shift[2]  & ~new_new_n284__;
  assign new_new_n286__ = ~\a[5]  & \shift[1] ;
  assign new_new_n287__ = ~\a[7]  & ~\shift[1] ;
  assign new_new_n288__ = ~new_new_n286__ & ~new_new_n287__;
  assign new_new_n289__ = \shift[0]  & ~new_new_n288__;
  assign new_new_n290__ = ~\a[8]  & ~\shift[1] ;
  assign new_new_n291__ = ~\a[6]  & \shift[1] ;
  assign new_new_n292__ = ~new_new_n290__ & ~new_new_n291__;
  assign new_new_n293__ = ~\shift[0]  & ~new_new_n292__;
  assign new_new_n294__ = ~new_new_n289__ & ~new_new_n293__;
  assign new_new_n295__ = \shift[3]  & ~new_new_n294__;
  assign new_new_n296__ = ~\a[13]  & \shift[1] ;
  assign new_new_n297__ = ~\a[15]  & ~\shift[1] ;
  assign new_new_n298__ = ~new_new_n296__ & ~new_new_n297__;
  assign new_new_n299__ = \shift[0]  & ~new_new_n298__;
  assign new_new_n300__ = ~\a[16]  & ~\shift[1] ;
  assign new_new_n301__ = ~\a[14]  & \shift[1] ;
  assign new_new_n302__ = ~new_new_n300__ & ~new_new_n301__;
  assign new_new_n303__ = ~\shift[0]  & ~new_new_n302__;
  assign new_new_n304__ = ~new_new_n299__ & ~new_new_n303__;
  assign new_new_n305__ = ~\shift[3]  & ~new_new_n304__;
  assign new_new_n306__ = ~new_new_n295__ & ~new_new_n305__;
  assign new_new_n307__ = ~\shift[2]  & ~new_new_n306__;
  assign new_new_n308__ = ~new_new_n285__ & ~new_new_n307__;
  assign new_new_n309__ = \shift[5]  & ~new_new_n308__;
  assign new_new_n310__ = ~\a[48]  & ~\shift[1] ;
  assign new_new_n311__ = ~\a[46]  & \shift[1] ;
  assign new_new_n312__ = ~new_new_n310__ & ~new_new_n311__;
  assign new_new_n313__ = ~\shift[0]  & new_new_n312__;
  assign new_new_n314__ = \a[47]  & ~\shift[1] ;
  assign new_new_n315__ = \a[45]  & \shift[1] ;
  assign new_new_n316__ = ~new_new_n314__ & ~new_new_n315__;
  assign new_new_n317__ = \shift[0]  & ~new_new_n316__;
  assign new_new_n318__ = ~new_new_n313__ & ~new_new_n317__;
  assign new_new_n319__ = ~\shift[3]  & new_new_n318__;
  assign new_new_n320__ = \a[40]  & ~\shift[1] ;
  assign new_new_n321__ = \a[38]  & \shift[1] ;
  assign new_new_n322__ = ~new_new_n320__ & ~new_new_n321__;
  assign new_new_n323__ = ~\shift[0]  & new_new_n322__;
  assign new_new_n324__ = ~\a[39]  & ~\shift[1] ;
  assign new_new_n325__ = ~\a[37]  & \shift[1] ;
  assign new_new_n326__ = ~new_new_n324__ & ~new_new_n325__;
  assign new_new_n327__ = \shift[0]  & ~new_new_n326__;
  assign new_new_n328__ = ~new_new_n323__ & ~new_new_n327__;
  assign new_new_n329__ = \shift[3]  & ~new_new_n328__;
  assign new_new_n330__ = ~new_new_n319__ & ~new_new_n329__;
  assign new_new_n331__ = ~\shift[2]  & ~new_new_n330__;
  assign new_new_n332__ = ~\a[33]  & \shift[1] ;
  assign new_new_n333__ = ~\a[35]  & ~\shift[1] ;
  assign new_new_n334__ = ~new_new_n332__ & ~new_new_n333__;
  assign new_new_n335__ = \shift[0]  & ~new_new_n334__;
  assign new_new_n336__ = ~\a[36]  & ~\shift[1] ;
  assign new_new_n337__ = ~\a[34]  & \shift[1] ;
  assign new_new_n338__ = ~new_new_n336__ & ~new_new_n337__;
  assign new_new_n339__ = ~\shift[0]  & ~new_new_n338__;
  assign new_new_n340__ = ~new_new_n335__ & ~new_new_n339__;
  assign new_new_n341__ = \shift[3]  & ~new_new_n340__;
  assign new_new_n342__ = ~\a[41]  & \shift[1] ;
  assign new_new_n343__ = ~\a[43]  & ~\shift[1] ;
  assign new_new_n344__ = ~new_new_n342__ & ~new_new_n343__;
  assign new_new_n345__ = \shift[0]  & ~new_new_n344__;
  assign new_new_n346__ = \a[44]  & ~\shift[1] ;
  assign new_new_n347__ = \a[42]  & \shift[1] ;
  assign new_new_n348__ = ~new_new_n346__ & ~new_new_n347__;
  assign new_new_n349__ = ~\shift[0]  & new_new_n348__;
  assign new_new_n350__ = ~new_new_n345__ & ~new_new_n349__;
  assign new_new_n351__ = ~\shift[3]  & ~new_new_n350__;
  assign new_new_n352__ = ~new_new_n341__ & ~new_new_n351__;
  assign new_new_n353__ = \shift[2]  & ~new_new_n352__;
  assign new_new_n354__ = ~new_new_n331__ & ~new_new_n353__;
  assign new_new_n355__ = ~\shift[5]  & ~new_new_n354__;
  assign new_new_n356__ = ~new_new_n309__ & ~new_new_n355__;
  assign new_new_n357__ = \shift[4]  & ~new_new_n356__;
  assign new_new_n358__ = ~\a[17]  & \shift[1] ;
  assign new_new_n359__ = ~\a[19]  & ~\shift[1] ;
  assign new_new_n360__ = ~new_new_n358__ & ~new_new_n359__;
  assign new_new_n361__ = \shift[0]  & ~new_new_n360__;
  assign new_new_n362__ = ~\a[20]  & ~\shift[1] ;
  assign new_new_n363__ = ~\a[18]  & \shift[1] ;
  assign new_new_n364__ = ~new_new_n362__ & ~new_new_n363__;
  assign new_new_n365__ = ~\shift[0]  & ~new_new_n364__;
  assign new_new_n366__ = ~new_new_n361__ & ~new_new_n365__;
  assign new_new_n367__ = \shift[3]  & ~new_new_n366__;
  assign new_new_n368__ = ~\a[25]  & \shift[1] ;
  assign new_new_n369__ = ~\a[27]  & ~\shift[1] ;
  assign new_new_n370__ = ~new_new_n368__ & ~new_new_n369__;
  assign new_new_n371__ = \shift[0]  & ~new_new_n370__;
  assign new_new_n372__ = ~\a[28]  & ~\shift[1] ;
  assign new_new_n373__ = ~\a[26]  & \shift[1] ;
  assign new_new_n374__ = ~new_new_n372__ & ~new_new_n373__;
  assign new_new_n375__ = ~\shift[0]  & ~new_new_n374__;
  assign new_new_n376__ = ~new_new_n371__ & ~new_new_n375__;
  assign new_new_n377__ = ~\shift[3]  & ~new_new_n376__;
  assign new_new_n378__ = ~new_new_n367__ & ~new_new_n377__;
  assign new_new_n379__ = \shift[2]  & ~new_new_n378__;
  assign new_new_n380__ = ~\a[21]  & \shift[1] ;
  assign new_new_n381__ = ~\a[23]  & ~\shift[1] ;
  assign new_new_n382__ = ~new_new_n380__ & ~new_new_n381__;
  assign new_new_n383__ = \shift[0]  & ~new_new_n382__;
  assign new_new_n384__ = ~\a[24]  & ~\shift[1] ;
  assign new_new_n385__ = ~\a[22]  & \shift[1] ;
  assign new_new_n386__ = ~new_new_n384__ & ~new_new_n385__;
  assign new_new_n387__ = ~\shift[0]  & ~new_new_n386__;
  assign new_new_n388__ = ~new_new_n383__ & ~new_new_n387__;
  assign new_new_n389__ = \shift[3]  & ~new_new_n388__;
  assign new_new_n390__ = ~\a[29]  & \shift[1] ;
  assign new_new_n391__ = ~\a[31]  & ~\shift[1] ;
  assign new_new_n392__ = ~new_new_n390__ & ~new_new_n391__;
  assign new_new_n393__ = \shift[0]  & ~new_new_n392__;
  assign new_new_n394__ = ~\a[32]  & ~\shift[1] ;
  assign new_new_n395__ = ~\a[30]  & \shift[1] ;
  assign new_new_n396__ = ~new_new_n394__ & ~new_new_n395__;
  assign new_new_n397__ = ~\shift[0]  & ~new_new_n396__;
  assign new_new_n398__ = ~new_new_n393__ & ~new_new_n397__;
  assign new_new_n399__ = ~\shift[3]  & ~new_new_n398__;
  assign new_new_n400__ = ~new_new_n389__ & ~new_new_n399__;
  assign new_new_n401__ = ~\shift[2]  & ~new_new_n400__;
  assign new_new_n402__ = ~new_new_n379__ & ~new_new_n401__;
  assign new_new_n403__ = \shift[5]  & ~new_new_n402__;
  assign new_new_n404__ = ~\a[49]  & \shift[1] ;
  assign new_new_n405__ = ~\a[51]  & ~\shift[1] ;
  assign new_new_n406__ = ~new_new_n404__ & ~new_new_n405__;
  assign new_new_n407__ = \shift[0]  & ~new_new_n406__;
  assign new_new_n408__ = ~\a[52]  & ~\shift[1] ;
  assign new_new_n409__ = ~\a[50]  & \shift[1] ;
  assign new_new_n410__ = ~new_new_n408__ & ~new_new_n409__;
  assign new_new_n411__ = ~\shift[0]  & ~new_new_n410__;
  assign new_new_n412__ = ~new_new_n407__ & ~new_new_n411__;
  assign new_new_n413__ = \shift[3]  & ~new_new_n412__;
  assign new_new_n414__ = ~\a[57]  & \shift[1] ;
  assign new_new_n415__ = ~\a[59]  & ~\shift[1] ;
  assign new_new_n416__ = ~new_new_n414__ & ~new_new_n415__;
  assign new_new_n417__ = \shift[0]  & ~new_new_n416__;
  assign new_new_n418__ = ~\a[60]  & ~\shift[1] ;
  assign new_new_n419__ = ~\a[58]  & \shift[1] ;
  assign new_new_n420__ = ~new_new_n418__ & ~new_new_n419__;
  assign new_new_n421__ = ~\shift[0]  & ~new_new_n420__;
  assign new_new_n422__ = ~new_new_n417__ & ~new_new_n421__;
  assign new_new_n423__ = ~\shift[3]  & ~new_new_n422__;
  assign new_new_n424__ = ~new_new_n413__ & ~new_new_n423__;
  assign new_new_n425__ = \shift[2]  & ~new_new_n424__;
  assign new_new_n426__ = ~\a[53]  & \shift[1] ;
  assign new_new_n427__ = ~\a[55]  & ~\shift[1] ;
  assign new_new_n428__ = ~new_new_n426__ & ~new_new_n427__;
  assign new_new_n429__ = \shift[0]  & ~new_new_n428__;
  assign new_new_n430__ = ~\a[56]  & ~\shift[1] ;
  assign new_new_n431__ = ~\a[54]  & \shift[1] ;
  assign new_new_n432__ = ~new_new_n430__ & ~new_new_n431__;
  assign new_new_n433__ = ~\shift[0]  & ~new_new_n432__;
  assign new_new_n434__ = ~new_new_n429__ & ~new_new_n433__;
  assign new_new_n435__ = \shift[3]  & ~new_new_n434__;
  assign new_new_n436__ = ~\a[61]  & \shift[1] ;
  assign new_new_n437__ = ~\a[63]  & ~\shift[1] ;
  assign new_new_n438__ = ~new_new_n436__ & ~new_new_n437__;
  assign new_new_n439__ = \shift[0]  & ~new_new_n438__;
  assign new_new_n440__ = ~\a[64]  & ~\shift[1] ;
  assign new_new_n441__ = ~\a[62]  & \shift[1] ;
  assign new_new_n442__ = ~new_new_n440__ & ~new_new_n441__;
  assign new_new_n443__ = ~\shift[0]  & ~new_new_n442__;
  assign new_new_n444__ = ~new_new_n439__ & ~new_new_n443__;
  assign new_new_n445__ = ~\shift[3]  & ~new_new_n444__;
  assign new_new_n446__ = ~new_new_n435__ & ~new_new_n445__;
  assign new_new_n447__ = ~\shift[2]  & ~new_new_n446__;
  assign new_new_n448__ = ~new_new_n425__ & ~new_new_n447__;
  assign new_new_n449__ = ~\shift[5]  & ~new_new_n448__;
  assign new_new_n450__ = ~new_new_n403__ & ~new_new_n449__;
  assign new_new_n451__ = ~\shift[4]  & ~new_new_n450__;
  assign new_new_n452__ = ~new_new_n357__ & ~new_new_n451__;
  assign new_new_n453__ = \shift[6]  & ~new_new_n452__;
  assign new_new_n454__ = ~\a[65]  & \shift[1] ;
  assign new_new_n455__ = ~\a[67]  & ~\shift[1] ;
  assign new_new_n456__ = ~new_new_n454__ & ~new_new_n455__;
  assign new_new_n457__ = \shift[0]  & ~new_new_n456__;
  assign new_new_n458__ = ~\a[68]  & ~\shift[1] ;
  assign new_new_n459__ = ~\a[66]  & \shift[1] ;
  assign new_new_n460__ = ~new_new_n458__ & ~new_new_n459__;
  assign new_new_n461__ = ~\shift[0]  & ~new_new_n460__;
  assign new_new_n462__ = ~new_new_n457__ & ~new_new_n461__;
  assign new_new_n463__ = \shift[3]  & ~new_new_n462__;
  assign new_new_n464__ = ~\a[73]  & \shift[1] ;
  assign new_new_n465__ = ~\a[75]  & ~\shift[1] ;
  assign new_new_n466__ = ~new_new_n464__ & ~new_new_n465__;
  assign new_new_n467__ = \shift[0]  & ~new_new_n466__;
  assign new_new_n468__ = ~\a[76]  & ~\shift[1] ;
  assign new_new_n469__ = ~\a[74]  & \shift[1] ;
  assign new_new_n470__ = ~new_new_n468__ & ~new_new_n469__;
  assign new_new_n471__ = ~\shift[0]  & ~new_new_n470__;
  assign new_new_n472__ = ~new_new_n467__ & ~new_new_n471__;
  assign new_new_n473__ = ~\shift[3]  & ~new_new_n472__;
  assign new_new_n474__ = ~new_new_n463__ & ~new_new_n473__;
  assign new_new_n475__ = \shift[2]  & ~new_new_n474__;
  assign new_new_n476__ = ~\a[69]  & \shift[1] ;
  assign new_new_n477__ = ~\a[71]  & ~\shift[1] ;
  assign new_new_n478__ = ~new_new_n476__ & ~new_new_n477__;
  assign new_new_n479__ = \shift[0]  & ~new_new_n478__;
  assign new_new_n480__ = ~\a[72]  & ~\shift[1] ;
  assign new_new_n481__ = ~\a[70]  & \shift[1] ;
  assign new_new_n482__ = ~new_new_n480__ & ~new_new_n481__;
  assign new_new_n483__ = ~\shift[0]  & ~new_new_n482__;
  assign new_new_n484__ = ~new_new_n479__ & ~new_new_n483__;
  assign new_new_n485__ = \shift[3]  & ~new_new_n484__;
  assign new_new_n486__ = ~\a[77]  & \shift[1] ;
  assign new_new_n487__ = ~\a[79]  & ~\shift[1] ;
  assign new_new_n488__ = ~new_new_n486__ & ~new_new_n487__;
  assign new_new_n489__ = \shift[0]  & ~new_new_n488__;
  assign new_new_n490__ = ~\a[80]  & ~\shift[1] ;
  assign new_new_n491__ = ~\a[78]  & \shift[1] ;
  assign new_new_n492__ = ~new_new_n490__ & ~new_new_n491__;
  assign new_new_n493__ = ~\shift[0]  & ~new_new_n492__;
  assign new_new_n494__ = ~new_new_n489__ & ~new_new_n493__;
  assign new_new_n495__ = ~\shift[3]  & ~new_new_n494__;
  assign new_new_n496__ = ~new_new_n485__ & ~new_new_n495__;
  assign new_new_n497__ = ~\shift[2]  & ~new_new_n496__;
  assign new_new_n498__ = ~new_new_n475__ & ~new_new_n497__;
  assign new_new_n499__ = \shift[5]  & ~new_new_n498__;
  assign new_new_n500__ = ~\a[97]  & \shift[1] ;
  assign new_new_n501__ = ~\a[99]  & ~\shift[1] ;
  assign new_new_n502__ = ~new_new_n500__ & ~new_new_n501__;
  assign new_new_n503__ = \shift[0]  & ~new_new_n502__;
  assign new_new_n504__ = ~\a[100]  & ~\shift[1] ;
  assign new_new_n505__ = ~\a[98]  & \shift[1] ;
  assign new_new_n506__ = ~new_new_n504__ & ~new_new_n505__;
  assign new_new_n507__ = ~\shift[0]  & ~new_new_n506__;
  assign new_new_n508__ = ~new_new_n503__ & ~new_new_n507__;
  assign new_new_n509__ = \shift[3]  & ~new_new_n508__;
  assign new_new_n510__ = ~\a[105]  & \shift[1] ;
  assign new_new_n511__ = ~\a[107]  & ~\shift[1] ;
  assign new_new_n512__ = ~new_new_n510__ & ~new_new_n511__;
  assign new_new_n513__ = \shift[0]  & ~new_new_n512__;
  assign new_new_n514__ = ~\a[108]  & ~\shift[1] ;
  assign new_new_n515__ = ~\a[106]  & \shift[1] ;
  assign new_new_n516__ = ~new_new_n514__ & ~new_new_n515__;
  assign new_new_n517__ = ~\shift[0]  & ~new_new_n516__;
  assign new_new_n518__ = ~new_new_n513__ & ~new_new_n517__;
  assign new_new_n519__ = ~\shift[3]  & ~new_new_n518__;
  assign new_new_n520__ = ~new_new_n509__ & ~new_new_n519__;
  assign new_new_n521__ = \shift[2]  & ~new_new_n520__;
  assign new_new_n522__ = ~\a[101]  & \shift[1] ;
  assign new_new_n523__ = ~\a[103]  & ~\shift[1] ;
  assign new_new_n524__ = ~new_new_n522__ & ~new_new_n523__;
  assign new_new_n525__ = \shift[0]  & ~new_new_n524__;
  assign new_new_n526__ = ~\a[104]  & ~\shift[1] ;
  assign new_new_n527__ = ~\a[102]  & \shift[1] ;
  assign new_new_n528__ = ~new_new_n526__ & ~new_new_n527__;
  assign new_new_n529__ = ~\shift[0]  & ~new_new_n528__;
  assign new_new_n530__ = ~new_new_n525__ & ~new_new_n529__;
  assign new_new_n531__ = \shift[3]  & ~new_new_n530__;
  assign new_new_n532__ = ~\a[109]  & \shift[1] ;
  assign new_new_n533__ = ~\a[111]  & ~\shift[1] ;
  assign new_new_n534__ = ~new_new_n532__ & ~new_new_n533__;
  assign new_new_n535__ = \shift[0]  & ~new_new_n534__;
  assign new_new_n536__ = ~\a[112]  & ~\shift[1] ;
  assign new_new_n537__ = ~\a[110]  & \shift[1] ;
  assign new_new_n538__ = ~new_new_n536__ & ~new_new_n537__;
  assign new_new_n539__ = ~\shift[0]  & ~new_new_n538__;
  assign new_new_n540__ = ~new_new_n535__ & ~new_new_n539__;
  assign new_new_n541__ = ~\shift[3]  & ~new_new_n540__;
  assign new_new_n542__ = ~new_new_n531__ & ~new_new_n541__;
  assign new_new_n543__ = ~\shift[2]  & ~new_new_n542__;
  assign new_new_n544__ = ~new_new_n521__ & ~new_new_n543__;
  assign new_new_n545__ = ~\shift[5]  & ~new_new_n544__;
  assign new_new_n546__ = ~new_new_n499__ & ~new_new_n545__;
  assign new_new_n547__ = \shift[4]  & ~new_new_n546__;
  assign new_new_n548__ = ~\a[81]  & \shift[1] ;
  assign new_new_n549__ = ~\a[83]  & ~\shift[1] ;
  assign new_new_n550__ = ~new_new_n548__ & ~new_new_n549__;
  assign new_new_n551__ = \shift[0]  & ~new_new_n550__;
  assign new_new_n552__ = ~\a[84]  & ~\shift[1] ;
  assign new_new_n553__ = ~\a[82]  & \shift[1] ;
  assign new_new_n554__ = ~new_new_n552__ & ~new_new_n553__;
  assign new_new_n555__ = ~\shift[0]  & ~new_new_n554__;
  assign new_new_n556__ = ~new_new_n551__ & ~new_new_n555__;
  assign new_new_n557__ = \shift[3]  & ~new_new_n556__;
  assign new_new_n558__ = ~\a[89]  & \shift[1] ;
  assign new_new_n559__ = ~\a[91]  & ~\shift[1] ;
  assign new_new_n560__ = ~new_new_n558__ & ~new_new_n559__;
  assign new_new_n561__ = \shift[0]  & ~new_new_n560__;
  assign new_new_n562__ = ~\a[92]  & ~\shift[1] ;
  assign new_new_n563__ = ~\a[90]  & \shift[1] ;
  assign new_new_n564__ = ~new_new_n562__ & ~new_new_n563__;
  assign new_new_n565__ = ~\shift[0]  & ~new_new_n564__;
  assign new_new_n566__ = ~new_new_n561__ & ~new_new_n565__;
  assign new_new_n567__ = ~\shift[3]  & ~new_new_n566__;
  assign new_new_n568__ = ~new_new_n557__ & ~new_new_n567__;
  assign new_new_n569__ = \shift[2]  & ~new_new_n568__;
  assign new_new_n570__ = ~\a[85]  & \shift[1] ;
  assign new_new_n571__ = ~\a[87]  & ~\shift[1] ;
  assign new_new_n572__ = ~new_new_n570__ & ~new_new_n571__;
  assign new_new_n573__ = \shift[0]  & ~new_new_n572__;
  assign new_new_n574__ = ~\a[88]  & ~\shift[1] ;
  assign new_new_n575__ = ~\a[86]  & \shift[1] ;
  assign new_new_n576__ = ~new_new_n574__ & ~new_new_n575__;
  assign new_new_n577__ = ~\shift[0]  & ~new_new_n576__;
  assign new_new_n578__ = ~new_new_n573__ & ~new_new_n577__;
  assign new_new_n579__ = \shift[3]  & ~new_new_n578__;
  assign new_new_n580__ = ~\a[93]  & \shift[1] ;
  assign new_new_n581__ = ~\a[95]  & ~\shift[1] ;
  assign new_new_n582__ = ~new_new_n580__ & ~new_new_n581__;
  assign new_new_n583__ = \shift[0]  & ~new_new_n582__;
  assign new_new_n584__ = ~\a[96]  & ~\shift[1] ;
  assign new_new_n585__ = ~\a[94]  & \shift[1] ;
  assign new_new_n586__ = ~new_new_n584__ & ~new_new_n585__;
  assign new_new_n587__ = ~\shift[0]  & ~new_new_n586__;
  assign new_new_n588__ = ~new_new_n583__ & ~new_new_n587__;
  assign new_new_n589__ = ~\shift[3]  & ~new_new_n588__;
  assign new_new_n590__ = ~new_new_n579__ & ~new_new_n589__;
  assign new_new_n591__ = ~\shift[2]  & ~new_new_n590__;
  assign new_new_n592__ = ~new_new_n569__ & ~new_new_n591__;
  assign new_new_n593__ = \shift[5]  & ~new_new_n592__;
  assign new_new_n594__ = ~\a[113]  & \shift[1] ;
  assign new_new_n595__ = ~\a[115]  & ~\shift[1] ;
  assign new_new_n596__ = ~new_new_n594__ & ~new_new_n595__;
  assign new_new_n597__ = \shift[0]  & ~new_new_n596__;
  assign new_new_n598__ = ~\a[116]  & ~\shift[1] ;
  assign new_new_n599__ = ~\a[114]  & \shift[1] ;
  assign new_new_n600__ = ~new_new_n598__ & ~new_new_n599__;
  assign new_new_n601__ = ~\shift[0]  & ~new_new_n600__;
  assign new_new_n602__ = ~new_new_n597__ & ~new_new_n601__;
  assign new_new_n603__ = \shift[3]  & ~new_new_n602__;
  assign new_new_n604__ = ~\a[121]  & \shift[1] ;
  assign new_new_n605__ = ~\a[123]  & ~\shift[1] ;
  assign new_new_n606__ = ~new_new_n604__ & ~new_new_n605__;
  assign new_new_n607__ = \shift[0]  & ~new_new_n606__;
  assign new_new_n608__ = ~\a[124]  & ~\shift[1] ;
  assign new_new_n609__ = ~\a[122]  & \shift[1] ;
  assign new_new_n610__ = ~new_new_n608__ & ~new_new_n609__;
  assign new_new_n611__ = ~\shift[0]  & ~new_new_n610__;
  assign new_new_n612__ = ~new_new_n607__ & ~new_new_n611__;
  assign new_new_n613__ = ~\shift[3]  & ~new_new_n612__;
  assign new_new_n614__ = ~new_new_n603__ & ~new_new_n613__;
  assign new_new_n615__ = \shift[2]  & ~new_new_n614__;
  assign new_new_n616__ = ~\a[117]  & \shift[1] ;
  assign new_new_n617__ = ~\a[119]  & ~\shift[1] ;
  assign new_new_n618__ = ~new_new_n616__ & ~new_new_n617__;
  assign new_new_n619__ = \shift[0]  & ~new_new_n618__;
  assign new_new_n620__ = ~\a[120]  & ~\shift[1] ;
  assign new_new_n621__ = ~\a[118]  & \shift[1] ;
  assign new_new_n622__ = ~new_new_n620__ & ~new_new_n621__;
  assign new_new_n623__ = ~\shift[0]  & ~new_new_n622__;
  assign new_new_n624__ = ~new_new_n619__ & ~new_new_n623__;
  assign new_new_n625__ = \shift[3]  & ~new_new_n624__;
  assign new_new_n626__ = ~\a[125]  & \shift[1] ;
  assign new_new_n627__ = ~\a[127]  & ~\shift[1] ;
  assign new_new_n628__ = ~new_new_n626__ & ~new_new_n627__;
  assign new_new_n629__ = \shift[0]  & ~new_new_n628__;
  assign new_new_n630__ = ~\a[0]  & ~\shift[1] ;
  assign new_new_n631__ = ~\a[126]  & \shift[1] ;
  assign new_new_n632__ = ~new_new_n630__ & ~new_new_n631__;
  assign new_new_n633__ = ~\shift[0]  & ~new_new_n632__;
  assign new_new_n634__ = ~new_new_n629__ & ~new_new_n633__;
  assign new_new_n635__ = ~\shift[3]  & ~new_new_n634__;
  assign new_new_n636__ = ~new_new_n625__ & ~new_new_n635__;
  assign new_new_n637__ = ~\shift[2]  & ~new_new_n636__;
  assign new_new_n638__ = ~new_new_n615__ & ~new_new_n637__;
  assign new_new_n639__ = ~\shift[5]  & ~new_new_n638__;
  assign new_new_n640__ = ~new_new_n593__ & ~new_new_n639__;
  assign new_new_n641__ = ~\shift[4]  & ~new_new_n640__;
  assign new_new_n642__ = ~new_new_n547__ & ~new_new_n641__;
  assign new_new_n643__ = ~\shift[6]  & ~new_new_n642__;
  assign \result[0]  = ~new_new_n453__ & ~new_new_n643__;
  assign new_new_n645__ = \a[1]  & ~\shift[1] ;
  assign new_new_n646__ = \a[127]  & \shift[1] ;
  assign new_new_n647__ = ~new_new_n645__ & ~new_new_n646__;
  assign new_new_n648__ = ~\shift[0]  & ~new_new_n647__;
  assign new_new_n649__ = \shift[0]  & new_new_n632__;
  assign new_new_n650__ = ~new_new_n648__ & ~new_new_n649__;
  assign new_new_n651__ = ~\shift[3]  & ~new_new_n650__;
  assign new_new_n652__ = \a[121]  & ~\shift[1] ;
  assign new_new_n653__ = \a[119]  & \shift[1] ;
  assign new_new_n654__ = ~new_new_n652__ & ~new_new_n653__;
  assign new_new_n655__ = ~\shift[0]  & ~new_new_n654__;
  assign new_new_n656__ = \shift[0]  & new_new_n622__;
  assign new_new_n657__ = ~new_new_n655__ & ~new_new_n656__;
  assign new_new_n658__ = \shift[3]  & ~new_new_n657__;
  assign new_new_n659__ = ~new_new_n651__ & ~new_new_n658__;
  assign new_new_n660__ = ~\shift[2]  & ~new_new_n659__;
  assign new_new_n661__ = \a[125]  & ~\shift[1] ;
  assign new_new_n662__ = \a[123]  & \shift[1] ;
  assign new_new_n663__ = ~new_new_n661__ & ~new_new_n662__;
  assign new_new_n664__ = ~\shift[0]  & ~new_new_n663__;
  assign new_new_n665__ = \shift[0]  & new_new_n610__;
  assign new_new_n666__ = ~new_new_n664__ & ~new_new_n665__;
  assign new_new_n667__ = ~\shift[3]  & ~new_new_n666__;
  assign new_new_n668__ = \a[117]  & ~\shift[1] ;
  assign new_new_n669__ = \a[115]  & \shift[1] ;
  assign new_new_n670__ = ~new_new_n668__ & ~new_new_n669__;
  assign new_new_n671__ = ~\shift[0]  & ~new_new_n670__;
  assign new_new_n672__ = \shift[0]  & new_new_n600__;
  assign new_new_n673__ = ~new_new_n671__ & ~new_new_n672__;
  assign new_new_n674__ = \shift[3]  & ~new_new_n673__;
  assign new_new_n675__ = ~new_new_n667__ & ~new_new_n674__;
  assign new_new_n676__ = \shift[2]  & ~new_new_n675__;
  assign new_new_n677__ = ~new_new_n660__ & ~new_new_n676__;
  assign new_new_n678__ = ~\shift[5]  & ~new_new_n677__;
  assign new_new_n679__ = \a[97]  & ~\shift[1] ;
  assign new_new_n680__ = \a[95]  & \shift[1] ;
  assign new_new_n681__ = ~new_new_n679__ & ~new_new_n680__;
  assign new_new_n682__ = ~\shift[0]  & ~new_new_n681__;
  assign new_new_n683__ = \shift[0]  & new_new_n586__;
  assign new_new_n684__ = ~new_new_n682__ & ~new_new_n683__;
  assign new_new_n685__ = ~\shift[3]  & ~new_new_n684__;
  assign new_new_n686__ = \a[89]  & ~\shift[1] ;
  assign new_new_n687__ = \a[87]  & \shift[1] ;
  assign new_new_n688__ = ~new_new_n686__ & ~new_new_n687__;
  assign new_new_n689__ = ~\shift[0]  & ~new_new_n688__;
  assign new_new_n690__ = \shift[0]  & new_new_n576__;
  assign new_new_n691__ = ~new_new_n689__ & ~new_new_n690__;
  assign new_new_n692__ = \shift[3]  & ~new_new_n691__;
  assign new_new_n693__ = ~new_new_n685__ & ~new_new_n692__;
  assign new_new_n694__ = ~\shift[2]  & ~new_new_n693__;
  assign new_new_n695__ = \a[93]  & ~\shift[1] ;
  assign new_new_n696__ = \a[91]  & \shift[1] ;
  assign new_new_n697__ = ~new_new_n695__ & ~new_new_n696__;
  assign new_new_n698__ = ~\shift[0]  & ~new_new_n697__;
  assign new_new_n699__ = \shift[0]  & new_new_n564__;
  assign new_new_n700__ = ~new_new_n698__ & ~new_new_n699__;
  assign new_new_n701__ = ~\shift[3]  & ~new_new_n700__;
  assign new_new_n702__ = \a[85]  & ~\shift[1] ;
  assign new_new_n703__ = \a[83]  & \shift[1] ;
  assign new_new_n704__ = ~new_new_n702__ & ~new_new_n703__;
  assign new_new_n705__ = ~\shift[0]  & ~new_new_n704__;
  assign new_new_n706__ = \shift[0]  & new_new_n554__;
  assign new_new_n707__ = ~new_new_n705__ & ~new_new_n706__;
  assign new_new_n708__ = \shift[3]  & ~new_new_n707__;
  assign new_new_n709__ = ~new_new_n701__ & ~new_new_n708__;
  assign new_new_n710__ = \shift[2]  & ~new_new_n709__;
  assign new_new_n711__ = ~new_new_n694__ & ~new_new_n710__;
  assign new_new_n712__ = \shift[5]  & ~new_new_n711__;
  assign new_new_n713__ = ~new_new_n678__ & ~new_new_n712__;
  assign new_new_n714__ = ~\shift[4]  & ~new_new_n713__;
  assign new_new_n715__ = \a[113]  & ~\shift[1] ;
  assign new_new_n716__ = \a[111]  & \shift[1] ;
  assign new_new_n717__ = ~new_new_n715__ & ~new_new_n716__;
  assign new_new_n718__ = ~\shift[0]  & ~new_new_n717__;
  assign new_new_n719__ = \shift[0]  & new_new_n538__;
  assign new_new_n720__ = ~new_new_n718__ & ~new_new_n719__;
  assign new_new_n721__ = ~\shift[3]  & ~new_new_n720__;
  assign new_new_n722__ = \a[105]  & ~\shift[1] ;
  assign new_new_n723__ = \a[103]  & \shift[1] ;
  assign new_new_n724__ = ~new_new_n722__ & ~new_new_n723__;
  assign new_new_n725__ = ~\shift[0]  & ~new_new_n724__;
  assign new_new_n726__ = \shift[0]  & new_new_n528__;
  assign new_new_n727__ = ~new_new_n725__ & ~new_new_n726__;
  assign new_new_n728__ = \shift[3]  & ~new_new_n727__;
  assign new_new_n729__ = ~new_new_n721__ & ~new_new_n728__;
  assign new_new_n730__ = ~\shift[2]  & ~new_new_n729__;
  assign new_new_n731__ = \a[109]  & ~\shift[1] ;
  assign new_new_n732__ = \a[107]  & \shift[1] ;
  assign new_new_n733__ = ~new_new_n731__ & ~new_new_n732__;
  assign new_new_n734__ = ~\shift[0]  & ~new_new_n733__;
  assign new_new_n735__ = \shift[0]  & new_new_n516__;
  assign new_new_n736__ = ~new_new_n734__ & ~new_new_n735__;
  assign new_new_n737__ = ~\shift[3]  & ~new_new_n736__;
  assign new_new_n738__ = \a[101]  & ~\shift[1] ;
  assign new_new_n739__ = \a[99]  & \shift[1] ;
  assign new_new_n740__ = ~new_new_n738__ & ~new_new_n739__;
  assign new_new_n741__ = ~\shift[0]  & ~new_new_n740__;
  assign new_new_n742__ = \shift[0]  & new_new_n506__;
  assign new_new_n743__ = ~new_new_n741__ & ~new_new_n742__;
  assign new_new_n744__ = \shift[3]  & ~new_new_n743__;
  assign new_new_n745__ = ~new_new_n737__ & ~new_new_n744__;
  assign new_new_n746__ = \shift[2]  & ~new_new_n745__;
  assign new_new_n747__ = ~new_new_n730__ & ~new_new_n746__;
  assign new_new_n748__ = ~\shift[5]  & ~new_new_n747__;
  assign new_new_n749__ = \a[81]  & ~\shift[1] ;
  assign new_new_n750__ = \a[79]  & \shift[1] ;
  assign new_new_n751__ = ~new_new_n749__ & ~new_new_n750__;
  assign new_new_n752__ = ~\shift[0]  & ~new_new_n751__;
  assign new_new_n753__ = \shift[0]  & new_new_n492__;
  assign new_new_n754__ = ~new_new_n752__ & ~new_new_n753__;
  assign new_new_n755__ = ~\shift[3]  & ~new_new_n754__;
  assign new_new_n756__ = \a[73]  & ~\shift[1] ;
  assign new_new_n757__ = \a[71]  & \shift[1] ;
  assign new_new_n758__ = ~new_new_n756__ & ~new_new_n757__;
  assign new_new_n759__ = ~\shift[0]  & ~new_new_n758__;
  assign new_new_n760__ = \shift[0]  & new_new_n482__;
  assign new_new_n761__ = ~new_new_n759__ & ~new_new_n760__;
  assign new_new_n762__ = \shift[3]  & ~new_new_n761__;
  assign new_new_n763__ = ~new_new_n755__ & ~new_new_n762__;
  assign new_new_n764__ = ~\shift[2]  & ~new_new_n763__;
  assign new_new_n765__ = \a[77]  & ~\shift[1] ;
  assign new_new_n766__ = \a[75]  & \shift[1] ;
  assign new_new_n767__ = ~new_new_n765__ & ~new_new_n766__;
  assign new_new_n768__ = ~\shift[0]  & ~new_new_n767__;
  assign new_new_n769__ = \shift[0]  & new_new_n470__;
  assign new_new_n770__ = ~new_new_n768__ & ~new_new_n769__;
  assign new_new_n771__ = ~\shift[3]  & ~new_new_n770__;
  assign new_new_n772__ = \a[69]  & ~\shift[1] ;
  assign new_new_n773__ = \a[67]  & \shift[1] ;
  assign new_new_n774__ = ~new_new_n772__ & ~new_new_n773__;
  assign new_new_n775__ = ~\shift[0]  & ~new_new_n774__;
  assign new_new_n776__ = \shift[0]  & new_new_n460__;
  assign new_new_n777__ = ~new_new_n775__ & ~new_new_n776__;
  assign new_new_n778__ = \shift[3]  & ~new_new_n777__;
  assign new_new_n779__ = ~new_new_n771__ & ~new_new_n778__;
  assign new_new_n780__ = \shift[2]  & ~new_new_n779__;
  assign new_new_n781__ = ~new_new_n764__ & ~new_new_n780__;
  assign new_new_n782__ = \shift[5]  & ~new_new_n781__;
  assign new_new_n783__ = ~new_new_n748__ & ~new_new_n782__;
  assign new_new_n784__ = \shift[4]  & ~new_new_n783__;
  assign new_new_n785__ = ~new_new_n714__ & ~new_new_n784__;
  assign new_new_n786__ = ~\shift[6]  & ~new_new_n785__;
  assign new_new_n787__ = \a[49]  & ~\shift[1] ;
  assign new_new_n788__ = \a[47]  & \shift[1] ;
  assign new_new_n789__ = ~new_new_n787__ & ~new_new_n788__;
  assign new_new_n790__ = ~\shift[0]  & ~new_new_n789__;
  assign new_new_n791__ = \shift[0]  & new_new_n312__;
  assign new_new_n792__ = ~new_new_n790__ & ~new_new_n791__;
  assign new_new_n793__ = ~\shift[3]  & ~new_new_n792__;
  assign new_new_n794__ = \shift[0]  & ~new_new_n322__;
  assign new_new_n795__ = \a[41]  & ~\shift[1] ;
  assign new_new_n796__ = \a[39]  & \shift[1] ;
  assign new_new_n797__ = ~new_new_n795__ & ~new_new_n796__;
  assign new_new_n798__ = ~\shift[0]  & ~new_new_n797__;
  assign new_new_n799__ = ~new_new_n794__ & ~new_new_n798__;
  assign new_new_n800__ = \shift[3]  & ~new_new_n799__;
  assign new_new_n801__ = ~new_new_n793__ & ~new_new_n800__;
  assign new_new_n802__ = ~\shift[2]  & ~new_new_n801__;
  assign new_new_n803__ = \a[37]  & ~\shift[1] ;
  assign new_new_n804__ = \a[35]  & \shift[1] ;
  assign new_new_n805__ = ~new_new_n803__ & ~new_new_n804__;
  assign new_new_n806__ = ~\shift[0]  & ~new_new_n805__;
  assign new_new_n807__ = \shift[0]  & new_new_n338__;
  assign new_new_n808__ = ~new_new_n806__ & ~new_new_n807__;
  assign new_new_n809__ = \shift[3]  & ~new_new_n808__;
  assign new_new_n810__ = \shift[0]  & ~new_new_n348__;
  assign new_new_n811__ = \a[45]  & ~\shift[1] ;
  assign new_new_n812__ = \a[43]  & \shift[1] ;
  assign new_new_n813__ = ~new_new_n811__ & ~new_new_n812__;
  assign new_new_n814__ = ~\shift[0]  & ~new_new_n813__;
  assign new_new_n815__ = ~new_new_n810__ & ~new_new_n814__;
  assign new_new_n816__ = ~\shift[3]  & ~new_new_n815__;
  assign new_new_n817__ = ~new_new_n809__ & ~new_new_n816__;
  assign new_new_n818__ = \shift[2]  & ~new_new_n817__;
  assign new_new_n819__ = ~new_new_n802__ & ~new_new_n818__;
  assign new_new_n820__ = ~\shift[5]  & ~new_new_n819__;
  assign new_new_n821__ = \a[17]  & ~\shift[1] ;
  assign new_new_n822__ = \a[15]  & \shift[1] ;
  assign new_new_n823__ = ~new_new_n821__ & ~new_new_n822__;
  assign new_new_n824__ = ~\shift[0]  & ~new_new_n823__;
  assign new_new_n825__ = \shift[0]  & new_new_n302__;
  assign new_new_n826__ = ~new_new_n824__ & ~new_new_n825__;
  assign new_new_n827__ = ~\shift[3]  & ~new_new_n826__;
  assign new_new_n828__ = \a[9]  & ~\shift[1] ;
  assign new_new_n829__ = \a[7]  & \shift[1] ;
  assign new_new_n830__ = ~new_new_n828__ & ~new_new_n829__;
  assign new_new_n831__ = ~\shift[0]  & ~new_new_n830__;
  assign new_new_n832__ = \shift[0]  & new_new_n292__;
  assign new_new_n833__ = ~new_new_n831__ & ~new_new_n832__;
  assign new_new_n834__ = \shift[3]  & ~new_new_n833__;
  assign new_new_n835__ = ~new_new_n827__ & ~new_new_n834__;
  assign new_new_n836__ = ~\shift[2]  & ~new_new_n835__;
  assign new_new_n837__ = \a[13]  & ~\shift[1] ;
  assign new_new_n838__ = \a[11]  & \shift[1] ;
  assign new_new_n839__ = ~new_new_n837__ & ~new_new_n838__;
  assign new_new_n840__ = ~\shift[0]  & ~new_new_n839__;
  assign new_new_n841__ = \shift[0]  & new_new_n280__;
  assign new_new_n842__ = ~new_new_n840__ & ~new_new_n841__;
  assign new_new_n843__ = ~\shift[3]  & ~new_new_n842__;
  assign new_new_n844__ = \a[5]  & ~\shift[1] ;
  assign new_new_n845__ = \a[3]  & \shift[1] ;
  assign new_new_n846__ = ~new_new_n844__ & ~new_new_n845__;
  assign new_new_n847__ = ~\shift[0]  & ~new_new_n846__;
  assign new_new_n848__ = \shift[0]  & new_new_n270__;
  assign new_new_n849__ = ~new_new_n847__ & ~new_new_n848__;
  assign new_new_n850__ = \shift[3]  & ~new_new_n849__;
  assign new_new_n851__ = ~new_new_n843__ & ~new_new_n850__;
  assign new_new_n852__ = \shift[2]  & ~new_new_n851__;
  assign new_new_n853__ = ~new_new_n836__ & ~new_new_n852__;
  assign new_new_n854__ = \shift[5]  & ~new_new_n853__;
  assign new_new_n855__ = ~new_new_n820__ & ~new_new_n854__;
  assign new_new_n856__ = \shift[4]  & ~new_new_n855__;
  assign new_new_n857__ = \a[65]  & ~\shift[1] ;
  assign new_new_n858__ = \a[63]  & \shift[1] ;
  assign new_new_n859__ = ~new_new_n857__ & ~new_new_n858__;
  assign new_new_n860__ = ~\shift[0]  & ~new_new_n859__;
  assign new_new_n861__ = \shift[0]  & new_new_n442__;
  assign new_new_n862__ = ~new_new_n860__ & ~new_new_n861__;
  assign new_new_n863__ = ~\shift[3]  & ~new_new_n862__;
  assign new_new_n864__ = \a[57]  & ~\shift[1] ;
  assign new_new_n865__ = \a[55]  & \shift[1] ;
  assign new_new_n866__ = ~new_new_n864__ & ~new_new_n865__;
  assign new_new_n867__ = ~\shift[0]  & ~new_new_n866__;
  assign new_new_n868__ = \shift[0]  & new_new_n432__;
  assign new_new_n869__ = ~new_new_n867__ & ~new_new_n868__;
  assign new_new_n870__ = \shift[3]  & ~new_new_n869__;
  assign new_new_n871__ = ~new_new_n863__ & ~new_new_n870__;
  assign new_new_n872__ = ~\shift[2]  & ~new_new_n871__;
  assign new_new_n873__ = \a[61]  & ~\shift[1] ;
  assign new_new_n874__ = \a[59]  & \shift[1] ;
  assign new_new_n875__ = ~new_new_n873__ & ~new_new_n874__;
  assign new_new_n876__ = ~\shift[0]  & ~new_new_n875__;
  assign new_new_n877__ = \shift[0]  & new_new_n420__;
  assign new_new_n878__ = ~new_new_n876__ & ~new_new_n877__;
  assign new_new_n879__ = ~\shift[3]  & ~new_new_n878__;
  assign new_new_n880__ = \a[53]  & ~\shift[1] ;
  assign new_new_n881__ = \a[51]  & \shift[1] ;
  assign new_new_n882__ = ~new_new_n880__ & ~new_new_n881__;
  assign new_new_n883__ = ~\shift[0]  & ~new_new_n882__;
  assign new_new_n884__ = \shift[0]  & new_new_n410__;
  assign new_new_n885__ = ~new_new_n883__ & ~new_new_n884__;
  assign new_new_n886__ = \shift[3]  & ~new_new_n885__;
  assign new_new_n887__ = ~new_new_n879__ & ~new_new_n886__;
  assign new_new_n888__ = \shift[2]  & ~new_new_n887__;
  assign new_new_n889__ = ~new_new_n872__ & ~new_new_n888__;
  assign new_new_n890__ = ~\shift[5]  & ~new_new_n889__;
  assign new_new_n891__ = \a[33]  & ~\shift[1] ;
  assign new_new_n892__ = \a[31]  & \shift[1] ;
  assign new_new_n893__ = ~new_new_n891__ & ~new_new_n892__;
  assign new_new_n894__ = ~\shift[0]  & ~new_new_n893__;
  assign new_new_n895__ = \shift[0]  & new_new_n396__;
  assign new_new_n896__ = ~new_new_n894__ & ~new_new_n895__;
  assign new_new_n897__ = ~\shift[3]  & ~new_new_n896__;
  assign new_new_n898__ = \a[25]  & ~\shift[1] ;
  assign new_new_n899__ = \a[23]  & \shift[1] ;
  assign new_new_n900__ = ~new_new_n898__ & ~new_new_n899__;
  assign new_new_n901__ = ~\shift[0]  & ~new_new_n900__;
  assign new_new_n902__ = \shift[0]  & new_new_n386__;
  assign new_new_n903__ = ~new_new_n901__ & ~new_new_n902__;
  assign new_new_n904__ = \shift[3]  & ~new_new_n903__;
  assign new_new_n905__ = ~new_new_n897__ & ~new_new_n904__;
  assign new_new_n906__ = ~\shift[2]  & ~new_new_n905__;
  assign new_new_n907__ = \a[29]  & ~\shift[1] ;
  assign new_new_n908__ = \a[27]  & \shift[1] ;
  assign new_new_n909__ = ~new_new_n907__ & ~new_new_n908__;
  assign new_new_n910__ = ~\shift[0]  & ~new_new_n909__;
  assign new_new_n911__ = \shift[0]  & new_new_n374__;
  assign new_new_n912__ = ~new_new_n910__ & ~new_new_n911__;
  assign new_new_n913__ = ~\shift[3]  & ~new_new_n912__;
  assign new_new_n914__ = \a[21]  & ~\shift[1] ;
  assign new_new_n915__ = \a[19]  & \shift[1] ;
  assign new_new_n916__ = ~new_new_n914__ & ~new_new_n915__;
  assign new_new_n917__ = ~\shift[0]  & ~new_new_n916__;
  assign new_new_n918__ = \shift[0]  & new_new_n364__;
  assign new_new_n919__ = ~new_new_n917__ & ~new_new_n918__;
  assign new_new_n920__ = \shift[3]  & ~new_new_n919__;
  assign new_new_n921__ = ~new_new_n913__ & ~new_new_n920__;
  assign new_new_n922__ = \shift[2]  & ~new_new_n921__;
  assign new_new_n923__ = ~new_new_n906__ & ~new_new_n922__;
  assign new_new_n924__ = \shift[5]  & ~new_new_n923__;
  assign new_new_n925__ = ~new_new_n890__ & ~new_new_n924__;
  assign new_new_n926__ = ~\shift[4]  & ~new_new_n925__;
  assign new_new_n927__ = ~new_new_n856__ & ~new_new_n926__;
  assign new_new_n928__ = \shift[6]  & ~new_new_n927__;
  assign \result[1]  = new_new_n786__ | new_new_n928__;
  assign new_new_n930__ = ~\a[22]  & ~\shift[1] ;
  assign new_new_n931__ = ~\a[20]  & \shift[1] ;
  assign new_new_n932__ = ~new_new_n930__ & ~new_new_n931__;
  assign new_new_n933__ = ~\shift[0]  & ~new_new_n932__;
  assign new_new_n934__ = \shift[0]  & new_new_n916__;
  assign new_new_n935__ = ~new_new_n933__ & ~new_new_n934__;
  assign new_new_n936__ = \shift[3]  & ~new_new_n935__;
  assign new_new_n937__ = ~\a[30]  & ~\shift[1] ;
  assign new_new_n938__ = ~\a[28]  & \shift[1] ;
  assign new_new_n939__ = ~new_new_n937__ & ~new_new_n938__;
  assign new_new_n940__ = ~\shift[0]  & ~new_new_n939__;
  assign new_new_n941__ = \shift[0]  & new_new_n909__;
  assign new_new_n942__ = ~new_new_n940__ & ~new_new_n941__;
  assign new_new_n943__ = ~\shift[3]  & ~new_new_n942__;
  assign new_new_n944__ = ~new_new_n936__ & ~new_new_n943__;
  assign new_new_n945__ = \shift[2]  & ~new_new_n944__;
  assign new_new_n946__ = ~\a[26]  & ~\shift[1] ;
  assign new_new_n947__ = ~\a[24]  & \shift[1] ;
  assign new_new_n948__ = ~new_new_n946__ & ~new_new_n947__;
  assign new_new_n949__ = ~\shift[0]  & ~new_new_n948__;
  assign new_new_n950__ = \shift[0]  & new_new_n900__;
  assign new_new_n951__ = ~new_new_n949__ & ~new_new_n950__;
  assign new_new_n952__ = \shift[3]  & ~new_new_n951__;
  assign new_new_n953__ = ~\a[34]  & ~\shift[1] ;
  assign new_new_n954__ = ~\a[32]  & \shift[1] ;
  assign new_new_n955__ = ~new_new_n953__ & ~new_new_n954__;
  assign new_new_n956__ = ~\shift[0]  & ~new_new_n955__;
  assign new_new_n957__ = \shift[0]  & new_new_n893__;
  assign new_new_n958__ = ~new_new_n956__ & ~new_new_n957__;
  assign new_new_n959__ = ~\shift[3]  & ~new_new_n958__;
  assign new_new_n960__ = ~new_new_n952__ & ~new_new_n959__;
  assign new_new_n961__ = ~\shift[2]  & ~new_new_n960__;
  assign new_new_n962__ = ~new_new_n945__ & ~new_new_n961__;
  assign new_new_n963__ = \shift[5]  & ~new_new_n962__;
  assign new_new_n964__ = ~\a[54]  & ~\shift[1] ;
  assign new_new_n965__ = ~\a[52]  & \shift[1] ;
  assign new_new_n966__ = ~new_new_n964__ & ~new_new_n965__;
  assign new_new_n967__ = ~\shift[0]  & ~new_new_n966__;
  assign new_new_n968__ = \shift[0]  & new_new_n882__;
  assign new_new_n969__ = ~new_new_n967__ & ~new_new_n968__;
  assign new_new_n970__ = \shift[3]  & ~new_new_n969__;
  assign new_new_n971__ = ~\a[62]  & ~\shift[1] ;
  assign new_new_n972__ = ~\a[60]  & \shift[1] ;
  assign new_new_n973__ = ~new_new_n971__ & ~new_new_n972__;
  assign new_new_n974__ = ~\shift[0]  & ~new_new_n973__;
  assign new_new_n975__ = \shift[0]  & new_new_n875__;
  assign new_new_n976__ = ~new_new_n974__ & ~new_new_n975__;
  assign new_new_n977__ = ~\shift[3]  & ~new_new_n976__;
  assign new_new_n978__ = ~new_new_n970__ & ~new_new_n977__;
  assign new_new_n979__ = \shift[2]  & ~new_new_n978__;
  assign new_new_n980__ = ~\a[58]  & ~\shift[1] ;
  assign new_new_n981__ = ~\a[56]  & \shift[1] ;
  assign new_new_n982__ = ~new_new_n980__ & ~new_new_n981__;
  assign new_new_n983__ = ~\shift[0]  & ~new_new_n982__;
  assign new_new_n984__ = \shift[0]  & new_new_n866__;
  assign new_new_n985__ = ~new_new_n983__ & ~new_new_n984__;
  assign new_new_n986__ = \shift[3]  & ~new_new_n985__;
  assign new_new_n987__ = ~\a[66]  & ~\shift[1] ;
  assign new_new_n988__ = ~\a[64]  & \shift[1] ;
  assign new_new_n989__ = ~new_new_n987__ & ~new_new_n988__;
  assign new_new_n990__ = ~\shift[0]  & ~new_new_n989__;
  assign new_new_n991__ = \shift[0]  & new_new_n859__;
  assign new_new_n992__ = ~new_new_n990__ & ~new_new_n991__;
  assign new_new_n993__ = ~\shift[3]  & ~new_new_n992__;
  assign new_new_n994__ = ~new_new_n986__ & ~new_new_n993__;
  assign new_new_n995__ = ~\shift[2]  & ~new_new_n994__;
  assign new_new_n996__ = ~new_new_n979__ & ~new_new_n995__;
  assign new_new_n997__ = ~\shift[5]  & ~new_new_n996__;
  assign new_new_n998__ = ~new_new_n963__ & ~new_new_n997__;
  assign new_new_n999__ = ~\shift[4]  & ~new_new_n998__;
  assign new_new_n1000__ = ~\a[6]  & ~\shift[1] ;
  assign new_new_n1001__ = ~\a[4]  & \shift[1] ;
  assign new_new_n1002__ = ~new_new_n1000__ & ~new_new_n1001__;
  assign new_new_n1003__ = ~\shift[0]  & ~new_new_n1002__;
  assign new_new_n1004__ = \shift[0]  & new_new_n846__;
  assign new_new_n1005__ = ~new_new_n1003__ & ~new_new_n1004__;
  assign new_new_n1006__ = \shift[3]  & ~new_new_n1005__;
  assign new_new_n1007__ = ~\a[14]  & ~\shift[1] ;
  assign new_new_n1008__ = ~\a[12]  & \shift[1] ;
  assign new_new_n1009__ = ~new_new_n1007__ & ~new_new_n1008__;
  assign new_new_n1010__ = ~\shift[0]  & ~new_new_n1009__;
  assign new_new_n1011__ = \shift[0]  & new_new_n839__;
  assign new_new_n1012__ = ~new_new_n1010__ & ~new_new_n1011__;
  assign new_new_n1013__ = ~\shift[3]  & ~new_new_n1012__;
  assign new_new_n1014__ = ~new_new_n1006__ & ~new_new_n1013__;
  assign new_new_n1015__ = \shift[2]  & ~new_new_n1014__;
  assign new_new_n1016__ = ~\a[10]  & ~\shift[1] ;
  assign new_new_n1017__ = ~\a[8]  & \shift[1] ;
  assign new_new_n1018__ = ~new_new_n1016__ & ~new_new_n1017__;
  assign new_new_n1019__ = ~\shift[0]  & ~new_new_n1018__;
  assign new_new_n1020__ = \shift[0]  & new_new_n830__;
  assign new_new_n1021__ = ~new_new_n1019__ & ~new_new_n1020__;
  assign new_new_n1022__ = \shift[3]  & ~new_new_n1021__;
  assign new_new_n1023__ = ~\a[18]  & ~\shift[1] ;
  assign new_new_n1024__ = ~\a[16]  & \shift[1] ;
  assign new_new_n1025__ = ~new_new_n1023__ & ~new_new_n1024__;
  assign new_new_n1026__ = ~\shift[0]  & ~new_new_n1025__;
  assign new_new_n1027__ = \shift[0]  & new_new_n823__;
  assign new_new_n1028__ = ~new_new_n1026__ & ~new_new_n1027__;
  assign new_new_n1029__ = ~\shift[3]  & ~new_new_n1028__;
  assign new_new_n1030__ = ~new_new_n1022__ & ~new_new_n1029__;
  assign new_new_n1031__ = ~\shift[2]  & ~new_new_n1030__;
  assign new_new_n1032__ = ~new_new_n1015__ & ~new_new_n1031__;
  assign new_new_n1033__ = \shift[5]  & ~new_new_n1032__;
  assign new_new_n1034__ = ~\a[38]  & ~\shift[1] ;
  assign new_new_n1035__ = ~\a[36]  & \shift[1] ;
  assign new_new_n1036__ = ~new_new_n1034__ & ~new_new_n1035__;
  assign new_new_n1037__ = ~\shift[0]  & ~new_new_n1036__;
  assign new_new_n1038__ = \shift[0]  & new_new_n805__;
  assign new_new_n1039__ = ~new_new_n1037__ & ~new_new_n1038__;
  assign new_new_n1040__ = \shift[3]  & ~new_new_n1039__;
  assign new_new_n1041__ = \shift[0]  & ~new_new_n813__;
  assign new_new_n1042__ = \a[46]  & ~\shift[1] ;
  assign new_new_n1043__ = \a[44]  & \shift[1] ;
  assign new_new_n1044__ = ~new_new_n1042__ & ~new_new_n1043__;
  assign new_new_n1045__ = ~\shift[0]  & ~new_new_n1044__;
  assign new_new_n1046__ = ~new_new_n1041__ & ~new_new_n1045__;
  assign new_new_n1047__ = ~\shift[3]  & new_new_n1046__;
  assign new_new_n1048__ = ~new_new_n1040__ & ~new_new_n1047__;
  assign new_new_n1049__ = \shift[2]  & ~new_new_n1048__;
  assign new_new_n1050__ = ~\a[42]  & ~\shift[1] ;
  assign new_new_n1051__ = ~\a[40]  & \shift[1] ;
  assign new_new_n1052__ = ~new_new_n1050__ & ~new_new_n1051__;
  assign new_new_n1053__ = ~\shift[0]  & ~new_new_n1052__;
  assign new_new_n1054__ = \shift[0]  & new_new_n797__;
  assign new_new_n1055__ = ~new_new_n1053__ & ~new_new_n1054__;
  assign new_new_n1056__ = \shift[3]  & ~new_new_n1055__;
  assign new_new_n1057__ = ~\a[50]  & ~\shift[1] ;
  assign new_new_n1058__ = ~\a[48]  & \shift[1] ;
  assign new_new_n1059__ = ~new_new_n1057__ & ~new_new_n1058__;
  assign new_new_n1060__ = ~\shift[0]  & ~new_new_n1059__;
  assign new_new_n1061__ = \shift[0]  & new_new_n789__;
  assign new_new_n1062__ = ~new_new_n1060__ & ~new_new_n1061__;
  assign new_new_n1063__ = ~\shift[3]  & ~new_new_n1062__;
  assign new_new_n1064__ = ~new_new_n1056__ & ~new_new_n1063__;
  assign new_new_n1065__ = ~\shift[2]  & ~new_new_n1064__;
  assign new_new_n1066__ = ~new_new_n1049__ & ~new_new_n1065__;
  assign new_new_n1067__ = ~\shift[5]  & ~new_new_n1066__;
  assign new_new_n1068__ = ~new_new_n1033__ & ~new_new_n1067__;
  assign new_new_n1069__ = \shift[4]  & ~new_new_n1068__;
  assign new_new_n1070__ = ~new_new_n999__ & ~new_new_n1069__;
  assign new_new_n1071__ = \shift[6]  & ~new_new_n1070__;
  assign new_new_n1072__ = ~\a[70]  & ~\shift[1] ;
  assign new_new_n1073__ = ~\a[68]  & \shift[1] ;
  assign new_new_n1074__ = ~new_new_n1072__ & ~new_new_n1073__;
  assign new_new_n1075__ = ~\shift[0]  & ~new_new_n1074__;
  assign new_new_n1076__ = \shift[0]  & new_new_n774__;
  assign new_new_n1077__ = ~new_new_n1075__ & ~new_new_n1076__;
  assign new_new_n1078__ = \shift[3]  & ~new_new_n1077__;
  assign new_new_n1079__ = ~\a[78]  & ~\shift[1] ;
  assign new_new_n1080__ = ~\a[76]  & \shift[1] ;
  assign new_new_n1081__ = ~new_new_n1079__ & ~new_new_n1080__;
  assign new_new_n1082__ = ~\shift[0]  & ~new_new_n1081__;
  assign new_new_n1083__ = \shift[0]  & new_new_n767__;
  assign new_new_n1084__ = ~new_new_n1082__ & ~new_new_n1083__;
  assign new_new_n1085__ = ~\shift[3]  & ~new_new_n1084__;
  assign new_new_n1086__ = ~new_new_n1078__ & ~new_new_n1085__;
  assign new_new_n1087__ = \shift[2]  & ~new_new_n1086__;
  assign new_new_n1088__ = ~\a[74]  & ~\shift[1] ;
  assign new_new_n1089__ = ~\a[72]  & \shift[1] ;
  assign new_new_n1090__ = ~new_new_n1088__ & ~new_new_n1089__;
  assign new_new_n1091__ = ~\shift[0]  & ~new_new_n1090__;
  assign new_new_n1092__ = \shift[0]  & new_new_n758__;
  assign new_new_n1093__ = ~new_new_n1091__ & ~new_new_n1092__;
  assign new_new_n1094__ = \shift[3]  & ~new_new_n1093__;
  assign new_new_n1095__ = ~\a[82]  & ~\shift[1] ;
  assign new_new_n1096__ = ~\a[80]  & \shift[1] ;
  assign new_new_n1097__ = ~new_new_n1095__ & ~new_new_n1096__;
  assign new_new_n1098__ = ~\shift[0]  & ~new_new_n1097__;
  assign new_new_n1099__ = \shift[0]  & new_new_n751__;
  assign new_new_n1100__ = ~new_new_n1098__ & ~new_new_n1099__;
  assign new_new_n1101__ = ~\shift[3]  & ~new_new_n1100__;
  assign new_new_n1102__ = ~new_new_n1094__ & ~new_new_n1101__;
  assign new_new_n1103__ = ~\shift[2]  & ~new_new_n1102__;
  assign new_new_n1104__ = ~new_new_n1087__ & ~new_new_n1103__;
  assign new_new_n1105__ = \shift[5]  & ~new_new_n1104__;
  assign new_new_n1106__ = ~\a[102]  & ~\shift[1] ;
  assign new_new_n1107__ = ~\a[100]  & \shift[1] ;
  assign new_new_n1108__ = ~new_new_n1106__ & ~new_new_n1107__;
  assign new_new_n1109__ = ~\shift[0]  & ~new_new_n1108__;
  assign new_new_n1110__ = \shift[0]  & new_new_n740__;
  assign new_new_n1111__ = ~new_new_n1109__ & ~new_new_n1110__;
  assign new_new_n1112__ = \shift[3]  & ~new_new_n1111__;
  assign new_new_n1113__ = ~\a[110]  & ~\shift[1] ;
  assign new_new_n1114__ = ~\a[108]  & \shift[1] ;
  assign new_new_n1115__ = ~new_new_n1113__ & ~new_new_n1114__;
  assign new_new_n1116__ = ~\shift[0]  & ~new_new_n1115__;
  assign new_new_n1117__ = \shift[0]  & new_new_n733__;
  assign new_new_n1118__ = ~new_new_n1116__ & ~new_new_n1117__;
  assign new_new_n1119__ = ~\shift[3]  & ~new_new_n1118__;
  assign new_new_n1120__ = ~new_new_n1112__ & ~new_new_n1119__;
  assign new_new_n1121__ = \shift[2]  & ~new_new_n1120__;
  assign new_new_n1122__ = ~\a[106]  & ~\shift[1] ;
  assign new_new_n1123__ = ~\a[104]  & \shift[1] ;
  assign new_new_n1124__ = ~new_new_n1122__ & ~new_new_n1123__;
  assign new_new_n1125__ = ~\shift[0]  & ~new_new_n1124__;
  assign new_new_n1126__ = \shift[0]  & new_new_n724__;
  assign new_new_n1127__ = ~new_new_n1125__ & ~new_new_n1126__;
  assign new_new_n1128__ = \shift[3]  & ~new_new_n1127__;
  assign new_new_n1129__ = ~\a[114]  & ~\shift[1] ;
  assign new_new_n1130__ = ~\a[112]  & \shift[1] ;
  assign new_new_n1131__ = ~new_new_n1129__ & ~new_new_n1130__;
  assign new_new_n1132__ = ~\shift[0]  & ~new_new_n1131__;
  assign new_new_n1133__ = \shift[0]  & new_new_n717__;
  assign new_new_n1134__ = ~new_new_n1132__ & ~new_new_n1133__;
  assign new_new_n1135__ = ~\shift[3]  & ~new_new_n1134__;
  assign new_new_n1136__ = ~new_new_n1128__ & ~new_new_n1135__;
  assign new_new_n1137__ = ~\shift[2]  & ~new_new_n1136__;
  assign new_new_n1138__ = ~new_new_n1121__ & ~new_new_n1137__;
  assign new_new_n1139__ = ~\shift[5]  & ~new_new_n1138__;
  assign new_new_n1140__ = ~new_new_n1105__ & ~new_new_n1139__;
  assign new_new_n1141__ = \shift[4]  & ~new_new_n1140__;
  assign new_new_n1142__ = ~\a[86]  & ~\shift[1] ;
  assign new_new_n1143__ = ~\a[84]  & \shift[1] ;
  assign new_new_n1144__ = ~new_new_n1142__ & ~new_new_n1143__;
  assign new_new_n1145__ = ~\shift[0]  & ~new_new_n1144__;
  assign new_new_n1146__ = \shift[0]  & new_new_n704__;
  assign new_new_n1147__ = ~new_new_n1145__ & ~new_new_n1146__;
  assign new_new_n1148__ = \shift[3]  & ~new_new_n1147__;
  assign new_new_n1149__ = ~\a[94]  & ~\shift[1] ;
  assign new_new_n1150__ = ~\a[92]  & \shift[1] ;
  assign new_new_n1151__ = ~new_new_n1149__ & ~new_new_n1150__;
  assign new_new_n1152__ = ~\shift[0]  & ~new_new_n1151__;
  assign new_new_n1153__ = \shift[0]  & new_new_n697__;
  assign new_new_n1154__ = ~new_new_n1152__ & ~new_new_n1153__;
  assign new_new_n1155__ = ~\shift[3]  & ~new_new_n1154__;
  assign new_new_n1156__ = ~new_new_n1148__ & ~new_new_n1155__;
  assign new_new_n1157__ = \shift[2]  & ~new_new_n1156__;
  assign new_new_n1158__ = ~\a[90]  & ~\shift[1] ;
  assign new_new_n1159__ = ~\a[88]  & \shift[1] ;
  assign new_new_n1160__ = ~new_new_n1158__ & ~new_new_n1159__;
  assign new_new_n1161__ = ~\shift[0]  & ~new_new_n1160__;
  assign new_new_n1162__ = \shift[0]  & new_new_n688__;
  assign new_new_n1163__ = ~new_new_n1161__ & ~new_new_n1162__;
  assign new_new_n1164__ = \shift[3]  & ~new_new_n1163__;
  assign new_new_n1165__ = ~\a[98]  & ~\shift[1] ;
  assign new_new_n1166__ = ~\a[96]  & \shift[1] ;
  assign new_new_n1167__ = ~new_new_n1165__ & ~new_new_n1166__;
  assign new_new_n1168__ = ~\shift[0]  & ~new_new_n1167__;
  assign new_new_n1169__ = \shift[0]  & new_new_n681__;
  assign new_new_n1170__ = ~new_new_n1168__ & ~new_new_n1169__;
  assign new_new_n1171__ = ~\shift[3]  & ~new_new_n1170__;
  assign new_new_n1172__ = ~new_new_n1164__ & ~new_new_n1171__;
  assign new_new_n1173__ = ~\shift[2]  & ~new_new_n1172__;
  assign new_new_n1174__ = ~new_new_n1157__ & ~new_new_n1173__;
  assign new_new_n1175__ = \shift[5]  & ~new_new_n1174__;
  assign new_new_n1176__ = ~\a[118]  & ~\shift[1] ;
  assign new_new_n1177__ = ~\a[116]  & \shift[1] ;
  assign new_new_n1178__ = ~new_new_n1176__ & ~new_new_n1177__;
  assign new_new_n1179__ = ~\shift[0]  & ~new_new_n1178__;
  assign new_new_n1180__ = \shift[0]  & new_new_n670__;
  assign new_new_n1181__ = ~new_new_n1179__ & ~new_new_n1180__;
  assign new_new_n1182__ = \shift[3]  & ~new_new_n1181__;
  assign new_new_n1183__ = ~\a[126]  & ~\shift[1] ;
  assign new_new_n1184__ = ~\a[124]  & \shift[1] ;
  assign new_new_n1185__ = ~new_new_n1183__ & ~new_new_n1184__;
  assign new_new_n1186__ = ~\shift[0]  & ~new_new_n1185__;
  assign new_new_n1187__ = \shift[0]  & new_new_n663__;
  assign new_new_n1188__ = ~new_new_n1186__ & ~new_new_n1187__;
  assign new_new_n1189__ = ~\shift[3]  & ~new_new_n1188__;
  assign new_new_n1190__ = ~new_new_n1182__ & ~new_new_n1189__;
  assign new_new_n1191__ = \shift[2]  & ~new_new_n1190__;
  assign new_new_n1192__ = ~\a[122]  & ~\shift[1] ;
  assign new_new_n1193__ = ~\a[120]  & \shift[1] ;
  assign new_new_n1194__ = ~new_new_n1192__ & ~new_new_n1193__;
  assign new_new_n1195__ = ~\shift[0]  & ~new_new_n1194__;
  assign new_new_n1196__ = \shift[0]  & new_new_n654__;
  assign new_new_n1197__ = ~new_new_n1195__ & ~new_new_n1196__;
  assign new_new_n1198__ = \shift[3]  & ~new_new_n1197__;
  assign new_new_n1199__ = ~\a[2]  & ~\shift[1] ;
  assign new_new_n1200__ = ~\a[0]  & \shift[1] ;
  assign new_new_n1201__ = ~new_new_n1199__ & ~new_new_n1200__;
  assign new_new_n1202__ = ~\shift[0]  & ~new_new_n1201__;
  assign new_new_n1203__ = \shift[0]  & new_new_n647__;
  assign new_new_n1204__ = ~new_new_n1202__ & ~new_new_n1203__;
  assign new_new_n1205__ = ~\shift[3]  & ~new_new_n1204__;
  assign new_new_n1206__ = ~new_new_n1198__ & ~new_new_n1205__;
  assign new_new_n1207__ = ~\shift[2]  & ~new_new_n1206__;
  assign new_new_n1208__ = ~new_new_n1191__ & ~new_new_n1207__;
  assign new_new_n1209__ = ~\shift[5]  & ~new_new_n1208__;
  assign new_new_n1210__ = ~new_new_n1175__ & ~new_new_n1209__;
  assign new_new_n1211__ = ~\shift[4]  & ~new_new_n1210__;
  assign new_new_n1212__ = ~new_new_n1141__ & ~new_new_n1211__;
  assign new_new_n1213__ = ~\shift[6]  & ~new_new_n1212__;
  assign \result[2]  = ~new_new_n1071__ & ~new_new_n1213__;
  assign new_new_n1215__ = \shift[0]  & ~new_new_n1002__;
  assign new_new_n1216__ = ~\shift[0]  & ~new_new_n288__;
  assign new_new_n1217__ = ~new_new_n1215__ & ~new_new_n1216__;
  assign new_new_n1218__ = \shift[3]  & ~new_new_n1217__;
  assign new_new_n1219__ = \shift[0]  & ~new_new_n1009__;
  assign new_new_n1220__ = ~\shift[0]  & ~new_new_n298__;
  assign new_new_n1221__ = ~new_new_n1219__ & ~new_new_n1220__;
  assign new_new_n1222__ = ~\shift[3]  & ~new_new_n1221__;
  assign new_new_n1223__ = ~new_new_n1218__ & ~new_new_n1222__;
  assign new_new_n1224__ = \shift[2]  & ~new_new_n1223__;
  assign new_new_n1225__ = \shift[0]  & ~new_new_n1018__;
  assign new_new_n1226__ = ~\shift[0]  & ~new_new_n276__;
  assign new_new_n1227__ = ~new_new_n1225__ & ~new_new_n1226__;
  assign new_new_n1228__ = \shift[3]  & ~new_new_n1227__;
  assign new_new_n1229__ = \shift[0]  & ~new_new_n1025__;
  assign new_new_n1230__ = ~\shift[0]  & ~new_new_n360__;
  assign new_new_n1231__ = ~new_new_n1229__ & ~new_new_n1230__;
  assign new_new_n1232__ = ~\shift[3]  & ~new_new_n1231__;
  assign new_new_n1233__ = ~new_new_n1228__ & ~new_new_n1232__;
  assign new_new_n1234__ = ~\shift[2]  & ~new_new_n1233__;
  assign new_new_n1235__ = ~new_new_n1224__ & ~new_new_n1234__;
  assign new_new_n1236__ = \shift[5]  & ~new_new_n1235__;
  assign new_new_n1237__ = \shift[0]  & ~new_new_n1052__;
  assign new_new_n1238__ = ~\shift[0]  & ~new_new_n344__;
  assign new_new_n1239__ = ~new_new_n1237__ & ~new_new_n1238__;
  assign new_new_n1240__ = \shift[3]  & ~new_new_n1239__;
  assign new_new_n1241__ = \shift[0]  & ~new_new_n1059__;
  assign new_new_n1242__ = ~\shift[0]  & ~new_new_n406__;
  assign new_new_n1243__ = ~new_new_n1241__ & ~new_new_n1242__;
  assign new_new_n1244__ = ~\shift[3]  & ~new_new_n1243__;
  assign new_new_n1245__ = ~new_new_n1240__ & ~new_new_n1244__;
  assign new_new_n1246__ = ~\shift[2]  & ~new_new_n1245__;
  assign new_new_n1247__ = \shift[0]  & ~new_new_n1036__;
  assign new_new_n1248__ = ~\shift[0]  & ~new_new_n326__;
  assign new_new_n1249__ = ~new_new_n1247__ & ~new_new_n1248__;
  assign new_new_n1250__ = \shift[3]  & ~new_new_n1249__;
  assign new_new_n1251__ = \shift[0]  & ~new_new_n1044__;
  assign new_new_n1252__ = ~\shift[0]  & ~new_new_n316__;
  assign new_new_n1253__ = ~new_new_n1251__ & ~new_new_n1252__;
  assign new_new_n1254__ = ~\shift[3]  & new_new_n1253__;
  assign new_new_n1255__ = ~new_new_n1250__ & ~new_new_n1254__;
  assign new_new_n1256__ = \shift[2]  & ~new_new_n1255__;
  assign new_new_n1257__ = ~new_new_n1246__ & ~new_new_n1256__;
  assign new_new_n1258__ = ~\shift[5]  & ~new_new_n1257__;
  assign new_new_n1259__ = ~new_new_n1236__ & ~new_new_n1258__;
  assign new_new_n1260__ = \shift[4]  & ~new_new_n1259__;
  assign new_new_n1261__ = \shift[0]  & ~new_new_n932__;
  assign new_new_n1262__ = ~\shift[0]  & ~new_new_n382__;
  assign new_new_n1263__ = ~new_new_n1261__ & ~new_new_n1262__;
  assign new_new_n1264__ = \shift[3]  & ~new_new_n1263__;
  assign new_new_n1265__ = \shift[0]  & ~new_new_n939__;
  assign new_new_n1266__ = ~\shift[0]  & ~new_new_n392__;
  assign new_new_n1267__ = ~new_new_n1265__ & ~new_new_n1266__;
  assign new_new_n1268__ = ~\shift[3]  & ~new_new_n1267__;
  assign new_new_n1269__ = ~new_new_n1264__ & ~new_new_n1268__;
  assign new_new_n1270__ = \shift[2]  & ~new_new_n1269__;
  assign new_new_n1271__ = \shift[0]  & ~new_new_n948__;
  assign new_new_n1272__ = ~\shift[0]  & ~new_new_n370__;
  assign new_new_n1273__ = ~new_new_n1271__ & ~new_new_n1272__;
  assign new_new_n1274__ = \shift[3]  & ~new_new_n1273__;
  assign new_new_n1275__ = \shift[0]  & ~new_new_n955__;
  assign new_new_n1276__ = ~\shift[0]  & ~new_new_n334__;
  assign new_new_n1277__ = ~new_new_n1275__ & ~new_new_n1276__;
  assign new_new_n1278__ = ~\shift[3]  & ~new_new_n1277__;
  assign new_new_n1279__ = ~new_new_n1274__ & ~new_new_n1278__;
  assign new_new_n1280__ = ~\shift[2]  & ~new_new_n1279__;
  assign new_new_n1281__ = ~new_new_n1270__ & ~new_new_n1280__;
  assign new_new_n1282__ = \shift[5]  & ~new_new_n1281__;
  assign new_new_n1283__ = \shift[0]  & ~new_new_n966__;
  assign new_new_n1284__ = ~\shift[0]  & ~new_new_n428__;
  assign new_new_n1285__ = ~new_new_n1283__ & ~new_new_n1284__;
  assign new_new_n1286__ = \shift[3]  & ~new_new_n1285__;
  assign new_new_n1287__ = \shift[0]  & ~new_new_n973__;
  assign new_new_n1288__ = ~\shift[0]  & ~new_new_n438__;
  assign new_new_n1289__ = ~new_new_n1287__ & ~new_new_n1288__;
  assign new_new_n1290__ = ~\shift[3]  & ~new_new_n1289__;
  assign new_new_n1291__ = ~new_new_n1286__ & ~new_new_n1290__;
  assign new_new_n1292__ = \shift[2]  & ~new_new_n1291__;
  assign new_new_n1293__ = \shift[0]  & ~new_new_n982__;
  assign new_new_n1294__ = ~\shift[0]  & ~new_new_n416__;
  assign new_new_n1295__ = ~new_new_n1293__ & ~new_new_n1294__;
  assign new_new_n1296__ = \shift[3]  & ~new_new_n1295__;
  assign new_new_n1297__ = \shift[0]  & ~new_new_n989__;
  assign new_new_n1298__ = ~\shift[0]  & ~new_new_n456__;
  assign new_new_n1299__ = ~new_new_n1297__ & ~new_new_n1298__;
  assign new_new_n1300__ = ~\shift[3]  & ~new_new_n1299__;
  assign new_new_n1301__ = ~new_new_n1296__ & ~new_new_n1300__;
  assign new_new_n1302__ = ~\shift[2]  & ~new_new_n1301__;
  assign new_new_n1303__ = ~new_new_n1292__ & ~new_new_n1302__;
  assign new_new_n1304__ = ~\shift[5]  & ~new_new_n1303__;
  assign new_new_n1305__ = ~new_new_n1282__ & ~new_new_n1304__;
  assign new_new_n1306__ = ~\shift[4]  & ~new_new_n1305__;
  assign new_new_n1307__ = ~new_new_n1260__ & ~new_new_n1306__;
  assign new_new_n1308__ = \shift[6]  & ~new_new_n1307__;
  assign new_new_n1309__ = \shift[0]  & ~new_new_n1144__;
  assign new_new_n1310__ = ~\shift[0]  & ~new_new_n572__;
  assign new_new_n1311__ = ~new_new_n1309__ & ~new_new_n1310__;
  assign new_new_n1312__ = \shift[3]  & ~new_new_n1311__;
  assign new_new_n1313__ = \shift[0]  & ~new_new_n1151__;
  assign new_new_n1314__ = ~\shift[0]  & ~new_new_n582__;
  assign new_new_n1315__ = ~new_new_n1313__ & ~new_new_n1314__;
  assign new_new_n1316__ = ~\shift[3]  & ~new_new_n1315__;
  assign new_new_n1317__ = ~new_new_n1312__ & ~new_new_n1316__;
  assign new_new_n1318__ = \shift[2]  & ~new_new_n1317__;
  assign new_new_n1319__ = \shift[0]  & ~new_new_n1160__;
  assign new_new_n1320__ = ~\shift[0]  & ~new_new_n560__;
  assign new_new_n1321__ = ~new_new_n1319__ & ~new_new_n1320__;
  assign new_new_n1322__ = \shift[3]  & ~new_new_n1321__;
  assign new_new_n1323__ = \shift[0]  & ~new_new_n1167__;
  assign new_new_n1324__ = ~\shift[0]  & ~new_new_n502__;
  assign new_new_n1325__ = ~new_new_n1323__ & ~new_new_n1324__;
  assign new_new_n1326__ = ~\shift[3]  & ~new_new_n1325__;
  assign new_new_n1327__ = ~new_new_n1322__ & ~new_new_n1326__;
  assign new_new_n1328__ = ~\shift[2]  & ~new_new_n1327__;
  assign new_new_n1329__ = ~new_new_n1318__ & ~new_new_n1328__;
  assign new_new_n1330__ = \shift[5]  & ~new_new_n1329__;
  assign new_new_n1331__ = \shift[0]  & ~new_new_n1178__;
  assign new_new_n1332__ = ~\shift[0]  & ~new_new_n618__;
  assign new_new_n1333__ = ~new_new_n1331__ & ~new_new_n1332__;
  assign new_new_n1334__ = \shift[3]  & ~new_new_n1333__;
  assign new_new_n1335__ = \shift[0]  & ~new_new_n1185__;
  assign new_new_n1336__ = ~\shift[0]  & ~new_new_n628__;
  assign new_new_n1337__ = ~new_new_n1335__ & ~new_new_n1336__;
  assign new_new_n1338__ = ~\shift[3]  & ~new_new_n1337__;
  assign new_new_n1339__ = ~new_new_n1334__ & ~new_new_n1338__;
  assign new_new_n1340__ = \shift[2]  & ~new_new_n1339__;
  assign new_new_n1341__ = \shift[0]  & ~new_new_n1194__;
  assign new_new_n1342__ = ~\shift[0]  & ~new_new_n606__;
  assign new_new_n1343__ = ~new_new_n1341__ & ~new_new_n1342__;
  assign new_new_n1344__ = \shift[3]  & ~new_new_n1343__;
  assign new_new_n1345__ = \shift[0]  & ~new_new_n1201__;
  assign new_new_n1346__ = ~\shift[0]  & ~new_new_n266__;
  assign new_new_n1347__ = ~new_new_n1345__ & ~new_new_n1346__;
  assign new_new_n1348__ = ~\shift[3]  & ~new_new_n1347__;
  assign new_new_n1349__ = ~new_new_n1344__ & ~new_new_n1348__;
  assign new_new_n1350__ = ~\shift[2]  & ~new_new_n1349__;
  assign new_new_n1351__ = ~new_new_n1340__ & ~new_new_n1350__;
  assign new_new_n1352__ = ~\shift[5]  & ~new_new_n1351__;
  assign new_new_n1353__ = ~new_new_n1330__ & ~new_new_n1352__;
  assign new_new_n1354__ = ~\shift[4]  & ~new_new_n1353__;
  assign new_new_n1355__ = \shift[0]  & ~new_new_n1074__;
  assign new_new_n1356__ = ~\shift[0]  & ~new_new_n478__;
  assign new_new_n1357__ = ~new_new_n1355__ & ~new_new_n1356__;
  assign new_new_n1358__ = \shift[3]  & ~new_new_n1357__;
  assign new_new_n1359__ = \shift[0]  & ~new_new_n1081__;
  assign new_new_n1360__ = ~\shift[0]  & ~new_new_n488__;
  assign new_new_n1361__ = ~new_new_n1359__ & ~new_new_n1360__;
  assign new_new_n1362__ = ~\shift[3]  & ~new_new_n1361__;
  assign new_new_n1363__ = ~new_new_n1358__ & ~new_new_n1362__;
  assign new_new_n1364__ = \shift[2]  & ~new_new_n1363__;
  assign new_new_n1365__ = \shift[0]  & ~new_new_n1090__;
  assign new_new_n1366__ = ~\shift[0]  & ~new_new_n466__;
  assign new_new_n1367__ = ~new_new_n1365__ & ~new_new_n1366__;
  assign new_new_n1368__ = \shift[3]  & ~new_new_n1367__;
  assign new_new_n1369__ = \shift[0]  & ~new_new_n1097__;
  assign new_new_n1370__ = ~\shift[0]  & ~new_new_n550__;
  assign new_new_n1371__ = ~new_new_n1369__ & ~new_new_n1370__;
  assign new_new_n1372__ = ~\shift[3]  & ~new_new_n1371__;
  assign new_new_n1373__ = ~new_new_n1368__ & ~new_new_n1372__;
  assign new_new_n1374__ = ~\shift[2]  & ~new_new_n1373__;
  assign new_new_n1375__ = ~new_new_n1364__ & ~new_new_n1374__;
  assign new_new_n1376__ = \shift[5]  & ~new_new_n1375__;
  assign new_new_n1377__ = \shift[0]  & ~new_new_n1108__;
  assign new_new_n1378__ = ~\shift[0]  & ~new_new_n524__;
  assign new_new_n1379__ = ~new_new_n1377__ & ~new_new_n1378__;
  assign new_new_n1380__ = \shift[3]  & ~new_new_n1379__;
  assign new_new_n1381__ = \shift[0]  & ~new_new_n1115__;
  assign new_new_n1382__ = ~\shift[0]  & ~new_new_n534__;
  assign new_new_n1383__ = ~new_new_n1381__ & ~new_new_n1382__;
  assign new_new_n1384__ = ~\shift[3]  & ~new_new_n1383__;
  assign new_new_n1385__ = ~new_new_n1380__ & ~new_new_n1384__;
  assign new_new_n1386__ = \shift[2]  & ~new_new_n1385__;
  assign new_new_n1387__ = \shift[0]  & ~new_new_n1124__;
  assign new_new_n1388__ = ~\shift[0]  & ~new_new_n512__;
  assign new_new_n1389__ = ~new_new_n1387__ & ~new_new_n1388__;
  assign new_new_n1390__ = \shift[3]  & ~new_new_n1389__;
  assign new_new_n1391__ = \shift[0]  & ~new_new_n1131__;
  assign new_new_n1392__ = ~\shift[0]  & ~new_new_n596__;
  assign new_new_n1393__ = ~new_new_n1391__ & ~new_new_n1392__;
  assign new_new_n1394__ = ~\shift[3]  & ~new_new_n1393__;
  assign new_new_n1395__ = ~new_new_n1390__ & ~new_new_n1394__;
  assign new_new_n1396__ = ~\shift[2]  & ~new_new_n1395__;
  assign new_new_n1397__ = ~new_new_n1386__ & ~new_new_n1396__;
  assign new_new_n1398__ = ~\shift[5]  & ~new_new_n1397__;
  assign new_new_n1399__ = ~new_new_n1376__ & ~new_new_n1398__;
  assign new_new_n1400__ = \shift[4]  & ~new_new_n1399__;
  assign new_new_n1401__ = ~new_new_n1354__ & ~new_new_n1400__;
  assign new_new_n1402__ = ~\shift[6]  & ~new_new_n1401__;
  assign \result[3]  = ~new_new_n1308__ & ~new_new_n1402__;
  assign new_new_n1404__ = ~\shift[3]  & ~new_new_n366__;
  assign new_new_n1405__ = \shift[3]  & ~new_new_n282__;
  assign new_new_n1406__ = ~new_new_n1404__ & ~new_new_n1405__;
  assign new_new_n1407__ = ~\shift[2]  & ~new_new_n1406__;
  assign new_new_n1408__ = \shift[2]  & ~new_new_n306__;
  assign new_new_n1409__ = ~new_new_n1407__ & ~new_new_n1408__;
  assign new_new_n1410__ = \shift[5]  & ~new_new_n1409__;
  assign new_new_n1411__ = \shift[2]  & ~new_new_n330__;
  assign new_new_n1412__ = \shift[3]  & ~new_new_n350__;
  assign new_new_n1413__ = ~\shift[3]  & ~new_new_n412__;
  assign new_new_n1414__ = ~new_new_n1412__ & ~new_new_n1413__;
  assign new_new_n1415__ = ~\shift[2]  & ~new_new_n1414__;
  assign new_new_n1416__ = ~new_new_n1411__ & ~new_new_n1415__;
  assign new_new_n1417__ = ~\shift[5]  & ~new_new_n1416__;
  assign new_new_n1418__ = ~new_new_n1410__ & ~new_new_n1417__;
  assign new_new_n1419__ = \shift[4]  & ~new_new_n1418__;
  assign new_new_n1420__ = ~\shift[3]  & ~new_new_n340__;
  assign new_new_n1421__ = \shift[3]  & ~new_new_n376__;
  assign new_new_n1422__ = ~new_new_n1420__ & ~new_new_n1421__;
  assign new_new_n1423__ = ~\shift[2]  & ~new_new_n1422__;
  assign new_new_n1424__ = \shift[2]  & ~new_new_n400__;
  assign new_new_n1425__ = ~new_new_n1423__ & ~new_new_n1424__;
  assign new_new_n1426__ = \shift[5]  & ~new_new_n1425__;
  assign new_new_n1427__ = ~\shift[3]  & ~new_new_n462__;
  assign new_new_n1428__ = \shift[3]  & ~new_new_n422__;
  assign new_new_n1429__ = ~new_new_n1427__ & ~new_new_n1428__;
  assign new_new_n1430__ = ~\shift[2]  & ~new_new_n1429__;
  assign new_new_n1431__ = \shift[2]  & ~new_new_n446__;
  assign new_new_n1432__ = ~new_new_n1430__ & ~new_new_n1431__;
  assign new_new_n1433__ = ~\shift[5]  & ~new_new_n1432__;
  assign new_new_n1434__ = ~new_new_n1426__ & ~new_new_n1433__;
  assign new_new_n1435__ = ~\shift[4]  & ~new_new_n1434__;
  assign new_new_n1436__ = ~new_new_n1419__ & ~new_new_n1435__;
  assign new_new_n1437__ = \shift[6]  & ~new_new_n1436__;
  assign new_new_n1438__ = ~\shift[3]  & ~new_new_n556__;
  assign new_new_n1439__ = \shift[3]  & ~new_new_n472__;
  assign new_new_n1440__ = ~new_new_n1438__ & ~new_new_n1439__;
  assign new_new_n1441__ = ~\shift[2]  & ~new_new_n1440__;
  assign new_new_n1442__ = \shift[2]  & ~new_new_n496__;
  assign new_new_n1443__ = ~new_new_n1441__ & ~new_new_n1442__;
  assign new_new_n1444__ = \shift[5]  & ~new_new_n1443__;
  assign new_new_n1445__ = \shift[3]  & ~new_new_n518__;
  assign new_new_n1446__ = ~\shift[3]  & ~new_new_n602__;
  assign new_new_n1447__ = ~new_new_n1445__ & ~new_new_n1446__;
  assign new_new_n1448__ = ~\shift[2]  & ~new_new_n1447__;
  assign new_new_n1449__ = \shift[2]  & ~new_new_n542__;
  assign new_new_n1450__ = ~new_new_n1448__ & ~new_new_n1449__;
  assign new_new_n1451__ = ~\shift[5]  & ~new_new_n1450__;
  assign new_new_n1452__ = ~new_new_n1444__ & ~new_new_n1451__;
  assign new_new_n1453__ = \shift[4]  & ~new_new_n1452__;
  assign new_new_n1454__ = ~\shift[3]  & ~new_new_n508__;
  assign new_new_n1455__ = \shift[3]  & ~new_new_n566__;
  assign new_new_n1456__ = ~new_new_n1454__ & ~new_new_n1455__;
  assign new_new_n1457__ = ~\shift[2]  & ~new_new_n1456__;
  assign new_new_n1458__ = \shift[2]  & ~new_new_n590__;
  assign new_new_n1459__ = ~new_new_n1457__ & ~new_new_n1458__;
  assign new_new_n1460__ = \shift[5]  & ~new_new_n1459__;
  assign new_new_n1461__ = \shift[3]  & ~new_new_n612__;
  assign new_new_n1462__ = ~\shift[3]  & ~new_new_n272__;
  assign new_new_n1463__ = ~new_new_n1461__ & ~new_new_n1462__;
  assign new_new_n1464__ = ~\shift[2]  & ~new_new_n1463__;
  assign new_new_n1465__ = \shift[2]  & ~new_new_n636__;
  assign new_new_n1466__ = ~new_new_n1464__ & ~new_new_n1465__;
  assign new_new_n1467__ = ~\shift[5]  & ~new_new_n1466__;
  assign new_new_n1468__ = ~new_new_n1460__ & ~new_new_n1467__;
  assign new_new_n1469__ = ~\shift[4]  & ~new_new_n1468__;
  assign new_new_n1470__ = ~new_new_n1453__ & ~new_new_n1469__;
  assign new_new_n1471__ = ~\shift[6]  & ~new_new_n1470__;
  assign \result[4]  = ~new_new_n1437__ & ~new_new_n1471__;
  assign new_new_n1473__ = \shift[2]  & ~new_new_n659__;
  assign new_new_n1474__ = ~\shift[3]  & ~new_new_n849__;
  assign new_new_n1475__ = \shift[3]  & ~new_new_n666__;
  assign new_new_n1476__ = ~new_new_n1474__ & ~new_new_n1475__;
  assign new_new_n1477__ = ~\shift[2]  & ~new_new_n1476__;
  assign new_new_n1478__ = ~new_new_n1473__ & ~new_new_n1477__;
  assign new_new_n1479__ = ~\shift[5]  & ~new_new_n1478__;
  assign new_new_n1480__ = \shift[2]  & ~new_new_n693__;
  assign new_new_n1481__ = ~\shift[3]  & ~new_new_n743__;
  assign new_new_n1482__ = \shift[3]  & ~new_new_n700__;
  assign new_new_n1483__ = ~new_new_n1481__ & ~new_new_n1482__;
  assign new_new_n1484__ = ~\shift[2]  & ~new_new_n1483__;
  assign new_new_n1485__ = ~new_new_n1480__ & ~new_new_n1484__;
  assign new_new_n1486__ = \shift[5]  & ~new_new_n1485__;
  assign new_new_n1487__ = ~new_new_n1479__ & ~new_new_n1486__;
  assign new_new_n1488__ = ~\shift[4]  & ~new_new_n1487__;
  assign new_new_n1489__ = \shift[2]  & ~new_new_n729__;
  assign new_new_n1490__ = ~\shift[3]  & ~new_new_n673__;
  assign new_new_n1491__ = \shift[3]  & ~new_new_n736__;
  assign new_new_n1492__ = ~new_new_n1490__ & ~new_new_n1491__;
  assign new_new_n1493__ = ~\shift[2]  & ~new_new_n1492__;
  assign new_new_n1494__ = ~new_new_n1489__ & ~new_new_n1493__;
  assign new_new_n1495__ = ~\shift[5]  & ~new_new_n1494__;
  assign new_new_n1496__ = \shift[2]  & ~new_new_n763__;
  assign new_new_n1497__ = ~\shift[3]  & ~new_new_n707__;
  assign new_new_n1498__ = \shift[3]  & ~new_new_n770__;
  assign new_new_n1499__ = ~new_new_n1497__ & ~new_new_n1498__;
  assign new_new_n1500__ = ~\shift[2]  & ~new_new_n1499__;
  assign new_new_n1501__ = ~new_new_n1496__ & ~new_new_n1500__;
  assign new_new_n1502__ = \shift[5]  & ~new_new_n1501__;
  assign new_new_n1503__ = ~new_new_n1495__ & ~new_new_n1502__;
  assign new_new_n1504__ = \shift[4]  & ~new_new_n1503__;
  assign new_new_n1505__ = ~new_new_n1488__ & ~new_new_n1504__;
  assign new_new_n1506__ = ~\shift[6]  & ~new_new_n1505__;
  assign new_new_n1507__ = \shift[2]  & ~new_new_n871__;
  assign new_new_n1508__ = ~\shift[3]  & ~new_new_n777__;
  assign new_new_n1509__ = \shift[3]  & ~new_new_n878__;
  assign new_new_n1510__ = ~new_new_n1508__ & ~new_new_n1509__;
  assign new_new_n1511__ = ~\shift[2]  & ~new_new_n1510__;
  assign new_new_n1512__ = ~new_new_n1507__ & ~new_new_n1511__;
  assign new_new_n1513__ = ~\shift[5]  & ~new_new_n1512__;
  assign new_new_n1514__ = \shift[2]  & ~new_new_n905__;
  assign new_new_n1515__ = ~\shift[3]  & ~new_new_n808__;
  assign new_new_n1516__ = \shift[3]  & ~new_new_n912__;
  assign new_new_n1517__ = ~new_new_n1515__ & ~new_new_n1516__;
  assign new_new_n1518__ = ~\shift[2]  & ~new_new_n1517__;
  assign new_new_n1519__ = ~new_new_n1514__ & ~new_new_n1518__;
  assign new_new_n1520__ = \shift[5]  & ~new_new_n1519__;
  assign new_new_n1521__ = ~new_new_n1513__ & ~new_new_n1520__;
  assign new_new_n1522__ = ~\shift[4]  & ~new_new_n1521__;
  assign new_new_n1523__ = ~\shift[3]  & ~new_new_n885__;
  assign new_new_n1524__ = \shift[3]  & ~new_new_n815__;
  assign new_new_n1525__ = ~new_new_n1523__ & ~new_new_n1524__;
  assign new_new_n1526__ = ~\shift[2]  & ~new_new_n1525__;
  assign new_new_n1527__ = \shift[2]  & ~new_new_n801__;
  assign new_new_n1528__ = ~new_new_n1526__ & ~new_new_n1527__;
  assign new_new_n1529__ = ~\shift[5]  & ~new_new_n1528__;
  assign new_new_n1530__ = \shift[2]  & ~new_new_n835__;
  assign new_new_n1531__ = ~\shift[3]  & ~new_new_n919__;
  assign new_new_n1532__ = \shift[3]  & ~new_new_n842__;
  assign new_new_n1533__ = ~new_new_n1531__ & ~new_new_n1532__;
  assign new_new_n1534__ = ~\shift[2]  & ~new_new_n1533__;
  assign new_new_n1535__ = ~new_new_n1530__ & ~new_new_n1534__;
  assign new_new_n1536__ = \shift[5]  & ~new_new_n1535__;
  assign new_new_n1537__ = ~new_new_n1529__ & ~new_new_n1536__;
  assign new_new_n1538__ = \shift[4]  & ~new_new_n1537__;
  assign new_new_n1539__ = ~new_new_n1522__ & ~new_new_n1538__;
  assign new_new_n1540__ = \shift[6]  & ~new_new_n1539__;
  assign \result[5]  = new_new_n1506__ | new_new_n1540__;
  assign new_new_n1542__ = ~\shift[3]  & ~new_new_n935__;
  assign new_new_n1543__ = \shift[3]  & ~new_new_n1012__;
  assign new_new_n1544__ = ~new_new_n1542__ & ~new_new_n1543__;
  assign new_new_n1545__ = ~\shift[2]  & ~new_new_n1544__;
  assign new_new_n1546__ = \shift[2]  & ~new_new_n1030__;
  assign new_new_n1547__ = ~new_new_n1545__ & ~new_new_n1546__;
  assign new_new_n1548__ = \shift[5]  & ~new_new_n1547__;
  assign new_new_n1549__ = ~\shift[3]  & ~new_new_n969__;
  assign new_new_n1550__ = \shift[3]  & new_new_n1046__;
  assign new_new_n1551__ = ~new_new_n1549__ & ~new_new_n1550__;
  assign new_new_n1552__ = ~\shift[2]  & ~new_new_n1551__;
  assign new_new_n1553__ = \shift[2]  & ~new_new_n1064__;
  assign new_new_n1554__ = ~new_new_n1552__ & ~new_new_n1553__;
  assign new_new_n1555__ = ~\shift[5]  & ~new_new_n1554__;
  assign new_new_n1556__ = ~new_new_n1548__ & ~new_new_n1555__;
  assign new_new_n1557__ = \shift[4]  & ~new_new_n1556__;
  assign new_new_n1558__ = \shift[3]  & ~new_new_n942__;
  assign new_new_n1559__ = ~\shift[3]  & ~new_new_n1039__;
  assign new_new_n1560__ = ~new_new_n1558__ & ~new_new_n1559__;
  assign new_new_n1561__ = ~\shift[2]  & ~new_new_n1560__;
  assign new_new_n1562__ = \shift[2]  & ~new_new_n960__;
  assign new_new_n1563__ = ~new_new_n1561__ & ~new_new_n1562__;
  assign new_new_n1564__ = \shift[5]  & ~new_new_n1563__;
  assign new_new_n1565__ = ~\shift[3]  & ~new_new_n1077__;
  assign new_new_n1566__ = \shift[3]  & ~new_new_n976__;
  assign new_new_n1567__ = ~new_new_n1565__ & ~new_new_n1566__;
  assign new_new_n1568__ = ~\shift[2]  & ~new_new_n1567__;
  assign new_new_n1569__ = \shift[2]  & ~new_new_n994__;
  assign new_new_n1570__ = ~new_new_n1568__ & ~new_new_n1569__;
  assign new_new_n1571__ = ~\shift[5]  & ~new_new_n1570__;
  assign new_new_n1572__ = ~new_new_n1564__ & ~new_new_n1571__;
  assign new_new_n1573__ = ~\shift[4]  & ~new_new_n1572__;
  assign new_new_n1574__ = ~new_new_n1557__ & ~new_new_n1573__;
  assign new_new_n1575__ = \shift[6]  & ~new_new_n1574__;
  assign new_new_n1576__ = ~\shift[3]  & ~new_new_n1147__;
  assign new_new_n1577__ = \shift[3]  & ~new_new_n1084__;
  assign new_new_n1578__ = ~new_new_n1576__ & ~new_new_n1577__;
  assign new_new_n1579__ = ~\shift[2]  & ~new_new_n1578__;
  assign new_new_n1580__ = \shift[2]  & ~new_new_n1102__;
  assign new_new_n1581__ = ~new_new_n1579__ & ~new_new_n1580__;
  assign new_new_n1582__ = \shift[5]  & ~new_new_n1581__;
  assign new_new_n1583__ = \shift[3]  & ~new_new_n1118__;
  assign new_new_n1584__ = ~\shift[3]  & ~new_new_n1181__;
  assign new_new_n1585__ = ~new_new_n1583__ & ~new_new_n1584__;
  assign new_new_n1586__ = ~\shift[2]  & ~new_new_n1585__;
  assign new_new_n1587__ = \shift[2]  & ~new_new_n1136__;
  assign new_new_n1588__ = ~new_new_n1586__ & ~new_new_n1587__;
  assign new_new_n1589__ = ~\shift[5]  & ~new_new_n1588__;
  assign new_new_n1590__ = ~new_new_n1582__ & ~new_new_n1589__;
  assign new_new_n1591__ = \shift[4]  & ~new_new_n1590__;
  assign new_new_n1592__ = ~\shift[3]  & ~new_new_n1111__;
  assign new_new_n1593__ = \shift[3]  & ~new_new_n1154__;
  assign new_new_n1594__ = ~new_new_n1592__ & ~new_new_n1593__;
  assign new_new_n1595__ = ~\shift[2]  & ~new_new_n1594__;
  assign new_new_n1596__ = \shift[2]  & ~new_new_n1172__;
  assign new_new_n1597__ = ~new_new_n1595__ & ~new_new_n1596__;
  assign new_new_n1598__ = \shift[5]  & ~new_new_n1597__;
  assign new_new_n1599__ = \shift[3]  & ~new_new_n1188__;
  assign new_new_n1600__ = ~\shift[3]  & ~new_new_n1005__;
  assign new_new_n1601__ = ~new_new_n1599__ & ~new_new_n1600__;
  assign new_new_n1602__ = ~\shift[2]  & ~new_new_n1601__;
  assign new_new_n1603__ = \shift[2]  & ~new_new_n1206__;
  assign new_new_n1604__ = ~new_new_n1602__ & ~new_new_n1603__;
  assign new_new_n1605__ = ~\shift[5]  & ~new_new_n1604__;
  assign new_new_n1606__ = ~new_new_n1598__ & ~new_new_n1605__;
  assign new_new_n1607__ = ~\shift[4]  & ~new_new_n1606__;
  assign new_new_n1608__ = ~new_new_n1591__ & ~new_new_n1607__;
  assign new_new_n1609__ = ~\shift[6]  & ~new_new_n1608__;
  assign \result[6]  = ~new_new_n1575__ & ~new_new_n1609__;
  assign new_new_n1611__ = \shift[3]  & ~new_new_n1221__;
  assign new_new_n1612__ = ~\shift[3]  & ~new_new_n1263__;
  assign new_new_n1613__ = ~new_new_n1611__ & ~new_new_n1612__;
  assign new_new_n1614__ = ~\shift[2]  & ~new_new_n1613__;
  assign new_new_n1615__ = \shift[2]  & ~new_new_n1233__;
  assign new_new_n1616__ = ~new_new_n1614__ & ~new_new_n1615__;
  assign new_new_n1617__ = \shift[5]  & ~new_new_n1616__;
  assign new_new_n1618__ = \shift[2]  & ~new_new_n1245__;
  assign new_new_n1619__ = ~\shift[3]  & new_new_n1285__;
  assign new_new_n1620__ = \shift[3]  & ~new_new_n1253__;
  assign new_new_n1621__ = ~new_new_n1619__ & ~new_new_n1620__;
  assign new_new_n1622__ = ~\shift[2]  & new_new_n1621__;
  assign new_new_n1623__ = ~new_new_n1618__ & ~new_new_n1622__;
  assign new_new_n1624__ = ~\shift[5]  & ~new_new_n1623__;
  assign new_new_n1625__ = ~new_new_n1617__ & ~new_new_n1624__;
  assign new_new_n1626__ = \shift[4]  & ~new_new_n1625__;
  assign new_new_n1627__ = \shift[3]  & ~new_new_n1267__;
  assign new_new_n1628__ = ~\shift[3]  & ~new_new_n1249__;
  assign new_new_n1629__ = ~new_new_n1627__ & ~new_new_n1628__;
  assign new_new_n1630__ = ~\shift[2]  & ~new_new_n1629__;
  assign new_new_n1631__ = \shift[2]  & ~new_new_n1279__;
  assign new_new_n1632__ = ~new_new_n1630__ & ~new_new_n1631__;
  assign new_new_n1633__ = \shift[5]  & ~new_new_n1632__;
  assign new_new_n1634__ = \shift[3]  & ~new_new_n1289__;
  assign new_new_n1635__ = ~\shift[3]  & ~new_new_n1357__;
  assign new_new_n1636__ = ~new_new_n1634__ & ~new_new_n1635__;
  assign new_new_n1637__ = ~\shift[2]  & ~new_new_n1636__;
  assign new_new_n1638__ = \shift[2]  & ~new_new_n1301__;
  assign new_new_n1639__ = ~new_new_n1637__ & ~new_new_n1638__;
  assign new_new_n1640__ = ~\shift[5]  & ~new_new_n1639__;
  assign new_new_n1641__ = ~new_new_n1633__ & ~new_new_n1640__;
  assign new_new_n1642__ = ~\shift[4]  & ~new_new_n1641__;
  assign new_new_n1643__ = ~new_new_n1626__ & ~new_new_n1642__;
  assign new_new_n1644__ = \shift[6]  & ~new_new_n1643__;
  assign new_new_n1645__ = \shift[3]  & ~new_new_n1361__;
  assign new_new_n1646__ = ~\shift[3]  & ~new_new_n1311__;
  assign new_new_n1647__ = ~new_new_n1645__ & ~new_new_n1646__;
  assign new_new_n1648__ = ~\shift[2]  & ~new_new_n1647__;
  assign new_new_n1649__ = \shift[2]  & ~new_new_n1373__;
  assign new_new_n1650__ = ~new_new_n1648__ & ~new_new_n1649__;
  assign new_new_n1651__ = \shift[5]  & ~new_new_n1650__;
  assign new_new_n1652__ = \shift[3]  & ~new_new_n1383__;
  assign new_new_n1653__ = ~\shift[3]  & ~new_new_n1333__;
  assign new_new_n1654__ = ~new_new_n1652__ & ~new_new_n1653__;
  assign new_new_n1655__ = ~\shift[2]  & ~new_new_n1654__;
  assign new_new_n1656__ = \shift[2]  & ~new_new_n1395__;
  assign new_new_n1657__ = ~new_new_n1655__ & ~new_new_n1656__;
  assign new_new_n1658__ = ~\shift[5]  & ~new_new_n1657__;
  assign new_new_n1659__ = ~new_new_n1651__ & ~new_new_n1658__;
  assign new_new_n1660__ = \shift[4]  & ~new_new_n1659__;
  assign new_new_n1661__ = \shift[3]  & ~new_new_n1315__;
  assign new_new_n1662__ = ~\shift[3]  & ~new_new_n1379__;
  assign new_new_n1663__ = ~new_new_n1661__ & ~new_new_n1662__;
  assign new_new_n1664__ = ~\shift[2]  & ~new_new_n1663__;
  assign new_new_n1665__ = \shift[2]  & ~new_new_n1327__;
  assign new_new_n1666__ = ~new_new_n1664__ & ~new_new_n1665__;
  assign new_new_n1667__ = \shift[5]  & ~new_new_n1666__;
  assign new_new_n1668__ = \shift[3]  & ~new_new_n1337__;
  assign new_new_n1669__ = ~\shift[3]  & ~new_new_n1217__;
  assign new_new_n1670__ = ~new_new_n1668__ & ~new_new_n1669__;
  assign new_new_n1671__ = ~\shift[2]  & ~new_new_n1670__;
  assign new_new_n1672__ = \shift[2]  & ~new_new_n1349__;
  assign new_new_n1673__ = ~new_new_n1671__ & ~new_new_n1672__;
  assign new_new_n1674__ = ~\shift[5]  & ~new_new_n1673__;
  assign new_new_n1675__ = ~new_new_n1667__ & ~new_new_n1674__;
  assign new_new_n1676__ = ~\shift[4]  & ~new_new_n1675__;
  assign new_new_n1677__ = ~new_new_n1660__ & ~new_new_n1676__;
  assign new_new_n1678__ = ~\shift[6]  & ~new_new_n1677__;
  assign \result[7]  = ~new_new_n1644__ & ~new_new_n1678__;
  assign new_new_n1680__ = \shift[2]  & ~new_new_n1406__;
  assign new_new_n1681__ = \shift[3]  & ~new_new_n304__;
  assign new_new_n1682__ = ~\shift[3]  & ~new_new_n388__;
  assign new_new_n1683__ = ~new_new_n1681__ & ~new_new_n1682__;
  assign new_new_n1684__ = ~\shift[2]  & ~new_new_n1683__;
  assign new_new_n1685__ = ~new_new_n1680__ & ~new_new_n1684__;
  assign new_new_n1686__ = \shift[5]  & ~new_new_n1685__;
  assign new_new_n1687__ = \shift[2]  & ~new_new_n1414__;
  assign new_new_n1688__ = ~\shift[3]  & new_new_n434__;
  assign new_new_n1689__ = \shift[3]  & ~new_new_n318__;
  assign new_new_n1690__ = ~new_new_n1688__ & ~new_new_n1689__;
  assign new_new_n1691__ = ~\shift[2]  & new_new_n1690__;
  assign new_new_n1692__ = ~new_new_n1687__ & ~new_new_n1691__;
  assign new_new_n1693__ = ~\shift[5]  & ~new_new_n1692__;
  assign new_new_n1694__ = ~new_new_n1686__ & ~new_new_n1693__;
  assign new_new_n1695__ = \shift[4]  & ~new_new_n1694__;
  assign new_new_n1696__ = \shift[2]  & ~new_new_n1422__;
  assign new_new_n1697__ = ~\shift[3]  & ~new_new_n328__;
  assign new_new_n1698__ = \shift[3]  & ~new_new_n398__;
  assign new_new_n1699__ = ~new_new_n1697__ & ~new_new_n1698__;
  assign new_new_n1700__ = ~\shift[2]  & ~new_new_n1699__;
  assign new_new_n1701__ = ~new_new_n1696__ & ~new_new_n1700__;
  assign new_new_n1702__ = \shift[5]  & ~new_new_n1701__;
  assign new_new_n1703__ = \shift[2]  & ~new_new_n1429__;
  assign new_new_n1704__ = \shift[3]  & ~new_new_n444__;
  assign new_new_n1705__ = ~\shift[3]  & ~new_new_n484__;
  assign new_new_n1706__ = ~new_new_n1704__ & ~new_new_n1705__;
  assign new_new_n1707__ = ~\shift[2]  & ~new_new_n1706__;
  assign new_new_n1708__ = ~new_new_n1703__ & ~new_new_n1707__;
  assign new_new_n1709__ = ~\shift[5]  & ~new_new_n1708__;
  assign new_new_n1710__ = ~new_new_n1702__ & ~new_new_n1709__;
  assign new_new_n1711__ = ~\shift[4]  & ~new_new_n1710__;
  assign new_new_n1712__ = ~new_new_n1695__ & ~new_new_n1711__;
  assign new_new_n1713__ = \shift[6]  & ~new_new_n1712__;
  assign new_new_n1714__ = \shift[2]  & ~new_new_n1440__;
  assign new_new_n1715__ = \shift[3]  & ~new_new_n494__;
  assign new_new_n1716__ = ~\shift[3]  & ~new_new_n578__;
  assign new_new_n1717__ = ~new_new_n1715__ & ~new_new_n1716__;
  assign new_new_n1718__ = ~\shift[2]  & ~new_new_n1717__;
  assign new_new_n1719__ = ~new_new_n1714__ & ~new_new_n1718__;
  assign new_new_n1720__ = \shift[5]  & ~new_new_n1719__;
  assign new_new_n1721__ = \shift[2]  & ~new_new_n1447__;
  assign new_new_n1722__ = \shift[3]  & ~new_new_n540__;
  assign new_new_n1723__ = ~\shift[3]  & ~new_new_n624__;
  assign new_new_n1724__ = ~new_new_n1722__ & ~new_new_n1723__;
  assign new_new_n1725__ = ~\shift[2]  & ~new_new_n1724__;
  assign new_new_n1726__ = ~new_new_n1721__ & ~new_new_n1725__;
  assign new_new_n1727__ = ~\shift[5]  & ~new_new_n1726__;
  assign new_new_n1728__ = ~new_new_n1720__ & ~new_new_n1727__;
  assign new_new_n1729__ = \shift[4]  & ~new_new_n1728__;
  assign new_new_n1730__ = \shift[2]  & ~new_new_n1456__;
  assign new_new_n1731__ = \shift[3]  & ~new_new_n588__;
  assign new_new_n1732__ = ~\shift[3]  & ~new_new_n530__;
  assign new_new_n1733__ = ~new_new_n1731__ & ~new_new_n1732__;
  assign new_new_n1734__ = ~\shift[2]  & ~new_new_n1733__;
  assign new_new_n1735__ = ~new_new_n1730__ & ~new_new_n1734__;
  assign new_new_n1736__ = \shift[5]  & ~new_new_n1735__;
  assign new_new_n1737__ = \shift[2]  & ~new_new_n1463__;
  assign new_new_n1738__ = \shift[3]  & ~new_new_n634__;
  assign new_new_n1739__ = ~\shift[3]  & ~new_new_n294__;
  assign new_new_n1740__ = ~new_new_n1738__ & ~new_new_n1739__;
  assign new_new_n1741__ = ~\shift[2]  & ~new_new_n1740__;
  assign new_new_n1742__ = ~new_new_n1737__ & ~new_new_n1741__;
  assign new_new_n1743__ = ~\shift[5]  & ~new_new_n1742__;
  assign new_new_n1744__ = ~new_new_n1736__ & ~new_new_n1743__;
  assign new_new_n1745__ = ~\shift[4]  & ~new_new_n1744__;
  assign new_new_n1746__ = ~new_new_n1729__ & ~new_new_n1745__;
  assign new_new_n1747__ = ~\shift[6]  & ~new_new_n1746__;
  assign \result[8]  = ~new_new_n1713__ & ~new_new_n1747__;
  assign new_new_n1749__ = \shift[2]  & ~new_new_n1476__;
  assign new_new_n1750__ = ~\shift[3]  & ~new_new_n833__;
  assign new_new_n1751__ = \shift[3]  & ~new_new_n650__;
  assign new_new_n1752__ = ~new_new_n1750__ & ~new_new_n1751__;
  assign new_new_n1753__ = ~\shift[2]  & ~new_new_n1752__;
  assign new_new_n1754__ = ~new_new_n1749__ & ~new_new_n1753__;
  assign new_new_n1755__ = ~\shift[5]  & ~new_new_n1754__;
  assign new_new_n1756__ = ~\shift[3]  & ~new_new_n727__;
  assign new_new_n1757__ = \shift[3]  & ~new_new_n684__;
  assign new_new_n1758__ = ~new_new_n1756__ & ~new_new_n1757__;
  assign new_new_n1759__ = ~\shift[2]  & ~new_new_n1758__;
  assign new_new_n1760__ = \shift[2]  & ~new_new_n1483__;
  assign new_new_n1761__ = ~new_new_n1759__ & ~new_new_n1760__;
  assign new_new_n1762__ = \shift[5]  & ~new_new_n1761__;
  assign new_new_n1763__ = ~new_new_n1755__ & ~new_new_n1762__;
  assign new_new_n1764__ = ~\shift[4]  & ~new_new_n1763__;
  assign new_new_n1765__ = \shift[2]  & ~new_new_n1492__;
  assign new_new_n1766__ = ~\shift[3]  & ~new_new_n657__;
  assign new_new_n1767__ = \shift[3]  & ~new_new_n720__;
  assign new_new_n1768__ = ~new_new_n1766__ & ~new_new_n1767__;
  assign new_new_n1769__ = ~\shift[2]  & ~new_new_n1768__;
  assign new_new_n1770__ = ~new_new_n1765__ & ~new_new_n1769__;
  assign new_new_n1771__ = ~\shift[5]  & ~new_new_n1770__;
  assign new_new_n1772__ = ~\shift[3]  & ~new_new_n691__;
  assign new_new_n1773__ = \shift[3]  & ~new_new_n754__;
  assign new_new_n1774__ = ~new_new_n1772__ & ~new_new_n1773__;
  assign new_new_n1775__ = ~\shift[2]  & ~new_new_n1774__;
  assign new_new_n1776__ = \shift[2]  & ~new_new_n1499__;
  assign new_new_n1777__ = ~new_new_n1775__ & ~new_new_n1776__;
  assign new_new_n1778__ = \shift[5]  & ~new_new_n1777__;
  assign new_new_n1779__ = ~new_new_n1771__ & ~new_new_n1778__;
  assign new_new_n1780__ = \shift[4]  & ~new_new_n1779__;
  assign new_new_n1781__ = ~new_new_n1764__ & ~new_new_n1780__;
  assign new_new_n1782__ = ~\shift[6]  & ~new_new_n1781__;
  assign new_new_n1783__ = ~\shift[3]  & ~new_new_n761__;
  assign new_new_n1784__ = \shift[3]  & ~new_new_n862__;
  assign new_new_n1785__ = ~new_new_n1783__ & ~new_new_n1784__;
  assign new_new_n1786__ = ~\shift[2]  & ~new_new_n1785__;
  assign new_new_n1787__ = \shift[2]  & ~new_new_n1510__;
  assign new_new_n1788__ = ~new_new_n1786__ & ~new_new_n1787__;
  assign new_new_n1789__ = ~\shift[5]  & ~new_new_n1788__;
  assign new_new_n1790__ = \shift[3]  & ~new_new_n896__;
  assign new_new_n1791__ = ~\shift[3]  & ~new_new_n799__;
  assign new_new_n1792__ = ~new_new_n1790__ & ~new_new_n1791__;
  assign new_new_n1793__ = ~\shift[2]  & ~new_new_n1792__;
  assign new_new_n1794__ = \shift[2]  & ~new_new_n1517__;
  assign new_new_n1795__ = ~new_new_n1793__ & ~new_new_n1794__;
  assign new_new_n1796__ = \shift[5]  & ~new_new_n1795__;
  assign new_new_n1797__ = ~new_new_n1789__ & ~new_new_n1796__;
  assign new_new_n1798__ = ~\shift[4]  & ~new_new_n1797__;
  assign new_new_n1799__ = ~\shift[3]  & ~new_new_n869__;
  assign new_new_n1800__ = \shift[3]  & ~new_new_n792__;
  assign new_new_n1801__ = ~new_new_n1799__ & ~new_new_n1800__;
  assign new_new_n1802__ = ~\shift[2]  & ~new_new_n1801__;
  assign new_new_n1803__ = \shift[2]  & ~new_new_n1525__;
  assign new_new_n1804__ = ~new_new_n1802__ & ~new_new_n1803__;
  assign new_new_n1805__ = ~\shift[5]  & ~new_new_n1804__;
  assign new_new_n1806__ = ~\shift[3]  & ~new_new_n903__;
  assign new_new_n1807__ = \shift[3]  & ~new_new_n826__;
  assign new_new_n1808__ = ~new_new_n1806__ & ~new_new_n1807__;
  assign new_new_n1809__ = ~\shift[2]  & ~new_new_n1808__;
  assign new_new_n1810__ = \shift[2]  & ~new_new_n1533__;
  assign new_new_n1811__ = ~new_new_n1809__ & ~new_new_n1810__;
  assign new_new_n1812__ = \shift[5]  & ~new_new_n1811__;
  assign new_new_n1813__ = ~new_new_n1805__ & ~new_new_n1812__;
  assign new_new_n1814__ = \shift[4]  & ~new_new_n1813__;
  assign new_new_n1815__ = ~new_new_n1798__ & ~new_new_n1814__;
  assign new_new_n1816__ = \shift[6]  & ~new_new_n1815__;
  assign \result[9]  = new_new_n1782__ | new_new_n1816__;
  assign new_new_n1818__ = \shift[2]  & ~new_new_n1544__;
  assign new_new_n1819__ = \shift[3]  & ~new_new_n1028__;
  assign new_new_n1820__ = ~\shift[3]  & ~new_new_n951__;
  assign new_new_n1821__ = ~new_new_n1819__ & ~new_new_n1820__;
  assign new_new_n1822__ = ~\shift[2]  & ~new_new_n1821__;
  assign new_new_n1823__ = ~new_new_n1818__ & ~new_new_n1822__;
  assign new_new_n1824__ = \shift[5]  & ~new_new_n1823__;
  assign new_new_n1825__ = \shift[2]  & ~new_new_n1551__;
  assign new_new_n1826__ = \shift[3]  & ~new_new_n1062__;
  assign new_new_n1827__ = ~\shift[3]  & ~new_new_n985__;
  assign new_new_n1828__ = ~new_new_n1826__ & ~new_new_n1827__;
  assign new_new_n1829__ = ~\shift[2]  & ~new_new_n1828__;
  assign new_new_n1830__ = ~new_new_n1825__ & ~new_new_n1829__;
  assign new_new_n1831__ = ~\shift[5]  & ~new_new_n1830__;
  assign new_new_n1832__ = ~new_new_n1824__ & ~new_new_n1831__;
  assign new_new_n1833__ = \shift[4]  & ~new_new_n1832__;
  assign new_new_n1834__ = \shift[2]  & ~new_new_n1560__;
  assign new_new_n1835__ = \shift[3]  & ~new_new_n958__;
  assign new_new_n1836__ = ~\shift[3]  & ~new_new_n1055__;
  assign new_new_n1837__ = ~new_new_n1835__ & ~new_new_n1836__;
  assign new_new_n1838__ = ~\shift[2]  & ~new_new_n1837__;
  assign new_new_n1839__ = ~new_new_n1834__ & ~new_new_n1838__;
  assign new_new_n1840__ = \shift[5]  & ~new_new_n1839__;
  assign new_new_n1841__ = \shift[2]  & ~new_new_n1567__;
  assign new_new_n1842__ = \shift[3]  & ~new_new_n992__;
  assign new_new_n1843__ = ~\shift[3]  & ~new_new_n1093__;
  assign new_new_n1844__ = ~new_new_n1842__ & ~new_new_n1843__;
  assign new_new_n1845__ = ~\shift[2]  & ~new_new_n1844__;
  assign new_new_n1846__ = ~new_new_n1841__ & ~new_new_n1845__;
  assign new_new_n1847__ = ~\shift[5]  & ~new_new_n1846__;
  assign new_new_n1848__ = ~new_new_n1840__ & ~new_new_n1847__;
  assign new_new_n1849__ = ~\shift[4]  & ~new_new_n1848__;
  assign new_new_n1850__ = ~new_new_n1833__ & ~new_new_n1849__;
  assign new_new_n1851__ = \shift[6]  & ~new_new_n1850__;
  assign new_new_n1852__ = \shift[2]  & ~new_new_n1578__;
  assign new_new_n1853__ = \shift[3]  & ~new_new_n1100__;
  assign new_new_n1854__ = ~\shift[3]  & ~new_new_n1163__;
  assign new_new_n1855__ = ~new_new_n1853__ & ~new_new_n1854__;
  assign new_new_n1856__ = ~\shift[2]  & ~new_new_n1855__;
  assign new_new_n1857__ = ~new_new_n1852__ & ~new_new_n1856__;
  assign new_new_n1858__ = \shift[5]  & ~new_new_n1857__;
  assign new_new_n1859__ = \shift[2]  & ~new_new_n1585__;
  assign new_new_n1860__ = \shift[3]  & ~new_new_n1134__;
  assign new_new_n1861__ = ~\shift[3]  & ~new_new_n1197__;
  assign new_new_n1862__ = ~new_new_n1860__ & ~new_new_n1861__;
  assign new_new_n1863__ = ~\shift[2]  & ~new_new_n1862__;
  assign new_new_n1864__ = ~new_new_n1859__ & ~new_new_n1863__;
  assign new_new_n1865__ = ~\shift[5]  & ~new_new_n1864__;
  assign new_new_n1866__ = ~new_new_n1858__ & ~new_new_n1865__;
  assign new_new_n1867__ = \shift[4]  & ~new_new_n1866__;
  assign new_new_n1868__ = \shift[2]  & ~new_new_n1594__;
  assign new_new_n1869__ = \shift[3]  & ~new_new_n1170__;
  assign new_new_n1870__ = ~\shift[3]  & ~new_new_n1127__;
  assign new_new_n1871__ = ~new_new_n1869__ & ~new_new_n1870__;
  assign new_new_n1872__ = ~\shift[2]  & ~new_new_n1871__;
  assign new_new_n1873__ = ~new_new_n1868__ & ~new_new_n1872__;
  assign new_new_n1874__ = \shift[5]  & ~new_new_n1873__;
  assign new_new_n1875__ = \shift[2]  & ~new_new_n1601__;
  assign new_new_n1876__ = \shift[3]  & ~new_new_n1204__;
  assign new_new_n1877__ = ~\shift[3]  & ~new_new_n1021__;
  assign new_new_n1878__ = ~new_new_n1876__ & ~new_new_n1877__;
  assign new_new_n1879__ = ~\shift[2]  & ~new_new_n1878__;
  assign new_new_n1880__ = ~new_new_n1875__ & ~new_new_n1879__;
  assign new_new_n1881__ = ~\shift[5]  & ~new_new_n1880__;
  assign new_new_n1882__ = ~new_new_n1874__ & ~new_new_n1881__;
  assign new_new_n1883__ = ~\shift[4]  & ~new_new_n1882__;
  assign new_new_n1884__ = ~new_new_n1867__ & ~new_new_n1883__;
  assign new_new_n1885__ = ~\shift[6]  & ~new_new_n1884__;
  assign \result[10]  = ~new_new_n1851__ & ~new_new_n1885__;
  assign new_new_n1887__ = \shift[2]  & ~new_new_n1613__;
  assign new_new_n1888__ = \shift[3]  & ~new_new_n1231__;
  assign new_new_n1889__ = ~\shift[3]  & ~new_new_n1273__;
  assign new_new_n1890__ = ~new_new_n1888__ & ~new_new_n1889__;
  assign new_new_n1891__ = ~\shift[2]  & ~new_new_n1890__;
  assign new_new_n1892__ = ~new_new_n1887__ & ~new_new_n1891__;
  assign new_new_n1893__ = \shift[5]  & ~new_new_n1892__;
  assign new_new_n1894__ = \shift[3]  & ~new_new_n1243__;
  assign new_new_n1895__ = ~\shift[3]  & ~new_new_n1295__;
  assign new_new_n1896__ = ~new_new_n1894__ & ~new_new_n1895__;
  assign new_new_n1897__ = ~\shift[2]  & ~new_new_n1896__;
  assign new_new_n1898__ = \shift[2]  & new_new_n1621__;
  assign new_new_n1899__ = ~new_new_n1897__ & ~new_new_n1898__;
  assign new_new_n1900__ = ~\shift[5]  & ~new_new_n1899__;
  assign new_new_n1901__ = ~new_new_n1893__ & ~new_new_n1900__;
  assign new_new_n1902__ = \shift[4]  & ~new_new_n1901__;
  assign new_new_n1903__ = \shift[3]  & ~new_new_n1277__;
  assign new_new_n1904__ = ~\shift[3]  & ~new_new_n1239__;
  assign new_new_n1905__ = ~new_new_n1903__ & ~new_new_n1904__;
  assign new_new_n1906__ = ~\shift[2]  & ~new_new_n1905__;
  assign new_new_n1907__ = \shift[2]  & ~new_new_n1629__;
  assign new_new_n1908__ = ~new_new_n1906__ & ~new_new_n1907__;
  assign new_new_n1909__ = \shift[5]  & ~new_new_n1908__;
  assign new_new_n1910__ = \shift[2]  & ~new_new_n1636__;
  assign new_new_n1911__ = \shift[3]  & ~new_new_n1299__;
  assign new_new_n1912__ = ~\shift[3]  & ~new_new_n1367__;
  assign new_new_n1913__ = ~new_new_n1911__ & ~new_new_n1912__;
  assign new_new_n1914__ = ~\shift[2]  & ~new_new_n1913__;
  assign new_new_n1915__ = ~new_new_n1910__ & ~new_new_n1914__;
  assign new_new_n1916__ = ~\shift[5]  & ~new_new_n1915__;
  assign new_new_n1917__ = ~new_new_n1909__ & ~new_new_n1916__;
  assign new_new_n1918__ = ~\shift[4]  & ~new_new_n1917__;
  assign new_new_n1919__ = ~new_new_n1902__ & ~new_new_n1918__;
  assign new_new_n1920__ = \shift[6]  & ~new_new_n1919__;
  assign new_new_n1921__ = \shift[3]  & ~new_new_n1371__;
  assign new_new_n1922__ = ~\shift[3]  & ~new_new_n1321__;
  assign new_new_n1923__ = ~new_new_n1921__ & ~new_new_n1922__;
  assign new_new_n1924__ = ~\shift[2]  & ~new_new_n1923__;
  assign new_new_n1925__ = \shift[2]  & ~new_new_n1647__;
  assign new_new_n1926__ = ~new_new_n1924__ & ~new_new_n1925__;
  assign new_new_n1927__ = \shift[5]  & ~new_new_n1926__;
  assign new_new_n1928__ = \shift[2]  & ~new_new_n1654__;
  assign new_new_n1929__ = \shift[3]  & ~new_new_n1393__;
  assign new_new_n1930__ = ~\shift[3]  & ~new_new_n1343__;
  assign new_new_n1931__ = ~new_new_n1929__ & ~new_new_n1930__;
  assign new_new_n1932__ = ~\shift[2]  & ~new_new_n1931__;
  assign new_new_n1933__ = ~new_new_n1928__ & ~new_new_n1932__;
  assign new_new_n1934__ = ~\shift[5]  & ~new_new_n1933__;
  assign new_new_n1935__ = ~new_new_n1927__ & ~new_new_n1934__;
  assign new_new_n1936__ = \shift[4]  & ~new_new_n1935__;
  assign new_new_n1937__ = \shift[3]  & ~new_new_n1325__;
  assign new_new_n1938__ = ~\shift[3]  & ~new_new_n1389__;
  assign new_new_n1939__ = ~new_new_n1937__ & ~new_new_n1938__;
  assign new_new_n1940__ = ~\shift[2]  & ~new_new_n1939__;
  assign new_new_n1941__ = \shift[2]  & ~new_new_n1663__;
  assign new_new_n1942__ = ~new_new_n1940__ & ~new_new_n1941__;
  assign new_new_n1943__ = \shift[5]  & ~new_new_n1942__;
  assign new_new_n1944__ = \shift[3]  & ~new_new_n1347__;
  assign new_new_n1945__ = ~\shift[3]  & ~new_new_n1227__;
  assign new_new_n1946__ = ~new_new_n1944__ & ~new_new_n1945__;
  assign new_new_n1947__ = ~\shift[2]  & ~new_new_n1946__;
  assign new_new_n1948__ = \shift[2]  & ~new_new_n1670__;
  assign new_new_n1949__ = ~new_new_n1947__ & ~new_new_n1948__;
  assign new_new_n1950__ = ~\shift[5]  & ~new_new_n1949__;
  assign new_new_n1951__ = ~new_new_n1943__ & ~new_new_n1950__;
  assign new_new_n1952__ = ~\shift[4]  & ~new_new_n1951__;
  assign new_new_n1953__ = ~new_new_n1936__ & ~new_new_n1952__;
  assign new_new_n1954__ = ~\shift[6]  & ~new_new_n1953__;
  assign \result[11]  = ~new_new_n1920__ & ~new_new_n1954__;
  assign new_new_n1956__ = \shift[2]  & ~new_new_n1683__;
  assign new_new_n1957__ = ~\shift[2]  & ~new_new_n378__;
  assign new_new_n1958__ = ~new_new_n1956__ & ~new_new_n1957__;
  assign new_new_n1959__ = \shift[5]  & ~new_new_n1958__;
  assign new_new_n1960__ = ~\shift[2]  & ~new_new_n424__;
  assign new_new_n1961__ = \shift[2]  & new_new_n1690__;
  assign new_new_n1962__ = ~new_new_n1960__ & ~new_new_n1961__;
  assign new_new_n1963__ = ~\shift[5]  & ~new_new_n1962__;
  assign new_new_n1964__ = ~new_new_n1959__ & ~new_new_n1963__;
  assign new_new_n1965__ = \shift[4]  & ~new_new_n1964__;
  assign new_new_n1966__ = ~\shift[2]  & ~new_new_n352__;
  assign new_new_n1967__ = \shift[2]  & ~new_new_n1699__;
  assign new_new_n1968__ = ~new_new_n1966__ & ~new_new_n1967__;
  assign new_new_n1969__ = \shift[5]  & ~new_new_n1968__;
  assign new_new_n1970__ = \shift[2]  & ~new_new_n1706__;
  assign new_new_n1971__ = ~\shift[2]  & ~new_new_n474__;
  assign new_new_n1972__ = ~new_new_n1970__ & ~new_new_n1971__;
  assign new_new_n1973__ = ~\shift[5]  & ~new_new_n1972__;
  assign new_new_n1974__ = ~new_new_n1969__ & ~new_new_n1973__;
  assign new_new_n1975__ = ~\shift[4]  & ~new_new_n1974__;
  assign new_new_n1976__ = ~new_new_n1965__ & ~new_new_n1975__;
  assign new_new_n1977__ = \shift[6]  & ~new_new_n1976__;
  assign new_new_n1978__ = \shift[2]  & ~new_new_n1717__;
  assign new_new_n1979__ = ~\shift[2]  & ~new_new_n568__;
  assign new_new_n1980__ = ~new_new_n1978__ & ~new_new_n1979__;
  assign new_new_n1981__ = \shift[5]  & ~new_new_n1980__;
  assign new_new_n1982__ = \shift[2]  & ~new_new_n1724__;
  assign new_new_n1983__ = ~\shift[2]  & ~new_new_n614__;
  assign new_new_n1984__ = ~new_new_n1982__ & ~new_new_n1983__;
  assign new_new_n1985__ = ~\shift[5]  & ~new_new_n1984__;
  assign new_new_n1986__ = ~new_new_n1981__ & ~new_new_n1985__;
  assign new_new_n1987__ = \shift[4]  & ~new_new_n1986__;
  assign new_new_n1988__ = \shift[2]  & ~new_new_n1733__;
  assign new_new_n1989__ = ~\shift[2]  & ~new_new_n520__;
  assign new_new_n1990__ = ~new_new_n1988__ & ~new_new_n1989__;
  assign new_new_n1991__ = \shift[5]  & ~new_new_n1990__;
  assign new_new_n1992__ = \shift[2]  & ~new_new_n1740__;
  assign new_new_n1993__ = ~\shift[2]  & ~new_new_n284__;
  assign new_new_n1994__ = ~new_new_n1992__ & ~new_new_n1993__;
  assign new_new_n1995__ = ~\shift[5]  & ~new_new_n1994__;
  assign new_new_n1996__ = ~new_new_n1991__ & ~new_new_n1995__;
  assign new_new_n1997__ = ~\shift[4]  & ~new_new_n1996__;
  assign new_new_n1998__ = ~new_new_n1987__ & ~new_new_n1997__;
  assign new_new_n1999__ = ~\shift[6]  & ~new_new_n1998__;
  assign \result[12]  = ~new_new_n1977__ & ~new_new_n1999__;
  assign new_new_n2001__ = ~\shift[2]  & ~new_new_n851__;
  assign new_new_n2002__ = \shift[2]  & ~new_new_n1752__;
  assign new_new_n2003__ = ~new_new_n2001__ & ~new_new_n2002__;
  assign new_new_n2004__ = ~\shift[5]  & ~new_new_n2003__;
  assign new_new_n2005__ = \shift[2]  & ~new_new_n1758__;
  assign new_new_n2006__ = ~\shift[2]  & ~new_new_n745__;
  assign new_new_n2007__ = ~new_new_n2005__ & ~new_new_n2006__;
  assign new_new_n2008__ = \shift[5]  & ~new_new_n2007__;
  assign new_new_n2009__ = ~new_new_n2004__ & ~new_new_n2008__;
  assign new_new_n2010__ = ~\shift[4]  & ~new_new_n2009__;
  assign new_new_n2011__ = ~\shift[2]  & ~new_new_n675__;
  assign new_new_n2012__ = \shift[2]  & ~new_new_n1768__;
  assign new_new_n2013__ = ~new_new_n2011__ & ~new_new_n2012__;
  assign new_new_n2014__ = ~\shift[5]  & ~new_new_n2013__;
  assign new_new_n2015__ = \shift[2]  & ~new_new_n1774__;
  assign new_new_n2016__ = ~\shift[2]  & ~new_new_n709__;
  assign new_new_n2017__ = ~new_new_n2015__ & ~new_new_n2016__;
  assign new_new_n2018__ = \shift[5]  & ~new_new_n2017__;
  assign new_new_n2019__ = ~new_new_n2014__ & ~new_new_n2018__;
  assign new_new_n2020__ = \shift[4]  & ~new_new_n2019__;
  assign new_new_n2021__ = ~new_new_n2010__ & ~new_new_n2020__;
  assign new_new_n2022__ = ~\shift[6]  & ~new_new_n2021__;
  assign new_new_n2023__ = \shift[2]  & ~new_new_n1785__;
  assign new_new_n2024__ = ~\shift[2]  & ~new_new_n779__;
  assign new_new_n2025__ = ~new_new_n2023__ & ~new_new_n2024__;
  assign new_new_n2026__ = ~\shift[5]  & ~new_new_n2025__;
  assign new_new_n2027__ = ~\shift[2]  & ~new_new_n817__;
  assign new_new_n2028__ = \shift[2]  & ~new_new_n1792__;
  assign new_new_n2029__ = ~new_new_n2027__ & ~new_new_n2028__;
  assign new_new_n2030__ = \shift[5]  & ~new_new_n2029__;
  assign new_new_n2031__ = ~new_new_n2026__ & ~new_new_n2030__;
  assign new_new_n2032__ = ~\shift[4]  & ~new_new_n2031__;
  assign new_new_n2033__ = ~\shift[2]  & ~new_new_n887__;
  assign new_new_n2034__ = \shift[2]  & ~new_new_n1801__;
  assign new_new_n2035__ = ~new_new_n2033__ & ~new_new_n2034__;
  assign new_new_n2036__ = ~\shift[5]  & ~new_new_n2035__;
  assign new_new_n2037__ = \shift[2]  & ~new_new_n1808__;
  assign new_new_n2038__ = ~\shift[2]  & ~new_new_n921__;
  assign new_new_n2039__ = ~new_new_n2037__ & ~new_new_n2038__;
  assign new_new_n2040__ = \shift[5]  & ~new_new_n2039__;
  assign new_new_n2041__ = ~new_new_n2036__ & ~new_new_n2040__;
  assign new_new_n2042__ = \shift[4]  & ~new_new_n2041__;
  assign new_new_n2043__ = ~new_new_n2032__ & ~new_new_n2042__;
  assign new_new_n2044__ = \shift[6]  & ~new_new_n2043__;
  assign \result[13]  = new_new_n2022__ | new_new_n2044__;
  assign new_new_n2046__ = \shift[2]  & ~new_new_n1821__;
  assign new_new_n2047__ = ~\shift[2]  & ~new_new_n944__;
  assign new_new_n2048__ = ~new_new_n2046__ & ~new_new_n2047__;
  assign new_new_n2049__ = \shift[5]  & ~new_new_n2048__;
  assign new_new_n2050__ = \shift[2]  & ~new_new_n1828__;
  assign new_new_n2051__ = ~\shift[2]  & ~new_new_n978__;
  assign new_new_n2052__ = ~new_new_n2050__ & ~new_new_n2051__;
  assign new_new_n2053__ = ~\shift[5]  & ~new_new_n2052__;
  assign new_new_n2054__ = ~new_new_n2049__ & ~new_new_n2053__;
  assign new_new_n2055__ = \shift[4]  & ~new_new_n2054__;
  assign new_new_n2056__ = \shift[2]  & ~new_new_n1837__;
  assign new_new_n2057__ = ~\shift[2]  & ~new_new_n1048__;
  assign new_new_n2058__ = ~new_new_n2056__ & ~new_new_n2057__;
  assign new_new_n2059__ = \shift[5]  & ~new_new_n2058__;
  assign new_new_n2060__ = \shift[2]  & ~new_new_n1844__;
  assign new_new_n2061__ = ~\shift[2]  & ~new_new_n1086__;
  assign new_new_n2062__ = ~new_new_n2060__ & ~new_new_n2061__;
  assign new_new_n2063__ = ~\shift[5]  & ~new_new_n2062__;
  assign new_new_n2064__ = ~new_new_n2059__ & ~new_new_n2063__;
  assign new_new_n2065__ = ~\shift[4]  & ~new_new_n2064__;
  assign new_new_n2066__ = ~new_new_n2055__ & ~new_new_n2065__;
  assign new_new_n2067__ = \shift[6]  & ~new_new_n2066__;
  assign new_new_n2068__ = \shift[2]  & ~new_new_n1855__;
  assign new_new_n2069__ = ~\shift[2]  & ~new_new_n1156__;
  assign new_new_n2070__ = ~new_new_n2068__ & ~new_new_n2069__;
  assign new_new_n2071__ = \shift[5]  & ~new_new_n2070__;
  assign new_new_n2072__ = \shift[2]  & ~new_new_n1862__;
  assign new_new_n2073__ = ~\shift[2]  & ~new_new_n1190__;
  assign new_new_n2074__ = ~new_new_n2072__ & ~new_new_n2073__;
  assign new_new_n2075__ = ~\shift[5]  & ~new_new_n2074__;
  assign new_new_n2076__ = ~new_new_n2071__ & ~new_new_n2075__;
  assign new_new_n2077__ = \shift[4]  & ~new_new_n2076__;
  assign new_new_n2078__ = \shift[2]  & ~new_new_n1871__;
  assign new_new_n2079__ = ~\shift[2]  & ~new_new_n1120__;
  assign new_new_n2080__ = ~new_new_n2078__ & ~new_new_n2079__;
  assign new_new_n2081__ = \shift[5]  & ~new_new_n2080__;
  assign new_new_n2082__ = \shift[2]  & ~new_new_n1878__;
  assign new_new_n2083__ = ~\shift[2]  & ~new_new_n1014__;
  assign new_new_n2084__ = ~new_new_n2082__ & ~new_new_n2083__;
  assign new_new_n2085__ = ~\shift[5]  & ~new_new_n2084__;
  assign new_new_n2086__ = ~new_new_n2081__ & ~new_new_n2085__;
  assign new_new_n2087__ = ~\shift[4]  & ~new_new_n2086__;
  assign new_new_n2088__ = ~new_new_n2077__ & ~new_new_n2087__;
  assign new_new_n2089__ = ~\shift[6]  & ~new_new_n2088__;
  assign \result[14]  = ~new_new_n2067__ & ~new_new_n2089__;
  assign new_new_n2091__ = ~\shift[2]  & ~new_new_n1269__;
  assign new_new_n2092__ = \shift[2]  & ~new_new_n1890__;
  assign new_new_n2093__ = ~new_new_n2091__ & ~new_new_n2092__;
  assign new_new_n2094__ = \shift[5]  & ~new_new_n2093__;
  assign new_new_n2095__ = \shift[2]  & ~new_new_n1896__;
  assign new_new_n2096__ = ~\shift[2]  & ~new_new_n1291__;
  assign new_new_n2097__ = ~new_new_n2095__ & ~new_new_n2096__;
  assign new_new_n2098__ = ~\shift[5]  & ~new_new_n2097__;
  assign new_new_n2099__ = ~new_new_n2094__ & ~new_new_n2098__;
  assign new_new_n2100__ = \shift[4]  & ~new_new_n2099__;
  assign new_new_n2101__ = \shift[2]  & ~new_new_n1905__;
  assign new_new_n2102__ = ~\shift[2]  & ~new_new_n1255__;
  assign new_new_n2103__ = ~new_new_n2101__ & ~new_new_n2102__;
  assign new_new_n2104__ = \shift[5]  & ~new_new_n2103__;
  assign new_new_n2105__ = ~\shift[2]  & ~new_new_n1363__;
  assign new_new_n2106__ = \shift[2]  & ~new_new_n1913__;
  assign new_new_n2107__ = ~new_new_n2105__ & ~new_new_n2106__;
  assign new_new_n2108__ = ~\shift[5]  & ~new_new_n2107__;
  assign new_new_n2109__ = ~new_new_n2104__ & ~new_new_n2108__;
  assign new_new_n2110__ = ~\shift[4]  & ~new_new_n2109__;
  assign new_new_n2111__ = ~new_new_n2100__ & ~new_new_n2110__;
  assign new_new_n2112__ = \shift[6]  & ~new_new_n2111__;
  assign new_new_n2113__ = \shift[2]  & ~new_new_n1923__;
  assign new_new_n2114__ = ~\shift[2]  & ~new_new_n1317__;
  assign new_new_n2115__ = ~new_new_n2113__ & ~new_new_n2114__;
  assign new_new_n2116__ = \shift[5]  & ~new_new_n2115__;
  assign new_new_n2117__ = ~\shift[2]  & ~new_new_n1339__;
  assign new_new_n2118__ = \shift[2]  & ~new_new_n1931__;
  assign new_new_n2119__ = ~new_new_n2117__ & ~new_new_n2118__;
  assign new_new_n2120__ = ~\shift[5]  & ~new_new_n2119__;
  assign new_new_n2121__ = ~new_new_n2116__ & ~new_new_n2120__;
  assign new_new_n2122__ = \shift[4]  & ~new_new_n2121__;
  assign new_new_n2123__ = \shift[2]  & ~new_new_n1939__;
  assign new_new_n2124__ = ~\shift[2]  & ~new_new_n1385__;
  assign new_new_n2125__ = ~new_new_n2123__ & ~new_new_n2124__;
  assign new_new_n2126__ = \shift[5]  & ~new_new_n2125__;
  assign new_new_n2127__ = \shift[2]  & ~new_new_n1946__;
  assign new_new_n2128__ = ~\shift[2]  & ~new_new_n1223__;
  assign new_new_n2129__ = ~new_new_n2127__ & ~new_new_n2128__;
  assign new_new_n2130__ = ~\shift[5]  & ~new_new_n2129__;
  assign new_new_n2131__ = ~new_new_n2126__ & ~new_new_n2130__;
  assign new_new_n2132__ = ~\shift[4]  & ~new_new_n2131__;
  assign new_new_n2133__ = ~new_new_n2122__ & ~new_new_n2132__;
  assign new_new_n2134__ = ~\shift[6]  & ~new_new_n2133__;
  assign \result[15]  = ~new_new_n2112__ & ~new_new_n2134__;
  assign new_new_n2136__ = \shift[4]  & ~new_new_n450__;
  assign new_new_n2137__ = ~\shift[5]  & ~new_new_n498__;
  assign new_new_n2138__ = \shift[5]  & ~new_new_n354__;
  assign new_new_n2139__ = ~new_new_n2137__ & ~new_new_n2138__;
  assign new_new_n2140__ = ~\shift[4]  & ~new_new_n2139__;
  assign new_new_n2141__ = ~new_new_n2136__ & ~new_new_n2140__;
  assign new_new_n2142__ = \shift[6]  & ~new_new_n2141__;
  assign new_new_n2143__ = \shift[5]  & ~new_new_n544__;
  assign new_new_n2144__ = ~\shift[5]  & ~new_new_n308__;
  assign new_new_n2145__ = ~new_new_n2143__ & ~new_new_n2144__;
  assign new_new_n2146__ = ~\shift[4]  & ~new_new_n2145__;
  assign new_new_n2147__ = \shift[4]  & ~new_new_n640__;
  assign new_new_n2148__ = ~new_new_n2146__ & ~new_new_n2147__;
  assign new_new_n2149__ = ~\shift[6]  & ~new_new_n2148__;
  assign \result[16]  = ~new_new_n2142__ & ~new_new_n2149__;
  assign new_new_n2151__ = \shift[4]  & ~new_new_n713__;
  assign new_new_n2152__ = ~\shift[5]  & ~new_new_n853__;
  assign new_new_n2153__ = \shift[5]  & ~new_new_n747__;
  assign new_new_n2154__ = ~new_new_n2152__ & ~new_new_n2153__;
  assign new_new_n2155__ = ~\shift[4]  & ~new_new_n2154__;
  assign new_new_n2156__ = ~new_new_n2151__ & ~new_new_n2155__;
  assign new_new_n2157__ = ~\shift[6]  & ~new_new_n2156__;
  assign new_new_n2158__ = \shift[4]  & ~new_new_n925__;
  assign new_new_n2159__ = \shift[5]  & ~new_new_n819__;
  assign new_new_n2160__ = ~\shift[5]  & ~new_new_n781__;
  assign new_new_n2161__ = ~new_new_n2159__ & ~new_new_n2160__;
  assign new_new_n2162__ = ~\shift[4]  & ~new_new_n2161__;
  assign new_new_n2163__ = ~new_new_n2158__ & ~new_new_n2162__;
  assign new_new_n2164__ = \shift[6]  & ~new_new_n2163__;
  assign \result[17]  = new_new_n2157__ | new_new_n2164__;
  assign new_new_n2166__ = ~\shift[5]  & ~new_new_n1104__;
  assign new_new_n2167__ = \shift[5]  & ~new_new_n1066__;
  assign new_new_n2168__ = ~new_new_n2166__ & ~new_new_n2167__;
  assign new_new_n2169__ = ~\shift[4]  & ~new_new_n2168__;
  assign new_new_n2170__ = \shift[4]  & ~new_new_n998__;
  assign new_new_n2171__ = ~new_new_n2169__ & ~new_new_n2170__;
  assign new_new_n2172__ = \shift[6]  & ~new_new_n2171__;
  assign new_new_n2173__ = \shift[5]  & ~new_new_n1138__;
  assign new_new_n2174__ = ~\shift[5]  & ~new_new_n1032__;
  assign new_new_n2175__ = ~new_new_n2173__ & ~new_new_n2174__;
  assign new_new_n2176__ = ~\shift[4]  & ~new_new_n2175__;
  assign new_new_n2177__ = \shift[4]  & ~new_new_n1210__;
  assign new_new_n2178__ = ~new_new_n2176__ & ~new_new_n2177__;
  assign new_new_n2179__ = ~\shift[6]  & ~new_new_n2178__;
  assign \result[18]  = ~new_new_n2172__ & ~new_new_n2179__;
  assign new_new_n2181__ = ~\shift[5]  & ~new_new_n1375__;
  assign new_new_n2182__ = \shift[5]  & ~new_new_n1257__;
  assign new_new_n2183__ = ~new_new_n2181__ & ~new_new_n2182__;
  assign new_new_n2184__ = ~\shift[4]  & ~new_new_n2183__;
  assign new_new_n2185__ = \shift[4]  & ~new_new_n1305__;
  assign new_new_n2186__ = ~new_new_n2184__ & ~new_new_n2185__;
  assign new_new_n2187__ = \shift[6]  & ~new_new_n2186__;
  assign new_new_n2188__ = \shift[5]  & ~new_new_n1397__;
  assign new_new_n2189__ = ~\shift[5]  & ~new_new_n1235__;
  assign new_new_n2190__ = ~new_new_n2188__ & ~new_new_n2189__;
  assign new_new_n2191__ = ~\shift[4]  & ~new_new_n2190__;
  assign new_new_n2192__ = \shift[4]  & ~new_new_n1353__;
  assign new_new_n2193__ = ~new_new_n2191__ & ~new_new_n2192__;
  assign new_new_n2194__ = ~\shift[6]  & ~new_new_n2193__;
  assign \result[19]  = ~new_new_n2187__ & ~new_new_n2194__;
  assign new_new_n2196__ = \shift[4]  & ~new_new_n1434__;
  assign new_new_n2197__ = \shift[5]  & ~new_new_n1416__;
  assign new_new_n2198__ = ~\shift[5]  & ~new_new_n1443__;
  assign new_new_n2199__ = ~new_new_n2197__ & ~new_new_n2198__;
  assign new_new_n2200__ = ~\shift[4]  & ~new_new_n2199__;
  assign new_new_n2201__ = ~new_new_n2196__ & ~new_new_n2200__;
  assign new_new_n2202__ = \shift[6]  & ~new_new_n2201__;
  assign new_new_n2203__ = \shift[5]  & ~new_new_n1450__;
  assign new_new_n2204__ = ~\shift[5]  & ~new_new_n1409__;
  assign new_new_n2205__ = ~new_new_n2203__ & ~new_new_n2204__;
  assign new_new_n2206__ = ~\shift[4]  & ~new_new_n2205__;
  assign new_new_n2207__ = \shift[4]  & ~new_new_n1468__;
  assign new_new_n2208__ = ~new_new_n2206__ & ~new_new_n2207__;
  assign new_new_n2209__ = ~\shift[6]  & ~new_new_n2208__;
  assign \result[20]  = ~new_new_n2202__ & ~new_new_n2209__;
  assign new_new_n2211__ = \shift[4]  & ~new_new_n1487__;
  assign new_new_n2212__ = ~\shift[5]  & ~new_new_n1535__;
  assign new_new_n2213__ = \shift[5]  & ~new_new_n1494__;
  assign new_new_n2214__ = ~new_new_n2212__ & ~new_new_n2213__;
  assign new_new_n2215__ = ~\shift[4]  & ~new_new_n2214__;
  assign new_new_n2216__ = ~new_new_n2211__ & ~new_new_n2215__;
  assign new_new_n2217__ = ~\shift[6]  & ~new_new_n2216__;
  assign new_new_n2218__ = ~\shift[5]  & ~new_new_n1501__;
  assign new_new_n2219__ = \shift[5]  & ~new_new_n1528__;
  assign new_new_n2220__ = ~new_new_n2218__ & ~new_new_n2219__;
  assign new_new_n2221__ = ~\shift[4]  & ~new_new_n2220__;
  assign new_new_n2222__ = \shift[4]  & ~new_new_n1521__;
  assign new_new_n2223__ = ~new_new_n2221__ & ~new_new_n2222__;
  assign new_new_n2224__ = \shift[6]  & ~new_new_n2223__;
  assign \result[21]  = new_new_n2217__ | new_new_n2224__;
  assign new_new_n2226__ = \shift[4]  & ~new_new_n1572__;
  assign new_new_n2227__ = \shift[5]  & ~new_new_n1554__;
  assign new_new_n2228__ = ~\shift[5]  & ~new_new_n1581__;
  assign new_new_n2229__ = ~new_new_n2227__ & ~new_new_n2228__;
  assign new_new_n2230__ = ~\shift[4]  & ~new_new_n2229__;
  assign new_new_n2231__ = ~new_new_n2226__ & ~new_new_n2230__;
  assign new_new_n2232__ = \shift[6]  & ~new_new_n2231__;
  assign new_new_n2233__ = \shift[5]  & ~new_new_n1588__;
  assign new_new_n2234__ = ~\shift[5]  & ~new_new_n1547__;
  assign new_new_n2235__ = ~new_new_n2233__ & ~new_new_n2234__;
  assign new_new_n2236__ = ~\shift[4]  & ~new_new_n2235__;
  assign new_new_n2237__ = \shift[4]  & ~new_new_n1606__;
  assign new_new_n2238__ = ~new_new_n2236__ & ~new_new_n2237__;
  assign new_new_n2239__ = ~\shift[6]  & ~new_new_n2238__;
  assign \result[22]  = ~new_new_n2232__ & ~new_new_n2239__;
  assign new_new_n2241__ = \shift[4]  & ~new_new_n1641__;
  assign new_new_n2242__ = \shift[5]  & ~new_new_n1623__;
  assign new_new_n2243__ = ~\shift[5]  & ~new_new_n1650__;
  assign new_new_n2244__ = ~new_new_n2242__ & ~new_new_n2243__;
  assign new_new_n2245__ = ~\shift[4]  & ~new_new_n2244__;
  assign new_new_n2246__ = ~new_new_n2241__ & ~new_new_n2245__;
  assign new_new_n2247__ = \shift[6]  & ~new_new_n2246__;
  assign new_new_n2248__ = \shift[5]  & ~new_new_n1657__;
  assign new_new_n2249__ = ~\shift[5]  & ~new_new_n1616__;
  assign new_new_n2250__ = ~new_new_n2248__ & ~new_new_n2249__;
  assign new_new_n2251__ = ~\shift[4]  & ~new_new_n2250__;
  assign new_new_n2252__ = \shift[4]  & ~new_new_n1675__;
  assign new_new_n2253__ = ~new_new_n2251__ & ~new_new_n2252__;
  assign new_new_n2254__ = ~\shift[6]  & ~new_new_n2253__;
  assign \result[23]  = ~new_new_n2247__ & ~new_new_n2254__;
  assign new_new_n2256__ = \shift[4]  & ~new_new_n1710__;
  assign new_new_n2257__ = \shift[5]  & ~new_new_n1692__;
  assign new_new_n2258__ = ~\shift[5]  & ~new_new_n1719__;
  assign new_new_n2259__ = ~new_new_n2257__ & ~new_new_n2258__;
  assign new_new_n2260__ = ~\shift[4]  & ~new_new_n2259__;
  assign new_new_n2261__ = ~new_new_n2256__ & ~new_new_n2260__;
  assign new_new_n2262__ = \shift[6]  & ~new_new_n2261__;
  assign new_new_n2263__ = \shift[5]  & ~new_new_n1726__;
  assign new_new_n2264__ = ~\shift[5]  & ~new_new_n1685__;
  assign new_new_n2265__ = ~new_new_n2263__ & ~new_new_n2264__;
  assign new_new_n2266__ = ~\shift[4]  & ~new_new_n2265__;
  assign new_new_n2267__ = \shift[4]  & ~new_new_n1744__;
  assign new_new_n2268__ = ~new_new_n2266__ & ~new_new_n2267__;
  assign new_new_n2269__ = ~\shift[6]  & ~new_new_n2268__;
  assign \result[24]  = ~new_new_n2262__ & ~new_new_n2269__;
  assign new_new_n2271__ = \shift[4]  & ~new_new_n1763__;
  assign new_new_n2272__ = ~\shift[5]  & ~new_new_n1811__;
  assign new_new_n2273__ = \shift[5]  & ~new_new_n1770__;
  assign new_new_n2274__ = ~new_new_n2272__ & ~new_new_n2273__;
  assign new_new_n2275__ = ~\shift[4]  & ~new_new_n2274__;
  assign new_new_n2276__ = ~new_new_n2271__ & ~new_new_n2275__;
  assign new_new_n2277__ = ~\shift[6]  & ~new_new_n2276__;
  assign new_new_n2278__ = ~\shift[5]  & ~new_new_n1777__;
  assign new_new_n2279__ = \shift[5]  & ~new_new_n1804__;
  assign new_new_n2280__ = ~new_new_n2278__ & ~new_new_n2279__;
  assign new_new_n2281__ = ~\shift[4]  & ~new_new_n2280__;
  assign new_new_n2282__ = \shift[4]  & ~new_new_n1797__;
  assign new_new_n2283__ = ~new_new_n2281__ & ~new_new_n2282__;
  assign new_new_n2284__ = \shift[6]  & ~new_new_n2283__;
  assign \result[25]  = new_new_n2277__ | new_new_n2284__;
  assign new_new_n2286__ = \shift[4]  & ~new_new_n1848__;
  assign new_new_n2287__ = \shift[5]  & ~new_new_n1830__;
  assign new_new_n2288__ = ~\shift[5]  & ~new_new_n1857__;
  assign new_new_n2289__ = ~new_new_n2287__ & ~new_new_n2288__;
  assign new_new_n2290__ = ~\shift[4]  & ~new_new_n2289__;
  assign new_new_n2291__ = ~new_new_n2286__ & ~new_new_n2290__;
  assign new_new_n2292__ = \shift[6]  & ~new_new_n2291__;
  assign new_new_n2293__ = \shift[5]  & ~new_new_n1864__;
  assign new_new_n2294__ = ~\shift[5]  & ~new_new_n1823__;
  assign new_new_n2295__ = ~new_new_n2293__ & ~new_new_n2294__;
  assign new_new_n2296__ = ~\shift[4]  & ~new_new_n2295__;
  assign new_new_n2297__ = \shift[4]  & ~new_new_n1882__;
  assign new_new_n2298__ = ~new_new_n2296__ & ~new_new_n2297__;
  assign new_new_n2299__ = ~\shift[6]  & ~new_new_n2298__;
  assign \result[26]  = ~new_new_n2292__ & ~new_new_n2299__;
  assign new_new_n2301__ = \shift[4]  & ~new_new_n1917__;
  assign new_new_n2302__ = \shift[5]  & ~new_new_n1899__;
  assign new_new_n2303__ = ~\shift[5]  & ~new_new_n1926__;
  assign new_new_n2304__ = ~new_new_n2302__ & ~new_new_n2303__;
  assign new_new_n2305__ = ~\shift[4]  & ~new_new_n2304__;
  assign new_new_n2306__ = ~new_new_n2301__ & ~new_new_n2305__;
  assign new_new_n2307__ = \shift[6]  & ~new_new_n2306__;
  assign new_new_n2308__ = \shift[5]  & ~new_new_n1933__;
  assign new_new_n2309__ = ~\shift[5]  & ~new_new_n1892__;
  assign new_new_n2310__ = ~new_new_n2308__ & ~new_new_n2309__;
  assign new_new_n2311__ = ~\shift[4]  & ~new_new_n2310__;
  assign new_new_n2312__ = \shift[4]  & ~new_new_n1951__;
  assign new_new_n2313__ = ~new_new_n2311__ & ~new_new_n2312__;
  assign new_new_n2314__ = ~\shift[6]  & ~new_new_n2313__;
  assign \result[27]  = ~new_new_n2307__ & ~new_new_n2314__;
  assign new_new_n2316__ = \shift[4]  & ~new_new_n1974__;
  assign new_new_n2317__ = \shift[5]  & ~new_new_n1962__;
  assign new_new_n2318__ = ~\shift[5]  & ~new_new_n1980__;
  assign new_new_n2319__ = ~new_new_n2317__ & ~new_new_n2318__;
  assign new_new_n2320__ = ~\shift[4]  & ~new_new_n2319__;
  assign new_new_n2321__ = ~new_new_n2316__ & ~new_new_n2320__;
  assign new_new_n2322__ = \shift[6]  & ~new_new_n2321__;
  assign new_new_n2323__ = \shift[5]  & ~new_new_n1984__;
  assign new_new_n2324__ = ~\shift[5]  & ~new_new_n1958__;
  assign new_new_n2325__ = ~new_new_n2323__ & ~new_new_n2324__;
  assign new_new_n2326__ = ~\shift[4]  & ~new_new_n2325__;
  assign new_new_n2327__ = \shift[4]  & ~new_new_n1996__;
  assign new_new_n2328__ = ~new_new_n2326__ & ~new_new_n2327__;
  assign new_new_n2329__ = ~\shift[6]  & ~new_new_n2328__;
  assign \result[28]  = ~new_new_n2322__ & ~new_new_n2329__;
  assign new_new_n2331__ = \shift[4]  & ~new_new_n2009__;
  assign new_new_n2332__ = ~\shift[5]  & ~new_new_n2039__;
  assign new_new_n2333__ = \shift[5]  & ~new_new_n2013__;
  assign new_new_n2334__ = ~new_new_n2332__ & ~new_new_n2333__;
  assign new_new_n2335__ = ~\shift[4]  & ~new_new_n2334__;
  assign new_new_n2336__ = ~new_new_n2331__ & ~new_new_n2335__;
  assign new_new_n2337__ = ~\shift[6]  & ~new_new_n2336__;
  assign new_new_n2338__ = ~\shift[5]  & ~new_new_n2017__;
  assign new_new_n2339__ = \shift[5]  & ~new_new_n2035__;
  assign new_new_n2340__ = ~new_new_n2338__ & ~new_new_n2339__;
  assign new_new_n2341__ = ~\shift[4]  & ~new_new_n2340__;
  assign new_new_n2342__ = \shift[4]  & ~new_new_n2031__;
  assign new_new_n2343__ = ~new_new_n2341__ & ~new_new_n2342__;
  assign new_new_n2344__ = \shift[6]  & ~new_new_n2343__;
  assign \result[29]  = new_new_n2337__ | new_new_n2344__;
  assign new_new_n2346__ = \shift[4]  & ~new_new_n2064__;
  assign new_new_n2347__ = \shift[5]  & ~new_new_n2052__;
  assign new_new_n2348__ = ~\shift[5]  & ~new_new_n2070__;
  assign new_new_n2349__ = ~new_new_n2347__ & ~new_new_n2348__;
  assign new_new_n2350__ = ~\shift[4]  & ~new_new_n2349__;
  assign new_new_n2351__ = ~new_new_n2346__ & ~new_new_n2350__;
  assign new_new_n2352__ = \shift[6]  & ~new_new_n2351__;
  assign new_new_n2353__ = \shift[5]  & ~new_new_n2074__;
  assign new_new_n2354__ = ~\shift[5]  & ~new_new_n2048__;
  assign new_new_n2355__ = ~new_new_n2353__ & ~new_new_n2354__;
  assign new_new_n2356__ = ~\shift[4]  & ~new_new_n2355__;
  assign new_new_n2357__ = \shift[4]  & ~new_new_n2086__;
  assign new_new_n2358__ = ~new_new_n2356__ & ~new_new_n2357__;
  assign new_new_n2359__ = ~\shift[6]  & ~new_new_n2358__;
  assign \result[30]  = ~new_new_n2352__ & ~new_new_n2359__;
  assign new_new_n2361__ = \shift[4]  & ~new_new_n2109__;
  assign new_new_n2362__ = \shift[5]  & ~new_new_n2097__;
  assign new_new_n2363__ = ~\shift[5]  & ~new_new_n2115__;
  assign new_new_n2364__ = ~new_new_n2362__ & ~new_new_n2363__;
  assign new_new_n2365__ = ~\shift[4]  & ~new_new_n2364__;
  assign new_new_n2366__ = ~new_new_n2361__ & ~new_new_n2365__;
  assign new_new_n2367__ = \shift[6]  & ~new_new_n2366__;
  assign new_new_n2368__ = \shift[5]  & ~new_new_n2119__;
  assign new_new_n2369__ = ~\shift[5]  & ~new_new_n2093__;
  assign new_new_n2370__ = ~new_new_n2368__ & ~new_new_n2369__;
  assign new_new_n2371__ = ~\shift[4]  & ~new_new_n2370__;
  assign new_new_n2372__ = \shift[4]  & ~new_new_n2131__;
  assign new_new_n2373__ = ~new_new_n2371__ & ~new_new_n2372__;
  assign new_new_n2374__ = ~\shift[6]  & ~new_new_n2373__;
  assign \result[31]  = ~new_new_n2367__ & ~new_new_n2374__;
  assign new_new_n2376__ = \shift[4]  & ~new_new_n2139__;
  assign new_new_n2377__ = \shift[5]  & ~new_new_n448__;
  assign new_new_n2378__ = ~\shift[5]  & ~new_new_n592__;
  assign new_new_n2379__ = ~new_new_n2377__ & ~new_new_n2378__;
  assign new_new_n2380__ = ~\shift[4]  & ~new_new_n2379__;
  assign new_new_n2381__ = ~new_new_n2376__ & ~new_new_n2380__;
  assign new_new_n2382__ = \shift[6]  & ~new_new_n2381__;
  assign new_new_n2383__ = \shift[4]  & ~new_new_n2145__;
  assign new_new_n2384__ = \shift[5]  & ~new_new_n638__;
  assign new_new_n2385__ = ~\shift[5]  & ~new_new_n402__;
  assign new_new_n2386__ = ~new_new_n2384__ & ~new_new_n2385__;
  assign new_new_n2387__ = ~\shift[4]  & ~new_new_n2386__;
  assign new_new_n2388__ = ~new_new_n2383__ & ~new_new_n2387__;
  assign new_new_n2389__ = ~\shift[6]  & ~new_new_n2388__;
  assign \result[32]  = ~new_new_n2382__ & ~new_new_n2389__;
  assign new_new_n2391__ = ~\shift[5]  & ~new_new_n923__;
  assign new_new_n2392__ = \shift[5]  & ~new_new_n677__;
  assign new_new_n2393__ = ~new_new_n2391__ & ~new_new_n2392__;
  assign new_new_n2394__ = ~\shift[4]  & ~new_new_n2393__;
  assign new_new_n2395__ = \shift[4]  & ~new_new_n2154__;
  assign new_new_n2396__ = ~new_new_n2394__ & ~new_new_n2395__;
  assign new_new_n2397__ = ~\shift[6]  & ~new_new_n2396__;
  assign new_new_n2398__ = ~\shift[5]  & ~new_new_n711__;
  assign new_new_n2399__ = \shift[5]  & ~new_new_n889__;
  assign new_new_n2400__ = ~new_new_n2398__ & ~new_new_n2399__;
  assign new_new_n2401__ = ~\shift[4]  & ~new_new_n2400__;
  assign new_new_n2402__ = \shift[4]  & ~new_new_n2161__;
  assign new_new_n2403__ = ~new_new_n2401__ & ~new_new_n2402__;
  assign new_new_n2404__ = \shift[6]  & ~new_new_n2403__;
  assign \result[33]  = new_new_n2397__ | new_new_n2404__;
  assign new_new_n2406__ = \shift[4]  & ~new_new_n2168__;
  assign new_new_n2407__ = \shift[5]  & ~new_new_n996__;
  assign new_new_n2408__ = ~\shift[5]  & ~new_new_n1174__;
  assign new_new_n2409__ = ~new_new_n2407__ & ~new_new_n2408__;
  assign new_new_n2410__ = ~\shift[4]  & ~new_new_n2409__;
  assign new_new_n2411__ = ~new_new_n2406__ & ~new_new_n2410__;
  assign new_new_n2412__ = \shift[6]  & ~new_new_n2411__;
  assign new_new_n2413__ = \shift[4]  & ~new_new_n2175__;
  assign new_new_n2414__ = \shift[5]  & ~new_new_n1208__;
  assign new_new_n2415__ = ~\shift[5]  & ~new_new_n962__;
  assign new_new_n2416__ = ~new_new_n2414__ & ~new_new_n2415__;
  assign new_new_n2417__ = ~\shift[4]  & ~new_new_n2416__;
  assign new_new_n2418__ = ~new_new_n2413__ & ~new_new_n2417__;
  assign new_new_n2419__ = ~\shift[6]  & ~new_new_n2418__;
  assign \result[34]  = ~new_new_n2412__ & ~new_new_n2419__;
  assign new_new_n2421__ = \shift[4]  & ~new_new_n2183__;
  assign new_new_n2422__ = \shift[5]  & ~new_new_n1303__;
  assign new_new_n2423__ = ~\shift[5]  & ~new_new_n1329__;
  assign new_new_n2424__ = ~new_new_n2422__ & ~new_new_n2423__;
  assign new_new_n2425__ = ~\shift[4]  & ~new_new_n2424__;
  assign new_new_n2426__ = ~new_new_n2421__ & ~new_new_n2425__;
  assign new_new_n2427__ = \shift[6]  & ~new_new_n2426__;
  assign new_new_n2428__ = \shift[4]  & ~new_new_n2190__;
  assign new_new_n2429__ = ~\shift[5]  & ~new_new_n1281__;
  assign new_new_n2430__ = \shift[5]  & ~new_new_n1351__;
  assign new_new_n2431__ = ~new_new_n2429__ & ~new_new_n2430__;
  assign new_new_n2432__ = ~\shift[4]  & ~new_new_n2431__;
  assign new_new_n2433__ = ~new_new_n2428__ & ~new_new_n2432__;
  assign new_new_n2434__ = ~\shift[6]  & ~new_new_n2433__;
  assign \result[35]  = ~new_new_n2427__ & ~new_new_n2434__;
  assign new_new_n2436__ = \shift[4]  & ~new_new_n2199__;
  assign new_new_n2437__ = ~\shift[5]  & ~new_new_n1459__;
  assign new_new_n2438__ = \shift[5]  & ~new_new_n1432__;
  assign new_new_n2439__ = ~new_new_n2437__ & ~new_new_n2438__;
  assign new_new_n2440__ = ~\shift[4]  & ~new_new_n2439__;
  assign new_new_n2441__ = ~new_new_n2436__ & ~new_new_n2440__;
  assign new_new_n2442__ = \shift[6]  & ~new_new_n2441__;
  assign new_new_n2443__ = \shift[5]  & ~new_new_n1466__;
  assign new_new_n2444__ = ~\shift[5]  & ~new_new_n1425__;
  assign new_new_n2445__ = ~new_new_n2443__ & ~new_new_n2444__;
  assign new_new_n2446__ = ~\shift[4]  & ~new_new_n2445__;
  assign new_new_n2447__ = \shift[4]  & ~new_new_n2205__;
  assign new_new_n2448__ = ~new_new_n2446__ & ~new_new_n2447__;
  assign new_new_n2449__ = ~\shift[6]  & ~new_new_n2448__;
  assign \result[36]  = ~new_new_n2442__ & ~new_new_n2449__;
  assign new_new_n2451__ = \shift[4]  & ~new_new_n2214__;
  assign new_new_n2452__ = ~\shift[5]  & ~new_new_n1519__;
  assign new_new_n2453__ = \shift[5]  & ~new_new_n1478__;
  assign new_new_n2454__ = ~new_new_n2452__ & ~new_new_n2453__;
  assign new_new_n2455__ = ~\shift[4]  & ~new_new_n2454__;
  assign new_new_n2456__ = ~new_new_n2451__ & ~new_new_n2455__;
  assign new_new_n2457__ = ~\shift[6]  & ~new_new_n2456__;
  assign new_new_n2458__ = \shift[5]  & ~new_new_n1512__;
  assign new_new_n2459__ = ~\shift[5]  & ~new_new_n1485__;
  assign new_new_n2460__ = ~new_new_n2458__ & ~new_new_n2459__;
  assign new_new_n2461__ = ~\shift[4]  & ~new_new_n2460__;
  assign new_new_n2462__ = \shift[4]  & ~new_new_n2220__;
  assign new_new_n2463__ = ~new_new_n2461__ & ~new_new_n2462__;
  assign new_new_n2464__ = \shift[6]  & ~new_new_n2463__;
  assign \result[37]  = new_new_n2457__ | new_new_n2464__;
  assign new_new_n2466__ = \shift[4]  & ~new_new_n2229__;
  assign new_new_n2467__ = ~\shift[5]  & ~new_new_n1597__;
  assign new_new_n2468__ = \shift[5]  & ~new_new_n1570__;
  assign new_new_n2469__ = ~new_new_n2467__ & ~new_new_n2468__;
  assign new_new_n2470__ = ~\shift[4]  & ~new_new_n2469__;
  assign new_new_n2471__ = ~new_new_n2466__ & ~new_new_n2470__;
  assign new_new_n2472__ = \shift[6]  & ~new_new_n2471__;
  assign new_new_n2473__ = \shift[5]  & ~new_new_n1604__;
  assign new_new_n2474__ = ~\shift[5]  & ~new_new_n1563__;
  assign new_new_n2475__ = ~new_new_n2473__ & ~new_new_n2474__;
  assign new_new_n2476__ = ~\shift[4]  & ~new_new_n2475__;
  assign new_new_n2477__ = \shift[4]  & ~new_new_n2235__;
  assign new_new_n2478__ = ~new_new_n2476__ & ~new_new_n2477__;
  assign new_new_n2479__ = ~\shift[6]  & ~new_new_n2478__;
  assign \result[38]  = ~new_new_n2472__ & ~new_new_n2479__;
  assign new_new_n2481__ = \shift[4]  & ~new_new_n2244__;
  assign new_new_n2482__ = ~\shift[5]  & ~new_new_n1666__;
  assign new_new_n2483__ = \shift[5]  & ~new_new_n1639__;
  assign new_new_n2484__ = ~new_new_n2482__ & ~new_new_n2483__;
  assign new_new_n2485__ = ~\shift[4]  & ~new_new_n2484__;
  assign new_new_n2486__ = ~new_new_n2481__ & ~new_new_n2485__;
  assign new_new_n2487__ = \shift[6]  & ~new_new_n2486__;
  assign new_new_n2488__ = \shift[5]  & ~new_new_n1673__;
  assign new_new_n2489__ = ~\shift[5]  & ~new_new_n1632__;
  assign new_new_n2490__ = ~new_new_n2488__ & ~new_new_n2489__;
  assign new_new_n2491__ = ~\shift[4]  & ~new_new_n2490__;
  assign new_new_n2492__ = \shift[4]  & ~new_new_n2250__;
  assign new_new_n2493__ = ~new_new_n2491__ & ~new_new_n2492__;
  assign new_new_n2494__ = ~\shift[6]  & ~new_new_n2493__;
  assign \result[39]  = ~new_new_n2487__ & ~new_new_n2494__;
  assign new_new_n2496__ = \shift[4]  & ~new_new_n2259__;
  assign new_new_n2497__ = ~\shift[5]  & ~new_new_n1735__;
  assign new_new_n2498__ = \shift[5]  & ~new_new_n1708__;
  assign new_new_n2499__ = ~new_new_n2497__ & ~new_new_n2498__;
  assign new_new_n2500__ = ~\shift[4]  & ~new_new_n2499__;
  assign new_new_n2501__ = ~new_new_n2496__ & ~new_new_n2500__;
  assign new_new_n2502__ = \shift[6]  & ~new_new_n2501__;
  assign new_new_n2503__ = \shift[5]  & ~new_new_n1742__;
  assign new_new_n2504__ = ~\shift[5]  & ~new_new_n1701__;
  assign new_new_n2505__ = ~new_new_n2503__ & ~new_new_n2504__;
  assign new_new_n2506__ = ~\shift[4]  & ~new_new_n2505__;
  assign new_new_n2507__ = \shift[4]  & ~new_new_n2265__;
  assign new_new_n2508__ = ~new_new_n2506__ & ~new_new_n2507__;
  assign new_new_n2509__ = ~\shift[6]  & ~new_new_n2508__;
  assign \result[40]  = ~new_new_n2502__ & ~new_new_n2509__;
  assign new_new_n2511__ = \shift[4]  & ~new_new_n2274__;
  assign new_new_n2512__ = ~\shift[5]  & ~new_new_n1795__;
  assign new_new_n2513__ = \shift[5]  & ~new_new_n1754__;
  assign new_new_n2514__ = ~new_new_n2512__ & ~new_new_n2513__;
  assign new_new_n2515__ = ~\shift[4]  & ~new_new_n2514__;
  assign new_new_n2516__ = ~new_new_n2511__ & ~new_new_n2515__;
  assign new_new_n2517__ = ~\shift[6]  & ~new_new_n2516__;
  assign new_new_n2518__ = \shift[5]  & ~new_new_n1788__;
  assign new_new_n2519__ = ~\shift[5]  & ~new_new_n1761__;
  assign new_new_n2520__ = ~new_new_n2518__ & ~new_new_n2519__;
  assign new_new_n2521__ = ~\shift[4]  & ~new_new_n2520__;
  assign new_new_n2522__ = \shift[4]  & ~new_new_n2280__;
  assign new_new_n2523__ = ~new_new_n2521__ & ~new_new_n2522__;
  assign new_new_n2524__ = \shift[6]  & ~new_new_n2523__;
  assign \result[41]  = new_new_n2517__ | new_new_n2524__;
  assign new_new_n2526__ = \shift[4]  & ~new_new_n2289__;
  assign new_new_n2527__ = ~\shift[5]  & ~new_new_n1873__;
  assign new_new_n2528__ = \shift[5]  & ~new_new_n1846__;
  assign new_new_n2529__ = ~new_new_n2527__ & ~new_new_n2528__;
  assign new_new_n2530__ = ~\shift[4]  & ~new_new_n2529__;
  assign new_new_n2531__ = ~new_new_n2526__ & ~new_new_n2530__;
  assign new_new_n2532__ = \shift[6]  & ~new_new_n2531__;
  assign new_new_n2533__ = \shift[5]  & ~new_new_n1880__;
  assign new_new_n2534__ = ~\shift[5]  & ~new_new_n1839__;
  assign new_new_n2535__ = ~new_new_n2533__ & ~new_new_n2534__;
  assign new_new_n2536__ = ~\shift[4]  & ~new_new_n2535__;
  assign new_new_n2537__ = \shift[4]  & ~new_new_n2295__;
  assign new_new_n2538__ = ~new_new_n2536__ & ~new_new_n2537__;
  assign new_new_n2539__ = ~\shift[6]  & ~new_new_n2538__;
  assign \result[42]  = ~new_new_n2532__ & ~new_new_n2539__;
  assign new_new_n2541__ = \shift[4]  & ~new_new_n2304__;
  assign new_new_n2542__ = ~\shift[5]  & ~new_new_n1942__;
  assign new_new_n2543__ = \shift[5]  & ~new_new_n1915__;
  assign new_new_n2544__ = ~new_new_n2542__ & ~new_new_n2543__;
  assign new_new_n2545__ = ~\shift[4]  & ~new_new_n2544__;
  assign new_new_n2546__ = ~new_new_n2541__ & ~new_new_n2545__;
  assign new_new_n2547__ = \shift[6]  & ~new_new_n2546__;
  assign new_new_n2548__ = \shift[5]  & ~new_new_n1949__;
  assign new_new_n2549__ = ~\shift[5]  & ~new_new_n1908__;
  assign new_new_n2550__ = ~new_new_n2548__ & ~new_new_n2549__;
  assign new_new_n2551__ = ~\shift[4]  & ~new_new_n2550__;
  assign new_new_n2552__ = \shift[4]  & ~new_new_n2310__;
  assign new_new_n2553__ = ~new_new_n2551__ & ~new_new_n2552__;
  assign new_new_n2554__ = ~\shift[6]  & ~new_new_n2553__;
  assign \result[43]  = ~new_new_n2547__ & ~new_new_n2554__;
  assign new_new_n2556__ = \shift[4]  & ~new_new_n2319__;
  assign new_new_n2557__ = ~\shift[5]  & ~new_new_n1990__;
  assign new_new_n2558__ = \shift[5]  & ~new_new_n1972__;
  assign new_new_n2559__ = ~new_new_n2557__ & ~new_new_n2558__;
  assign new_new_n2560__ = ~\shift[4]  & ~new_new_n2559__;
  assign new_new_n2561__ = ~new_new_n2556__ & ~new_new_n2560__;
  assign new_new_n2562__ = \shift[6]  & ~new_new_n2561__;
  assign new_new_n2563__ = \shift[5]  & ~new_new_n1994__;
  assign new_new_n2564__ = ~\shift[5]  & ~new_new_n1968__;
  assign new_new_n2565__ = ~new_new_n2563__ & ~new_new_n2564__;
  assign new_new_n2566__ = ~\shift[4]  & ~new_new_n2565__;
  assign new_new_n2567__ = \shift[4]  & ~new_new_n2325__;
  assign new_new_n2568__ = ~new_new_n2566__ & ~new_new_n2567__;
  assign new_new_n2569__ = ~\shift[6]  & ~new_new_n2568__;
  assign \result[44]  = ~new_new_n2562__ & ~new_new_n2569__;
  assign new_new_n2571__ = \shift[4]  & ~new_new_n2334__;
  assign new_new_n2572__ = ~\shift[5]  & ~new_new_n2029__;
  assign new_new_n2573__ = \shift[5]  & ~new_new_n2003__;
  assign new_new_n2574__ = ~new_new_n2572__ & ~new_new_n2573__;
  assign new_new_n2575__ = ~\shift[4]  & ~new_new_n2574__;
  assign new_new_n2576__ = ~new_new_n2571__ & ~new_new_n2575__;
  assign new_new_n2577__ = ~\shift[6]  & ~new_new_n2576__;
  assign new_new_n2578__ = \shift[5]  & ~new_new_n2025__;
  assign new_new_n2579__ = ~\shift[5]  & ~new_new_n2007__;
  assign new_new_n2580__ = ~new_new_n2578__ & ~new_new_n2579__;
  assign new_new_n2581__ = ~\shift[4]  & ~new_new_n2580__;
  assign new_new_n2582__ = \shift[4]  & ~new_new_n2340__;
  assign new_new_n2583__ = ~new_new_n2581__ & ~new_new_n2582__;
  assign new_new_n2584__ = \shift[6]  & ~new_new_n2583__;
  assign \result[45]  = new_new_n2577__ | new_new_n2584__;
  assign new_new_n2586__ = \shift[4]  & ~new_new_n2349__;
  assign new_new_n2587__ = ~\shift[5]  & ~new_new_n2080__;
  assign new_new_n2588__ = \shift[5]  & ~new_new_n2062__;
  assign new_new_n2589__ = ~new_new_n2587__ & ~new_new_n2588__;
  assign new_new_n2590__ = ~\shift[4]  & ~new_new_n2589__;
  assign new_new_n2591__ = ~new_new_n2586__ & ~new_new_n2590__;
  assign new_new_n2592__ = \shift[6]  & ~new_new_n2591__;
  assign new_new_n2593__ = \shift[5]  & ~new_new_n2084__;
  assign new_new_n2594__ = ~\shift[5]  & ~new_new_n2058__;
  assign new_new_n2595__ = ~new_new_n2593__ & ~new_new_n2594__;
  assign new_new_n2596__ = ~\shift[4]  & ~new_new_n2595__;
  assign new_new_n2597__ = \shift[4]  & ~new_new_n2355__;
  assign new_new_n2598__ = ~new_new_n2596__ & ~new_new_n2597__;
  assign new_new_n2599__ = ~\shift[6]  & ~new_new_n2598__;
  assign \result[46]  = ~new_new_n2592__ & ~new_new_n2599__;
  assign new_new_n2601__ = \shift[4]  & ~new_new_n2364__;
  assign new_new_n2602__ = ~\shift[5]  & ~new_new_n2125__;
  assign new_new_n2603__ = \shift[5]  & ~new_new_n2107__;
  assign new_new_n2604__ = ~new_new_n2602__ & ~new_new_n2603__;
  assign new_new_n2605__ = ~\shift[4]  & ~new_new_n2604__;
  assign new_new_n2606__ = ~new_new_n2601__ & ~new_new_n2605__;
  assign new_new_n2607__ = \shift[6]  & ~new_new_n2606__;
  assign new_new_n2608__ = \shift[5]  & ~new_new_n2129__;
  assign new_new_n2609__ = ~\shift[5]  & ~new_new_n2103__;
  assign new_new_n2610__ = ~new_new_n2608__ & ~new_new_n2609__;
  assign new_new_n2611__ = ~\shift[4]  & ~new_new_n2610__;
  assign new_new_n2612__ = \shift[4]  & ~new_new_n2370__;
  assign new_new_n2613__ = ~new_new_n2611__ & ~new_new_n2612__;
  assign new_new_n2614__ = ~\shift[6]  & ~new_new_n2613__;
  assign \result[47]  = ~new_new_n2607__ & ~new_new_n2614__;
  assign new_new_n2616__ = \shift[4]  & ~new_new_n2379__;
  assign new_new_n2617__ = ~\shift[4]  & ~new_new_n546__;
  assign new_new_n2618__ = ~new_new_n2616__ & ~new_new_n2617__;
  assign new_new_n2619__ = \shift[6]  & ~new_new_n2618__;
  assign new_new_n2620__ = \shift[4]  & ~new_new_n2386__;
  assign new_new_n2621__ = ~\shift[4]  & ~new_new_n356__;
  assign new_new_n2622__ = ~new_new_n2620__ & ~new_new_n2621__;
  assign new_new_n2623__ = ~\shift[6]  & ~new_new_n2622__;
  assign \result[48]  = ~new_new_n2619__ & ~new_new_n2623__;
  assign new_new_n2625__ = ~\shift[4]  & ~new_new_n855__;
  assign new_new_n2626__ = \shift[4]  & ~new_new_n2393__;
  assign new_new_n2627__ = ~new_new_n2625__ & ~new_new_n2626__;
  assign new_new_n2628__ = ~\shift[6]  & ~new_new_n2627__;
  assign new_new_n2629__ = ~\shift[4]  & ~new_new_n783__;
  assign new_new_n2630__ = \shift[4]  & ~new_new_n2400__;
  assign new_new_n2631__ = ~new_new_n2629__ & ~new_new_n2630__;
  assign new_new_n2632__ = \shift[6]  & ~new_new_n2631__;
  assign \result[49]  = new_new_n2628__ | new_new_n2632__;
  assign new_new_n2634__ = \shift[4]  & ~new_new_n2409__;
  assign new_new_n2635__ = ~\shift[4]  & ~new_new_n1140__;
  assign new_new_n2636__ = ~new_new_n2634__ & ~new_new_n2635__;
  assign new_new_n2637__ = \shift[6]  & ~new_new_n2636__;
  assign new_new_n2638__ = \shift[4]  & ~new_new_n2416__;
  assign new_new_n2639__ = ~\shift[4]  & ~new_new_n1068__;
  assign new_new_n2640__ = ~new_new_n2638__ & ~new_new_n2639__;
  assign new_new_n2641__ = ~\shift[6]  & ~new_new_n2640__;
  assign \result[50]  = ~new_new_n2637__ & ~new_new_n2641__;
  assign new_new_n2643__ = \shift[4]  & ~new_new_n2424__;
  assign new_new_n2644__ = ~\shift[4]  & ~new_new_n1399__;
  assign new_new_n2645__ = ~new_new_n2643__ & ~new_new_n2644__;
  assign new_new_n2646__ = \shift[6]  & ~new_new_n2645__;
  assign new_new_n2647__ = \shift[4]  & ~new_new_n2431__;
  assign new_new_n2648__ = ~\shift[4]  & ~new_new_n1259__;
  assign new_new_n2649__ = ~new_new_n2647__ & ~new_new_n2648__;
  assign new_new_n2650__ = ~\shift[6]  & ~new_new_n2649__;
  assign \result[51]  = ~new_new_n2646__ & ~new_new_n2650__;
  assign new_new_n2652__ = \shift[4]  & ~new_new_n2439__;
  assign new_new_n2653__ = ~\shift[4]  & ~new_new_n1452__;
  assign new_new_n2654__ = ~new_new_n2652__ & ~new_new_n2653__;
  assign new_new_n2655__ = \shift[6]  & ~new_new_n2654__;
  assign new_new_n2656__ = ~\shift[4]  & ~new_new_n1418__;
  assign new_new_n2657__ = \shift[4]  & ~new_new_n2445__;
  assign new_new_n2658__ = ~new_new_n2656__ & ~new_new_n2657__;
  assign new_new_n2659__ = ~\shift[6]  & ~new_new_n2658__;
  assign \result[52]  = ~new_new_n2655__ & ~new_new_n2659__;
  assign new_new_n2661__ = \shift[4]  & ~new_new_n2454__;
  assign new_new_n2662__ = ~\shift[4]  & ~new_new_n1537__;
  assign new_new_n2663__ = ~new_new_n2661__ & ~new_new_n2662__;
  assign new_new_n2664__ = ~\shift[6]  & ~new_new_n2663__;
  assign new_new_n2665__ = ~\shift[4]  & ~new_new_n1503__;
  assign new_new_n2666__ = \shift[4]  & ~new_new_n2460__;
  assign new_new_n2667__ = ~new_new_n2665__ & ~new_new_n2666__;
  assign new_new_n2668__ = \shift[6]  & ~new_new_n2667__;
  assign \result[53]  = new_new_n2664__ | new_new_n2668__;
  assign new_new_n2670__ = \shift[4]  & ~new_new_n2469__;
  assign new_new_n2671__ = ~\shift[4]  & ~new_new_n1590__;
  assign new_new_n2672__ = ~new_new_n2670__ & ~new_new_n2671__;
  assign new_new_n2673__ = \shift[6]  & ~new_new_n2672__;
  assign new_new_n2674__ = ~\shift[4]  & ~new_new_n1556__;
  assign new_new_n2675__ = \shift[4]  & ~new_new_n2475__;
  assign new_new_n2676__ = ~new_new_n2674__ & ~new_new_n2675__;
  assign new_new_n2677__ = ~\shift[6]  & ~new_new_n2676__;
  assign \result[54]  = ~new_new_n2673__ & ~new_new_n2677__;
  assign new_new_n2679__ = \shift[4]  & ~new_new_n2484__;
  assign new_new_n2680__ = ~\shift[4]  & ~new_new_n1659__;
  assign new_new_n2681__ = ~new_new_n2679__ & ~new_new_n2680__;
  assign new_new_n2682__ = \shift[6]  & ~new_new_n2681__;
  assign new_new_n2683__ = ~\shift[4]  & ~new_new_n1625__;
  assign new_new_n2684__ = \shift[4]  & ~new_new_n2490__;
  assign new_new_n2685__ = ~new_new_n2683__ & ~new_new_n2684__;
  assign new_new_n2686__ = ~\shift[6]  & ~new_new_n2685__;
  assign \result[55]  = ~new_new_n2682__ & ~new_new_n2686__;
  assign new_new_n2688__ = \shift[4]  & ~new_new_n2499__;
  assign new_new_n2689__ = ~\shift[4]  & ~new_new_n1728__;
  assign new_new_n2690__ = ~new_new_n2688__ & ~new_new_n2689__;
  assign new_new_n2691__ = \shift[6]  & ~new_new_n2690__;
  assign new_new_n2692__ = ~\shift[4]  & ~new_new_n1694__;
  assign new_new_n2693__ = \shift[4]  & ~new_new_n2505__;
  assign new_new_n2694__ = ~new_new_n2692__ & ~new_new_n2693__;
  assign new_new_n2695__ = ~\shift[6]  & ~new_new_n2694__;
  assign \result[56]  = ~new_new_n2691__ & ~new_new_n2695__;
  assign new_new_n2697__ = \shift[4]  & ~new_new_n2514__;
  assign new_new_n2698__ = ~\shift[4]  & ~new_new_n1813__;
  assign new_new_n2699__ = ~new_new_n2697__ & ~new_new_n2698__;
  assign new_new_n2700__ = ~\shift[6]  & ~new_new_n2699__;
  assign new_new_n2701__ = ~\shift[4]  & ~new_new_n1779__;
  assign new_new_n2702__ = \shift[4]  & ~new_new_n2520__;
  assign new_new_n2703__ = ~new_new_n2701__ & ~new_new_n2702__;
  assign new_new_n2704__ = \shift[6]  & ~new_new_n2703__;
  assign \result[57]  = new_new_n2700__ | new_new_n2704__;
  assign new_new_n2706__ = \shift[4]  & ~new_new_n2529__;
  assign new_new_n2707__ = ~\shift[4]  & ~new_new_n1866__;
  assign new_new_n2708__ = ~new_new_n2706__ & ~new_new_n2707__;
  assign new_new_n2709__ = \shift[6]  & ~new_new_n2708__;
  assign new_new_n2710__ = ~\shift[4]  & ~new_new_n1832__;
  assign new_new_n2711__ = \shift[4]  & ~new_new_n2535__;
  assign new_new_n2712__ = ~new_new_n2710__ & ~new_new_n2711__;
  assign new_new_n2713__ = ~\shift[6]  & ~new_new_n2712__;
  assign \result[58]  = ~new_new_n2709__ & ~new_new_n2713__;
  assign new_new_n2715__ = \shift[4]  & ~new_new_n2544__;
  assign new_new_n2716__ = ~\shift[4]  & ~new_new_n1935__;
  assign new_new_n2717__ = ~new_new_n2715__ & ~new_new_n2716__;
  assign new_new_n2718__ = \shift[6]  & ~new_new_n2717__;
  assign new_new_n2719__ = ~\shift[4]  & ~new_new_n1901__;
  assign new_new_n2720__ = \shift[4]  & ~new_new_n2550__;
  assign new_new_n2721__ = ~new_new_n2719__ & ~new_new_n2720__;
  assign new_new_n2722__ = ~\shift[6]  & ~new_new_n2721__;
  assign \result[59]  = ~new_new_n2718__ & ~new_new_n2722__;
  assign new_new_n2724__ = \shift[4]  & ~new_new_n2559__;
  assign new_new_n2725__ = ~\shift[4]  & ~new_new_n1986__;
  assign new_new_n2726__ = ~new_new_n2724__ & ~new_new_n2725__;
  assign new_new_n2727__ = \shift[6]  & ~new_new_n2726__;
  assign new_new_n2728__ = ~\shift[4]  & ~new_new_n1964__;
  assign new_new_n2729__ = \shift[4]  & ~new_new_n2565__;
  assign new_new_n2730__ = ~new_new_n2728__ & ~new_new_n2729__;
  assign new_new_n2731__ = ~\shift[6]  & ~new_new_n2730__;
  assign \result[60]  = ~new_new_n2727__ & ~new_new_n2731__;
  assign new_new_n2733__ = \shift[4]  & ~new_new_n2574__;
  assign new_new_n2734__ = ~\shift[4]  & ~new_new_n2041__;
  assign new_new_n2735__ = ~new_new_n2733__ & ~new_new_n2734__;
  assign new_new_n2736__ = ~\shift[6]  & ~new_new_n2735__;
  assign new_new_n2737__ = ~\shift[4]  & ~new_new_n2019__;
  assign new_new_n2738__ = \shift[4]  & ~new_new_n2580__;
  assign new_new_n2739__ = ~new_new_n2737__ & ~new_new_n2738__;
  assign new_new_n2740__ = \shift[6]  & ~new_new_n2739__;
  assign \result[61]  = new_new_n2736__ | new_new_n2740__;
  assign new_new_n2742__ = \shift[4]  & ~new_new_n2589__;
  assign new_new_n2743__ = ~\shift[4]  & ~new_new_n2076__;
  assign new_new_n2744__ = ~new_new_n2742__ & ~new_new_n2743__;
  assign new_new_n2745__ = \shift[6]  & ~new_new_n2744__;
  assign new_new_n2746__ = ~\shift[4]  & ~new_new_n2054__;
  assign new_new_n2747__ = \shift[4]  & ~new_new_n2595__;
  assign new_new_n2748__ = ~new_new_n2746__ & ~new_new_n2747__;
  assign new_new_n2749__ = ~\shift[6]  & ~new_new_n2748__;
  assign \result[62]  = ~new_new_n2745__ & ~new_new_n2749__;
  assign new_new_n2751__ = \shift[4]  & ~new_new_n2604__;
  assign new_new_n2752__ = ~\shift[4]  & ~new_new_n2121__;
  assign new_new_n2753__ = ~new_new_n2751__ & ~new_new_n2752__;
  assign new_new_n2754__ = \shift[6]  & ~new_new_n2753__;
  assign new_new_n2755__ = ~\shift[4]  & ~new_new_n2099__;
  assign new_new_n2756__ = \shift[4]  & ~new_new_n2610__;
  assign new_new_n2757__ = ~new_new_n2755__ & ~new_new_n2756__;
  assign new_new_n2758__ = ~\shift[6]  & ~new_new_n2757__;
  assign \result[63]  = ~new_new_n2754__ & ~new_new_n2758__;
  assign new_new_n2760__ = \shift[6]  & ~new_new_n642__;
  assign new_new_n2761__ = ~\shift[6]  & ~new_new_n452__;
  assign \result[64]  = ~new_new_n2760__ & ~new_new_n2761__;
  assign new_new_n2763__ = ~\shift[6]  & ~new_new_n927__;
  assign new_new_n2764__ = \shift[6]  & ~new_new_n785__;
  assign \result[65]  = new_new_n2763__ | new_new_n2764__;
  assign new_new_n2766__ = \shift[6]  & ~new_new_n1212__;
  assign new_new_n2767__ = ~\shift[6]  & ~new_new_n1070__;
  assign \result[66]  = ~new_new_n2766__ & ~new_new_n2767__;
  assign new_new_n2769__ = \shift[6]  & ~new_new_n1401__;
  assign new_new_n2770__ = ~\shift[6]  & ~new_new_n1307__;
  assign \result[67]  = ~new_new_n2769__ & ~new_new_n2770__;
  assign new_new_n2772__ = \shift[6]  & ~new_new_n1470__;
  assign new_new_n2773__ = ~\shift[6]  & ~new_new_n1436__;
  assign \result[68]  = ~new_new_n2772__ & ~new_new_n2773__;
  assign new_new_n2775__ = ~\shift[6]  & ~new_new_n1539__;
  assign new_new_n2776__ = \shift[6]  & ~new_new_n1505__;
  assign \result[69]  = new_new_n2775__ | new_new_n2776__;
  assign new_new_n2778__ = \shift[6]  & ~new_new_n1608__;
  assign new_new_n2779__ = ~\shift[6]  & ~new_new_n1574__;
  assign \result[70]  = ~new_new_n2778__ & ~new_new_n2779__;
  assign new_new_n2781__ = \shift[6]  & ~new_new_n1677__;
  assign new_new_n2782__ = ~\shift[6]  & ~new_new_n1643__;
  assign \result[71]  = ~new_new_n2781__ & ~new_new_n2782__;
  assign new_new_n2784__ = \shift[6]  & ~new_new_n1746__;
  assign new_new_n2785__ = ~\shift[6]  & ~new_new_n1712__;
  assign \result[72]  = ~new_new_n2784__ & ~new_new_n2785__;
  assign new_new_n2787__ = ~\shift[6]  & ~new_new_n1815__;
  assign new_new_n2788__ = \shift[6]  & ~new_new_n1781__;
  assign \result[73]  = new_new_n2787__ | new_new_n2788__;
  assign new_new_n2790__ = \shift[6]  & ~new_new_n1884__;
  assign new_new_n2791__ = ~\shift[6]  & ~new_new_n1850__;
  assign \result[74]  = ~new_new_n2790__ & ~new_new_n2791__;
  assign new_new_n2793__ = \shift[6]  & ~new_new_n1953__;
  assign new_new_n2794__ = ~\shift[6]  & ~new_new_n1919__;
  assign \result[75]  = ~new_new_n2793__ & ~new_new_n2794__;
  assign new_new_n2796__ = \shift[6]  & ~new_new_n1998__;
  assign new_new_n2797__ = ~\shift[6]  & ~new_new_n1976__;
  assign \result[76]  = ~new_new_n2796__ & ~new_new_n2797__;
  assign new_new_n2799__ = ~\shift[6]  & ~new_new_n2043__;
  assign new_new_n2800__ = \shift[6]  & ~new_new_n2021__;
  assign \result[77]  = new_new_n2799__ | new_new_n2800__;
  assign new_new_n2802__ = \shift[6]  & ~new_new_n2088__;
  assign new_new_n2803__ = ~\shift[6]  & ~new_new_n2066__;
  assign \result[78]  = ~new_new_n2802__ & ~new_new_n2803__;
  assign new_new_n2805__ = \shift[6]  & ~new_new_n2133__;
  assign new_new_n2806__ = ~\shift[6]  & ~new_new_n2111__;
  assign \result[79]  = ~new_new_n2805__ & ~new_new_n2806__;
  assign new_new_n2808__ = \shift[6]  & ~new_new_n2148__;
  assign new_new_n2809__ = ~\shift[6]  & ~new_new_n2141__;
  assign \result[80]  = ~new_new_n2808__ & ~new_new_n2809__;
  assign new_new_n2811__ = ~\shift[6]  & ~new_new_n2163__;
  assign new_new_n2812__ = \shift[6]  & ~new_new_n2156__;
  assign \result[81]  = new_new_n2811__ | new_new_n2812__;
  assign new_new_n2814__ = \shift[6]  & ~new_new_n2178__;
  assign new_new_n2815__ = ~\shift[6]  & ~new_new_n2171__;
  assign \result[82]  = ~new_new_n2814__ & ~new_new_n2815__;
  assign new_new_n2817__ = \shift[6]  & ~new_new_n2193__;
  assign new_new_n2818__ = ~\shift[6]  & ~new_new_n2186__;
  assign \result[83]  = ~new_new_n2817__ & ~new_new_n2818__;
  assign new_new_n2820__ = \shift[6]  & ~new_new_n2208__;
  assign new_new_n2821__ = ~\shift[6]  & ~new_new_n2201__;
  assign \result[84]  = ~new_new_n2820__ & ~new_new_n2821__;
  assign new_new_n2823__ = ~\shift[6]  & ~new_new_n2223__;
  assign new_new_n2824__ = \shift[6]  & ~new_new_n2216__;
  assign \result[85]  = new_new_n2823__ | new_new_n2824__;
  assign new_new_n2826__ = \shift[6]  & ~new_new_n2238__;
  assign new_new_n2827__ = ~\shift[6]  & ~new_new_n2231__;
  assign \result[86]  = ~new_new_n2826__ & ~new_new_n2827__;
  assign new_new_n2829__ = \shift[6]  & ~new_new_n2253__;
  assign new_new_n2830__ = ~\shift[6]  & ~new_new_n2246__;
  assign \result[87]  = ~new_new_n2829__ & ~new_new_n2830__;
  assign new_new_n2832__ = \shift[6]  & ~new_new_n2268__;
  assign new_new_n2833__ = ~\shift[6]  & ~new_new_n2261__;
  assign \result[88]  = ~new_new_n2832__ & ~new_new_n2833__;
  assign new_new_n2835__ = ~\shift[6]  & ~new_new_n2283__;
  assign new_new_n2836__ = \shift[6]  & ~new_new_n2276__;
  assign \result[89]  = new_new_n2835__ | new_new_n2836__;
  assign new_new_n2838__ = \shift[6]  & ~new_new_n2298__;
  assign new_new_n2839__ = ~\shift[6]  & ~new_new_n2291__;
  assign \result[90]  = ~new_new_n2838__ & ~new_new_n2839__;
  assign new_new_n2841__ = \shift[6]  & ~new_new_n2313__;
  assign new_new_n2842__ = ~\shift[6]  & ~new_new_n2306__;
  assign \result[91]  = ~new_new_n2841__ & ~new_new_n2842__;
  assign new_new_n2844__ = \shift[6]  & ~new_new_n2328__;
  assign new_new_n2845__ = ~\shift[6]  & ~new_new_n2321__;
  assign \result[92]  = ~new_new_n2844__ & ~new_new_n2845__;
  assign new_new_n2847__ = ~\shift[6]  & ~new_new_n2343__;
  assign new_new_n2848__ = \shift[6]  & ~new_new_n2336__;
  assign \result[93]  = new_new_n2847__ | new_new_n2848__;
  assign new_new_n2850__ = \shift[6]  & ~new_new_n2358__;
  assign new_new_n2851__ = ~\shift[6]  & ~new_new_n2351__;
  assign \result[94]  = ~new_new_n2850__ & ~new_new_n2851__;
  assign new_new_n2853__ = \shift[6]  & ~new_new_n2373__;
  assign new_new_n2854__ = ~\shift[6]  & ~new_new_n2366__;
  assign \result[95]  = ~new_new_n2853__ & ~new_new_n2854__;
  assign new_new_n2856__ = \shift[6]  & ~new_new_n2388__;
  assign new_new_n2857__ = ~\shift[6]  & ~new_new_n2381__;
  assign \result[96]  = ~new_new_n2856__ & ~new_new_n2857__;
  assign new_new_n2859__ = ~\shift[6]  & ~new_new_n2403__;
  assign new_new_n2860__ = \shift[6]  & ~new_new_n2396__;
  assign \result[97]  = new_new_n2859__ | new_new_n2860__;
  assign new_new_n2862__ = \shift[6]  & ~new_new_n2418__;
  assign new_new_n2863__ = ~\shift[6]  & ~new_new_n2411__;
  assign \result[98]  = ~new_new_n2862__ & ~new_new_n2863__;
  assign new_new_n2865__ = \shift[6]  & ~new_new_n2433__;
  assign new_new_n2866__ = ~\shift[6]  & ~new_new_n2426__;
  assign \result[99]  = ~new_new_n2865__ & ~new_new_n2866__;
  assign new_new_n2868__ = \shift[6]  & ~new_new_n2448__;
  assign new_new_n2869__ = ~\shift[6]  & ~new_new_n2441__;
  assign \result[100]  = ~new_new_n2868__ & ~new_new_n2869__;
  assign new_new_n2871__ = ~\shift[6]  & ~new_new_n2463__;
  assign new_new_n2872__ = \shift[6]  & ~new_new_n2456__;
  assign \result[101]  = new_new_n2871__ | new_new_n2872__;
  assign new_new_n2874__ = \shift[6]  & ~new_new_n2478__;
  assign new_new_n2875__ = ~\shift[6]  & ~new_new_n2471__;
  assign \result[102]  = ~new_new_n2874__ & ~new_new_n2875__;
  assign new_new_n2877__ = \shift[6]  & ~new_new_n2493__;
  assign new_new_n2878__ = ~\shift[6]  & ~new_new_n2486__;
  assign \result[103]  = ~new_new_n2877__ & ~new_new_n2878__;
  assign new_new_n2880__ = \shift[6]  & ~new_new_n2508__;
  assign new_new_n2881__ = ~\shift[6]  & ~new_new_n2501__;
  assign \result[104]  = ~new_new_n2880__ & ~new_new_n2881__;
  assign new_new_n2883__ = ~\shift[6]  & ~new_new_n2523__;
  assign new_new_n2884__ = \shift[6]  & ~new_new_n2516__;
  assign \result[105]  = new_new_n2883__ | new_new_n2884__;
  assign new_new_n2886__ = \shift[6]  & ~new_new_n2538__;
  assign new_new_n2887__ = ~\shift[6]  & ~new_new_n2531__;
  assign \result[106]  = ~new_new_n2886__ & ~new_new_n2887__;
  assign new_new_n2889__ = \shift[6]  & ~new_new_n2553__;
  assign new_new_n2890__ = ~\shift[6]  & ~new_new_n2546__;
  assign \result[107]  = ~new_new_n2889__ & ~new_new_n2890__;
  assign new_new_n2892__ = \shift[6]  & ~new_new_n2568__;
  assign new_new_n2893__ = ~\shift[6]  & ~new_new_n2561__;
  assign \result[108]  = ~new_new_n2892__ & ~new_new_n2893__;
  assign new_new_n2895__ = ~\shift[6]  & ~new_new_n2583__;
  assign new_new_n2896__ = \shift[6]  & ~new_new_n2576__;
  assign \result[109]  = new_new_n2895__ | new_new_n2896__;
  assign new_new_n2898__ = \shift[6]  & ~new_new_n2598__;
  assign new_new_n2899__ = ~\shift[6]  & ~new_new_n2591__;
  assign \result[110]  = ~new_new_n2898__ & ~new_new_n2899__;
  assign new_new_n2901__ = \shift[6]  & ~new_new_n2613__;
  assign new_new_n2902__ = ~\shift[6]  & ~new_new_n2606__;
  assign \result[111]  = ~new_new_n2901__ & ~new_new_n2902__;
  assign new_new_n2904__ = \shift[6]  & ~new_new_n2622__;
  assign new_new_n2905__ = ~\shift[6]  & ~new_new_n2618__;
  assign \result[112]  = ~new_new_n2904__ & ~new_new_n2905__;
  assign new_new_n2907__ = ~\shift[6]  & ~new_new_n2631__;
  assign new_new_n2908__ = \shift[6]  & ~new_new_n2627__;
  assign \result[113]  = new_new_n2907__ | new_new_n2908__;
  assign new_new_n2910__ = \shift[6]  & ~new_new_n2640__;
  assign new_new_n2911__ = ~\shift[6]  & ~new_new_n2636__;
  assign \result[114]  = ~new_new_n2910__ & ~new_new_n2911__;
  assign new_new_n2913__ = \shift[6]  & ~new_new_n2649__;
  assign new_new_n2914__ = ~\shift[6]  & ~new_new_n2645__;
  assign \result[115]  = ~new_new_n2913__ & ~new_new_n2914__;
  assign new_new_n2916__ = \shift[6]  & ~new_new_n2658__;
  assign new_new_n2917__ = ~\shift[6]  & ~new_new_n2654__;
  assign \result[116]  = ~new_new_n2916__ & ~new_new_n2917__;
  assign new_new_n2919__ = ~\shift[6]  & ~new_new_n2667__;
  assign new_new_n2920__ = \shift[6]  & ~new_new_n2663__;
  assign \result[117]  = new_new_n2919__ | new_new_n2920__;
  assign new_new_n2922__ = \shift[6]  & ~new_new_n2676__;
  assign new_new_n2923__ = ~\shift[6]  & ~new_new_n2672__;
  assign \result[118]  = ~new_new_n2922__ & ~new_new_n2923__;
  assign new_new_n2925__ = \shift[6]  & ~new_new_n2685__;
  assign new_new_n2926__ = ~\shift[6]  & ~new_new_n2681__;
  assign \result[119]  = ~new_new_n2925__ & ~new_new_n2926__;
  assign new_new_n2928__ = \shift[6]  & ~new_new_n2694__;
  assign new_new_n2929__ = ~\shift[6]  & ~new_new_n2690__;
  assign \result[120]  = ~new_new_n2928__ & ~new_new_n2929__;
  assign new_new_n2931__ = ~\shift[6]  & ~new_new_n2703__;
  assign new_new_n2932__ = \shift[6]  & ~new_new_n2699__;
  assign \result[121]  = new_new_n2931__ | new_new_n2932__;
  assign new_new_n2934__ = \shift[6]  & ~new_new_n2712__;
  assign new_new_n2935__ = ~\shift[6]  & ~new_new_n2708__;
  assign \result[122]  = ~new_new_n2934__ & ~new_new_n2935__;
  assign new_new_n2937__ = \shift[6]  & ~new_new_n2721__;
  assign new_new_n2938__ = ~\shift[6]  & ~new_new_n2717__;
  assign \result[123]  = ~new_new_n2937__ & ~new_new_n2938__;
  assign new_new_n2940__ = \shift[6]  & ~new_new_n2730__;
  assign new_new_n2941__ = ~\shift[6]  & ~new_new_n2726__;
  assign \result[124]  = ~new_new_n2940__ & ~new_new_n2941__;
  assign new_new_n2943__ = ~\shift[6]  & ~new_new_n2739__;
  assign new_new_n2944__ = \shift[6]  & ~new_new_n2735__;
  assign \result[125]  = new_new_n2943__ | new_new_n2944__;
  assign new_new_n2946__ = \shift[6]  & ~new_new_n2748__;
  assign new_new_n2947__ = ~\shift[6]  & ~new_new_n2744__;
  assign \result[126]  = ~new_new_n2946__ & ~new_new_n2947__;
  assign new_new_n2949__ = \shift[6]  & ~new_new_n2757__;
  assign new_new_n2950__ = ~\shift[6]  & ~new_new_n2753__;
  assign \result[127]  = ~new_new_n2949__ & ~new_new_n2950__;
endmodule


